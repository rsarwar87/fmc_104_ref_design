`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "XILINX"
`pragma protect encrypt_agent_info = "Xilinx Encryption Tool 2015"
`pragma protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`pragma protect key_block
Hh9mLrxAUJcIbXQpft7WyV47P9aViqoaS94GUQZBJMKIArARgBgQc1WFNWCsVxnWTpoRM4Q802VD
KHcn8rDNdQ==

`pragma protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-1", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
qW2mxZDr8+IjkBqgd6E1jQTj/H1HLIzxOoIVvUUx7vdIlmtataFUiII4JtuulWdxbcpTthe5+sJ5
VWF8NMqxnfP5oWAtXoV9HqP1gRHGHx2J+KUlW6DZ7GIU/WyqWs3qNQWXHxs7LTcVJVae7H1lmgRN
SBi80coo3C7mis9oxeQ=

`pragma protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
t4hz3Ob5qw0EXJS4gVKhwysffp6z2c7Ih85mnavXdlK6D503iiCd6rB4ze+hdNSttlhN8OtLFq44
wrFkilzS8VthRdI44iVz72YX52H2DcA6y9Yqu4zThZrXxdWqlDvevFx0MwbXSs0zyMyhVvmtOrPK
L2Pd6K4YIT0CB2nc7caRkaYgx7byc/MTJX85Q3R0SgpOjrsaMgWK/r+dSdMadTCosrZPdkdgy9eB
21xnY9YuXhFZmw6rRFBh28/VMNIEvNGx6bES/R8geeUbnGPNGod+VU/W4UpCDHQ82G5HZStN9MjI
O/roEuQsAfz1j+p5P6Z9ZG3QJGAquX8A2uwRSA==

`pragma protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
ps6cFpBLd+D5dON+Ptem3RLEOImhhkkhXBuAnjwn5nZ5oLTtAp22FCmw4Urq+uXxyv/xxqTaFfL8
BUNthoX5gipGphaR9SB9Yd+VFSqNPLtxUeJHyOi8KGGMd6P+126a9KGqTn9EKGyjbXdfu8wN+vNh
wiOwqbXy46T9jR01erhzQfw8uP5RLx0FU19GWONhgXhpdy/vVnBQvJDqzphOC0mrbDRaSfHpwgSy
cmo0Urq4QvOoXeAmRyBD0dUNRXJl3OYQ9jCsSGMHoDM2OXY7Ya+I1M1UxzvKmpzIM4u4HQrf4Nvd
vEpjCJYEdqly86zplVG78Upl1if0gYlfPE7OWw==

`pragma protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2017_05", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
Y3cOH7Z+DibqmubiJsOOQQjDdkakLXPknDx1DgseouUjaeVy/kn3bUDWCynRqkehtwUXxZv05Tym
4PkTlkz3Huxek39b28/vpDAszh1BqCjM2ZMB+sAOzpphihvxptW0q1G6TM3LdAeUbiRA01Hg0/4j
qyTePjJEYnq77hxSn1SFvocjy4dvbStbvAO0l2aiuqSitxMctlsCro6J0MjJCuZw9iIlAYvqqC/Z
ptKGJIU8oLtyoHYEblGvKwLDF35CuvbpBwiOCvq/pvi/8zeASIIxwyaVIAVEk0dQwiOXL8kMrZCQ
U8uYHcSJJEwyFSTqIBtaZNTrEeAQEMH0LRlJdw==

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`pragma protect key_block
lIEO9V+mMmOA3vniDmXxjOhUWLLhqWAhx/DmboPDf38dhnoR4b3igTC+cFc+reyYNTm1Dxo+p1cB
QvdxLGGDXwXhPHhAd9QMKUUnMABO18VAZGikoLBwlJH95VwPhudWnwFWcC4gu38gIEIjy9+pmsWD
iUzkZTtHsHtmg7cQuyA=

`pragma protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`pragma protect key_block
DJO2eFD4TbRVLdxCKXGkwvXrrkDDbe7jcSnV7Myqdd/QMMIxZMOL2apyMhk4gcKcPtHJy8zBb4Yh
NSAb4J6LBJdhMxZXOeHcniylZq4xX6k8zWW1N3qAZeBYRewNcP3j6zmToNwfBiqQ87So8C0qqYNW
uwEoHOtKpN2vwvvXsMiRHGeEHMBSwFzapolFGwKjLgiGmUCQzrB96Mu3wrbBsR9Fm87zx+reChel
2quaOyT63CPr80m4hsvEjgPPZv7XzF0bxu8XsqAnM9k3UsTx+JtAsaB9VlA8LWZVKPoRrJyZ0hTd
AVmPE7MNv/LRiSBeTmQA0kN3N8MCWX8K2kFwCg==

`pragma protect data_method = "AES128-CBC"
`pragma protect encoding = (enctype = "BASE64", line_length = 76, bytes = 2578496)
`pragma protect data_block
bYV8svsYLMrJ90pm+GgL6lzB8Cri3wA8yx20G0NvFvB4vL8rIlg7JOR/+6LgqYnHQs8HgpuWO8jR
QgxAmQLsQ7l98yX43cmvDjDDY+JZT7WIUEDN/C15CkiUU1YFdGxXI7gl41bwwS5wFPpzQDbhyq0m
i5mvyYKGqfAGmyyT0QA+kI9g3RN65CB+tiDj/0brfzqnoR1AyUpUIZQzqSlFQ298Y8H8Pc+4Cd3F
ClANOzj2NBw4zb6SAechRaAXJ30msUjdQN5vsomRjfdroi/JHHc8RAEImt9MAHZN68RPMQbfoQaW
btsX1rOBllGkNCU5bFt33Cg1FaUVz8kog1VRIt7zMBrpnUxZ3GRrn48TymB19rwDfwLtws3GqUQT
8fMV31p/dojWB10L07XMRWnni+4LWrfqrRusVoLbW3DU6SWh+Qq1wopiklSp9Vrww5ggv+NbhHk4
WEvO1sgbyhfmhN1uEttE/gN0ALCmTCccT57oo+EJvo58nSrPd2sFeHwvBeJuaw9qhOEwdLclDLxj
JDdFkOoJTOjgBDK+O2wF9n/ER5RbI9J7apCxJd9WQ62WlpETlpy6KOPW0MJd/PXWkjrFBwxMOYVD
fTktCHhCdgu2RYv1vkRwDUk+OtHlZoW8ToNCZGT5nSxBfVPgfMvYRx1tSyGvfZdThCe6xaSbv3pt
N74o+ce92cX8VgQQxTNKkXsgb4JRMNFfWC0oeuIAGUSrL5bJ37jCI8R3d5F8PxTU5qSk/0Ml8S1U
0tWt+M1IIE1aN1YFto5BzJvjY6y2D7p4ojiAX5jZmcei2La0Aw83RnrEPrSjy4Q5IL3vFXALg+Hg
sU/iWGwIcoVugFiatlKVTAuvaCnRo6taGLdVOnglhT5Lrj9ZpTdHoYaCN0PHhucKWchbxX1yS6DH
osw6z1N38R+O8/9WOez/etS1W/JCiR/oOWwbOe2b7h8KMTVWsELIyOe+sWCL+Y8m5x/H9F3NhPef
jar75k1XKx0fbAHzimvAp55XHw32AQ9lxLGSgZ0lQp9lF26Y/78LBdH0TWNdjnhPS2zsfNtUn4Is
HjpN+yi9QS65t7KLhAdlZ/1dy8eGjP1fiWU3phLcA+HglWBPd5ys8bTwRS7jLx/hdNvzDIiLQuwj
k9wPnjKgUiK65LIEkwwTmz+RDQr6tWN5KJS3pkL2++cyqPDnAArur1E838Dz6FBw8EJUKtCBIgCk
U++cQpXCqYPZT2Pwf0f78wLaZ+9dvv5vih/QD+TvWrc2gacVCm6Wx0cRXT9eycFuih9Gm2CwOtwr
XYnhuHgjIMOAteiEE+cVPIhBBiJyEV46eMaj/vZTKSSKz78JintmVdaf5j/5vH+lBHjg7YAkLWvi
N4kUT2rQo1QcIcCpCcvD5J1vn5tG5mq+LA1fdaWUfZ9MYydb2Q1t3Fc94/IchCZ+Xe6AdBQNCx3P
uKcQ/X/9X+D4m0veb39UYG1RD1oohU3/GfblYldVAtV4DyuueFGJ0zmHXNlJZ8oLd1BlppxWx/Mu
xPay1aJzFQYpMP+EA3wYUehugtbPUyItQ8PZpdpS13I99TeoxynRTkAK00G6OunIlZAj3b7K7neB
9cP1kZ4JfmIebyt+MBkQFh9Dli1+ofk4RUxT74oXnktRcLlkTKGotWTOlNjGRQugrR9OS9OsYQrM
dHWzat4SUGfpVeC0JqBlKF4PdVxbL8Zo5ISv6lDPAcIBL3iH90XFkxYbzJ6x8kELlMqlYo5HH9ac
ymGwXhLG9RK/2mzQ0JDSuY8OHdQ9vuBf4oFbiBvJAP2rJ/8jP/rr6qoJ7D9MHbWIXRn04guGGKqx
CZaaakDikjx1EvFtCjZWsatAJMHVtZVoiPfMhNevSjSg4IA8ZZ82KC+769qWY3Z1Gw56O/OTj7Nt
54kPeLlZtB9Rj6kpp7RJSlOyULslkt3ntnVbT7VJAQdE9oeKYQkEnQ8gPLfdQOmXzHnKv38XS/d9
9aH3zlleL2TYAcOlvr24WzmbY3F8dCLmz8XBw+0IKvvLeX29pzcJiuguaAmsI4ic0d+x8E1Xj4pL
eneR7iccxT/t4uZmOwjogrcN4VdilFTTiu8M8CxuKC1U4Jbx5rd0oosSD8H2EhWOx/iUl8Utub7A
No9eqABv1712FZElACiNtsbzeNHOBD+j8Q2LuJpatmcEUBJrfIE2+5L8CDrGoBkcr45ds26wAgyt
tvsYpb7eS/1FTK130rOdHxTGEvbG95CY1jkGgOoyrSBwMmWvoA8k69MZPNHX1P+LXB9huomh8bN4
FG/Fpv7AqoyBaM96AW9tPdCKXOFImGiLwXQmzZQYuecXwT3hxz9+CPBEfQakMsWlc3TIBhj5mzaE
oG2wOaqff+dOupDK/Zi4A+4tY3Efe31Hc/EgY1IZbAFnRt1Kis0Pb30uMEShOPUpBgPhZzwCc7AX
KxsUUxcy2YZ7a1DoftHCmME9EArZ5fgJU7cICLJA3pG1gJd14SRHp15kBqG+rjnbafm9O1JwvC/T
aVnPesKUpjzWVuy/yV6E388Q5HMqnOx5BM0A3zqFC2IA4YZKtPWcESuco1Ur3jl7kK7yi1XMnwoh
dbHmDGN0QkLkfShViSovxY9A6RzEf7R4J2OovhzQijOXzPHpOOEwHVUqAy7nW8VXGLbN43aVW6Ei
n0+7eWRtp/nrmpgb6uO51AF0AzWRCTFwR+OJYRzraLzUMdXDKYcKFFmtLS3gl39rT3qhccaFDU1F
cCVdrQF5lkJRFHXeg4sYZxXDob/aZ5clbNva56oMN97ubqc7+hlmdjvHeZbdfy7wGvKy76nqEC7G
QREmjb1Kwq86ZHP4IwXtXrPPdE1UfDUP6nVHw0/SyEcClwLvOEyiuTi07x/v9f9K+QNkflayiMwV
11uQQX7y6OacriMomrHbriRKJWqJrcHI1TZuKiq5c92hNrhCwWRwR3Ay7RieLwEy/MLTX0gxfvYb
GNMpP6GZuyvr6nCoPe7cUjz2/tw2YHvyjRehfsRp0h8A89lzF6bJ2jQXsXdnXiBbjRkQoJNJoiP2
3UWPEijJRbtVnMnUmkuosA7hZmHtlA+DPpZTIeifGks6PfqxXT0ZaUR2MBaL7TzNkWBC3Iu3SArb
paP0+4fbATMZdqv9ZTPsgTp9gvIBtKuqfFT+E6te9/2dnCVcjSiURyoEDljYmZce7kyeT+2s1Qsn
JTKkDElorjJrdh66HQxfFQ5k74XndE9qNXrMY2rKB52ydAeTFyBwYf3WNaLAUlUowtMa29yUuZM+
KPEm1AxN+QLodS7vFW2GXmwmvNUq5sBHWy8pQciqsMKVpoYjTawV9Y0G05Gq2xyFDx9grJMeRp/7
ArqP2WHY+Yed8C66ILl/2V9k79MWv3ll2c8/MxWMgIjvBnNM3ra2WZ/Bohl4ZI5v2V2oU11WEDeR
o9D8sN5AJSaP99WHJkOJGCg/NfZBJsCioKlNUV9+899+SQSKxteJ4xjpWL2QdfL0vqewZjILAFv9
aJMq9EYJnU3BWXPVxMpAwOtHUSoaGsChxB7CEz0CQ/a8OBK8kXzLWBtbkrMAlwMGAdPCd2MxJ3PR
ADXgeIwxFXRRGZQG51Unhyq8siDaz66L7Km2Xx95er6QFOUAAhGJLcz/KCWLKjKu+fKbsPKX7BYG
cmEgfPO1gXBlFcxYgyxSR9Vmp6MNYz+JvXeiB5x/ctdW5zCilnA3Z82n6wPUSLlrLLJMgvVmnQIC
02uXUv0DPc3CDdh4kopwQkoN4th90vUPRBlre/wGTPXfKgRpZEhQFx+vN7C84wn7ngL3V8KRbCjr
j9LvcO9hcU9aqNVhYaZMtF+hK4wczcLk4yY50at1miiXIZ5fh9FG4V/dPc0+Hy0dQ/SFYJl6Sp7w
L6k6D61WEj8YFIL8KkiE6cPWnZcsW55Um3T9f2qKkYNWvc3pUzKlPfHr1laAFgeKc550U6OdA8DJ
3AQYO1SU1+x2APMo997nBmNz8Mxw+cAh6XIE8exPHBi2ebejLjvTJOnPoderQTYEOSnjrzdChT34
5TjUnrxuvz/aVhwSmkeHvIN0ihhzAelFOnKBAI+XHa0ibJVDyEu+3tmTak+f+x+Y9smuit0N0Pxt
1osohRJEEF9AtNu2u9D50JncmiCvMoNTy0jiTLd9YOQoFMpgLGizszGsthPCl4ndDQU8bAvIfYQx
UNaQJDsL11MykhErfK3c9rxE7PIPDCIRwnFlVOyXvUADOCeTUHvNs9hSzRlyIQVOx9eJde+vUQXw
1T8KD7GzbCeS2RlsHAJ1h6Cg+EXD+X/WpkTlo5Wi2C5D8Zh/Oe5EclNWJ3kSW6V/DY315dA6A+5B
rnNPwKsMs8fs+5AgEtTqXN+9qv1cKmTyLzYF8eYdXcX85etDclSZkVWFqFhGIGCbdFr4Afn6wEWX
ajGCgpm2SeDZcPgyqEcgShkZabR/lonNxVOz7+2ECqN54ZnDM4eXOk7TRfymuXGwmZruh1R67wMH
Jl+LLFi6MMDCb4+n+EVRfXQPqtY4u1JsBUqrs4/BqnkZtJz9ZSShYyLfeFAUxotJLOS8llK2Y5su
LW/gbW2SbIG0doe340M98L6Cfe4asa+gfOvfAQuVTQdSV9+sjldzSlDx+dD9PuMBzf0+Z3nHDF/4
sle7cIpwP5kjBOP+JDQjxg2gnO11/GOHLQw36oNhgHNXWHyCTE/bh2WbZWX6cWNYMKr9CBEv90zf
PfkdZB4hgFCUIZeTiMsULvN72K0zYCmE4v8Co6VjBTTZDkeNfXjnItHe8FkPdHhYFGeodbFH0zUp
S/ZkB+AfW17Q5kyAp605CcKm5K0ClgyUejAsyEex7hDEezjT/IqzqCwgtBqesi8+lKhz2WZ45+NQ
DR7fCfzx2WPCX2Ypz8FsxbbGZRIslmjLkkwNVgbc2qR4RrIEXXDTVrrn43CLy/7o/KG+Zjfxg3ES
tlAtF3Dp3rEYINri8TnpEvjDvMhnILDJ8EYSO2y8RvHLCYLt6rDFS8Uhn4qIxn6T0f4KCC4I8eZq
Eow2R1Be/VKcoq353YV9F8wDo5Yh0vybLstR4HGgoy0eqwqvv/qOParglTvGdCzS+dgYo+NsKdyb
Z/b8Ux2+Ll5Q0d9mpaeA9nT+jl3XTzpRLml1qjgONmNwTFCnFOlFN8gfPyYuXBO/2cxuuXqHNfj0
GeSwvz7jURds8gp/D7g4JAIqCrXVf47NcCqxSlBW7JPnP4bTvYkOZPwJQeLRexE+E1BjT/HNRlzA
BmNpwTsVYC9oTBtNxHcvQ68yMFNJElTUR/YfRa/InADPktZRVNNbsj8MULf+tCDL7TO72SoOmjzS
F5O9drnDxxEvPcvJva/l5GuWp2oagZ2cGpQUc+ZU3NKH1wgLzLB0DyNpXBErd915rAiAMLHmSKTo
7GKyqfJlIV3J0cvr8aAVddtNrJ9Ll5Q27W/amSq7TqH6yVAyV4e1hV5ccgadXCDTOdyQSGou/EGn
Dkb63/+1fOrbDq+o/nKenVcRiC2fteeVAGS+hRIoQ7bBBYbeH0qcMUSRRzJEt44rRfFVTnNZZQ/L
2nOUwO0lYbFDbGNNtkKELhGHyy0nMCdorZ8vTrUrr4PYyyUWtLi1ZzFRuTuzEXqJa9P1x6ri82eA
ZIFiIl1lROm1ABXmp02G4+Rk/TkA8pafYYjJtkIDq+jkdXerLiQiBKMa4z+tRq37JMm4yo2RwT3s
z1gsnOMkOsYy7m9w0p3p5CY+/Fcr51XiqVNgzbLf31Fj8Ex67JHvQUZ4jNJBz3O+wABE41iyQzAc
4ElGCUdsOzAT8SiG5lwQUZQzo7sHnrNaCs0fvAt3hbvslKm4Zu7SNheR3S79L71qzwPY3IKsHngM
nwYD/StjJHnodolMr43drOrsQKSyQy+yNll/wqGzUdAi6beyERnQlCpwJZW36/9JiJTdFvVUpM5h
IC7a7/ucGXSpIw5w+pqfaCfHSG4tYN+zUK7/Q60l0cq9MZj5JJDe6LATjhLJx/x108eMpdSkcgCT
2d4QBmPOsjuWQgiVW85oaaWz1loG9mNtFp8DKoFjg2YYaKeZWSF9R4qh/SpFroudK6aulfCUKD6E
2pYYBiayZpi8G1mJju8jwSCF29RIVMn8uNnJL5Q+8ppKjPsy/Dln21FLRX/V7GmYqO08ElqOOgMC
EO9HuXC6e9S7sIFw3+GalegEhg4wHSOe93k8JKCCoTdCMEx/ZaSIM4aZuVOf2bvMHdPE68opNT4K
Jp5wBBG7D2y8vw5qbGwC753WXrFaHrXzpg1dxt4A4JQf1K+DuzbwksijPH5KyB7AjOzWQXi8uWme
he1+TpgE9zifeypOm1uY4Hj3xJQFHUOesvSRUF7vdQh9t/LUKrE7FC3cMDRGcg85pS7Q+JPXTsnm
jl6Ywv7BHuTMiEs2/76SNwgLjiUSpKibXZQ0BqNZc1q3r5Vy/HOjoWlulkrc8oG+TeWI8VY7nIGQ
F3rTHU7YcG8sEqZFsaEbna0Y8usUrqw/HBITmuSBlNezJcwkOV0IHfyuw+HIzL1IDQSBE7yY8+of
wBxrvdftOLxadVJr3aKBobWsUVepU9WCFdjwSnRtqn/fq6G+jhNpmp4VwfB0iyJByeLMn5zGVL0e
2W4eMPvrVzvaIBXbVAu0ReNAQYeCKp2LIbdvdpfb1LZR6+YoBinARZr6pkyJtYJUmJ+HPy2qrqHf
LAJ8wJtIrQ2Hq28cvnjxBj29LgWoTWNUZPAKBuBsCDWRTza+9y9NH9ui5ho9UTmOj1MHxQiVUwia
3VAPbpJ5xbvSfq+0uVM6VXBG+yVgiFMN3LcDwN3ME7zQGheP8UupWIwSWVaX7v5u53mG7DGNxD7J
ErAsUMD564r9HjffSMRq8uUUWUqkoU5W6f90bBgOd5YzPOEYARzqDQbI31GxGqvPJCZJ6aoRQT/3
glETEV+rzo+pkv3T6jOKv8UhmJTlzTaM5ChcM6zvMuOeqDjIA6gz1GD+3YzC1EkgvrEKLX0fewvV
i08ryx+pDE/yCvX1rgtxxvhXxGSSM0Mnh4P+tC/QkzZ75RSz4jcxEoYn1qwgF2BGCyyQBFGe/Apa
8c2EKj1EBXrof/AQc6pn8gPxOEK+jFF/OF6w8NNUFN3CQ8Ha/BlcNY4/HhUKVOjIjnaDuAJlTv+T
s595NE+wr0sttTr5X9VsvlHAhSfN6vnvu2SvrbjiDylUhiTTycMHIz8ReaYbHCiqakrdqiXpPybV
jtPL08ynrwK1yCjW5Og1fSsDwr8o1fkYXhxhoKEiE5jU2IUSKpkUXZEnRVS8Eyq4whfL5Q39+fRm
nVE6OjVwebbJstWbpkOGk+bz3FEymT74KoMvnpp747YzT24lzR+3D6O693fV1imw8Ot9AS0a7pM5
nJ7EE2mvBQOxPVGLVnNIQddBBhQ0bT0u1mieMmgigM5/iYMWGBBGTtY0uM/AsBUCaQty1neas+/8
4dcE4O1tc5RGi08JBNcuvMMdRH7f/saIdRZAc5Dv10s4fbke1a5h6SQ1NEfW5x/nzQ1yaM3P62JA
1rA12C24Xso5oY14QwCf/0kjp9ZoEYTSJfGnPD0rHb1hqfUtYG51PiFRYXdsoQcYjj6AukJQg4Zl
s5C9r69fINDKsMy2YfJ4buiNryBfPmMLeav5zaKIW7I3mxbAwn5Yo7J40fN4VaLfCGpKNXqhAyxO
oqgoGyZQFKu0UiSxwGPprWZby0eZX2AfDHZjfiTctX3oiytnboYpOxUTXGnTO3kEUn58r/zn7L3K
N9rKLQkH7OXl5omp8kY0nT4OsfnYY/yHLGnjSlMSO+PR+7uf8SwQxPljjUm4hAPTjj+ShpIuwpwG
OXTvk0Tc35uKCdwKkvv4990zPQEF98tpi8kV9RYB0BRqcQU2b2WJscC4qf7bsSazTXsKdLpfV1uw
o6qHwwn1ISs7gX1CN5tBgspl1FQSHCzg6Btayan1uLZe3MTjhknJVQct76hF42H3v5+e4fpgQPq6
shhp0KRrEV6EAMOjFYLBJJWnx/ENEYjbXKHxheZmn6bjGNSAWTaUUGsKkFYvT9beA4w8msPngJBK
Hb0bpXgspVYzCbchALZ7uotLIKFBeG9onYhIxr7c0VBGPmIqWUtjG4pIUxizgzaN3TJuhLjN3370
tZeMXzIiTooYQ2zhL7MvJBEaP1/lvITvhSSLmVnVXKCzGTTmsegRKCpcI5ihZiOiBI/n8tdCA8fA
idfmcTBCtI7IA2R4C8JuJy8tUZwfSMNjm61e9rwPLbdk8RRZgRR40Cz/GRearMkIx/B1R70Fxl5r
xIlApYBkwKJjsnSoqGCjbvAmmGcSVEjYpo9E770saTo+zPtJVY6z7dhbsBGrWxl9/xabT8c7zxNJ
7adXyiE3cRyu8E3cGPPrT5XkdT7w/K/pAnsugaEjvVBSxI7qoTOltSo3PAUSv3IP48wNA8bgH7b6
kA2gyj1jNN79uAg1T18xjlMVYcO+Y8G+9EHAtY1Yw9kQNC4XnJZ+IJJv0EEQD4jrtd1gFvMYnK3j
me2+BEbGm5Y0yptrgxYmMOtt34VMuZL/hBgUJ8O0AEo8qZfmGUe0YDNiI3MOO3A0cF523uNvw/0n
A2jH6kOmWtuvm++4GDG+Bu1+KJLOpBNsXXCt3Q8IcV5U9AMCNvSqE3xvZ25xsa3UoUIRo/5qdV+j
P2RW+aXjtExzpiKh6LI9VaoO0j08QpbPSyEsR2bzF266MU3xYEL/r8jddVOems+6TLmv+vtCsQK8
yuAHDQt5saqiL1pNPoi9MzcB972JyX1CW5saQ0N/3o0kc7ab4SRkwqaAOBKMp6MDuJ2dakOlvGic
xpkeFLJnjJZVdAragIV80+eSDaciabEFpmIKFA6uwbsBJ52X7BjRHV/PG1+TMLv/7NSM45YddaSv
CbFLCAD7FWbYOQfAwjFOGMkytYyBm3+4HGgpfiA9qtOOdhymz7eqks0blr1k3RMwVXY7BBR5ogbI
4WU6Eoo4zQAnAE/Q1Z2QcoCg/qUmVqhGkbroz7+sS4H6tvD3jVc+mmIhVBMnaF8/+tihXctzJGqc
JKuHHVuB+mii2dnVbtbO5ITTSNRZTCHiNUe9WUb/4+90ohyEaHIgFLSvx0C/ysJzn4ngh2nVBiAu
zt3uXQwZ46sCqJiWNuP0259nvriZdMkEJz4Zqw/qe1mCKfZIo9cJxlPF/oY0Q3qRw3cLiPNlcRFe
REevXzLzu6OBX2LTS4rKm4h0x5MwYKdESMF7KEmM1nSTFZwaCr4FgQAalusYtsWkBccowixnbQoN
/uM/ST/Ha7o1UI/nk/7WHUKk27zU927B5VtRBYEbEciJo14q/kUewp0fiE6jthoWZYo4Zqf6ENF3
H72tSsV7MaGhK1m094jEgtKU/TxAXVawTrtPPmO2+gH/utsoo9x/gkyqOh4ldFQXKQi1mv/hZAn+
OEiMDpv+WrDdV+9StGA0qWi/2sLVHBBZa4qXAVovD7yYrWrtYLurXN7GrpNsZngLmk1TDntAx9Io
xfA0wpO6QW5qilG+Ejp0NnCs7avzqtZRlbB7AycN6pb7A1lbWRU2p/cBWzjCbgGUEkrO8hVOj5tZ
Tjv9XuSQDnf/91yjUpINiiYO2eJUaqozdGeiZv8Dzt5o1rICMXdSThOh8bFP4xxnLWEfxV/Vfwf4
heoPzQUudzEVDK+Ua2o9sRaJUhuKw7f4TkZv3W5uR/yOQfDK29/OPnvZpnm0WpuNNKRsvh7Btm40
dcfh2BSrHSwUAGKxMG4ojsV0B1IERnOI2+yOV400kz45MOuihLfDOoraRsHGqqGewIBFqP0gHZo2
78Jh8X0Y9DdHO167G5Zm3mh0E8T4VwLcxny6FzGyKY4Y2eOSJSjM3JNQHAXh4UMgYPqfUHXtaXWR
IYNirQPyU6loTDp4/GNl34nITRrly4a2ol33fqE2usNMvGefjyEltS/3K7Nyhjf7goz7hmuVc2uu
Szi7ozE0+Jxi/CPdR2gU1gcSbJB4a1HPIZnXgTe7YoVu26pnjSrKAuUvNfNh/OofgGGvfmF9CmAL
0iPzF31/VB2kvKfyLhMg086Y/fzUywGr+lAyYp1BxjW2e5E5Cflyn0VDfL29fo92YK7vSv9dvF+9
4xY7iTDIve4qlMENABX/m7x5BPQoff3W5tEX+OvJfYrUZe1p/XHqm3MxFQCnG4Ek7wWD7c9gZ+LO
rbYHqFRrqe6Hxz/XCyxysMHw36a9dcMQOtLd8/u0vWV2f6CBo7m+uUnbcPpE9N0/X5sR/HhlvjxD
u5/mm2FeaVFyQS64Du+kt82D9EXVak2d2L7jRs+3MG4HzPB/sgMDFE1vHrRqPgH17pubZ7MkJmo2
wYMWNfEgOLNQ19IrZYIf25zYrCNnRR2gYAzppuJ7/78OW1wylaG0/KyqYZRuMPRs6QA4S6MBsXZ9
hdOrT0RDBmyPHgyQkGezbsDOQJ5AsJHBf4i/0kMLE/bYDr5AWMLkdszj1vSK7LOB7aMzTkZfpxeg
s6jLUhPkfjuXcz6bYkATq6Q1Jys06tQbl/zIOmcla6PMxjV/KiaWyhkMxps6Ayok0gYL6dBIex3d
05qdJjHudr1xcCbXeJQR1cpCeZgqsjwlbSb4/OGiqoCV6cpROrKiTdI/hm51VqrSqK2zmk3UPfj9
/rJ/3TaHhuGvoXR9ld4RaiOCCbJ/d9G8BCYD9De5SR/aPUnbY/eQGB3Z571AVwp3PW8uKXmae0Kd
tukzkfG5trlLgEp4lbJ0hmZUMQ/rZsl563QpnmDHo+PA7N6kMIMwm6ycO8vvaYgE9TiH/b+vbFCR
unmgo9DvQnJNrtRI5SzQOtjzpG2BkCDCAg588ZdvslU3ICSGyyYKchjie4UpkSBEYXI/KsnB9tcc
3XcNB1j7HKKKv0egb0llHjhtpZPV9YfMkb7bgna2TQM3Dn1UQSOdqFArK98TVtazEgaRxaGiijOj
mq7A9yB9a8sFhoWKFbZvkRQH4j40Z/uHVhaBb3jtAVTWc+/XYfuY6bQHxpXYBWZg8h+KPFI5ASow
aTpVpWYKolDPIyvR5mqKBR3zUnKDhYCK50/er87GFuuqbbcXkuzIhPTvvjDQhLKpgFNWfklTyMf4
xLI/LgEmEC91MWRAFuM3hbaeTNZu4CrkBRMQplsNN4HJZBo8QSU5s/vBDyMmjAZd/5Lsg4/+pcsD
4m796kyjEINHUl8hwklnXdfA7fT6mpGUbUCI+WkmI0806PC24eS9xePS04TJAe0dtDLFpIO1TK2k
EsgFIqudE7wtl1PqKE4p9JtY1aIePZ1pYINWikDKrnfYa2aFQjYpTReRrm/G/36PCHpFuNlpWy3p
ycMvlfNxlBZVsKrX/PtTQ/eeygmjqVPNiHuIT4aSRBbzy9CCjRiw3sJ2ksRue7QHjoncu4spz0W0
gom3yP3rioUk6+7jOciPgNKombUGNW2dlyP+9YXlfDBi04aCKWQUtpY7VXr/Sen7h/LBTp+58gpr
iz4dgDwyKJ9AnFUctD9Mb//YmhDOnN9czshJM3weuz26/FwJc1PDgPjip0Je77w03mnL8frVGc9b
yVEzzCJBFtXzmL8MpykujRoyCxK8YU6IQDPQI0JxQzXsDoEiZYyj33sP/8/ycZ0dYSJSTerHfQpT
TVodlkIJB/H4P3JmztFdJ7OIsa1Soq980VAQLz9CEQq/0v+MzkdyeOlcTnHuKYfwizqBB7uyq8Qr
8qTBgubQ5+lsT8VsBQ/fI+NZgdRY+3lKPn2DP2vNjdGX+Ws0ahXWvI9Jq42osk23HHoITCzABd25
UARDGFZ7zTU1zxe9W/V9bUSklAf+FTruVvWInnhB80k3nAcsYO1L/S4eWoLdLDTY1eqEGXWy/ofH
dUAoOBWIndiciw1GVdVLyOyKbG5VTHY5V7BL+SzKIclNZA4agin9KtnRkO9o84FsXQszUJqBqn4/
ShhYSjJIENGP5kBdNy0F8Ipjr5UxixI6m3I7SC09zz+4j9M2iQwGd2PWLUJpSQoj6+5vF4FTVADV
DbSDwoBdiJVio3Vk0WIaA6bY/2wj/HEap+T4qsMHcrZHp4jbay5je+5SpheCcQNQ04LA9UR3WQFW
FWEGGSBJRt1vp4x/+ouaqPOoXNVuonOZHgKlQ44PUQQxa1NXEr5nghMDdm3d3hF3gIoG/zrHQiyC
+7xNhjT2yXpRaMqfToKhkOPUU5SF7sA3WiOSQfDuNW7pxgZgeoOLikjKL007bn/fizSMFfjDDk2U
1qEdVauJhDjROYVZZXeEj3X/RkzBeP6xUenhwfxC7tJ7zOTGA/I8CJq05sbEvoyqgRvBueLGrnqW
2vkIeRFEsmuZrFZGPLRdzfU+DheuIfqFSECIFJ9nRA6C5uciTq4iruPbiqhx4C5x1vPk7w4p+P1z
mKfTN+42WQ7QIzKsLnDCLVT2qsVNWupXWntPqXcoYaZqTdHCb0aTZK9JJNlRv8ers3993koNunBF
j/1lDfzkio3rqyH4e7HBt/Z8REToNtuumy74pOu0jjW6LiSMblnklIt7XBe3PunfWhzezD7BokFq
xgPAZHle8yWAHzbw68BvQaFtY+4yBfUMgPHGj6G/S5gkCNxAGUwwucXhEuCo/MgYtM+NmQ+2n6Id
dQPFulsXBComIr46cYF1/ah6kMFARdFZRuA2Cz9ILMoCQleNA/pz4JKOqfYxJw+qvupve+8l7zLl
P+tEFG7HXxY1SZXqkiwgUymz09EosgGV5yxGChy2lkYp/4Y7JrrUFWAbJXkqPynTF/alOYmxDsYT
IG4YTVJKPjOR5F14YbjsDiV2yXaYu2e9nQ7xNg8E6DhZ2bsB8wq4OdeHu2MkhTajRgwXSpqfsedP
MhpCIPlfX5pH8pQcaqY8cPHtbrJWLyRJh/LnvV2/ou122fVCs0N1MLNkPKfl+d10Jj329lMFYQWg
h0fJ8TDg0LiMxaxm5Jz4zJA6FIExRFhrE2v6ZmYGydc0c1y8F0JPwCZpEcFbiJzJL8P5ek3iVCNP
b3c9xgEa4OSZUymWaYIazevXzfpiMxD3FaR1FkS87U/tvn7KYRJyDDdWpfCDPnz+ZuNZxOGm4taD
W0lng2NBnl+R9HkDx1Nvlg9kaXY9hycThiDHnk1Jq9Ylt2KkKCTXtEM8x6iGlnOtvagKCuTiOt6T
CN2+w+y+Sit4ILvCGOZVykiPHa0bDabvhibjwOwBfnFGnLA8VrS8NIXkAqAe9Uz8YgBRVpG8IsFt
IJLfleoC6Fovdaqx6RcKpeES6Tdlji5gIrguL6GIg5x1ojaDsA1YSGEzsD5cDowQ50OFW2zDwrkj
U4n0jw96v5w+pSVYy4F9V5IxIS3n9mGizXQiMb4yIGD0W5r78xUsgPzkqj7kzXsz8Ki8RXQ1izwP
5l6fVa2PJfI6YncHUfZNSH/c0Tw/ZPN9Vy9ckzv4d/tEEUOPz04tyyyjCxKlCP7SnK+iVEzk72FV
orn2NP9Ikn8nFeOKaZkC+uot1wp1AIJW8dP2oWlvbY7XG5piSf3jm9TimhCYlnYCrPc9zxQLgx37
mm/wmGXmaAFiEy2KrlYM0ut8Xrj1bfrZ4Aq3uE9qW+PZ9B6hjgXC0ap559koI5qQmQ+IjDuIPURj
nP3rTsJgj7GYmLlXBxvPVx/CsO0wGylei/wn2b9SZUgV2ym3+HHM6UUrUqDlxDtdodGeAxVF8bZJ
K6mhMMRFE2HoX1D+wtcjDxHmj8J0/FZLvuRGENby4eV0pXAf6Cp+7PRxVzQAwnmJ/83mf6OSW7bD
/A3cSz+d6Bcp4isXdbNkSuPlsQF8kUNShEmFMen/ZRQgnaknuGKej9nJhhliWyXTeQRV1tBHj+Zs
sJclpQNW0ldg7na1nk8phsWTXKuhwJVnAdyb1UK6hPn1PUleWAvP4rcHh+nLWIEeZvwdCPXdhDqT
x0vhzTiSMzBrzrMTRhiTsz7ppNfeD3phk4GhCWjbfDNsHkGeZdaEDgpxeOOnz0Jkv/wvG36YoeYU
0jDY1snmGyXq91cA4FOBn5GLpTHOEnBWYCBwGNYa9fRAoFl6UCeiHdITVY3sG/6qpXNnYXGvNlIx
7b3NthF4urLQe0Lba0YB9moMMO/vIUsAEWolcof4rMK4YUx7wCITI/nkfeSh9gZu2KcvGN83jh7c
0TrE7C1LNxrMdLx0RatAFSsZct3Wp2mgnSLIyi+Li+yv8SeG/dszQldKsSNn/yl1xll4jAtybqH7
yhc99+mCVRJuSc7zbTHomdd4lMB2W6Ws29WF7mNj3jAlUifZ86zSjyN5WZghtyUbJmpihIlqHZOD
bHolsBEX+S6swxB99CktbLtNCGARU5Udh7jp6Y8uhb0SmVzTCDzyoGUkEfHowAeWW2l2nKKLRTL9
odXP6qlolvdW4pKVBQIvt0TPdxnVyNb2WeG0vXDeBtlVGtZjc5Nip+Ca23BLkVmdTjLjPN3QjtzS
VUuAP3yxeNX1QmcF7HCgEq45Ok03ghtDgDPKAuxa9XAgQQrYa7S6i7u22Gi/ZoOsCDb2kchNS+yE
ulVkdLbE4MjRoKtfvCpQGY1pHw6hY1Jgtvj2qmu9jDaLWU5sJzYh6WLp3Yz1cuQYKb81/deo3S4B
hXw82WsN01wzmHxLJ0c7aIPUKdv5CG8dRixvVovS41SoiWGYP1XDP71bdsM3yfp6fKqPMbAl5CVB
lOrdyVBLLg7v5hefTCKljz7oW2Qx2DffIxdFyOOGN/kLoFY/Z+Hic0QJy1cxHHrrxAvMy9h+nw7P
Jhlmg2LmaPWzqtVMdH7OiGVjJ/Ty86fVL1bKENIC91U5pTiOij7zuzbbZFPn5F0p4nu1xi17Lo7G
eRiTihefc1FebTUSok82VFG5lThyOZJ993l5NUDHkVUhqOAgzbHv6JGu87JTDriT5yzHzR73FCsW
A98ydjHNNB7CphHG9AdR4dOVXqKvVNSJ3BjZ1u4TryBq5+4BmIHjMIWzY7gh32YMRslA/RNFosKw
qzgw+fyMO0PZa58Wd60cX1hhRWGeJ5Z4yxdYKZO1Rcwgjhvb5WMtJytyDY+wldMFGh3pO2JNtlLn
LjmDfL3Nh4svci201p8xbO0Z9plxqr/p6EHDXZb+sLx301ClrEYIm3a+wYVw2Mssc7rPq2nEzD4I
sygSm5R75Et5tmeiuyrD6VBAkcinyvbH4fcn4JSLRaiggHma+ViirCBhhjlpPFVPswiLrt+LiNKW
TRkTeUm1O9WYtXn6caOEm49XhzUM88PWTWWRWfK/ARENulXUn+WtAd7C7dy5YJ8Pd3DvgO756pD8
RqgzrRd+F/1nFyObMvRwYzzKDEcgVE6ysMbxQ6qlv54Of+BOfPdKtNvgvZwm9YbDrjKg2iuGS2cH
RGl+EQ2/cmHZrRHvgC7K9gIwgxxgg+KNZ2o3rI+tIyolPpXCfWcRmzMIk79escM0BFmXZFpSFlrf
Rnkt7rDwk3ASEZXjZZ2AuTuClKxPKXSIGvkxmQKimLCWGREgW1mACW0M9Rv9lxytOs3boDnrD9pS
GyPraJQnnfjjLNdR6luR3fWrjljGaaQ8HRsgFV7Wa7FVb19VT39UCa6S8qVqoD2rvKDPutgYiKwc
t/b1ok3vx2OUl3bwv/V26//AItMswb4nLcfhX/rstNreDKYijAMYZU97ptXpzTX9xgyL83mINb9o
mKQJ00maPenI0eAaBjetJJSKAXWbmuI4Ula04ds+2XiOf9wWkkjF19iSQLyCML8jCPUc7bjrg36j
yDAcgBld8f1eMH54Fa4fV8AuAgo5p8loLmBLhfaVW3BRmdn9TOCzI7iG8z4EdVrOINO2mUoEGfWZ
1zAqECgf22vbWkwROHH3xyIiomoomPivaznHh1u0diBRvdqjNgk4ggKW5Sqomx4wbJ960OWZ1DoO
L6Y2RTawJt1zPYOExrnRF5Tsh5/OTUPUy58b6nSPPIafTTzRMVbZzMeyMQ7pb1dsn/Z938DURFmi
OzmTZfO+rU2U8z75eGGT5qvhBSy4tgXIRh3JbDXAcCT9lo3Sd1EXQJLLh2N4om/KlFtvWmvgs2fD
ueMyXTVA4zDztb1Jbbp1uaYw0GHBmh2wOCdYFNIJLP5zGLDi4yUL4xSQcIEMMG3e/ft3wt3jTcqL
IWsSKQPhupQHanlWhICG4g9QWflOhGLatm2Rauv5EKL3OqUvJuxi3hh8w4lwJXkMFrWVdyObrkPz
YxJKkFWEsPfH+IzA6KV1UbnqnXsxqGRbtvhRRXQqOlNVNa38KKEC1h+BiBeTG2NIl6xWxrL/PLtg
F9A6rKjVLHNLE6C4x5RqLkANoV/dF9P6T2nRjidW9Y3CURMweYmUr2xCW2VggxWMBWjdGzluUtJH
tM0ouySrf5UMY559yGtbDqxYUgXdmuJO3ClnCzJ7iBh/stWmiDNUtRn6ipNl+i+lplveVvPro0Sr
LS2giMh9JJXvbEdz3RhhyXIU5kzco+nzsLaorMJBDbjQFcXUL5dzzy9/Z70EodD9wcE6G/z2lxSK
rnrD+TJ+/6SOk4oP6KOjmrgQnYzvyOjX4h9jwGs1Oxzx9x4/aoiWSPmEdTRmgoAxjTMWdVp8Dc14
JpFU365bZiHXRmrP5LkOzrlD2luUdaLd9hxO07H5jrrENLamRyyOYHLswkEKhgZPH47I4NEVOzaJ
tRJwlwVp4fmRcpux5F2Bp7CYuopcV1cEP3AEeaLtpvmZyNDWaoC2HqaW2P36DZypEcxPt5MT2CKB
sGioGtVTNACw0VpXVADVsqVQa/sRhJD9c+1O1Fl+TxP/7Oyhef9J6glsVRmp/27TBnSVapZAtgyo
5nq375+LyfEPQqxgxHO0fgwBvzrSItLdih85gAG8XUrgUMkVNCX8jIALfXE2sHICCT4IvzjWTxyQ
hbRSky72fym3wFo94kXrT6nR+RUHNWSUuICaFzwfV78otzRJNs3Hh4V+OD1FzARja/0GzpopbSED
bL9PL5s8bHvWWReMuI8DWfLdrfGmp0BqQrmDdOMm/Y3/Q7Euvua4DcIqT++Ws7qHX5MVa14x6ETO
EfRViqnuaqy/5mkQWGEpO3wORx+Fips94p49T6deStF2kzYQ6fOt7AHo79rDb+wYiR2FYcgUk6Ur
Hn+LPmBlklhmNjrUA05J4vbnb5fNDu81RqEkh/J+6nq9CY3OFN6QI7iZR0VP6shmyVadouZttxFU
fvrqqMKkdNrlvwTJb6F2t4J1yLpKkNEHjWZU7ffdx2AQHY/m9vuUsNpuFjMu4++nd72ZiapHwCYL
bcVPYSaqDEjmx4+4wgI8kCh7iZfN8kTlqKo6VBLt8Op/y5fyVLbCMuq7pzy+RsCV2qhmqWUcPRn0
OtptdREXBMJ0wvR68v9+5wZiiHXWug06fvL6SSX3kTSNeKUUq00S5VaZTVHkJ2woulLcTKC+SmA8
20eWAq5Qj3FtkLe1leRdrE8pcrmd7OinLTpV1QGbVIP2GbNSXiVqLMD7pH33D+nwh3WI2N5VoneX
z79Py9fcLuFr4KGsHb6vqibyy004/CmIL5kNof9a97rExfENOeledPZ8zqJaO81J15jxbwJiDVch
5gvhKgNHyAq9XV62cScY+4FeVOfjJj49NZ+0Xt6o3rAH2ETXTn4la30zAIZeOUpGn6srWMs0dn2D
vfuL4lc7DvelxIXWCZ/fxxBoscN2X9/iysHZ4lSlsUrZPInjVKkKLFfA+x3RiO79SpBAh2yQRuo3
SaWbjsbFfFaHLKxVNrLPYGyy/J49y1UOWL4ZR3FSCmrgdNTCQbtpmJLvDEf2Lvlyd+WS4CJPAGl/
d+3SZ/WpPz2CzmgHBfwg3kmWaT8W9HBC/ZF9W/VCeBxByjaGdieQSijSUBCFhjwsKoyA9OwYW5I+
KsQS/NtgQZxzFk+OVGWSSiPHqcgMUUDuVfvvcRBV2ofSINOiAYSq+aWh59AVHCDeOEeSeIGevQ/l
ZlCZeBAvYD7ByfJnHnxdPoNde5cru+L7/grV8MWdDzB2Hg+srexHN//q23tTEU1q1pIB8Wu8GWQ8
GjXnm+V3bp8KtcCSJVPvv9D8Zmu/dlyM2RctYp+5Xasm+A4I17Z8TU4uufGL4AJFukq20Ds5zwB1
gryzdEU3SnrmtaDmXCP0fNu7uGOxL6XXcyPA0xb1POJjPI+Qut6sA+b8/MQGgzm1I9VMfAARLnxX
Aun/zUMnCa0G0HY2fyy0LpOTwOXNIuESHZFg16evsrHeDPwj5QNfFccm+6EngdeCZZ8RsGe+OpvY
5IqvFwu2lfXwuuAC6Hab2CuaSlVI6QwQIGSk5hETZnF1TpVr8+e+KbtZNlhIVz4vxyhf292rouI3
MBSX4WJT+4QuFHT//JDqlCqrKKt2AexEHKPeD8wc5/R+L3VFMGk+/CABwC0kcwaP8MXFQB01jiIJ
jpM9Z3iVqcYl6wH2jTAQHx7ytRvBFLFKwAUCExvZcIq56S6WQgZIOhYur81CNvtO1i5tOBBBAgWT
iD65pRQBc6xlaKCIMZ0TFjdZy6KCmTNaO6v0EeB/bRt49nkoC5J++Z3YD4iyK7Rprzl0ifjLaS3p
K9jzM08fdV1zN86M6jf2fdTaC4A7mREBmNqlFI9q7JSXQ/ApPh90My84J3S02swzatwkGg0TJ+ez
7Bo+5WnY5OlCduecNlzRyDhQn59JZm1W6+lOITPXnqCyD2OR1SYxH9H3f5XN068f5aV+aN1ZoC74
TDsCAksUqvHpQBNtkx0buwUuKFX7eiAsegU4Mgj23Gm52koQxzPTV1sp8+ASnu59aqYlgzBq7a07
YJprSXYTMagRgUbLh5cYqB3gw2T8G8s3FIez79VTkO4YgWLKXeTO54y/RDfL2oHlLDOywnfkdXHs
Qqsek7YIUb8fbxG1f6aDAGdNhL6Irjp6yrsxHKR6D/kR40ZevRrJkhfM2lgooApQ3W0l7i4vrl2N
WMI5U8nVhOHVZ+omi5qRWAJt7k/pa9McBJ7oNrOICMYoxlk+9ZWwamBBSHWL1mmeZWU8172EJcq/
smV8hwa6d+jfFW4ksj9B+b+HV0jyoo0QYVHS3mJgOPsSnPTcq1Weg7UgX+Z7oD/30di1lRx9t1iG
izhKQnyTyGrGnpi7v2QkUoZ0If3mvXecvu3BxwFHzMV1RS+uVv1APBMp3GJv7BQk0fhUnHOqtlU8
o14NCv4k84aPr0t+RXIIemUveMkkw5g4WRBLKzG+oxyAceBlAp4uNKua0rHzfm4Y/GnVoaXP991D
ylqodcXrSbgb6ldqkmFj3HoIipaYBJw7tfqp2AA69jbydJf11u3IGE6uxhavfVWcaT+95SkuDT86
jDdBmfEVHvQXU3Y840HLYzQscnXljku3bOZcFjEmRymXb9lPZBHB5/A3Wa2ImFxiqHXY+jc8TU6R
Lrwp9Lv1wFjzRdeMZmxjvqblmqSUeChZ0gBxxWMMLzNQgewLaJvNsa6t4B2kRo+oD+eFmFsvws2V
eihGhX3P3+CWuKMhAXQ3oWKbBObB7qakN3VHCaI42NaE5nM2Th2zKn2lH282X/QbRlHmWZCUEOZ0
er1kOHfoygZJ0KWZmWy24gK0XjO7mRS3+oOfPIsVLkXnxSxva/3XAAlQqbxbMn/AmkS7z2rlBy40
AQEaXxP0Z1d7KwcGeEnEGHk+y3E2AxgGyP4NFxrepEoA8Mb/BXn50DDD9FnqbVVrd9SL9J52KnOt
MKV8SKYRgNo2Hmc7oAiavmKN/Zf+2s2erh20c1S0cHIDhhvXa/JYPNMoMWkdzH9F8khEqOjP7Pky
R6xBBNdvJiIbzKAxSFab65l5Q79DFRzmIdm0WFT7ZkFXmo+XG9EVDLvXhscjfctiJ8dsiEaYblCK
KT+D5zRdzIu+sxkGYps8lmx5kJZzLzvCOrF+9OXPNrLFhJUjNVudY24B8BN7XHmFwh1GtTBwWbPf
MN15k79ROtHLRJOAYay0I4WhudUPN/x2BqH7AP5bOYaKt0b2vObyMNyLFcYvfkJ2GXCju1WcnibA
L5mXnAeX6W2XySEJw7ukBQ1Gca/fO65pNA2KBAu3yH40WlhTHnmFDLETL2UkAsTMMfv3YOvRbuYJ
ubOQ0a2btFp6QtaAb8eUEK9fv6/UZZ+4WHv/XcJNb09Tx/rPtiVySr9PrC+CptGubRrCIOmd6x67
r8dK29a/UiD1+RmdWg44IljdJqSWPjgCNVWVPQUx6tegGrixcAW4QBaB5VqXcnQG6xXBmFazF7iH
TMsXeW9pQQa4ao8neVTG7BV5pJw7GeLwgmm6oklJ9CjfCeQy7YJa2hjSmkCuiYdY8snrd4KPP301
b0urs1z7SSGVBJ4WD0cLQDGRHqItPVTy0frQqMUbxW+9GHbFusp4U0rfpqKnTfczwEvf+aEAls0g
DVzS6irVgnUJ2dQmq6M4dcEXaosw703qwVBsafce6CMbmA86gJfCoJVXGuIplLYRw9R7TrS/WGNH
i87ifNDINORr9XbsIP3YlWwJWYHidm9rbaNCaXdnVVIelpXmyFLEGzOG3+3Ow8ZTEHpG5CXNml1N
sGaYz9r81NQFPOaATFJAqB/9OwMfe4jhCsWlp/HZIhmkJ1rj38fkEtBhq/NZzH5AzREVVRAxiAF5
9mbmpRXhpWu9n/FHuJnRHrjN7AL7tbVq3K+RjEy4Id59LnhiA8H53z+3W5Tvsobd5WDLVbuJybuJ
LodYV51pNOk0Lqi7urfj+N949gCjhbh7qT/ZdELtqwXQPS5YJfzEKU5OCs5bGMFLs8arfzUm+GX0
0NRRwSMxdHjVRjeRaG7U2FweW0R2252un2QqQofUWbDuaW+39iQMRf0r1O4+9DQX0eEhHedfECQO
Dk82pzjH49wHavxETF+6y25Y/A2e0LCSYxBlY/67Qn5r7kraIJKUjiJiIDF1dDB1Cjwl1Rwe1tm4
0GarvclwEUXZz4bGD1LFsrL8nkowqF6rhkOtM3RqECAwq1YA0XHeWnGfS4lhjhaq1UDtrm2W32NX
UQ8ALQ2qaSbBOi2Olr3lORNecDNV7aJ/CqNB8rMSQM8oX6JxKNqNnhNmr8DUfPWwWG9klMwqyQqi
qCTt5+mGJTTtxKiGBmi5JfCi4iMnPlkHJDzM0812tKAqdwEb/d1nfoMCRhPYMAl5NKJDHTmvMMLE
CDKRl5fwcHcxrMFNzHVjj20L9iPpwfoV0skH8VqY/geWpsYj+rtnry208aNhBjih7b/kjFP1oUv1
lnym+xJPN5+v+2xLHAjXTl+B4aGMUysL3JsOtTUAwykGc8XGZXslU92vXKETn+PDXsth8Z8EDUX7
dxjETopmQ8KZGaz+c1OnNSmAHF581bkxQASR11i3P3zi4ylsxJFvDES7nOgLbvBUiJPcUQDqXWqT
CsWiPZgspcyb5XWAH2ATLu7KjBeUttps0ceVe0FssoPLI5jYAXCqZwmwxvz4AfnbVF5IDXrxYhCT
hXu+BccVlP7ShYEUQu60e0SGleeT7KNizjMSrwvF1ZUnuYPDrVjozVwKxfZkxMhjppQb/oZQLuaF
WmK2ccq1PMamj1FiziifrvUEfAOSgJCDnegxQt7rJXS81GuWG0uUPN7i92jcruLhsCX9Yv3bSP5h
TSad7sjnm5z6pL94icJO9sWkwB6mytrhOR2ZDEcP6zRlZQnbdYmQiXSVDjbHpsuoFBXV69QEN+bW
d8NREt+C03qUe/jKc3UmFJeHy5Xc7NA6He9SbMLdOAlBLlnPNvUGLwNkwv0J5DrIGBEMoFvljxnK
KwKjKahleGXNlgUnb4rgoAAftDeEiCNMML0x47rdYJ+LsW4M9yHnQNvMOr1q6td72nXGPNB/dspa
VempZ2mAzFboYA4FO/Hgn5m79inrmNdj1O8LjHqs8Pt2sOOnbglVmCaUXpTF/HPx/YJXr2bRa6PQ
j6xzKNSeyiCZ+gVbRHDqoYxDogHFtP5JMRo0NPp3btQig+8GFthpYid8DqxWCeDSHPsA+4Z/KpE0
sjHzZsfC+4MS//BYFThmzQ7Vft5aTpZU/dESJNTsDswXZlGfkEpTky/3vJNKjunep53byR/T+q2E
CdQWuwRqGo3angpCniqNuNvqNHLThxX1795+x8DpM1B3zpuLTh2CAj6uWGD1HqG9MJQb0+3jgkuT
QMbLVJ//eHSr9vT6tfxmL3ljLHSRap5aL2jNpUBiKmlOz+1AusGU043mXvVf9QhTuHcAkLAxBuIP
dvpftgEoS/fZXhfqBQfrup26X4HtxvddGHRruyuJvWhObTyLVwcLO/uqrvD6JR+NG/cPbkGZmuaL
6vsq1PUZZOUwN9UGQLoTPtHfeB5AeaEOOrklQ7lwu9l7Eg9qdE1X6Hnv9Y0eVbD2ljc/6InE36vJ
sIcpfe23WSd0NzfTvGbKzmw09cSt+tI0bVaTZMi6Vw3kaP/T5QsyFlzEleoooyF5LvLoFJ7JTu4Q
jyc1Ug3QmPxRv26osInZl+qk+mmKk2aXmIo4R2zdnjC5F/IhtSB4tC9EaUsVr1PoS/eJEjF6QPGQ
PVRiXG85s7wnWHejLMdQ65MjNGCt6mOMbkNaQ1JZkiyboObzegKtG8DXk/EM5P+QD76N/DcEBUgO
kGiBQdqHKw3QLwXrMjHr39jsy9ZlRDGlXlW7GVO6H9dNBmGpPP6AzTx2BLz4vfv/elGO4e38ntVf
zNwrLPsbCtWBF2lYUQd4RWQW6503ELpUVSNIlSGyo4dx/O7vEd12bUuvOcj2e3xEgsU1HszZn55y
ypZhOQYfrjF3ofDIPz3/X19Zvww0eTtAI5a3V+u+VxRhGlozlLmsbQtaVbKVxkar0/xdz12H55Zr
AfskMgConkeXM8GlBPg7b6D1tFtvM0TmRH+AsYp2DL+ptq6SZ6a1IRWqmaBDPaAoPCRHF++smmpY
kxNHttlY5sFjP72bqxnTMng3kHSy7pth92PomYgw3VWjsUYZsHks/gHkEV3Ya9+UI6wq3DZeY/h8
XXucK+09wHnQnWFce0Yvbh6x5UftV0Ur3MEjaNtPtu20nqpMhlyVe3M+zG0bncj6Cxtv0cOXkYis
o/pcpWN4LcWBUST8cidWZuR4fi56/hzoN9ugHkRryRwkbl6jQYfq7voTqUgwofVnbxTpRGC1b7ei
MN9gYBVNI2EeWgpREPE4qWt5diOEv4KWKE0NGkWGJ5LbHqfvqlXu5+5IgRNUpVczFWt4dVHVuMu8
kxlO9leol09haXAsWsO147K0vzd392u0KCQhls2vDl3pwWPaWPl5326cUHkja5RTvAFsEAqChAug
zOgJLVvareJf0cA0+KyrDOPhzWWS6wI+Dxox1mw+vZP9ZusZusHAZea2GY79J3tlE/dEm8TIxIkA
ol66eAUt0vAZEx91VBNGl+jLcScHs0BgZk86+fKRXTfpUgEFNE/aa2lQngDbxDqiwWhscaaIfUeF
dOMLwAsFTc4JB70VNXwu2JN1s/KDwMVf2ykMr6OPWFv+FTOtU8eSHhsNcPEGPZei0l/rjj4RLIpW
V+I20VcijebTjekEa5I4H17sJwQ1z1l70PHzfX0FEvouufptJ4j582cHbaWYjicpoHgK8TNGm5Z0
MTWZIC/sQvrZeOg31pCQXLmeqS08plPObynDTvFkBb9RQZM6qYIFz/wP307GUyq8qZtc1jN/dyVN
HSi9J6Vo5ebAg1CC3HSD86AW7Vdaghx8ti/XzV0KrYi20paGKaNnvOMdJiOjWTkxV+QlT45nrahT
LL4IEQqjyWq2chCGpmIa5+q3eRbh4wqHT2HivIW8pUH9a/eKOTEnLPgMfbIu49sFqvRfYbOjD788
2jHLmWjVcvjNCaTvgLA1F715q86c35uMjD/lQaxNPDHFrcg7DNHIuApbfT6WxfSpnNjf3eds5NzA
Z2uUe7988xbeyymnG9QHx1dAWLT9IK+7uciAx81OBRhaw+twEQ9Bsiw9dYFPCm7yHMC3rT5jVDsH
wqxpFIzCwCiPMAL4q2Myhjl45oUvgW5Kz392oNuuAxlKkDJqIpzIRa4+8ETuR2Q4Yk32kp2LgjxA
NTjNQw3/R+URQCivw7IEirrO8bOZ7+jzA71uR5EfCoI2Fp1FhZ2ruC48GPvDV8Wjs/nbAjaUn76X
QPbqMWqnVvcyoGrKpxXn2KHNjpUzMgJNV/H7lvxfdbV5DSRlEKjEsaNMchmuelu/Rq1NAXrOoMJZ
r0Ddp+8AZiC5yJJgoswEDZ4JS15YuOO/H9MXRrxGFXQzQWCgGMa8/Lqs3D7ap1y0c7AKtV1H9yi6
YxngHEewbLJ2hOgfhQzwtPK5P7g1qlHG07rdwjbFDW1kaaQNGsNuFV7b5VtLTADNgzM+HRkgV+I2
mEHS67XTO9B2lshE579WW8gWGcwO2zjOcGsSV8ewm53o8Vimlq8DtRptyzqInDiYDdLC53SxWjMb
ht8OH9xLEKtaajT5tdFszXzfB5F2KRPQvUXjcXjADC2HsKcDN9j+INNwGGMpoXGQ3SI3MUBiOdd1
Z9qzUCd7gDqtj4Z5Vw5RRCvQ8Jhk7+GWrL1GRJDhI15e68wnLcn/rvF4oOVoUTUtCGSAX3QJihuY
ErARe3mu2LQL/Cicg9zoBYmGFF5Cs8/MSDnQ06pFgQ/ixAhKCO+XjgQ7ZtxP+g5EUwG6Y5UBcZh2
z7dEM8yr8oie1ycAApVwaWPQRclgNXouNvsETYRPGC8avYMdvYzoPuEHSaRzU5eKi42otkCQ5bSu
Fq8W0UayxfMEw3O+c8CBxaP01sqO5JgyTmBU0fXdAyPjbmDsrp10dFflM5PdT9n5YWkzgPYYVR0a
YpWbsvDRGBrUaNURGvzB2jDTEZaL3o6mDow23LIzczOfDLSSkVlAahrpJM41mOKyHB2rwiCfgAWW
Wwcf/n+HgGGr+GEUBVkGl0+vpX/vS1eIP6hje+IiqaX7UUdqENN08eSbeN6PxWc5ERCeBmhjl+fS
eW7MPUMvMLXqYsieklUMSDAA6Pq+GsVq/jzg0FqHCnyEXna4x4ZMJUyyuZxCOvH7mQvVXmNVS/CV
dWROwS7OaArGb3h7r8jC6sS++3Livq/y574vuREyCWm72W4xn/QxW59FabWWW12GwW/3J/JxTQE5
jdmVlgAJRjNtHHcTxorvV5AUNSgyJJ6MsFXo0jR5qlUJhHhFPyuAG4s/S9WIEYA+EaQUwSnI2RmV
Kkj0cAduDUkxrVxgHpKHDGi2+xEKuHiVet8c8kMv68gr9Gpmw7suyeUhX+RHRjlEVRppK7Y18sZI
3x3ijdJN/QtcWVxOEGTaYD7qFUyNGFXxvryBoSUdG/guR35Hcoh4BZ9DvialAv3fr/QjgkDQDyXc
Vs8mNEIqRY65RjgHpa+WtPDIBGV72J31xOqzVwLeXMrG7MO9yhkcvD7ATWJ3xHF3MUUELUGGvkdI
tl1OpZXxBGuUaRgdPSZAMoXb5/K012t+bbj1QVjkcZoIZFksJyJLVrO48Y0dxaGp3YRwegFHfjKL
XfbmjVXQq+1lYv1OTWnO/5kNJZpW7PmpQxBecAkgoYieqCNUE1Clg7/OPCdFF75CXDNfCRLFtlCq
iNdWlHH4FDxIxJ9+M9ZRXVyBN8v6JZluRBPidnU7bx9v0BUbkB2dRUh2byLhVWJW8jeAas6dG7Kd
6jlL+DVbhkmsXoAibgy/XN8JbKU0J8IAcoTqgCRg4UCeWS14p+hTyLt0tvCf2pmYNVegX0rKUAlN
eUjn2Lumu4Ip5dW7H9mpJVLuJHqJLpUvh/PuBxkH+ev87keeQSbv/Zlj6OzXf72Vc+BKYJv6KCCe
mrvEAHUjYHNZTWcRWpbRPaEmzLFGCfvCLfRwmF6xJsLKEV4CUkMA+LDc67P00guAmN/XsL0L+F3+
GtOXhDOdKPrNksicUPohTMFh9jxABZFQcmTvjRjNHT1hGXQL25gSP+t1Wf4+/Vp2q/zIGThPO3ht
kvtskUrOwprJr3SBUGIV9yO7K+hi/kGm5AyyplB12JVeb/mhZDou7HB55kjC7ubjEJOGSJyNztWM
ctqMlq/nTcTh4LP0I7D038gZdG7n4B6hAwOw0EJSVpMFeaSCYQHQ5EazCkWM+3qs6EL3hWUL+fGH
p+YXM4IBKW2/eyNUMeOZdA+vufNxDFVVfQ1qf35Jz0D5woknO4SORXeW0osv1YRZMuRUbiYr1k9n
uZxpVTlQ+a17zW5qqFb0pB5bF3S1pZWZKexRf8bQR9v6Jzcto8emg0dJ+Mdqx2EjavIbAu/D7g6K
lu1QeSH1g65/rg/dJbyWdaQ2tm1gKIqZPHI/I8rMBahgvki77YrXxDfqfbJCsUCR4KNTTkWxS0X4
ERXp/N+TKQiU1osqjRRpUEgKEqgixV0arm3pcoae97ygDCttj48DzSWBhlY3iGX7o2yjNyDc+c2D
aQamcuystTZDHlqPBMPQM6VQcLL4KhfnaEPJD4KL+bq7xb/F7rm+kpkBwIhLGswzApAjXdH1bUeS
kOPgAS4MxoZf1bzoMYOsN/SaVEepzd6fy4THnphlNDhn4d9LAqDIKzNqZaElvJTjNicLNoHK6xAO
MBVO5TESG+ExpNoKXGIkkjnZa41qGpSC3+wN0hU3mxYEottMELEWOsC7ryoAq05KvA1OuZy/Mtr1
L5B+5JtXVuzOGNuQSAfm4220V3kBF0vjZ+/s+HXFupO3j2MVDPnRSoGuLm7XnbvUNYmVA5dofz7Z
AFtiAuUreNu0mPh+SvAdWBRUzyviZjTavuU+tOPGG22Edk7STktUKRxDu+jURHXYEBY3Frb+BbPo
Z+3cmw/AuKUCkYRnF373kkcp0ZKwBkpCE5Wt75rkQFot0I1AfluU5B0SbzHbPZ6joWwXThZUhdpE
X+yRs/yeUXpHkHYQiyhKLYmhiKTs1PZnAK1JmAc/WPiMaQfOiqxq9PZL8OW4vI/NXdVn5NIJZc1b
3JLICmixU7yIWv0GM2v22LrRqZCbqszpBrGeeWTiDnAElBoO0ghzMXSWopbz/SkDpornn+6u8MH1
dBhX3eu4vuDy5EIc2YuxuvEbpvPRKWyWDnM6V5z98qJrLMyYz/sgI8AqE+kjLMArK1guTWN5FaJZ
mjdJCT49w+/YEBdNgFdwngKhnYPfOgDldmQv2t6SO6PXMDpDtWrOGOiEfs9Cngz4/tyszWjNDMsj
rS7MPnWyTHoZFZxAU4+qBxE2ErOzXbEsD8AppNIb3dmaBCSf8So2MzM6dv/gKj6vcnbWIaQvI8wF
59kqSaRc6SYU9mR4lxSm29HRbzr8OTyS4g+w9qWy6pDLZT6RjNr55z8ovFlJzkzWcFUTlZUd02Sm
7g1B1u3imJApeOukAuQo2g/YJn2luSG8knUAgcq1RtG9dVGXvUHClsxOmvTwL0Kce+0AlnfqM8/m
s4cIpBhvfByUol/bYs+6VCN9vbeMAvoAe1zJ9CAR2lvNdH0f3bQHreqrNRhSvXNsz5C1775XQKZK
uwu0eRwV1m2Y54XtpqKC4ai+rEWSJckdsLGEhrZym8uspPOGoybdqeiMMP6mVCnUSyxHkYQ0TklE
beNq36Y4SxMaO1lGN+hlwtwufg2zK9r4Or94pfooy3gajSK2UM1bXB9pY/i367nSgogYSQjt+W2V
Fz4GFR3pEtrCIyqrtzIjjBaZPLtB2APsKlxs+ZvlClB0AOXERhWeQPKPbaxk6ZqPh6pcadcZcSn0
CKIWqwLVwj14f8r44rWggxFlPRb3JJ+6HnwDRDQXXA4ZIfwUgM9aLLnu2zxAM1XpvVFcEuf7KU/V
tPGFzrL/Go6yBYXTgGQvgOWGKdw2Xb7F6BjF3lFCQRwUpH0muHVvtETNjnR5QoUSo02tsIzHHpal
+ZgedHATd+OvGP7RuHfehyHEvJZMAfyF1HTnINFP5oPTPUk9KLBIPQL9vP1M7sBsKKgngdelj3cw
7GGJxCyFdL6hK6xZcWZfmd244t8EEDl8SUdoiCRv96wE68Y/4fYrtbalJcXIBDnIDkBwc0aHojUX
+Fyr2dxm2Kt2LyILeX9X5b99pvxlfdr7pJwnzIA3F8BUHnwAeWHIChtxAoE67hTh/BAn7pGS6K+s
ZBuJcqRBvFiGnLNNH+NSlmKhNkd9u4BWe9xnem1c2wQLOBuD4+TELWjv3c0O45bgbRF2m4pXyZfD
hAv8SJ+5eNH0HwVnJ72uqMYRW24Alk/p44ldif+UILAn/N2HyOZIR+UARdlRV2kzDKAL4sm1R8VD
M5aSXENO9kKhNUBpN9rmSOo82NEj87SFou4wY2DXNR9fks9hmMxGoGdDiTzYNWmkCLuc86Saa0k3
2I+hFiObW22Tu70EOFkR6/EcznVQ1bzYJ5BgLnEcc5luvphzTxb4GrlY77q3dnadX1qSQwQtbm9+
m9vXdlc1X1cgrlTpox2UrD6b6rgRBmbPvz3bcwvE6ddWznGJCryTFjXTVip9ZHK8NB/f4n4toIIM
evSHi101Syt9V13jRFpxo/N+zxLFXU/sk2fuHNSsE0qkmcvm6nNHRu31tE7rJvqywUSqsmNAM8Ra
JINs7/HkI+6Hrj2fn+ckTIvjRxD29IDKAgS5if9OPBItQt49sT3PBBkHIYud+MIak30HgQkRPJ1f
VADGpsjx0fuozOyIB31VEbhtPccet4wbikJWOeeaHJWLOQvRlRkdNJKTvM83p1FOo8OUJ1Y4Z0FZ
HzyV9X/YXuWSmeUuO8Ua9GLUW98ik8nnwOAe6WM2NWgw1V2t2S0OHB3SAaDIMFHVZ56nHirPosyK
XLgpc8kR7+wOEX3w8V+HJwGPDBW1sVfWG0oK4cCDO0xkIQVnzztF6lfFkNJLRnvc+yyMjMno/bqv
er7bV+ZGrTiZTaI0/GY+HPOLvqS3hjL+55X27JouWHDB8gGIHI6yoq25ctctvL538R3xZOzWGUig
aNIc0zaDmdCixHLiot403O2ZmuOQtaQysiu4ES1ionRLpsXMk2dvxJv5oxXy82zboCtSBCA+pScW
fPZg+OWHBM5B39iJV7PmHyjm4t7hqBN8HltHuNwDpXneg9Or2IjuiYLVhxtCIZPhX+LEWH+pNQTJ
1u2hRSduc+/EvKoK1KYi+leCG6NzLI1tWOplrjHvSqvdbSyfR7IuLcqy7FfxQQB5zS6FJA4pygMi
K2s3JhuCPOYbHBbt693Nh/qudh6IpfdGizp71PPrLEJLHfWHTOqcHbaWjTwew/po8PhIyf3PHV/B
SQEBCF6tqcbNNQoqWNV5PHmZIQRaqxGLyDBkGlNIxhO/Io5lxw/pOogMzkJPBzW62eLYlQuwwonB
bZ3xtzuz5xxF2742qdCM+ddVFgmTmaeVaHnmn98OryYpATf09MxVzVP0yVX5ILtnyNBXq8Pw7Kn9
msrhpnrIZ8wbpQk76mRgiXwEVxJaCYlMVf41kymaccwFO/lYpTmQVaxnLnP8ZNdT4GJdSARg7Z5y
2s6O+kSHxURXUQ7vvuKYgeyJz5fvU3n3mDVqykdfDCWClTSxn6W14wWy4w55PUMhq0/viK6/VFHm
awo+fVmnnSWVylsn5rQFNtZDlK81kdDxFPykSiCmB6jtbO6ORJaWOriXf7Kmyzd3BHonftQosK0g
uEaUgwrWm3cIVzJOlVhSKfpIXQ8mPjB2iQAqTYZrJ/biWAAw11iRBpJm5wHXYwmUENROSqvu3QK0
E1mDdubNECrF3q8pdXqZCoZQemlikb2NGghJIaJD0X7OiH5vxon4p7ROEyUheeo9ymc1fsUKRJRo
24DyPfPDGphalLRYauqUA8UrSBd8iT1FQbAhWY7xG5FJzd29BHImDx0Fr2uVK8sx+Mc0W7mrQRjo
kq6osrM4HEYoWsWnHe6hitQ/tC/RRowBtj8jMDSeNh71LbqfBJL8VLdcjcyGhA0jF5LnfPUizczv
NaD56PmCjDlZw2GKAdk381l1cDfzFUc5pMGzpZCc4imrs8ssqvdjkzFFTCcwnwmFKggmQdrPgvnt
6Lkym2bM24xaa43LQOxhWeslj+t8Z7luUsJ1SAdYpAtNIx7Uj8Tq8Lpj26Zkk9lPrkHjdjC9oPfm
sRriZvU0XbGrOZsLdaEeOjGionL4FEg54AE+OGWeYdjCWSI5AShNiWfFYS8NUyr2KfcWQLaoAzPI
Ygg6iqbmCsQb8kzE+LrdWryrvsiqok/klGFf3s8JGF5guadGzOBSNE0Ys3+M5QtOomO5L/WRGdYC
kFXOrgeF7kMVSIHoBBdebXLo0t8vg+Z2+cbEZG4jJEbiNJVtOFKR0ZdyAK/TOmNSuX1x5IBCQkNc
u4YnGMePCag6fJqkIF2IpayQioSxBaHJzIa2ZpVr1BXZ5jYnrfjtVOcnTZb87KQxgEfSEh2EbJ11
syc6gy7Csf741RBUb/QsBGcpdhnN1IoMLZsAQSDmF8pYOU6nCT++2ccnj6YJHoDD6htQNSR/LdLN
QRllXlZySecjpxHuUzOkI+RSC7Pip9Y6jVtxnSAZ9IC7Tg4nNqsGjWlDCWV2RizXPW1lSHk8UyXg
Y/JoN/xlW+sXO2YRelJ5toezE2mst578wDab6vR4Rlm2azPWG+osGflL8Bifx6ik3dOz9vPpf7EM
dtU695rxMO2hFNtGs5FiMAS18NwiX4M8TjLC/hv4BEi219b44ut4AKE9AuWQPR5fUHFMiu4He+MH
jNEFox8nwkmfiVbZHkGSjDxdvGzr+O/8wbT5FdNkqWkr30nh9UBH6pbwC7Ihw+bJ4lLQfuvwSubr
hYL0v8B9onkLLODb/O8Eu3MDKaAqF4CgWIXfXnRFCtXnLiD8/t/ntbMbJ+L+PoIVO0PqMAq3Xe3t
YKve30I9s7JlXPSwNZVabhIYxWz/451lgc/pSZ2sopknYecTlkUOPFAHPLzjvlNE/2HzMNgy9Kr4
zWi6AYsMzEeecTGtit4xLth9U5yGk5fVCzc5IDeE+nBliA7sWQFVsPxT+8m1dz5VCy9hY1pb02NW
2k4F+oicBzkslBxfISc2IBqMSvphn8VNgxA8Qty/IQc/n9ja1PbB31VzVq5z+r4C5gSdBEaqer/T
5K7RQXOt/+NPrtvzwymfHNeBk/WmSx/nlyKTxkjTLYi9d2B68jF+yLj+FKyteMUGqiRljeEf6C6c
e7kiVVTpNMPRDU2uDNuEWmJADOAFGROGfcHh4EYQvmNXvTDTT6bPTw7cGI61kP8S3KdrwuB95g3H
HbeeFGvHBVBS9Z2IWUy5KuPKH0gGdZGSSBPcyDNOnNNjEeFsr5UfEq+lGnTBC1SAsi6c8p+1gZY+
IhwmWgTeOi3IFBR4KQE+9vCqobkw0x6GazoQ22C5mJMrRnjJ/z5DaD87KcVe9sbWnFsRQkOzqa3W
vYdfNJzsaPtxLu0RS/wOg7Dvjyu+9L9AkBiCzDpVoiSLwLAxxaA16/UtAfVu8kJfce8RJ8xcgWD6
bFa0DnQq5UyX/0j8zPa47z+avXXh6NNmf/YxA7rp0wIR2VOi6kY7A9n6bacsY1jGRX7ZPVagCwDo
R4scYK8cjvLzDtlBT9GLg9QZVVwHo6ma/rCALYxLaWNvoY6e5g7Lww4EXi/UXYa8UMGLQk6meYro
5y/JPFsy78qUDyONHEq4PtuIJ3TPkzHtmfZ97TOFP8E6b6hjtuf/MrXhBxDGtR/r0yUzkt8f9YT7
+JBSPmB1e8TxbwLXQoiC4q9eg7HPWHywemtb4kilJmL47wYujPPwPLjSB84+UNSEM4767GjNWWAw
wJ4xtomNZ4MFYTkSejJtBo0BGoX7ca/ryUpbza9oV78XysLNsIX7K2iV5UMQijndAjMYCutZ7iQJ
EUdqZMhcp2O5l2LQfuHZAQ+J9Gr+2wZ7MtiyKkVpx4KQ790JPfPvZeEDMxJeGTxW7rqcUr0Vc7X6
h5FnrjOcdiXVhoMWyDSD51AwPsv9NVRYoahcfOJvB67ybrEIZ04yKgkrMOsBYaczGLe004wee3OK
9KA4NSDCbXYpux++ohkb6ToOQyNEyL7JcfSdJshlMGx0M6+wH3EDgg/+swETpFkPD/qbUQs/YC9h
72twR9P3/LF0R88jAlrcrZtzpNcKlZffo71mkbS+JyL4AJNQQBjPCLlSAv1Cj/++SbAOR/gnRZU2
vmCRbe9cLehduLjFOXeja5v8ywDWFYXyQUiY85TCWZRYZBfHkHKDdjnL8P1MRyLdp/chojmxAGHm
UgFrUgjv7ILKhEQoi8RfzOFDJLvYCQ2ym59o1uKQdDg4d1oL1mW6CfEEpnYrKBK9Yo6kKtzmdNlc
cgQRiuqTkGPkJO6inyI3+G6ybujOjMrdnxsc6oxl6yl4Er85z3U1Qbl+fU/VxJHbz3JDYMODbBnh
PH47x9AbfEbLAkweR36okjpzbN+dWjAS3j53lcJpTendJiftrOmZW2M3LNN5+jZAD516fAw8sALT
/P1iDFAbSoLSP6gWe9Qw1hnrcjoV3m1vKXNjLS26U3ZABGaso11zusssqW08WoUozPEEGfBd/Dmg
anqhtqQdRUymdXZhitDun1+yEGFfJ3YTu0t9YcL89u8XOrKL1ZAsd2fZ9Pv4/EmqeHXSiUTfWUO9
AF5Q9mbCEi15XN1jzepss9m9sTuUE79y/yeNQsdV8AGvjoKzfFRjwmeY0jEnTSmroBPLq6YYn95z
w1Rky/hJbADid4ybk0f9m2KHeTDJfr9iA3J9O+GyMK6wnRgt7zhRELmFQuWw73nz+5V5WgHdwtfD
+LeSVwqVBd/E7CqTAYyPMgFpKcNNBbIF5B+Mt0DCE3oc8iH5FJxvh0QZhKTvRMyhsbOtiQNpbshc
WRSyQlbenFQ9zH8xaW4An4cYUhlyJLRxny6D/E//8o0ls7OQ7ZIhOhQAuolBFEot2z6cG8tHcGVc
gqP5cb8l00hErGeYzm4ogZu14lh1Ld8Gt8P7Hvq2LRU9Eg2Wcd4ZZv+4Qg8fPWV46Yiu+636cimq
Gc8Uzir/uFcFpfuAQTlqX1fpYQNCOvVKnpBnGV6kI7v2nieBFmq2uXDWReUgSxCdePMJLMOwMK9U
acb0utaYmwL1mA9g1yGUe+9R2qNa5f/+QwPjiQ5cJXn7b2Z3rPwpoXNdhElkNZSaI4BezL9S592g
z6x8GcMZ3XgP4niwccXlRaE6pNiXT2ZjsoulSgrFFFbqVV5y9SDrpWXWgszhJmQSMeR0eR4NED0X
uOs3oQANv3dqNV5FW9YieXN5CtHPyf0NArO0Sy1Iw5NKbRY/KEuE0jX+ptDUATrjB3dl7avPcahw
RgGP0Mjdfv+ENYx71dmNSEHnerRs0m8hFQp7Iks9ntzhuOJ5OrglXYyEOW3IvKeVxTs2KdiP+Bqu
3o3WaJllqn+V6uBUz3BDpaQDUu5QPXUVR5TJpV+RoA3gZmNveeiy014vdX2cBfZeywcVb7DlU4Co
MS0SQqZv3JTIu7SVMOzXrVF4qhhJthexgKIAQKg48dVQfT0gFZKr0E4FmCPtKg12ypkQY5kEcErq
ogMJsLSIDAwdCreQUEoQiHahXnyTQ59ho7VMPCU7PDOpyG2lVC4oVum9WqBK6kU6c1417IvcduuQ
gMNf2WGZJR1IzEZs4wKUavb5uU/TjRrmYPOsCYwBffPw94fUXRJ6ULZ0JTa2bQ4dAy8MA0MAt6kd
Qa8TngJhrsPp3hWdNCM61MhboErVozSxygM7dhSV5Zpe2JBnFKhrwKCCOs2Tju7EZc412bYUrWLJ
FhZ2qdPpHv36SMulj/NQMtlL9/BkM4wQmJQM5t1vC+JMk/Vit8ZBjqWIeJd9d12i+9fIPCYMExb2
8LciTvxlZsAINvMSw3gTS0oyCHnGA5jzZFPKeeE2r9fBRegI6IZaResu30u6NyhP6mz2E3FNQbL3
VdxLeWThL0Ass6EQ7q8SQOyUBUw7K+xXSqZmz2+Yd58W1w4aQZUjuJMR2611v7fv3MR2N8AkUNK7
4ra2uFsqVuPBrc7eHxG3biRa4D+dPzPX8Q3DDSHSI5sG9MJJojGmvCTVfm6UY9krtDV7foxwNM+4
aC21SsoCcHB3Udp7fcBX+b3l/LoutqxhCYAlbAxJOlTgMXKtpb+Mo7ti9qonLTBbU+8Rl5djdeE0
KlzOPO8KvkHdnGh4JpuCIAo3oaHc7Vl4s34mDL6hbLiW/YtpnadGJ+CQ7tYedM3uEf2dDExofwIV
+IoIxb/7eNhuS0Kfsrls8LWV3TUm2CqbF4EqK89Likvyx5iw+IK8rFrOSGi0OJdzQMDAOiZ5qS+a
qfSwGggWD9gI9p/Cko8iypWuk4PRRQDghny18MrqGPzaK3trYjr9KTJVOHK5e2PxyGRGulbGytcR
qg/nCa6wFCS1do/7IxrVNhL5gZfB3WIHUNe5l281tHUL3vKDVbxHnlSAfwN5/gDGieRuWaJfyF2I
0zpZwkwnZLzgy1FI8j0RF1Qhmn/PdSzDrveK7qCVllAH52C9YvFHtsUbk3+LpjYS3J5vwZazOPrE
lUubfcLwcqkd1Mcek/NdZlqYAs8di14bH+bzBo9iw4qc/E+VwB/LlTcqIW7V9ENFGZsi003elLwN
AMlf8Avgs+x6QeNgY8jnhGVc7FiscBqDKvafO38s7IYf8plyxS7D+dIynUFvc2IABxhZCsug0YI2
WCx+2qsEkap98XmIKrBCvK2W7AEfTM+z+qtGrwyTLsXoODx2DEIZjvyXEYgHhjYvaaGxF7Dqpd0r
ArJSstWvtCDbzJmXADq1+4xVuvDU1WK/NfzEMbOW+mwoyJ5+GqY75xpmjLCmWNYUS+jYBWLpAXQs
6zbhbN0quqYmr6N1tulZD9aHbR14q9xeilY31IUvW9JRzaaAp9Q11TNFbWQ5BeW3mXjWUTMJv+aS
pvD7BcUkwOaORyqw0fNKruNLW3LUW36OjJBb5KM0kV55yRW6ZPmKzI+CDkciLrbIeZ52IOPPZpot
Mr4y07NHWI0l40oaip7+aC89z13W7vjo/EP4/cBcej6ysQabCIwTRQccqcPtIglgVHiBpS83/rwJ
ws/5tD04ipfcL7blA7Pf8icQW9UpIvKwY9EHLX4B07HteqjZytWIN8+wz90ynYXJRDdxZCSooL9P
+5fTk6WWc6Tkvaphycz5Yb62ATkrI6yKjABIjIM6XCA3LUHCY78vkLnFk1nyCHH5q7L42AhiXj/+
RMpjPZfC/KbCztp3F2QNTACYmGEG5Dzjqou+VjIYrx2y/LLqyWMn1dQfOkGdUX/9yrmz5ppjTyYL
LTK36GwUHhIKJchNvBSOS2/y36qT0oFqlKEoC+1HywG7HOJPENmQTkjpZhMW7bquWY1zHl/NtyFT
IHNiOwwegiNdWLPh5Pq6vde0ZhFpqJUgp4hp73FpQkSCtGMQSN8r1A5QKdoqsRIASZNpPxrna1Bc
hiLqTv/KJEMSDj8hLkAoTf/BD33KPIILsO7luAaJni/4KY2BE/UBGjwp/XBJr1LK4LKvM93BDa6E
Q1GZnYRNWALQbItKb6+06Xc5GZ1PZwuxEJAMWPp1DSUZTAgAaACGmOzoU3OzIVzhC8mDd6sgjn0o
Lz1tezAeb0XeprfuVGJ+A1/f0C0DmGWgjF9lvc5POLp7UPJWwZ3jbATV2Ucu0r336s2mVsqyL0Tu
3/jnn4QqZ7kVc2D0vQn5/Fu0JRTqcAZeiVPSsbXIBjJgUFgQi8CporBjlGBHK3Ms7+Ecqke6ogoG
kdHX4tLr+NLFJCOb1wsohY9FpoKZTBUb+3/T2GGezWlCWzwymOUPoy22soUTA5736cPy41k0EHtB
6PSm0vPEk/PEnt567Q3nQ9DwnG6oUeO5RU7AmsuCFuV0sYumK3MoQVOO/ExZHUjOnMxPRM53nfBI
7doGX33+99b17b/2tLo/KJlfRG+6TYs+S5kcS4d03UrVu+pnHdiS3zYlGrvPnhgZiMtu/xAJORfi
Teu74yXxzd/Z9q/CEPg0Vm/XWa4qtoUCQIT3AEwR1+Yf5sjNddYOyj7cobJFdFwxhWP1A3vM6y3M
Vcvdh2o8iZoLUqEZBekbBvblHpO//MCd2UC48/hWTP15HgqipMa5TW5bx4F23P3VyuVqjA+BhW2n
FdKi6qrjVxdyd7L2vlgEPP5zV6le6Z/aI8xBEovv5eXM8P+v7Xfpsh0h2rLF047/6WgF3fmxHBsJ
cqw88UA64Xe4fbFsJj6Pq0Hk5agCsSU/CEm4+noP/YxUIpccjY4nCzEGUZOTf6oeTE7K+6zBLbM2
PwaRO0ATCHLqfVtbUTf/qc4/b/CkQdWLlOzvuABRZ1+c/38d0baeA1RAyGW21TqL1e8UOV1UgKp4
6XPxOya+u36reHnNZ8Bp5TKji4Lg9VBXnkOPGDqf6R7XPfBhRlmhxBGYYGp6wNZx/ShGrK9L76LO
vNCfPLBQ/s7Fyr0RNXPUgbW+6aJVq4l3l4rma6VUQXj3gGQCqmNEGnvvMT1rfvmOF+FOhN3Z6b0+
Y80dfpR5cKTqFplNbHkVizITwJkcnmSacAVbgQCGgl/CClDeBaiHvVSxdVs0zbQM0nQX1Z9ykwmx
97bhs6zmZNUshm99D72tTRcS/ERqZj9pYqdErhViGnOP4ThQ7qg+bRJjjw6rTyAQ01f2O7KQ6kqw
JIklSJ2RaXg/0qxy5MSGrM/V5VYnoOx8xRhIpyANXsjUU3znhd252EQjiSd2+j1bKeFR1Pu7Ky/Z
pV9Gyy7KshnZMQyB3Kf+e20h2NSKpUEhyQlz+zn51rK+SoQB2XxTPmPouW4ohO1gaPahIXnD4qtM
qfj/YhnPUL8M/jsMc9YGxBGnGb1gLlU1bqJWzojhRpHjlkHnKSsmmBPPdPFZOye0nR22mArA25t8
9OMbWi/u1l4K9+qZrf/dHI92ol1A8H59TdjJuOeTNsim6TuFKyoWaPbKk/paHkKPOgYdWk9L5yep
qswfOjXCgG5zbaVjlSMj3PrELcq9ckmrDsbvZItWsEbuQdjQbYPy0LHq3Jl5inhgFSMuiVghiGvx
ilGKUT+mslQ6YwciFQ77VBLkec9H0b38LLhNWaa2tngaZf5aB7tUrrobK0514YA79vehzcEFFxLi
HNvbSbSNhCm3bTFDYzLJLdYhDT/l5ouqivAKAyPVj25Q8gDMWMqKFRk3+H63CoL9JpaqHaRKCZrO
wXPpCaXJeLu8TcXidX2XaiM4wtLGHuYDO+shFeY9W/LFekmG/OAeJi/OPmDO/bb/QWSzy3qPNSwN
/V+JFIfMVUdCAiHwAgqNRoXZgoOZ/+5v9gs5rDcx+E2WW2dIn7QTjltArb7HSOpsdAhSfe0YuKKT
TJxuSlHuGoa0txUb/bfG2Q4QeNpf0l1cdWm8FzGkeafBXk4uMcxFNaiYJyYDjFe770bmLV0utGDo
/PSiXCFmwfTupd6IsJrNT9aD3Zlf06GjaWJ5Cx6WMW04/Kpo3t3AYqgjKOwoMDkgP6nWDMAtDHPV
lGbK6R1Ag/Wii0iTJERPgIlnFyJWddmA6Qsy2gype3DfL9KHDHKNIY9Nd8SCj/2jEf9arpBYVPbc
uLkdNBsE8DRg25PILUVcmwYICLZM4a0N0gTRmZgvmb/C5YDGpJb0m7kgmfI/YJMM3TiIB1fHa3cx
luLQbAnoqySK25WAngk9QGwGMLS2hvCCf1vNhbMwD4hJq9RH7MxCCg9p6/s3cJpZz6beRjvKL6kI
3TOYPPo/YEyesNQOFd14tcXUBa8VrtG7iCLxwBrhg7DKN6SlzjAG73zGGPvR1w3G2iVgHrnYSUlg
tfstcBQBvSgUEY4xSnxxQcu3HGDu7g3WmXhtoMy2PR0C4Ep6HQ0zyqtMlUd5+ZsOR03c7pVTtq9i
696mSTWwga+Qmh0wnlPFJLzK+l85VsiwTH9QPN62bNI5HKDyjws6UobQ1sK4722SKbz7Ai4J4ovi
IdGyS++k9Fa41mmvwsXWbyBkTbj1nzo2kZbziRs6PhP8XXAE8Yyjcx4i/BNOnhuu47eS+HNg6RKk
zZFrss6pvIVPgfGZ6L0RBmluQDlM9FM1fB+5xZ6689XbHmdJhydOmpgo9bx3ZGimKWJBVAB+LeSa
+NlwB25xTidDN/YLtrle6iKVITcB6iHa5ayyxrH5jl5XT9tpO5ELGRFKfR/7QD5J3HxVZjI4Vf6F
NU7ipThIa4ed0SrQFPXXKP8hYvr8m6EEu8aqWBIHogEYvwfzmA6+1fcT2g9Y1GZ0LperkP65zooE
vF2yUXyHw54HJ6C2d14jM0Zxmyhz7ab7q1WDb9V+zBnJXHWUkxOHAxiww2WBVG9FYqaB4MfGocC3
gANFxFqxQZgxYsWnir6dN4vAVfMXckuAqcr0PsHhpcuPI/gnLEE+iM5+EiqKBW9ETIoAbEa02Pbb
l6aek1GtVv+sxvRFxvCT0ZtcsYEqgzu2MlpRj2HgrH7lCzPrmu2MYOPQUa6zI5RVzIvPTSO6Q98H
L+/58H7SGI4ATC+U5MY52oWNcqwyTYT/QxNU+J6XTocLxnmtyLrNZkOBKZ+6xADjtcfCY0P0EeeH
ZJk3xzDZ0ZV1cbbl9OFf3KmLh0NihAwwYSXGkfQJQ6NWlIHaDFNZ/TvMfy2azGW1YjT9ncwpKinW
k11QKdCouFTpAUoVFG9U11VY+TvtWmpdRvn20uI+lnW2uk4v2kJeDeBeqe4Ihm1Jo+vYtWV08bWn
vsrRqSFGmb6FeqDF0yl4PjS6sCt4QjMHz3oLARLeP95McYrKjnxp0oxIEJgxlTYRvPlKeXpK1YDT
ylCJaJPI66e2OEOwgKR8SLGTvIxmBCScDumvTTglt2t3fCB+7htF+uiFgHaXSG+N7SCMhO/K8sDg
MMtZVMPI73kqYFtCxCFzIdlApDlxOPKyR0kaCrgZGbXY2JDZcr9yV/Y+s3EEDfp+AczLbyQxcGzx
v0T6I8PHSjdYnpd89TsbvikgFJ07kWy2iwWT8I+z0dOGhUQyLiPujpcniGocN7qhO6fDpUb7Gvvt
/BQunKyNgFu9RpivJ9pBbPY/GThrwDcRswcOlLbMnlysvIlOQD8ShOoqAxYiE+4VnzW3DCra29bA
Hk0cclY4KE5J9ddFel9CIDtygmcfcYWVn2RQzCL1uoWmDbjhR/aE3C8XRtpPgUdoJOoPEBlmo1v9
0BsofFVbBwdLqsew0nsPnvcBVU5CiSj8YwVCmzyJUH9Cc1l5vNQ1WQySFx7gm2TjEbzfjEcZ8OoB
apyVTODjHWZSrXBOQRUvnpRqgoLtcV6wSdTVrPsRkBgo0NbTj9btCgTsYU3qDOjoMpWep96iYz+m
Pv4/MxTQJFKjVutiHVCtp7yg22GvHnuYXiTsORgKeRnyBGNkwPldBZn7j5JXZR4wLELCGIGOKg00
k0dFxv8+H9VpITeC15B0NVFkueGek6TYnZoO5xUAm4C0pdJi9iBPxT5rslfvzw1z9t0BHfFj7tgK
X08JI8WMXtMxD6cVtoGHbniW027z35Gq1uY5UHOGTXYemgF2nm5FH8pUF0SodSxq+TQvNSfd5Fxa
Vo4KgWh0Jz7FSZW5iY5aewCskI5Mhj63V9JAITSytcuPNOVO5q9SQQVRSQyIA3k8HcXOB2QeGigM
5IBdmXhrJEP4IiUvL+vURv0gUleRu0QVDQkHLJbYGOBZZmQNQBwFe6o9vMC3EAXrA2K5NEO4VUiO
PMoXicYUlKWdgRpHJe6+LaI8rHW9U1OiPh6951Ndg4ZRr7RHD0CEVyiLzpjh9zEyK+NOviKJUY+L
IGbIRxfbE2EC8LNDQs0R1VFs8WOZJRZy7jxExHo9U/OTw8NVRo5wV1DjmkvkMb9SsUR4+4Oyz8HW
2gmgQmec7YAi9d0x1Jz8p1MqrqLNc04ySGbBkYeT/53i6XuuFA574JxAw1efrMOYXLz2qijEqaPm
VfO1/AjeYDfPwCeYbnB51ongiQVnr9kj7jZ20hpCY5HuqmFAYE9qY4LhnKQrlohzfEBQeDpjPW/D
4biEl0Hz4y1h+jIMl2+dVhMAnGoU8Jdcf+NFekcl/CHDKx+f/f1ZJfTDZ72raDsH7rxDEqngvndi
R4IfPT15zqNc/lDrPN2g3fdkIk5IgyB3QcaGkxWk/i7qtvI+cbhsE+rudEN+aasTR47oOwaeHvfO
3GzUmGQ/vVS859k64sZPgpTfWGO7hF/QL7XmWlh5dBLC8pul0T4mpCjAAXPcdERFGYOxgQiuW11/
GSC+I/e1vKDpYhj5YkIMDs/l526PZSc55oREc+ZJosgnHhzFoUeSUlzp8HHX2xLJC1GZwFJV7O4E
15MlFf/O0X4T5+TIXRdblbbd1R+dJGAJQgrBkL/EvTicMWOrUkFpmNXoXIKoi19KQH99igD3UUTB
sI+33KnsWFbOjRiEfisUCxigygr87zS3/qQhpzvIL08hzYXPm2Q37WW7r7dLqX+g4TXls0jWvTIZ
jr2fx7vwLT7FD1VLWkmy6pJ70G2MXEh5TQHG8uGsD4DY6q1SM9iiaavMAANLpvBhQctNUF3tU4pN
54xGZBBwxpFhZXoYbXo+e7c+DqWwFajonW1jugth9hKBnQ559HB15KQTUOnt2BZS7UXluoMiow2u
cPNDC+kDPPxH8/aV6MyLGls9rsG9HQXoXz3wYVfSIyKxrzyJx27SeLSNiVxZl5H0tLzhzNzIxxJO
0ZWinPD0ajOB7N6NGfZx5KTy3V5ZXvOl+mrDIwgJG7KgTpCIWX0eEuTVTL3Sige1PoxACZBsozBp
6RtyIrxuwon3ocfw7Ktuuah8KyLG36iRTKKjl+E/U7B28VNaO9d/t4Bz23k5Fi8nPrbEaK+epaV4
00s2JsbSbsbQ0E/45P3RsRiSF+SsiMYxORjy8htwrKzKwS+1hPak6uTTs5bpGX4mEx1JzVT/wMo1
AUpDfYUFpAVTqccJZQqLyTWLEw1r+L9BIIQPusHYWzpLWngtt4IKZjROWrS1L0fzw6EI6U6tIl9M
GZS0kMZd7havDRs4sa4dRfAKEVt8vDfif+UyZVNOLZolf8TEKFkxzRsOsxRPUcbw2N0rddCZbQ4h
tEHOS3ov7kFLVMpZypRyjzMr+XNnaKKJluxLAxZJbDhHfs9lOEEdyIpzRo9l3DpLoi1uwSYPmMLP
qkQcdziAnqceIaBLm1v7YxinUlD1FNEZcGzsl4Yh99IUiow4y9/R+cZbhuAgkAFVF8vVvxHg0PKv
T0fDhOfu4eQAYO8kondjXfHJoqP7wu6f3+HWTXPu3fjcDJtciglPs75yGPYzIQkkASNLZjbt/cpV
LqYE9kRtf+J1Oc0uFSJvRyQw3bykr1urcTAKeanvUoOMmIir6YVxwuO+nT1NRsnxbfvoazQKagaX
+KKmp16aW+XtwXzjYGvTWDgMfyS/BI/1bQAiLnKJqh+p3zwL8z3X7P0WQy19fss30xnQv4Gugqj/
FszMd1phmNqIAkDUhQzy8W7rT90UP/EZZHCUt8k9Azw9PVI50xW5WtnihEXudMgNGwgI3hOhfrf4
4M+fsxubZDY8RXZEt3+4NAz6B/0DTOnhfJqH4TiZsC6BY1Muhc/vkOUnKpr7vkFL/RgKpyhs33/3
UUtwMoyffOiw700x3gW8mcsqRKqtl6bYT2m+YLKMuCxWSeGfS0M52/4FGg/M5mcslJOrIPLo+z7j
DvHvbZXQlHH6MhbBNRVKptoC9GFIDnwAIVUvdbfN79QwzH0el4o0di7f1PeqgDDNbNdnVde4o7+k
0E6V+tGETLQkgEP9NZC+mbiVwxtHQmnkV5GpRqZcZcNmnRU7w/PzTOW1AL9UII87vmSJ1U0RXuDr
HGhfheEyhbV2S8MhRWLStkJEYIEoB1zPPZ1eVD9owkum9B26w/L4N1tJq3pveNDL3wZi7Y/nZKL+
Nvw73nOQMaVAvR1OvyF7I3eVng/s7Un3fQqpLs8dQxS3i7GfSxaUqFmOICe/9RITMcDM4ZsC3lnr
fKUsTaNAIqI6jqG3qfdl5k3IpRm3o9wWEM7DT2JrHKQ5yPW8nrgh74HaH9CWLBomuYo2F9VOBXYC
WO4ocLeYOGdM56Ot1kLTLCBcJbQ4rZGBkzaJ9PRSEtGlrAP0y06ZRxZBtsD8J0cZ9cp9bLAFKbxi
ZErzF4Y0mxOctVnhNEWJoMwVwJYujmtuTFitJO1VaEeMY9KIWlDTpi+xHuj2YZnFCO2b8cL2PaUV
YIbbBU7rCHeQn9OtisxQqZMNLWR2gBVNMrNKl5XXBoOgKWj6SQYOebAQz9sSN/lHnmKXK57JmFXy
owbN8nlKpShpCgdKVvrWmERHE+S6gE68rjRSmRbAToPvRbfuWAOIaWM4opieieJj3bh8mLn010X+
yeZgNj7ZWLIAVrIpcwX8EzvC/F7RCg8BNjofzXsg03RtJbGwalOA5RCPnb4m7peQCDmuPA//BvvA
ZxtFuf8OLCdW1D57+Vu+iwUgwzmUZpe8jgZhZXhgVl+XpHNb7YwWpB8H+RT6sRWvAYK8+bph2WCQ
NyamGjQE2+MFg/4u/P3GjCqBM4W6205sq5MhioCNob7nOtnh+TFhEP3vmwV5slDWwyQlcqqAjwxT
QGFfnIEhClNqUJijqcJcaa/QhqDw6cx1B6tpRAWyGecYWKexXdnojg4I4q+7M+m1wZwPXATqJ4q9
mTzXWXwHQEyceb6juTIRqWRYZarL4QUllZAYPST3xbD7BgsBeuiuYeik4reu/dyHWwSU/5ZfdLKk
h1NY069YyB7GhytewdbPc55OH4vzy51ui1HLT7zfgSaW0l/ujZ7Z5+SrNKCt7s8khsDpiGBuXlL2
dNKiVzMjALxiPY4sS5Ub3Gok03SjrYeWun3h7FViCbVmWWV++dJvB7HoFQ8GJ770LVGG7olVTRj0
OQ0q0NJ2U4EgIgpWpJsB9jCHYgAslw2LyS58TPQ6k68RtmbrlEGjjK7W/t8mFcZ+ekpiPCwpymKn
piHwgkbXUrffvN097MG6kYjcopE6IV0Z6SOAbMFihGTt6CvW4EcAGaCyDWyGvt9DmiKve/3FLvPA
yCzlxAwqTRp8xLmiqiKd2e8ByLADs+6qDlSuGrPOdf4gVptojA7Dgb0AJIBKVpRNIKAoDiN9TGbb
wYlV0f6MOPiP0W6U+MRFi1H58WP3T8vTcMWQJMnlDNkfcO84Snb8+3W8PX3iofq6qeenAXmZieN6
bwtbFr0Zob9lJnx1u+/vj7yU5dxlzHEShX+BYmmyVGKbAcMtM6wYnOMxqG3BNP0h9+KtUUjXMl6m
VFrxFDxabqg/NK3y4/MSYuVAHDdJJ/DaXjTq35PPNTj4oYfdjIVvloptOWMKlZT2uELCG+N2b09Q
hli3Wxgfk6UDuybr/2q5eYIHPBEigsQjx4HW+OV+6T+FZ3lZGMUUtuuPceRgoQYWhPp/1jbldRU8
XRoG89XRiephzGvVIz+EfdLhM7srmwRZi3mFrRpUSEu2TZV9kZmshHwpNl9roOvAACAmwGULBtVZ
oIBbH46hWdqQ4c42E/sxmTTyxfYHL0sMbkvDuxkWBTlONYFyZrHYXYjtpjgMxbmYcqsz5Y5IWOb2
aK/MnHtDo6O9JiNHCUboLzzVzGcufsfWRhyl+kMAKRoBdmSoRD5q1ct3OiwnmarwQD0oMit0OU3j
J2QdVWQm/4ZHfuKMSe4Fe2vnaSqrC0XMHD0+CTP4aVyWghjDQKQAQ6ZV4P90LwCUOSXsvQfi5BE0
iNfMrqhh6CHizshGvCwZtUxXmgQCa3YwcukiwIFjU0rxsJCJOI0VIrM0eR+28S7aUaMWbeG74VNx
2pBd5zEvnRSoE0yVrUl2zmKe3jUD7H3z2kHH2c9rw7ouNUUNAB6O4pvFRsmd/tvAHnWrY5jJg6oI
AL3/yu+hTTKu3L5WhMJyytNUlO8MsT0Y+s2IYTtp6OcgybBxbLWVMQVW/x437DpFLbuF6+pvasbV
w3v96bESCuLAfZX8Hnu5IZF/y7ds5JDEo/o09YIoB7v8mZGVfq1ZrUaJrIh8SyYRX8CPYM8s7MvD
gdoueRbX+oMkDscdAoIPsSoAovOzfr+NOAp9/eFmhh3WFbNG2wluLZwJVhABAf/L21Q0bjOeobEH
4Yvezm5GrMyxJT78VOScgQTN0SD54obJW9l1LI/Z9EWrzGAzzIGHl8eDwhcJ5Il4B72XkwxMi/6k
QLufjJiYfZuxjWQA8t9KqkcCQcSMWZix+NLqzicDQ5umRanRftScVEz322r4gBeQMy0rdpd05EIt
/h95wXoc8pk8fFoAebTVlmHrhG95XjT8c0flixihpEuSSehaIjGnk5M9WkIEa0PUsAN/1FAWcLWf
XNC0TP7qlrOjVUtVKZfjrVrUGIbh6nUZmMH+DX7TosRo8oKQnEIkKq/kO1doEjtBtvUq2g+NSCIq
j0bYYJBqm2oavNw1P4rPq+zf9W9Eyv13a1C43qHARlzTbzDViJLh2g89Xwf1qmKzMTg1tUVUh/Oo
cj7MToXr2wvf9XjL5QkDzA3b6NIySvGHmRLiBVy5BHog+7Hc14Cg3N63uqqi3iVmLgJUZKHQd9S3
M/tnux9D8vTGLy/GZP7RBPJkqhZC2h7RvgcnRMBbBo2R2plAE9GtP1snzhphr7sL156x+DBuWjqy
pqYGDwvKk+4usrwV2RvhC6WWUUyKITIrQ2VpYw7Lu0cNWPS1jYIfnoSETBabdcbrAZu0bwRGLNUh
GhBwX0ChOdCBP4uwdWhLOFDMNXt+tkLIPgC1CWEVumPY+EWZZK8oYQ1Nfyb9XlbNNtfIwcyVJwke
AAF/zLUFjIKti6JEes8WGvnw0NcDKQ86v2x5cpSlpyQ0JHeo5RODAKmnCQ1ey5j2wKnx8Oq77ouv
cwGcPbzNVl2/0YRz9DmG9Vh2azJ+qK7UmJVahvnE8SJbO/k33joefjNXW+4/BQgD1GcPgpZPVn9o
NKigs3TMN0W2jqjc6cQPOoguiPct4oKcvUvcOXiqLXHt5m8g1RUbVFfrSPOENHfb36YjQjxUuo3G
22lOYX5v+2ES8Za+Dwc7VtE/kh7ginWUWIsR2SwDcpb/Xb4uXl0mjDrS1Z9SeZXy63KJ67pd5Nls
ujasEX/kRUzzGOiBrnff50HcsRxOIJ+sbAbwU7Zfp5fICSxHWJrqT/UHUx14hPumfkSlHyNfQW5N
d9R+sBccu8LM9w8ZOtxEurvwY7Qgp2Y5TXsZyTZi+/gtZRY3KT74/Ru4CcMc2Tjp0u3HetY0rEXT
+zZdCO6X4iSKx00WLEdX8AAN7yequNhMLjOzQ207pj5eqDhgxb0hGE8tMztLI9KDjNohmg3diCmB
x55KcIWMFfuVCbh/xR54agppcC3Y6kUp77y5hczVKTVdEhDqmBj8IBvMWZyILu5ZNfnaOAivtxaq
eJatoAJX/20DeuXoIB0lbSLFDynvVJJk4iRfkMf3WPt0Lu3/AI90152BbYIkNNVngH+QId+f4Uo0
eYwBTRhhM9vzN81HMQvM6jqCJHX6WPUwoCVS/K54QS6Zq9vO9U7tbbZ6h8mXukpCgdyEuXofGNoM
qKV567HKtwTF1mXR2G/NmndCe1tpnpQRYIvnAr0uS2uSAsUFAUarnqcN0mK7qg1+n6Igad2cGFC2
3dIdmcCAkdi3eieOjpAgwv1BFzFf1pZD8bbUH3YcriDOA1ozYYy+5HPc1DPpqG9F4e67Re8zbivy
fRTxou1pFZUCIjnYp6rxP9RoiINSeM8edcdj7rCNvsQEHQYpwnol5UArQqN1jN+7UpYoXWVb7BC8
YNVvaXtRSOC1T5+JLfHED4kMdu/eua59MOoR36T/LA+BZM5FD/pcjCPw1D4UkjnLu1r5sbnYTNgF
v0S9RWrxbpt7Uu9KOeLTtBGnU4wvNpqmHt+c3+A0SAeTpx8uK7Hg/I71r0mOZHdhD3PzUF5j5se3
L2J5R1hfeqjv8tu4TSYCmSndUFKMvkQIx+0RyICOpy2aCHxhVv7iKmlxfuwxVK9Jo+J9MYKKAWgD
ewqV8tEUQRzqplo5ciG8BunWkr2E/vJVYhcLQVt0Smax+EsrGpp8suL2iCv/tCUsizdapsOmOw5o
3G6o8IPd4Y3rVtyjDEe0V8+OFCeG5QyHFNqV7q122j09UwAg2ZprOchfOTuHLpR3BfhcNoX/UiDj
M2+YYhbLHAqDxIQZnf5lKLF0TJalf5XCu8dyXlA1O83rySTv3LC1O68T3d1Itf/PyTRjD83T8p2v
0iO0c7uMBeObmYpp3McFWOWS8npaCe74fks0xfjzLTSO82cVBsmYCYkRf0K1PCCn2S6StZq3UsEv
KF6C+tvira/xXvjtrBm4EtM6SDfHLM/QEUkg3e0yKr/LQchSv+LUwdroEefwgi7D7VqVjgggqYXE
IyStTAOYVrImvQvmA/zxrrEaeuKoOWekPRLZ5rv9qdNx7vVfmlAHtvnwwLbOL7t3cYgERTZugWTL
YW8rt77P5mLaD5uLywLNg8wWScWJbTYXO3oeer3rGaPqp/AuAwk/eADi5d1OObD9CWxugSqqYbTv
0OJfY27o6lVf4uM5u9cUvkqfwxOIglSFq9G5LMF9oDMbPfszUGBSfUHjEMlmfzjHkzrHtWAMgod4
5bKis/1pMrudKkUM4EFSyV1PzItRxJGlFX3GY5R8NK0oGgGumYBLTelAZsETBNC5AQxUzwMA/onT
mCtJwNKSum7nBTeZNGHdwnQrMqOdNNr8DCV0Qnwn7ItsYlPDS65iTLff2RxHq9LBTL+UqEYeiFXr
NcoQe8BnAPYM3AGAwkAu47q17qtCsdunb3To0JoJnNkyxxKvk8fZ772WLFSsmc6HkfW2/Ce587bO
T0dMnMfg9A1MXf64Q6B1HiyXQ6UPKHQiFBEEmkD0nqTFOOC+9iKPz+OTO0FPMAr3TyojCHqiEgys
aoJd8xKsIelb+GzVcnxXGDOiJ85TAGsVcSMlDZTPRDS24ohP9rGaXrmtECgUveWrCC6DXfRBiMH3
Ht9vjgN2b97CkaNlQKFkVFrxkRzgaNa4Z9Wdyg9S1Mnxiu6xZT/UirDHztZW7xpO6qm3wuKCdJjg
93BOG9++gBHc/U3zVQpINaA9rbpPd99zocGfMX2WAPwvbad5d1ymCBuoxPa2Qr3pHN1VFT0c6ccv
jP45Wamcmiaduc8XbyBoIEef3WNRxG7h9GIWuhCx/bAOBAMaN9rVV7Wc6fk4FxAPrI/52TZuKtfQ
TiLoxPE20M7mKflLDXWY3I+UtlOns3e7gmT1x4TyYwUfu5FRHvFAXJ3xwtMJZaCnfPa/wgkkEJ0/
qcLTrLGMoKyF5EMxkqffFJ6acNUIdSqFa6K7Wqf2jO++SJ2qVqUzFboQpHLyEhtiFLOkexmGhz8z
wU4MNQfT7MS7CJqLOyYVVHiC14PmpbObwFlTVQGpImVscOuVRvBEg8mSIgRmVWk5osIpJ0GP8xT7
+b3BP1qkWOsAXrlngplEu3YW/Ry4AxSxt4/XIIwW1SanXyllrv+uqYzzpSNxyA0LBGKBYfiT5QBy
6QStxtQGE4Rv9VVBQtecbey7bUsVq8V5KokFWuZ6FWNgRGYQ0DrYyfIbez9zML20rFt1YDrh/+Z8
V7I3Esb3Tky/bT4ZwT5QdIhGta5kFi0dMFbDiBWHCR1I/xk1JgoYvIhzoSNsiRjAFy2fQc8TSqdC
f9So2jWh6k3vhNhqyMLK4rorol4QCd/YqQ56Eo1G9ETbc013fZWSNZH50GDtCNCu4zQQlvCMqksE
ok88tr8HKjsjFkEOt6IbJtBVynvGsDWN8BLhk3StiImpmGR9m/0ipndaqli24HjlB3fEm77Kb80e
0JJy8aDUiQK+sSWD8NuuJezTfvb6tf2ialDni3/7IIdAFS8s+rHUrIc2zFFj+nywpiJniApkLHP3
vnF4F8Mmp+Bh+voktGOdUFkYwSqaPHUYfzZ8DbgI04fNndumjkhrzpeSsJt/prbFfCfNKJTUVC1G
PZC1ysNEazmRw17X2nYdIE6vBuYAg0wnmbUPv3w2EuDODCWppBeMM2rlEK0puRMKSt3vEwxK+d4g
VE4Z5rdOl/qE5yuAduI6Ts34yOBkYbJ+K5k4d5X3ZqirgUcb6fqVYvqFOfE41dBa68pBZiXg462o
i/KdM8KYjgCm9U5lY0Kx4r9+p+WOWQuplbRHcSsL8wCD4/1cF/IoBbc4fX5YBMbF2dFfDDSIHXiK
0gblpuAnSrJLycLaGth6uS/kE3Ps8U9p+aOc+z+w4Hcs8mk6d4xmP7zk8fdYc3eOJR1h3+TBzkxW
yWdoxWQYVj1lh5mIcHiOQE5a41Ce4+Klk3kFSWQZgfN5bWQNTMdSQIQ7SFTSX7OgXaeu0+fYJg8V
jPkXWwXMwImOt611Z42Ouwv764VLyW1ZQw69GWxTp/9LxU1e5tn2mJqfyTIt4t7YP/8wq7zZmlan
HOr3SrdVW/Cnsej040YGNFjDOUMq2donuK1uELSYOgF6uy5d/n120UZ5D3uQ5LRIrD3LILNK9uwG
BbjqKQA67CcUDO5bznL0iX6zEJt8j7UPxdRziiIVSjgTTl5R407/pEZOhC0+D+AbZzilHjTxgTaY
GFUjMJHRd7cdMqbJMKpkxfQsOwF2gMWJRCfSfYwkSxsLsl23yii+c8T+Uganlt4XVzw0WZxaGlah
LtvWlGM7wGnauzDzdvoKhNKl0+4kDI3Gd0ru1qu0BpDBkkP6a7QJBivzu3hhrc8MgtA3lbNortoj
BTLdYFgDBM59NL9NGoZCMGpEnWQ5DlyJYZfZPBEiYVJlfu8qxhH+cYw5uPqdRrpJ0hXe+rdgk0rp
E2v+Wc+nNsS6LQxzQgUCsKbV2pe+pX1dhvZAMvTBrtKmQ7PA4rNu1AYhZgmLvUgHvsM/+Tj/4zor
kTHv0uLtj0rI5fy7qBcYLxGS+Kd1zK0fuRNyGBGrb+rm/gUmSwRWQsc9zdJQCMDYyy9IFc+ln1kE
xg0Pwr0oBIO2BzsEHkHRJHYQDiaU/ljIPi4Xz8nsTkXQIeXzoFrGs3iZR1E3NyY9mCHvE11UQETy
r9X1a/jq1dG2AdiNbcdQAhPYI+/dU4HRMxGR1QTUU1t3pNBW6wcoOUtSM3cmsx6Ikkru35EcEGUD
p1wo2faZZhsR/fU2AWaSpnL/vNmLPxpxw6B+jmT9SMAmtZnVah5Bc+OB6GP1hQK39mWDnqCE3gLE
UnRzvRs4IyKEUZhGkxLQU1NWxhezuAgfIvmzxlMsr0vv3koV/HaYLF4qQ5eZubw2HVJbonFTb8YF
eJC4dEfvB1VCC60RJr5X9CtmI82iTaYrTkbnF/y5DbkVwgaHSFcbpXo0aiFEJ+jNlH6f/vg6OFuL
kh3N7ODkjtMQD+eAT9gA16Fui8DgaMYQ1/4ZQhtoJxvodHXH9E0xojGj0D1spYBl4adfYoZkPsQO
sBoETZGWz1qI2u6eTuYOOw8isAPNIYjP2GQFE1L1crhoJCXb40LBxJ5evSA1xkwyyXXebpftpE2o
wIaUjMnehPcmtGECsWj9I2LyJmhcH/1ZjDA4SxPtuMr8x1Jz1Fglk3ihz/AEk0UfJFCmVI1XAwx3
QB1Z3pXU/1XE08wJASEdpA96pZjJTb37G/bSJqvZLJoS4yQcC2eftV14DTMo5nbTyATTFdEKnICZ
8oVmBGELVRo6xF+xvgxaXnxOb3554z/0nfOP6jK/VyxaVbY7m2AjONhN1lTTinf68jHp5xhXUF4f
c3KysU59jndNybVrD6p3GokAYLv724HMXoLirFynO+lxEoinwfWkODSsHZXpCHcFr9aV+Kg7e7PJ
G6XMgcpfzVWmYWFfKcD+xERX+/E/MZIlUhoyUJYj78u4KeUDp/C3o9w2ddqTZ909cmNdQ9+ngBce
wBS8+iduh928jTclkfulv2saaaKQdW5SoxS7yO3oZYarA/HoYflRS2cUopj0mjxeG1JvISPe1F0u
Ia5ysn+R3RzsJ2wdzoxtwLDSvQgudkT3RPXEe1fCuhuEBB+/ygiW8F7baAvFlwAPjvvNsxaUdq5m
Tx5GCjXF8un0BWLeNh+hqwiHpqjL+NimiX0nkLtyRZh3ueLKEiLqn+DfK8CuUHAPA/4VEWE05u89
4AvQpMRsMrXO60804C9S9Y2C+mqukbjKXK1aeRfLcu38suVZZ0BPNFZyfUf5XHJ59MEEtg9sCzRK
MdFcgdXHWCRH2vnn5XyriAClzAdPon4RHeE77v7LOq3XcRwmdANmbRWECZpV05Gn47Bdp+GxOEp3
I4rkRJw+mWuxYcXeoY9TlVc4wq+EUB42OoTYoIiYG80WOePLyG0kagdn+j5GhmtSE9Bycx6Ypypb
bHWR2oeCeq2tGI772137KZUevVIXJdSEoIDkalPZMWYP57MU/XL1EzIcoHNKaYk1QPmno4JPFh0+
xrg7TnYeC+5zaR7a6iBdTLw8e5I2NvFIZvgSgfygOXgPGB3KP2yPxJQOcXeN6GptqoWBd8E/sF5Q
062kKmocKquH65zTSulGC+4bzLQw47yC73trfCF8zTVNbPuEp33dO0wy5SfYbCz1HIS5LJAZfaTD
412rTu4tFBxNUB/Yxjw9MMz1Z35U0H1UNiFaRcmJ8ym3fdYynBnG9MCcjm+5CFMFbGgmeF64LzYL
FsPuzAG+pGE4iJHtnyjcCJstx+U3nqdafiL6+YFjE82zM8EdyRCTBD7t9GFZBa3WSlvtIjBVfv30
RGtecJGU5K/Y+ZqEXXHvHLLb0cm5/zdIRnuBWj9/BITe1IciTiYmOQuzblF6knMSui+6TBS2KM8K
imF/OXddcrCe+7FmeAUs73DaFM2FYgAkhnwA1ad/+HPUbHUxaYnDte08ysCVrJye5qeYpI4Bn2mL
jzt2W39OU1E2GLith6qjcJnUfw5zRSuKXhHorh+eM+lzL9Bz6va9A+QSDDNwFT0e4EzzS88iP2MX
f9VLB+m16r0JwhUjn90fMPs5sQQKwF9hBRCYU87vUvIbmyOwdbHyG6WrxSlxgQCCUhgKKybEEo6i
/P26oeXeQFFTm/aAG4kY6aKW2YV/JFvDEMWWuTzjZnLHWiYxkXjRJyLBW4d5FSSZEeYCnOFnt6q8
o3xCcNcrFpDtLS786Hueu9snn82NUN2O0IjGeWLLBkaRwoxm0OCd7NtHPhvExD791FMK3xl7famW
2IPWJrGEydWHAHXHYOyj2+6RZHS58iKXqaA/ZfRNhMtdIcNY4Pypu2UOD0hXz3b4Id3iV2zTKF1Z
+CTOvUJt+oQ6q7f4xm33f7zRJIkGPAwdS/0/GRw5cHNOjekZTgPGi48lM8jxnUrwAwrwohIFEFEd
zBfsvi2dHBhSQr8PQy/SsYjG5DQO2qk5xDPX5KEe9yDspbaFwVPj3QxoYKOa/YN7S0xEsmwf4ZTu
40HMfGGYk1M4aiUFmvFODCUwKr3KYdJ2MkxC1GJUgJSKGo953CWdI/IlOuaFo9dVtFCIyYI/EjfZ
x+MN2hcPK8yaR/Eho0vNhKlapfExWMCwIngvhcO51Zs+3gB9+kq6rPo2XOtYy+aSuiS12LWAc/UP
LmwSzgOpeaSS25ovTL7etyvC7rgmucnuKARMlM6U3TPuqtdxJrlP+xWNwwZU/0IYz/cTUojGnYMX
u2kitpC3V9yIU/siiLmDs8rijuxUL3BZvzFdIiVDPo8nTQeiwY8HnDnKR+gpyvA66Z/wTzyVR31t
Sktvn0qxasKX2v+4PlJ9Y1WMulzRelA5JosQhumoS/2yCWzLtuxs9ZtyKwr+1zdJMh4tmoQ3kkHw
V4ltBhhuA/pVrjzqpggtXG0mqRkCz2G4+Ga2SxUtqTM4uweGnRmxvLZbBvvhNrPSpwC4I5hy/7x9
Q7ajNV1UHQZcOlazBHQoOR/oR3U8N+kWZ32GNTyX2jnoXjtWsQJOSI+/3AxYvUghsdyD8Lk6hzlb
xQVYgxeoVm4aTdPYI45k0st54tEDozpnQGWCDkFxOJfAhAnZaqeC0FmWynjeLfafCQ1Yn0Mwm/W0
bX11HukfBGHWzdmqnAZInTHffsltVQhuO4bKT+Kf0EWltwmyxxdhVfZSJWTbToDQ2DNc+mpdhJZG
9eHbeVEuOiTvBzCIdRVQQzJ6qci67pd1nLWGyvYV1wXc0XxnwANxwfRHhOjpi3V+tMhlQqk8B4Ax
iq/ebLu+UcxFFSdz5/x1y4i8y/ZweESVxo10oiESr65ltMKwORg7ypgGq2C8LrFuS7llCrmwhApV
gcM3Xal9aYmENgE4u1mCZv0ZSXN1MTorFfzAe85FGv2h4wG4bO1IaKFrIAiSXI0tYJnkV7hoSJ4B
Ybtur2tCUhJhje1iwZkkywxegr8An7j5uJqPLlAsdP6q6AjyjyhVWdJu3WP7rd39D0phDrfCPz8n
TdlXxJZ3BlhAWP2wpx0NgAvMMd1vWFZejoz6yxUTbCThQlWgn68LhYFETw+x6JLyEt2roFDVW45t
h7uObQTVmQO5gR3Q15fkL62/84LObWB1/7blI5cRT2m9T1kNRnm5U+YWJyWRbjHvWZIcvSEHLFnZ
+t+HqSPLVU7T7BNHSUcLkkw2eaKgFCYOmxLNXbsx7Js67avkSk/ZQjnhcGw3fszHivV6nuHIjGFK
h5yKLHsCQAgvcoV3/2fm8ht+agmUPzpDatktpAzsCbx2JF/I9/XBsdwTV4rsXJ8vPxT8/KVuTZ+z
VyAjPApF7VRqsi4aLGy4ACJjNc9K+9aW+lygdVFkDCz7dMKthSkEpePOuzb2eujmclwi2bnCITHp
xlVLifY+d+Dy3wCWTZEYqz36tVzB5jJaDNvVYt+BGS9PTyxeoRiEEYHXqgqIGCEq4X2i8wqhqGZq
A6dzw205u2zx9wkNL3hbl8SUBiVRTC/klT6U4EAyNuOupRit62Gwp7yyOwhP02EUMKb4q/RkexYJ
1HxS8yeDf2ltv4lMwB5ApyoYEi8RCXwF/9Yo3S6EvbjQJRwhgYD0WHpK83fCNLW9CiEeniSKc5jz
tR64BcAHZBF6aLoBS3qAx+KaJB3jtoYxmTKQB9dRTNTFzfle5Hf0EDr9LJhvlYKBmZn+KKxBlLwx
frEMlfaeY+G62m6yuifptCxlUHvWHNVWYPMta5FPryymLEU9IykQwQZprg6YqdUVVuV+s8Z0cy8Q
9lIqonxJCRC9ilLgCjNksGEHGgHV0ySCREp4JOum9txE19A1fUqanyaQvuswfsOGuA6F3KJwnU0k
hYQmCCEjPYtokewaCUH/tOiSH38iYJ8Il5Uq9wun7EOrqLawaE88Lcte5FM0NyAi0AeBJ2NByUhr
RmEx8J+6OGnRLgHCZ0+E4nbZq73v00JCA5WaMNyuD3x6RWxmMDgVqnypL5Slb7inBzlw8mb//9IU
6HZCVQVAE4AjJzOkJedRGNr8DtIedYWFJDzBYMFFKjNUyqs03rgHosA3CL/WCCna7dfOC1KuNV33
X2HZTzQElUzBDWywm77zf9ZrvM0iB62rMieSOhlFNrZ+m7UfkQt9Uhu+EuTObgPk1fbfQ/ykmGlk
T8ygoKsU1vPTrPY8RDhV0AxUIf/RHOsFm8ij0C/xff9lrAwB94WfkzyaW4SSmtPe36+U5hGRiOHX
y49lNDZ1mf59DfDQSqZBOlMmTZ643GQUVx+kRgeE003/oUGGWriLV9Z31IqnX1AsXfmq1dvwTL+7
xrDkla3f4qOzWp3bbtiG6e3lMVepuv7FgXUy53qW7+FHhnWYdHl3k8Zz3zjBkKpVHEUUVwqdzii4
adqN27lhYUMAa4vQTLNLgitEnzVfrfUR00k0jfLqqTtKMH4kyRARlH/p8ZTEalHfb+lPEIeb2Th3
swoh+mYmQ7qB0Jq4PVUgotNtfVfedOA+plo6VLjizaeb5HEPtyShAvDC8bxiGy5CuGTr7NFv8WR9
EKtiijnFCzDKu0TWsTEABkkWi29tUZnCP3ocDxjFweSAUqqDtQOOZxhvtoQ4rUBSoSwZAlMBTWet
K41hHpNovRSauZcbiPEwgi/ZVoHCHidt05OgVQPDsg2XLHT+U8bAoBH2l0Ra2gWdV6UAUbCGjhyk
F+62kLyaBXpzD5ivUb5kPhN7TwGkACrIevFEdDdQtuuzXrPkJbJJw3oBaFNhMhAo0XAq1298t9b+
XHKnUMR4+LlhpHveF0BfpvhTG4ZHujuO/BYTwo7Fu0neFnnIAWQ11zx+5+TX0r/GuM5AejYlhFX4
65vngunIYUxpsiVMzCR3DNcNXuo+AnO5LrHpQd7e6KbFE+IaGdBykAv9Z0Bzrz7yCpMhnJpQAUhh
fOD6VoptSpsz40E3vLrZBkYGFXgES7rtXnsYvN3tVlrRz67ecy0G31N3A5xN4jF5CNeT2CMWkD2v
ef61ftrvR7J3aHRT8BZqESmtAmp2ZavNcoCOm6oZTsdtvabPegd1lBD0FQ1/VOmhMhqNdwcpks7p
fk2OoRrCqca8mIHtilzuxYwo6AnsVHNUTUOhWtXXEz2FFRH1/+KtjCPVxVZIDXg8ORJZGfUpsyw3
qI7PA4ONl0Eqej+ughTJ3iOs4qzr6z702KlMB1nBj8nbCDUzzxrmeTmmbjM1dgBB8Cq2ZnuI3idc
wr2yKFa9SjEKPPMAbzUSFSSMmhBHQPiJXPix6AQY2Vg9nF3WbiIb11EnUEeZ5gwRfUjyaZnJRWNA
ahb4kuaXKXEanBfxHyFKDCEtHRvvVlGwUcQMm6yapMahyiAUeFhKIMIHjZMkmwWP7GjhiulpckfM
ulEjTRO1fJQaC2DD7NhbnuhCFCzOZYQ92omomXEjpRkuLgwjwk/oNs4qfitmgY270/vluugt1Zr8
I59x4mv+a8d4/v93J5zx97v/ljhlU+rm4D/f4mVYlKhGcxmyXnZzrAatSwapsU6JBAGQAeEdEHr6
HbczICXg7M/vGzT8IPMRTnFzSUFZKHpo9NmHZg2PV/RbSqs+p8Td0ByzHf7gTgvw9Wj6kyZKrZNX
3ehoARiI5V8+6tBijJhexUNshjKFN61PpPWbA/NpTnMszkp10lcLgHT+DDn5hVwclIhUAKcIX/8L
4B/+IEtBfLYNghSI9vXIuUr8zr0A5tXj2A+G1C2McJctp5eSZ+raqhbYZSW0C9aOQLba5+DCE5zD
a7kXg/tzz2JFOR0cpgkeXrGO9MkmRGbzEY0Mp7XojNs6PdEGQNPzPJw8ODKXrQln8Min6ul+E/5Q
aB0X3ZrMZUleZiWFIrPzBmAQUZE8M9WZuo/1eC0f02ni1r+spK+yfIrjALceZXtxyloFf8MSp25M
isvoKVX+qIccAGz1CDSwL15FWlYbSaJpiRAZHRtSP8qQb5vAiUUFVF77QATFtIP0AykLFvqPOmIu
9WfY9PMiPsF0CSUQz2G6tK/J/irZNEm1zcrRrkH75vnhoSM69YdRE3DJ/+s0BhaTcpZ1rirv4Chk
0kPlyaaV/RkQ7+mv+U+4Df7RMJyPLW8OpAayhfXxhP+btkgLK+LAGWL1K+tBUYYVFqhmQpcmNsQn
6ZAAF4szL701Ig6Ea0D/Qh2/wxTVZJrUOENIP9rQfCAgGZprowTFrw96Hty9sz+zW+Lg4HlBOEDM
FQGGjVn49aLqHJHA66tjtdJ6T5J+9qAbTdG7s5VxMm/xmVzXvD1pxlvWqDWEizEOO5FSVC0FKvy+
2t7cuN7wbyPGYVvqNE3EV3tUtNVuP8gZ4nxtoNhTjuv3mlvQ0rcD5nT02DE5anP35RMU48IDn82k
lwd3/Px35J9i/CkFcc4IbcY7jfsD46r2w/8andtP4C0UqmiI0nvWmt5j4PasdqNnFPpsX53D6h8G
iwRPFMVcs2meECN4NsYFtQ3a2L4cYYm4Bs3EXi6D3I0S+xx4MVQmtRdf0jNp/pYVZ0HKhbyP3QsZ
cesNAtQkcZYWR2uJZvf+0rjyK6LoEvQTS9tNa1kk9GRtigXJVP7Mk3n5ZETKMjJ13YMlduQ/Es3P
2vK/E0FSa/bdy4kLQ269Iz91TqQQA9o2efhO+Twd8Qki4z2QhvDXBFXfhoJNDlbjWwelLGTRJBmx
457LOr6Z6dR5EbeAaIABbJiisPQrM3ArbfabHRqpK4yWUH3vUlGl6o+yXVwQA06ijIIqebE8MUSC
1dt5jYPAETL8gcKECwNDkuB+y7XlYf3oFZ0dZ6myFQRj6Wdyp+QYJVxX7fYZ+xK5ZIEW267UhaMY
ZyVLSYetVZcKiulIJgiI4CjJrRu7mKTwONT2DQTyC70odzRuBPNF15FFIn87MmGKAiGLbA4NdTZa
lDxzYlt6MIwEb+jukYUqdqJRfIpmxF5S3IMe8GMYo3jigzrYKKi9Y1CWKkI/NLc8ap5vG39SFOff
Z8qXFL8JGBT+OMLTnf9uEGIIz+URfn7AZR0o/5T1JBSbfxiWJ1Kp/ninOxjzP/pJRVGpCPt4C6p6
EuDRglqLfxt+Xb3tfQGlGtcRG909cVL4dUZrKRdTw39wQQdu6qyUtfxrucdvke31tw8KmWPJIEyD
ebH7v5Gxbq79vEarDt4pm5TSAhlMMsdK2UZn/BimlEnN1vP3dfG6bRv/cUCehWIXSS5d8ssVtvW+
e4vO8n/y/Wrqb3er+xGBYzIxMyEbv9mbJCEfBjmSN4vWAKLZtjx0s/ZklMVK89gioRCMx2XETrh+
bNjdX3z8owcPhLcy4n29FKpG28jpWmWA7KO/T7vVYXHfjl4wV38Rg1CRniMnDKMaRBuYj6MlwBdv
sDGNk7CbfL8SrYVd2vRD4Ldq9ouahvO6hfkffk7pbn/1wJIOiwZUAR00T68IlYXbed8FPHvSQgIH
uVfZ0fR6Hce++5xGv5rCqkPMruDy02dN+W+FfexznIaRuq1qhCMK+lgErzgYYUsQ3RZIhqNyZQlu
gMd5M16hpf1b6kAVTlTQEEAupGf8MqMakw2zmkwnPaJbJwJgGgysNM1itrLSbsbycwwAuYCU2DON
Ye28S/S5umkUMkSqmNLyqQlxBuNk4Bzbt1iJEw96FIvdnzafO7z2ppCGa2m0zkJWYwyTeJO1ZTC0
leNHXqwD4LTlg9iubSS95gF516OxNKIIeME4WWMKLjLzX919EeIM1aOeDtDoGeCdZPJrJRPk7AkQ
zLkCg9RhJUI1Z1k9oCUuk+9LFW+ExBFMavdwTzDHM1aAOc0AQuw2938WsofmgDeLu9enN0DUGqb5
FTLkzN56Aek76EdBYMSjCjL7hUlrFcGW5Of+ho4yMqfQKDxr+28MlpbUFipoNB6QdRm1E0jKyI6P
9IUZXrK2/MWrCPp0CP8YfycpCiMJ7N6iL5Im+bc7apnPgokPTRnuXZiAVB60Rg6h9craGmE0MnRi
gXIptKVJUzeyJxDC8mBf/Yje9Ol4WLeK+H9FT2JwrQ5wLECGs4YINTW6/s/zbUdmJZRD30fdbhUm
GsKn17fpx9guwGH/Fetut0ulKkq6wyLwCYYZoDBRtVkT6h7xvPa3SJHvPXfTHoJZjGs0Qo11a/ra
Q4pxdIanYH8cWYCRVLIOmPgBxucmstM6YXRnjJ2DEV2SgHAP0oUN6tOLsicAwJ6gtOrcqM5jBLif
xwwGLryqfceYwZEZi/mJ7KQ5I48eLbNdzMWNzLye2v+Br1lgCz5KYUSWehoqINmaT70SHjQ2GBrs
8sDID6GqqYFHlP3PD5zAr/wKdNiwtBeSwZFFhh2lA0Q5KBHtMgmHblIUsmPzyO7VAKJKC/lJOkfg
wyfm0PvJpZa4gEPvf5OXRluD7mkdRi63V+gJKLDFa/MpCc7WNGcnBRP4FLCfftEVA9JVG8sBhgUV
L1BhSv95EjFAZFUA8b2ufCSBtWJxrDXzJ39Jyp9x4OBySfdBcaWhHC6OnKxT++Yj1GvHRRUYPfd9
Pz278LMF+lUx6u4Zm2fhR0LfWG90vaMf9/mYNQiOqsoIovM00bBo7xUjn8euMr1mNH/Nhz++R+s5
bEFKK8Z/KsnC6iffxQaFA516K+GuTUZ31oswZDFRo8kVjJhB2n53d3YnbiQdv47BZrUHGf3aCB+m
nBv9Q2DFJ5r3lR6PiLW3cK35lHyGeRALVCKUT83y8ZJHMqDTQfIjLMxl+5d72Y9l0y53xfuv+Sf2
vqUMa+JqZIRFvTMQ4cfw4nUdp6U3In5bI1Obmun1co3eAsodS47Yt5ppbG/ku6v3SToOtdhKTHH1
FWQn68zSNPSnglnXsJKBSJifpYW3FYAOQllTpZ2ZTiVaMR8dwf1n+4twOdqpHftu95lKBkyz1zh/
GiRWrsLkH8K1lJ0AeMG8q+1v7kkmAM5PhYy5y4cfcYSLEAokPYyoPa8/23ZYgO1zE4K9pyOW90E+
mGqMMLIPBLAsfsBEqa/rQ+KzFzITDcIijferOgs5BgU+64d1qnqNSGhlwnbtZd7v1ZeDP3jX3ZJf
2Q0wlpa1L7fWiDyFlh8ZfCuFNVboZdYhIKNgxoApICRU7GEa4VZ3jDnEAUB+qzGmYS0KyG8NXsSK
8JYGraD3saVQTGKuTXDdM8wFRHYYj1RtovvDTBDLCiqJulm8tJAVIspSLM5xNkJrPkebtlmYOe0N
DjAPAdKemjoJTn053ItLE4Py2Q/rkOMibEzwtKcuZNbA4TXh58QuSWHdgIQokKNwXDM7anQk0X4m
jS6IRq1gCmhs1+vi5Wxo662ZvyDeTdDjsn8eYRMyzV1RnfizO9fK8cP3yajNoYp8auXLxHcanwbp
5XQHrAcsruz5ELNllhX2Fif+r0fWIKnNSPN9Iv03c6DK0W+4GSPBVayTz0vx6yFi6gMs3xHBUiM7
twkaGBwMLy34n8EuepO0+u4HfpK2XrHUaY+1lYPIp7rqTXKtFs82AraK7KrV5/3zEF8tUDz3ELps
04jQuv/zoHxbVTx3t2YXVBTfHnrxHi3xxQCZz+rfnGnQtzTXR590lgciaEz0GO3PPRGXZVwMPAw3
383SrX60PB2p4XLZ0QJ2MXhbXBJlPID/wPBdTOKC2XJSzDs2hYxUAuVInS7pI+dqq1k0JVnwpc+5
bA6q9KuxM2i0PHqUnloKdx4rU77nPt0bNBRFL3lKtYGXBHlJHOXfflZbL9GL/bQGG1LRF4rrDixW
1Qk/A7aV9Xn02l4wJoP5nXL6zqSEIGrHPRYLgy5Kx7GbnCIdHL6U3tMM7DKsN+mT4lDNmMp0RjHH
WKzgE9zlztW7Nltf204WImEuwKbjonr0LaKVqlzUOCNASzCcyEnIGn9VcyTGeVVHfT08xVW+AJZL
g4Y7vPv63T9EcN8R/Zc9CT6UQmhN1yrbebOcYI1S7qTWyNm3nEbNio6sDgFSbcEhedRCNRlJzF25
MVkwmUuMiTK3IF27Gw+SHCez3IeIbW0cV35IQfVOK7+8/TVAbkk2FVEI9dI8X0i7gFIds7vlhggw
cVhW4yyAzITlh/QcqnlGs9zEFAQbUy2NsPynPtR4/+5gj0Q8uFmckMf8eF+LGjyg/FsGcQx6SHIp
qUqji9E9K1ZYUTTWdGGn+OIbUjU4xNHkwubJG5/bNOYpHTo/0W5B/31rjKPCQeI2M5OJuUjThDVh
qxmCCc6lbLWwKV+61JB4V/AUPkee344jY7en7Uu2LXR4o7848A+dWXHQHOo9SG5tWsMBHbKcuNj5
c1asRHHyw5HzdYJUpu5JJAlmALXfywocUYrsGM6QBIcwJCKFEQlBKJfowx2NvaEjoUZH3aIpy+c6
VG1ySq/eRvwbZLCBQd9WOvbEk0EspxOoe5RLy4dtFbgn6CfEfjuePy7w6GWZVXv/L8Qx7VRcu1xP
csvVc00kS58xPTWcsyAAWnsrkZQWvXU3OFt2CVsOQ1WrjShNeWfMDeKjxAndsld5BUJwUG7Gt/Ia
otlQG+CbLPg4gd8vqxuWqcBUoOrA0mWTQT7bqbCZv/tpIegkQeABcUeoe1BhIU0FmBnrS31AfITB
TkavcQIfAV5G3FzDRtHHkyqMV4A6a5lR1qTsIGJdqY5uddwNQvFLNiXxEsYGvOPNqiFeHfTdjaYC
51RhcFhANMIWIm3ebInWuMQyU6YoU6TLh4tcZFDKdVYMxJ7zsB9ffcWOH5b5B5J3Kgd7PQYaPLa9
bQYTtoR8s8Awd/Fx7kVgC1wBm8f1yGCWXUeaupqnaJepHy8VMQzD0olgGjwdz2itpiPoiL1ETZLd
UTPRVytd7NGC5f3iDn4yEJHmGL2y49iXagN96t8AyxlI96fp2GlIYqT5vacs5ASWycjC4q3DLLNW
HKbT6o7YHKHrcgHiNdMfp/7iwY8HGiH4uzlvp4Qxv4TlanUMF8c2fwk0Poa/PZbwDpXQG84Hy4Yi
/LcD9d9vsxtihYuRN5YX6lUG8oA9XHVBz5yrtaksq3WJ/fggWkkF++/VNu7i4JihKLq8ys/PzgMq
sJC/3V1QdLKdZLyUmOGb6nuipOt6UnWmpDoMd01cJsUnVwlHitzUgyzjGj5stC27PezJF2X6Axe/
KFX/mtl0s8hHZMLwy2HFtjFG/c5mEsBmaxaXTzaMjndOUo3XvMBpPoaRsnI/FIlO0iuckcCZd5Vg
QOCrUIY7mRwzzHwT+oX/gPqXlvaeGh0M8U5jdzJZPtaf5lLpEt7q/7kWZSn/Df0KC26KUc6LjAnS
8aMUn73+BD8mnz/bhhHI885/m6usweo4K38mKOZXsmTe0AcqWJoxOkENV/LFzXVOWd7TkTcFwI+S
u0IhL4otlbk1oaQiBYM4754i7AOgLM8kcRi1+uZ9Xb4ki/vwaL6egVHQEI9wz0J/s/eaTSeheWL7
qzdwDLzBKyc6cZXQ6nPF9gKht+D8BX+iDpX4eym97X/eRrgUW1pC+PzKgJ8tk4sAf0TTWIuqSWre
bbB59w48j1rdfZNMtmsfC/FVbWGk/Ga0CWrbZM9H6yX81zty0tfxh4dgzqpFVHM8dhP2gYrXxDQg
rIynMHS1KWk07SSTMGP9z6mQIUvvyxWljx38ghZhBVaSg3DNnzK8DBt0rAVYbgkk/qlF9FE/lcze
7QZY24JOS8AHcBQlLA6cCQ6C/UXuJZsibIHCZQfsVsAdYxtKmheaGtLiwevcig6XEgXGAR7f1U7+
WqzzhxT6jmFCy8af6bbfFvnScbaoYYQYCOCCD5g7CTGznE38gCbQZqKfxUeqJdQwKm6GP74nxNue
QvTbpjzP09UD28pw/P/hlWqXtHxELkZrfTDBj5g6bsCfn19hEjKPKliyRtV77chbpltMrd0Bfmz6
7Lw6Y3iQqIb3GcWWLdtfwFcIBj9+04zxoCnJ5xazVkRa6x8S58QpgsiLxwhGdNGU34d3nEU9dKpJ
YjbSnIzhisoNguzv1P6OxrDGsexEpQbeAs/+0j3sySj5ZuuRjs2Gqpl3RiewE8Qk05ryYjcSlb1j
xh6/W3Nld+CZxVGQKBSUdhPzzi1k5hwM3+4r5WPlyuglTXfGffE14K9HbrEPcbFWBdWknW+khmc4
QmgKVYJAhaIPn4QmaQu0CJ3s59sBZ0NzwcFWMAe+JHPrqrxbhe+r0+hi0kwTuc4Qdm0UZQw8IdFv
rlEm63kQzo8gF+vNbxFmRPtv3sHMHXDpiDWYhXaFkJhiQ/0CzNoRwHpwWF2I0E0rGU6KEGsxkf8k
a2+nYF6uokvoOqvRys572mudYLOFKrOF6QdIbeB/RkHyX+V2syglY1KKHmoOkAaFZJbMJh4BWijD
We4AM0C5RUjojBxdJKKH1FO4XN0S7EquNu/9IZDiOBZQ1B5E/OiylAhBDm/Ctv7lF0ZUZS3MH9Bd
bqvcxZWyPFzE4PydGQREhcVI+PKpkSvRl2g1EVjJYg58iBMbyuVjY7qjORi2npeCgeo8TWmktnGN
n2+t1eMtFBXPnvXVckWibiPpMeSzLgLRv7iPv6jQYqyuVPuVVb5VCmDZOE8Q8OHZGXE6r7ZLZbNw
USS3vpwTlozfTr6kgIZQYcoGWa6osBZFEuyg3vxRyJ4b/vIO6WtxIaG44xq/gJUAUuLLlLfnsVKA
MqVipsW+EHY2A2kGAXSr0Gcn/TKZatTlKXgLen1fMiLc4o8Udotkpfz50Q8XSZah57/0sAcJF8n9
WNcRg7tzZC78erEpWRHc9Tsdaj084Awa9O96T5NS9uZkFHMackc6BW0FyLchvlmRkpQOzrO2DfAf
ubKswrMrRaXQ7ofUXqyJnKlO7wY4mwuCcN6CBczODtb/aftovlegmdTVeq2TBk/+VXME7F+OHZWZ
sgcXgEQOy0EwqYPPDcodkSz5E4qv6AFxBCuJ/McXkxWJXNmCfDkSBDv72KlZITgEVnXbJvTOig5D
On3gjBS5/C/f3T4RwA4+i1EQQooId0Dm96V1LtnusAlkcriaKcb2KAoiEcOrHACF6tYHKWdvbFjh
S3sKhEFOVv3iURb0hTWRcKPr3JPfHYOtY2vVgMeyGuniXZiR3zlKdLU5ZAtlUD82R+V1MkU3+ofi
p+mb/kXhc/v/BOQ4uXdFUfAhWSx7fz7lzc1+v6AZeJDLlR67Sgq2NFgjzhjI/hMAlSEU4w2EnUuc
lSOwvDOm2IGKMbVuJAZPtY738qjOaIk3oR+aDu6spQTLAT4kbkmfN3T278RHKp0z3UBs597exn/s
kzef2ItTn91V+VgXWGxJWiGbI2ZqDdnkLHde1id2ayOP7jPb8Og4ewutuPw2myDzRnh+sf9oEtv9
rL2LuWx8NVTkj2h1zme9wEeEhhhMrRFN0y7n/qqinMRmWwN1ohV226rJdDzNbY4//oAP53i+EkEu
/CMciuL0NUBEbOKX5HAOnS+BU7UlRAur/z9xXr1PRJNpKRE7hLqQneoSfXqO22Bhs1ZBliJuw5uX
WZa6yjMaGYY49Ptpg4UNCQTo0wVINYO9NCvV60eouvZlOO/6Ao9z7lvUi/dtLl0zRCpE3QcFfSnB
P+8Q8UnHcRblN6ngyU6HQN+Ql0PzG5x0mMe8Cg0pv7Oqyi5Na+IKcHIOHh39vnREqGEsDDmqTvPV
x3/tzuAXIp8R85V8vVCAa4Li8NSEnkYum73pMVGd/3GeOYW8Gx2qsxTxPaNFZRbXUI5k5L/8O/g7
zDKYK7sdcp9ed810vw2bYKuCX4WDyYXOEk9wMqkks6U9o/ZMfhLIWvemCAvVr2IgTpPRV+A0ZYJG
91ypJyrUWKzNG5Byj+yhOChYDRs1/iBkU7YHhEDXsfsywnziZHt+gZw3WFlEeUmGDtNT5krG7H31
aQHo69y8KCL1x5z0qJaM8AKyw4DIYbUcQdXDkRMaz1jexrYWONIy7MUhJt1rySF/t8Au0yPuxuSs
2szzqRuzEb02N6UEH9/dXUmAGZosygLgQw/+nvXA6nFkKs6aWYab+gyAR7rsbLWiM0pddp5gGZ+j
hcX6Z/7uerCCyYpnQmLfGQvKl+XBMpPld2FdOvbksMlp5mv+iIqrhmH00Gg4CRIs4ygpldg6XH/0
Jmeho8cEJ7db90qS/MNJpVLlkpPeMGN6W2DDNxLnyk3Tc/NbnBPcLZseljET7tdw6bM2IAWWtr0i
xyuHyp4Mta40kLv/wr008LIIAzEMCPfXtke6GfQ3FFDKEt7GdYPI5d+CUM7wbiy1qam5U3wjQOFw
S+7ASjT2NaAhD6qlDXh10UyQbi4jYpP0Os9vqJ8B5jXWo88preIsG6sA+HgBrAoRZapgi0XuEQIT
ZczwUyvOxwytARFXrF0r7CWBWBdjXMwlGqBHAkN2u2zP3AZoJT19b0vs0m64sSVjcjt71KePTgcB
ZfI1N+vUPiWPz+Oux6p/cEm1XeC+S1wa0gCdSYJwces7kk2kA2nGxXMTMZ4EIDWmv4j5NFV/5TrB
o170mpqjbm02IbVsuWxIFlnnM0lZrS00072w8lCzrO7mljHwLneHWtWsyaAzXINtLTZ4xo0R4mnN
mIvfrgseprw/GtxKdb4FwwYUuOgecBLR3aoSXDk75eqcEnGfGWHgeTERxwU6PLuyyljM6V6sjA4g
+PPSc+gVYamZHB5kGdU7Dn8iyNlqnXLXLQPuKP0uQpMDg367o6VK4FW4g0ZcpWs9HyGW3B6VXx5x
qPNIWNz89/QVWjEidLneymSaPLzfmTszVbvInMq7lG4QHRm84y2wK78vAFQ/a4mwp7kMaT28xTPr
8KI3YzaQNHrCmOZWu0EFvpddEUBq4wKICxF30OkIJTKzTyHumrOC9AnGyK92Y56vPjqR89SoKjz6
F7Frz2m66AIhdw3L10yVdtQyVXYb6yVIEQbphFdwKXaVDo4Xli+kefal9qROSPn4Fq6riigWHMyU
v/gPGqXD/2tKeF52cF3BpgrEYPu4hs5Oz7DVk3pTJBUSHVoUKVuQ+b21yzA/oxVvRW36COcziX6O
sQ41y/3L20u5eMaYMbkSlSyPoIHPCgxU6X0cmJFEzANX9cMH91jwHW/CeXiLWTU9lcG1xowNCnHV
cxNBiagjVMw5h33zE9iya7Ker0NZLUE97gvaM5lNijeS+IgQZF3KaN6EKE3/FREhOdDzkCL9L4UF
365sY8AlgwAPd8fJJjqx0fHY3Z0jzv2tNYzCrywS+nHaxi8+xChVsTcwMUdh0BRMkEsoMv5EkJHP
SttKCVgefl4OtWxYcsN6wBtXyD6WVN/LkNLkINunOCKHiSMuxZzUk0gp0YC59S1G+FReLOIXyCsY
VUCPMPSkARmqnf39/LbHXvZ1D5M0plknTJFdF7/I7QQ/ZRBbOoWy2/BWdM8s4hSINhcub8eLfFi0
FpfVRCRrRyPaMIP9yexhbeP9McUhbgN8FuDWnoXyCnrlZlKWGhFVcvDw5cfqkWGZdL0kw74hJF9L
TDAMFewsRkQ9Q8p7/sjFMJ8/JqJFcjVVPcRaFl9Xvinl63hyRq/V5+SiyqCD/OsujoT4AWTLCNiF
jzFkY1iQBBsVbxbFZ+MzHWVU/ERCoEabdcIxIHvh+a4LHW4ISJuk75DU/VuNfDxAAKYX00mpiQtB
bobDu6PXDipy4NKG+v/LRE5a0GLw6VBW8KIkqAuJbwwYwf1AcBB86S6lgXoc4cF+DgR62WSwgnJW
6DTSko0pnARIFb2uqQwH7hMU6hEEE51muwqtJvOL9NOZbisBnOAUI/n69gXZpGb+pith+NwSDmVh
FeBZpemeGbock5NdBGjzBQJ3KGr82OeV6JAvxrbgQPMXaVsabMK317gv9U4V1MVfPormfQg1sFxY
h7tlXWLbFhMj78io5QHxNY6fzGwTg0VU0J3qX5cMObp4edaRGL4jBaRfEqgBok1S2YhpGuDjmMLi
gY6B+eb676nzOWjNjACqFN9fd6gwEwiznXKp11VXSd/5Ac2gOtinecJ8ZhVmn/eNoXRrAzcpREpU
4q/iMUHEY2+WA0DfK3rGXLurqG5ixWKp1SQqpk9d2wWHmq8GY00s3UPPCdFaRtGQZ6owLG+FFAR8
Yv3udkrByVxSnFE+pykDnVodISyO//pHrjxFRhwJY/FHkFrkzWIDnFg6i9WUub5MVVOxup3CSHJb
Rn7dwISNgNjiRsw6SbIB8izmvVIjMErbiI0zVE9Vq6sXYs50tRzQjubNQCQceyp489Vi3EG7KNV0
9iNHI9K0bDSsZtitqhTJzSz1rHRY2GGPgDlTlfeOA98tR33mTQ9JATXucJcGHcwN+3t1lNp+YujF
jzDFixbPMkP9rDdkv45kgOytU/Ti9t6I2iavqD4QMJlIWa41/7ppfl48bVc0IIPVe4bbGkE9K+Rk
G1DR8jrneOF8D7Gvg71MJMIJyb6ZFZ3puS5ITTm4hfki8NhR3CM3WqS4hb3Cg4FgQ6wqnDgVOAHs
BxQbr904GGKsOzzTGQIFxPTlHzp22pNh193Aza+Ari8c/aatfBMG9INQfLqwKBdiCBO9JJIT2SrX
LlSLQyfi9+pGuoR29FrJVOG6YI1j9NzhG5H5F+UKPQY+aDCyqEaaw4XITt3m42BR7VaxjHThZM1V
XjB0j4frNRsnWIX8wNKlgItrFR+XhE+94nOeodQbKbPTeZng64OpFW+e2KlZQeUs2t6RMcxMEpww
ZtQQIwzyTtJZc+Blt2eZ1y4lt98EIbFQIMzvdnmJTRuTgZfvJu+IskLheOMZ+50R7gs74jfVmTmF
hQisR8Jk/gTtU6cd3N/7CTeQ+cVzEHOBIRJB6nJnlKPQcYx+BBlzyF/Q+HTw805L9/Hwsu3x0fxX
6Z1j/G4FDlstAY4K37DEZ8p1Zu3bkJyPmqu0wv3v9bNzgAIsbAQ3NKf0sVDHi83Tnhv6vAf/Vqeh
vSq1U9eCnTzqI4NgMov5gFKHTGGxUIbfL6m43R6CWNMBoIgmu6uAoJGHawbxt3lDEBlYpPJnDSXc
HJ0kjuLqHmS++t2juTCEfU6Mcx7dL773b3PKGVmHYXCUrek3a32+vS3f5GKF2vBf+Zed52z9aEba
IS/1+r+ZC6lusqNGSv5MYYAN25+qTBSwI96I4i3eJyNXzTYZ9OKWnY4tLyeDBrqtQBNFHYmDa2L1
OeCroTNDIUIxHFeZ4ctedkJGCPgeUQg5nd5NXFQDzLu247HM9NkByOHBJLIju8ZmOCpCPL3wvF+o
7VCT/IENMoj6wkeESQetWLyTRSMSSHEojycsMAapAqEpWVYAXdmcYVHgWT6O4UwVKhWrSGZZKUl9
UxxcVN6lmYt3xgHv3lZ5/NVW1SmEoSt+7/P0BApPZvztcoAcGw9fxatXNisKIsUbCBxUVit7b73+
yBVYHxjLpWwE5bIoTVm9p/EpB+PrGEWZIu0kSJ4YsHaIbQiPcXLmrWe/fnZnfrtaf4SvBPt9GkXl
uQ0A+GLDf3I9FtKswj/vdDbu4ze3cCPRzL10PdxJkot7qDnItMqN56ffg9Vm/Lz0aoTzc4S7ElZe
+UON60JOgOXuoWV5r+Ecpj4/Xm8CEXEXxCes0fbgVfx0DpW1iv2pKPeumDydvPoLGc0pUaiI9bm2
2IEkQHG1MefpZZnFlTlaYtiMdqRpsWstJ1Zfk2B6euMiItfGB5fhNUDjyAxEXAumO5HXSicRj3hX
3NYE5ftOothdX5qg/DIOrV0Ca//k/8DvgrDwSduse4eEBhL74vHxj3NxTtkH/IhR8NZuWO3a+quh
+jxi2KhL+3CVrqH0I4KqUyAoUw7A6rZQPUqRirnTJmK9ZrtyX8yfUdJpLoC7b0eJuWASQbNOK+p2
xpFiv5O4wUik/zKI9Gp/HczNTrHOhRd31G7BnK/YMgwoDcXyT+l0z8ItgIM1y6mkE8QC8ZBvLWsV
GLDuvO5VySwcpiROWJfkmUukxGHoz+Y5TZ/k9HYcdIjunsh86t0RsyRTUPQU5Z67c7d/cH0pZBQs
hat2ksrhIhaGfZDcTlchxIB/mCzUhVo9rbGyscnuX9fvIxeGYeYo71BW6poIoULIts7wOGHCig87
CSYRn5Lxc5dMEEpeDAHTVwK3GphGqEYKfqPtVEi8umU4xi6zOO4X6Q/cmsruNHJ1ujGNP43qAZSg
YThZtm5JXi3dcMsuc/pCgMfQquAuDRCcSb8/nHY3eOVzNzpFS9WONxoSxDV1SMh46GPNV0g24nrb
5XXK084d+muRak4nIlpIuP/RE4ici72os46qiWqO1dFBJ26pV+2cBIc8RrNlnZ/NKPI7po3B1vTI
+BCKG/t5lTIxmjID+jjjRb7dfBs2C5cq7DIlJcZL2ZDBRF3xzyQKt4GoKsM1CStY/3vO6w//X8he
M8qpA3HCnJ873nvU45pqZ6pgA/H5opbKV65IVCkmpuBUQCLvMB/JKT8VXjWsFLY1XTYQMKZRAQOX
iX9TudEUE7a7BSS2fAxlZgeeN4RJNL1gPoaABGdwEbtNJcETYMuQqq8urGxA1NcVVsghN7AAwf9Z
6KUP69qJy1RicS/UNO56LT+3OrDnTFa9QgDSu/PDbBBSsVN8G1YF/ryk2R6ViZNLq/crkL1NJdSd
dA20o/Fy4eYK4cBUAhqF3BSPmtk15rTNumqXlCVt6i9+owYBMTeBC3BOZxyvredqPMODQLkbchHt
2h+MbQKDdzlUR/LdT7iVyAEH1j11GD4KQ+s6DzToO2Eg+e8dWUH++2pTimRSxPBYvobcgY+siw2z
pLuBuc7TWZ2w9TfskYQKbZkngwYoPcuzr4bC/IMH5fxv6xLHO7iiRUx5bAjX0plWsdGEjVmEnQJH
/4vCXc2NwhiD0wzoQuPmSWexBeuT2OtP/RWLLrIaNb1mqPENrc0MHUfCmVvUd0pIqclxDmZZkWBM
ByVZGfPxjvb/CYlAqVM+pBdCKnCHByFsOjEkPOCIZ1L8h7qaQNevgb0DAtCuoKT2bh5i0/5z7IxY
Gsil64DbOS9VUMXOX4vspw8KRMKzMm3zxOvYLuIQOqOq2x64qBjKJScfZiSnJeEjr0smCOalRvyo
L9WOuXZu4GacL1SqDCmE8TbQPfNDp+0PJOZPx1Q5AR0/7hLThW6xfxmDfDAyoHx8bEde7K45y0bW
KtUw01aqqz6OLPc8avwiYUZ8wUwLp+OLy2gKGVfacyFozGFJU7yPFUNKLscD0bipDDe383lQBY/z
FN2gGzV465ZP6Ohas1isjDe932gKzUEyckj19mm/4c3suSerEBHdQK7/D6HDM+ieUn9/cOlAWUNN
+j1ctOnjfzty8S0Ii5ZVP2ED690KbRklXVPYpKx2gnrJrLLleNnHvcORTZ0EcM9oQCg2wFeF8KYb
o3f2QPq5KP9oRMywgpUkMjKP1n2nbEP70Bdp087BkXKvl/X/Zjg0Zfia5+ppFgQZ0/nSWIy2xoqp
JDbWIiisrs5GvUXh1LIWe4RimA7g746TiIMSG+Mz30L92ElqfpqMuDV+HaLHrqrvT3kfZcXzPTB+
5AComqLCLeeaAzV6FJbzVvLpTgBJMYrb9dnsprL021X7pqOutVLjqUCxqu3zKSPQkMvMzzSV8MUX
zooTZppikBu6BmrcutU8qu2Yot1O9hZ3RTno1Mq55kSr1baQB5r4ZlmaGDZtei+APbzxWnJ2JHj/
6/79Fytc0KOFTvMWHHjIcoW3rmlXIaw7LcDKDW3uXJsXpOLryeaL9HRkafzBXvapfvTempeK7ehg
2vx2cP+2YZB/iukLEYxv/sqUNV8s/8212rCOUBS4Q9/GcYxUXpuDoeK6ICmZrx9btr1jrrfg1Ig0
LOTLR7eTHogyisc3F20qOw8IXaQq9CpV4j28lgbY/YuDMdeZfeHUHhUYtUQacMCRzKzIBWGg5ULe
vV+sypzmhompUqIO0J42u+5jCyhet89sIWuFZAA6GvP2JH0uMIY90+QbeX8p7VgyLFV0VqlUNr5e
nbB5srFn3yvEm77poEwABYFLSOAN2Bh7JIHJiRATJuORUQe+/CarSQSOt+qOy88E2uoeIJtcVPv8
OlMqt5dpuxoDwFb4ASL/TOwoTrMNjDzend7D+kxOJ3E3kVQ4v4hDTZjgJxTd98AnD1sSMCIVvT4G
9qi8R8upMh3FoCqX1bOi99VY+BvTmLXkF1CBOgy13K1wmxrXO0YCiAHwJxboUzHQHhBwjJ41vokL
pnXY3cIcv7ybionraZnAUpgIp4pUjoUtFDhR7biqar2sQc/Q2DYUL0m1i1aaaDIWqcdm9j2Jehmo
/tZhlq0IqDAdHQwIEM28NauIN6gpeS/XTFRRj4f+cOuFla2vF9QLrmpVN1UMyZwwzgsOtm2/DceX
qo/D7jFtVZ8UVwjYzJOz2Ypn9BWoFONCT+XPygNsb6CHLCKZ5qqU/WultvO8xJ+LG2HPvmpCQiw7
JFVrUZCTKOGou6z0s9RPJBlSjq01uxmFSeBmZbeRgpJ9q0gG3oU7mz+FfmOLpc/X6NVXbdpjSSiT
DruB/x1Uq74VTl6lQHmbKASBMOUs5dR9CvEdMEnQqSAQL1cIYnoZRXAk4eV1tgt9GJDp0c+qEgXD
XT7gHSU55Fkc0N/tDqyaZ0eU65wtTeCsBqQCGzHfy0vRVbTN29lUVy+yuYkR4GFM2qlYnjJ74h7H
yUHiP1Xy+NZewmuuSWPxm111lupjVtuwXoCUIwOKXox5dc9eoLXqbcX+LBtPLS/LLi56chHPUx7G
isAHTzSVvRTYWr4iDMjKHmj5WzlmoQH20W1LFbcyaXQIs0+4Xv98sNLxrYm/tWHskytTf0XXJDpl
iWK7A0xXSVc3AhTsg3C3JGpKKZstH/AiEBED5P2cvzDMuuBzxOlDI4W1B6mDIujymnwTFGRQ74xo
ekDmEv8lp/FyhkWfAombnVMxFz/OLZ2gTMDqtHxLJyFBc2e/gTZP7772PHsJFA0tFoLoCIWRK6hW
YwMlnGB/eHiR4pzxyZPJ5AAHuhH4n0R2Gz95EE5ZEKfrQ+KbDkmuHt+KtNsmtXcAyKuBmfs2PkPK
NAAOO1dnsoxpO98HT5TGi0i3g4aK3wyxjNlyO4tmvs2+7GgwHtwlRHFe04LYivA9EKguFfaBbWL+
grX3a/jYPVH+NNEOHFXTBWEfeTRErD1Q4OLOUVcfZdAZCi3JY+O1yqx/S4vIO53uGSu02x6pLSCE
zgfGR+srl4lJEBMH1PwPjtGWDurqEsD7UfN5xH1UD/n2BRjFpR50y2rOehzy25/pO2dHl2xIu9Pq
x587k0LSMBPo9TSh0GU0LTaA/r+giBQV7DZpRU4FXa7cv18JWO/SDLGLrq0MSUW1mUo30I6GrWpk
7ij2juEI9JHEkk6D32yLtybMFqLYKRs8MfjyOI4/LZpHwIip1OZcjldoACHJjoxbqL1l3+It4s96
4eVPkTju+gO7U/XjhN0XzVoZp1sNegX58gDLWB3mVjmTivSTssoiDWXDzqh7BSUg0I5zamp/jUE8
EMp8zDtUmYzuAQyJUUNO2QGeZI+AikNhNNYrwoiFN4gWXBFdhJpC6jgBoPHFHhHcJG69H+FRR9bt
aloVGAYkZ7mLWz4+1lzlxjSx/QrZAoeV2bWctGSzFlH0tIJ2PR0+YKzYpMu7KrbEEPlHQjzXKq3z
Tn/WM+idgRZT35x96mdG7TR96ydUxpGeuWfcTbCDt9/IQI0KRtIiuFwDEmUnK/tN8eqsNTbpYnkP
kEeaOV0dlFeDhGEjmMfOF91SfgXpRbVu/W/QbOruGJg71QDNyyPr7aFDKHqUXqeD0ReLmpd2kMRX
gXZoLLziLefZVh0v85HBbU8pAazMx9qFYqCxdM08Cl/Md98LxSFEaICkMtPPc+e9uvS2y/XXIhQr
0NGxyIx1tSpxdBrTY9lwU/tT8zD8nkSSF9Wp89c2/Uw2oWtx5lEx/s3oJOqCI1Mc3Zuqvo7E8aRu
opG8G9WLTM7R/uN0PFmqYRMVD7RLHw59bUY3orLJMaHF8UspCDeOfGueQN4fRuSjsOV2pRMqbAf5
bpZFA8Owvzzgcn9/EWeQM7hL5U5BiqzqdONNypoi/dZki9AnQc7dashH8WCNwdYh8pC3OBIZzuJ6
jNES/B32xoF/m5SK7GcpbfJhqq01I63tzJ+jXDMsmKg9EH3UtW8M0O0nvN8jRbrI44M9GYDoSygv
0GhlRPFe+Yi9nzXxG6COS+C/laJVijlgM5pQf5+ejpaZ4ouBFcqUv2S59XYdqozNyQceX9udHS20
65KsqzUbNGNLTrBq1Wx/xHEFsdinzGRTfwYvAGcllhpGxeVQQxVq/X9vd8OlY/0Yb41AKMOGrFv2
Qn1OyaJaa57JsEWHHBzcA6nSMrIp/qAVvinUOiDfxSQL4LljB8AVrF760PPLg+FPORQANLJE8Kmt
quSYw9DevcuPguzeCA0PLFEPbg6g36jFp5qRqUgCjcYdDQa5fXrS/JdDFq8CAZDltnpiQbbmITL4
KVi9gOQiuQHuZROuDoyBXJKawnf9+G+sR/o9hyI6dUt0FgYjuLI1d+0IVmzT8it8P7bwK8IKeyR4
2jLaHcLwFrae3Qgl12bYQ5DOEMa0jQdlRzOz6/aNWYj9AfhHO9KECqdN0n9wu/i9I6evdbQmzWpG
jHrQ8+Hv9hJ4judRGj0qP/C9IwJiBlFm9gAXT9PQLGkZ+pUe25teCihTkPVCe70Prk1e3w7/ADco
ZlBuWjOF5TK4XzGRn6Rar5ceeeDG9lhJksqb+KMy8rfJiJUSq4+Ugi0vb+zTfISF7iaBgHb5IQ9Z
kkBolKbcKEFd+xiCf2wGxIlPtq3AmHgIkcoNy2x3HUx1zbg1/ZpwqFpzU06IuEc51Mk/JqkwzzVv
yQBv2EDghHSljh26Wk4D1kxDKaJwjr6txnUbcC0Xi4WWWyh6p4QzY6jdKHHp/wGFZK6qcpTGrZDz
AaFfnIcz4MVa+8B+mMfzLbeZSpT1/eMTtwhG2TARH2vnx3/3pxHJwsFAYbvA9s29wgRxav2BjnAx
YSs7UYOvS9OL2SROBoydc4DszqETYrhZ0oZ9PjvDyaeoVwDB2iTUdryculD7SLBMgflbHuXdQxRB
aNwdWqdKFSQC7t323MzuD1IzcE5zp9oG4SaH/umNRWRpgci9VTJhzh6t+bV/UAT6wOqvouki38Xi
NXe7a91S3sdQChnu7fal8aEKnHeqxy/2KJPqefN/7l/1SlhOtgnaw33HCGHZ6Y+Bgm88sb3y5QHl
wRxy4APYSTyuHrOq9mzzz0/rVSzFUbdK1ih7qMGsHJ0Sl0CSyK+rdgc+jqNLAfst1n95NToRHAVt
k54R2GajUPjwWJS6bP22fAnt9BmEoLy/0xcPZQPEpqtk82fZP2VSQAJKYdYPtq4FuvCGDT+H5Qsw
0tulUQOcSzAARJqyQdEo7/yjIq/073Ixq42xTUg0iNEL6HIXxTA74IknNJ0a9D8Ilhdu0S1C+e4e
9qbLYPss3ne2sIs9BY6vaJjq212QLDYDVht2A6c+awrie3b4kHMs1xUfe27y+x+j5qK0uCMOY0aU
ek2kdhmnENEzX64Ctbeq+H1/1UqJUZyUljkhC4FMBl8GDZjBFA9WeRkuy147Q1CsMzpaIoeJ/wP3
bRClZvUgWG1XBMwvnX46Xw7M9CMRRgRL6iA5immgG7eyUf8f8iBjNvOee4u/dXf0Hg20zZSarOIE
ApFmGv01tczRhKP970yUge7P9L5E/kwoBRBucVpynlh4qno/UR7fBdCqfnW8xcxHDRZYdrE4ALcJ
NoekSLrl6ztVat2waTsRAXrcmO3BXDR2bTqJd4IU9GLH9UL8pi7Z7/03M4LbZ9TZ7ItKjYLVpYqH
4MM/NvZrd4cWZsPTQJIyCC3CkIJ/3ggAOm2Ax4MEjB1eXBSgNb/JXSjgFMX4eU2f79XDFI2mGFSH
h7c/PHsjXC25nf38L2dY760GVE3nCCsvYayQvdtQtTrrTVg+NqVh3ZOX2Bc+I0w5OMUW7Ye+XSrX
JoONdNAdyFMz+mjNMyQXlQsLaD4iE3FpCvFlGL4nXERnHBan+oa4LDUtS55YcRst8urJoUcOMFdV
6wQU5Szeoo0Y5TdeS67qrobQ6CKpak1ivPuxn7AbA8jgzoyuST0rp65ENFPWdrU3zZG9Ek2Wnmd7
29R5N/qTJepcJH2orZy3Nhkm4E7e+3QmxjaO/jmCxMzONV0c+PYNi5+J9CG18MtgbNnzyBAoT00d
YoaKbrgU8Og46jxLWuKZWyzkcEV9LD53Xi0QFn8qrFIYUWZzs7i0WWAHkQVUrnJQAJMJkgP6rZo1
UKfC21/dwrjG/mKou820esvzpsith3SxDEW2uetupsd/dmS3zPIKZdMkrdECRchtpk94H8bFc2wQ
yMXSBoCKIdEPb3dimXIX1udblEP1NiVqEOCNdkf/iCrSHDxSSHMZZw9d8gyTfM2SG3TtzkYVq//X
jd3hfMoSNz4n1OWHw787G1/12RX/CsKYoiQI5SqFljyWcXYFllgaYGUZOBIEQUX0k1Y6xZOKNTAJ
lH622lldYBVlMCXvPEwA4rpaV8VGelbrtiIkwppjye7tGPlPXQu+nZCd2BjCYyeulJJFmydtTW7G
pWSC33oZvhpiv7+ix6YkAhSjnsN7oWLEtYpz8as5rY0c1n7irHTZ3GqIK9uaHcl00tqZLnGr4tj2
Z4+lpntS1f1KnPjIhhdUQEIpRAAylEDOpCpqDo8WeLpSA099CCzKxml6iE94GRPexiMwodz9rBxk
nZQb2ZLoYoZXlfVFN6bDWN7ea+hBHepht5+W+ZUj5mUsPaHPRIFkI8uwKDvb0lSK1sDITnei1Pm0
+OcjCHLY/oLei515N2l18IqJmgGuXT78pS3cW2biMR6YA+7rjARgWc3SVtP7OCZPlQiyCfTAA4t2
HQuAUwnYdT4nh6eMxaSI8Wfz7wXdRdN4x3QBIU2FiwVGQSv9nLH8VgAoABCak0+XPZVTF3PZxN3i
SmBhvY95k1l29YsrFdnh7dfkLomgaWwAAeMTK7fMZ2prwpqmKLKu7S7m+Kov7CXf9lHyPnUNt6SP
8Z3K8eJEL0Akkl3bgc+N+xGghUu30OWMIuBWTdNxjs7ATirAWqBWbboZZ4pM1IZsLbJ27g66Fu/f
8KMkd32ddFOYg5YGeM+v6rCgil6Cm2VDccKGpwxWfFJU2DAuoHunSm+YNJUFQXuPa+QIMzrZWJkT
A1ZJpt0xKeR5T/wcssdHwXHMavMobYsxQo8xP3cgX0cz6pCSjWKFBF6jEbfUL6obpz+nemIbc94p
AaCl4Eg88Fo5cUYyGduEMLuSKacINIBa5suqx5i6O7uPCe98W1V2LVP2YtblT4gJ6jzQ56qg0xxY
J4FG7GCYu/+nPx+/W38yorllkJHyMhfhK9zGtS0kHE8y/Qu9RSSbPcvJ7iOJHoAgCOmXvo1yL35q
kXSZoca8R5yT8xO5GOqzhdSQJg9rmHnWYHfnQAyOYcoBvZur+Ql9LPWrfMYXrcpqiNjUFE6S3Vtt
pGXQzv/MHLykmtei3U7SIu09TBHX6RMo3FNEb42MvsYkYFJC81Q6dHHg7M72XfWsj/S9XTQo6SwC
XkMuZJTRWLALiai2JEvrlw2vkuyY6+TR7fj72b2NdSu5rn+panAlU1S1+A/TTvzh4Us7S8IyPDps
u3r4KxjR9xqW3SP54X+nwdglJYPO2jIPoxZVx00nR4BgC0UVqtSG4Fj3ZBqBQsg8MOhLPtC9x/L4
oTFZjy3K0rwmkyBiEqONmdYfEcRJLMp1ncO66tTj1AljbivtYptKpMKkyn6tz9eoa0fsm+LbY3MX
WXAmHJFJDKzP3fLLC96SBQC2eZR4PIb7F4Oe5Elkf9ZtJJkFeEAzOfhAIN2/BvTT6PMM2WCtDK0j
B1AaH/a24rpQBAaKoHTspxqbnYkxr4E+zFow7DoXSgiB1V5mpsefE959HuNgi+IivXCzw+CcF0Ef
mPcmRZgPz+eE035lIOKYrKW4NnfC1VbxNB6G4iFLhDQjeffmhZLu/hh7JRBDjeqgxR4Y+Z6e8iyI
nayq1JJgnX8TDqLTlfUS0ihWGedxo5rytY2E4ow3Hkyou1+ucg8gVz4bpIlUJ+fa9iXskMjxKmhd
9dHM4KeIeJQ+B6SOMvOMkVW0e9iRZhJferM2n8L1SVdyPF7MnIcTwuEtZRwapSeH/cl6WRyoDuKs
OJ0OCvylpvbxfrHtE1Q0i4NrBCn9AV20/QnWsmYSFjdD0WAmWulihs4KdUAcwNspY7RO0s5QHeyl
VFJ3Celc3CLzTLinXuBlyEx9iDfPkYx6x5Wd3iaBGuC9JwvF2fmpZB5eqkPTAlR045UQSVM7GVB4
pleiJzMfcMBanoGmF1NGNOq+9E4ZBVXpdvEz4N2BclhQaq8rzXSo2ijrktImDnnRZKs1oZRWomc9
XQik6eSyj36Z2dH9BAOMETEecRVpma5xZffwR9GAFPLRdjVBWDJGo/oKB4EQTWnw71G2vt567cgf
PQLFNrUEPbG48TvAeZ+iAroV0vRHJWUV8zoi4Om649z+JqqFTDQ8dsBsNeuaoS6rMNpcu7nX/Wl8
JWfSLFbNR2dJcicuRqyTGeVRq/ZjsQEevnfbWwW+jnfJq1bdRZ1KQ9EvZUGkeewgeHhEhpYXwGLP
04cBtmcIgOAbqzBXHCojcQ9o5QjZlA3/i1JiW7fpXrGqIvOUL4Vk92tM0ZqXy9wQpp5ekEApwXPk
zVGiyiVcmp0E4gRMszDUJL6wfkzlDYgUMW0crEr1tJvE6at9LkkpTwx3Ql+sihvVHuEQqY/VecmG
V5y7GLs3iHVz57KPNou66+cwSME6Zy5jxrFkzXkg0YUtwCFr1BHTgUpVQx8h6mtWz07QxrJdaIN3
yQ5leA1+KxeCLZ2bXSm2itaRFnJlIFDAAKAyqpEP06x2apcW4cYIYW+BUPBxMN1Ik1+p04335Og0
E/tu3V0H54UYSld+/osj/0oqU8BYTjzQtMOLUPI579Ad2pfDUHwY1F+66hnI3PwEczFnCyuC/NwY
v+I6g1L0IxzP43fp2YJd4YJMdNqkNE1tz/EZ6uwaEkmLn1G8Q111hpFCxjuzRA8GpT5q0HX91lP+
EvGLxuLocIWOeoFxDrTYGbeFbgSXmpyFPAaxe77vMvfl7PZ21HpsZBpTdNNe9yTkrqcJTTvavz3y
fd+1UQn845KKdYpgEV4NdX9jsePv4PQhFX889iVOz5djCNe1r7Me4izOeDC6ZIoN0daVAjTgE0C9
jsspQJ4Lk1IK1Cbi+j2Vfl0Kzjp68TJ46v499OKXQ3FPSow1NxraAjzucEu9ga/0JdgNRFXeMyTq
Uq7Jb4MpSkSwKMepQX+gLfhvb+soo0xla3ZdVH0PiLogVZ8ukhwrKwoPy32SvSiPcFX/apZ3wz8s
twKrlSfWcM2fBFExI0/w7xcAnvsqBko5t6gKH7XMfYr/7m1qLciUbbpEl0IPq3x6qYfLZqHfrGoE
aeq6g4z+wRNTJQUT5sFv3t1fL7yg0wfD9A6GEHWVp90Z2x8LQGJiZrvugOp5PycEvFyWoXOli0vQ
Lpe1IGokIgIdBOje00oAzVs3OvK5JDJlcHPsqjntjlo/VPl2CEamOptALZhLBuDUVLSENdOUlrbf
0l/ai1bQSRMh4fww0BYym3rRrq1PVcEafqXfMt8MN1ZhTYPkRtJvB4PQIlCGrh3DVVFuVQyxdaQZ
z9X9gC1wyMpK2/iTAgsQ23PxGX2JW6EEOj9d3fmNkdvUCaQoipnsK+S5GHW4Lk/gINmKK6oVYVnQ
C6Ym8PgO/iVxbddWnk9G8Z3R03hFQxXmhEIEDOUwsUcXnWqbNBZnqa3AivBbDIDj8wX6NF30t6Uq
ZhrpW4S1ca75maJl1bBBwyp7YxG8WDJGbzI8f2hWMBaoK65P3lxvREEWrb1jCPpGgjpgLb/MS7Wp
1MPJrR1ewYXWR75UQ8KFFQvT6ttfyFdaO4Ml+V+M30S4lm2t8w8yVL5RrkF0IZAb/XVOWAe3O58n
czjsr+yrInIA58svPma3PKKhZGzfWSrEgBj0e4SotgCryooZUAAry37I2BsKEwrIEzMgXN1zC3Ye
cFvbjTTx9CIhI1rFsxpndr2n5yfEIoZhElCRNKQnHkizCLQhenFPXSzcAW/siYIYiei2rXhVTJA9
Pyyc+glopg8LUSiLcd45c/pAhxBN9VY8mWQaiu7PoaLpjjcegKN2T6zjGWhu4vqA1G6ExieDq1oA
oVmMqtAkuhEa/Y7Ic3btVx6mpngd19a00vP8tdoG/X5pM/5ikXg8aKaAXOiQXCSEIrtQxBrz2xJ1
47f02bRdI3iIBAQ8YqaL0sc2SrmxXfty1DwgJy9KPbFk6G9VxXMMfELrcPJlTGdPng1sefwJode+
ZlzfG3ZblS0izAH69m8eKVQXjP1m14BWFzvNdmYAD1E7LUj2/ViNKA21l78YfpWb5SlTx3nJIPge
QNE8xSIWU7tioj58viMa1FgRc1x+IfwY1+C05TPdz3fkSqJTXVFLF8lJAd61NtK3Qti909/cFeoD
5+5QEZP9G+hC4QglmDVJrcsQKdBHoJc4vmQXSXEkY3oiLZQQG2/HMftLm5zjR1G6XpvI/mO2Eq5z
CHxt/IBDl2g66jQ7DMVb4hUxXNZuSucQULYX2EStKq/lMy81oFRbrzuScWTb1sL4G13z9sznW1VK
pLPoWBptyB8MzgmK1kyqD1Wv6rKyCfjRTEfvUEs+Ef16IEbq6NW7NzxGvrlK+G0idfl/lxWJKtrW
0xE7MGaZtpp/+XlZVu0o5GAstJX3HebZc1vBNngLjqrN8SZy6mk1C7RC5n90K41ukof8/2+fnTWj
O26s9M8TVtvQyqqnO0MAoOMXRVT0X3PrbkKmv0cmXvMJP6v9XiNPYMd0gFN9xF0HBKhbC+NePvSV
bRG0r19p0Q7OgKthlvM1OPNx2ayPqqPK3ywJ7KIwR+c36t1FAFk8QIdMdMRpnKoe7NUeIqUIGCtE
B1xzKqAvNydooGJKHA0XNatenFna3Fcy23gU+SF8r2eYAM+ErPt0jrp1G0PSRxrJTaF9kDfhsTEU
2blQvyreggdS+V8dMfeRJooq49g6dk1VjOnqon9Z0uIZjwTFO6lbB1kPl6MC5bM6Oebs9IC47sgz
ObqpJx9CkxIyuQpPgyk0zXmSslrO0FfzigffiM9KvNLmUomC0V4J69DSkVlk/ADfCTiE4J/EJSxW
D2o9rhHetWxJ2GUqbhcwKtnymRdnIZl83hvKOAcEDhBjJdcGaZM53JzOWUf5vguX+sJWNQz52Gsf
unbvBfMJm1f5A9LJLtZqpV2+y/jdr/2Lye0Qu/yK75HoOwmPfEbryfGSfJLikN7F4hUqiqVu9sb8
JvGTDdNSXf5Ciu13GdMTXZHcdpS2pFw1Kzgf87oYKMvnBEXVHvTaTKWf7c62sLj5hg7RGUECeys/
cCf0NTkvTJ7gcqcRR3lWYS6p6lqociYLNsRzd6jDX6DgfpmaZ96qj5I0B7nQGQy+OOQ1jtjOFn84
9lkcO2NMUt0NLLsL6AuzuMsW30bqAW3SRQ3SVD4mA7xIvmD9e6Zg7a6RTzOzeWPWLru5d3wcVaQp
LaWUbY+lNW2AQVOlw3kCxlseviFgmeTWONJvJDoB6A0KXIC7y0zdIk7/y6HLF4O+l/Z3yoDGkU8Y
JkUHoLytcC6v/UA3lGOi4OZ/1b+19ARHgzoR18Tk56FQEfbp4Y0NFb/zutDZD3gckDYegWHqoYxg
aPKBUmVliO+OlRintYp7FH4i4dybzZDTNJ7F2K3GyjxxAZYV0WRH4ce9FE8y+sMgLj/FobYBYyF4
rVuYkCmTZOIbQ7/HA2kSXB21+Uzq8mPHzo3bUQZZS9o3c362WaZ/0XjY4DmQxYTBNK06yPckSqji
DAy9DyKt9lCDjJftGWbg7OENQXR1vg+gXvDulXAbj82qg9CCBACU0xbNgMAZipeVSyGHPtDzwbjA
KXooxuk6j1vVccmPYfC7J0BzcKGBDQ44aO3zjAE35KbttgfaK0mOnvFb92vPz+pR8keaVui1vm5e
cIOCAtObj+vtbk+aM3859jd6KJubDkkpNUv0jUWbq/yr0DIpYJaxg58Vh+qkMoS505Jg3zQ3zidf
YtZhhhYIySn3o57+dEZ1VewL93sNymliNWkM+bBYncfVdxrbBLsrBEmIxoONxCV4dNrXqBY1EzXK
EZmh9XGa0B9PUzI+RWWB+aqal2LSeV8bImizykhi8LN1MCQHcJay+YoTJ/bJqgbUE2DAi2Uq/HpP
rOY87O/VIcOkEkF1jaYjDROAC2DvXlBOs/RMv1ahDf9i5JHI4wfysOcFVO+cT7qJjbkuN0OL1WlR
Qp/7SqEvwhapmdSfXGwPienvp7iPo6L+zokE1hD9s8llY9iZSv0lFH9sajICuXiw0wR4WwDA7ZGP
hFe2Vo+UsXEx2e/eFtO3yuComqZyJ3h1jBL+eYhwYbSVWdvPWOltKW1IhAo6JFLVbvmOgiEbPGZy
nd1kQHtrawYNdXraGDjdGeJ38MnplwW6qC0cNEBVYa6cKS/g9E14staa3AOCjWt9mrb+8Y2axGEA
HBUXscNEFOd9hOdfD7j5Ad81Uk4XIXCOwsXApCXSfNhJ9U31SoD130mVtLEFhpUjVUIIZoMhjzxS
xPfjHaY0S6OteDni2xrICPPhTNVocqTTOume8aSJMgzFO6ZQttMMu6+JZ0uRVpozsxa39HhjLQtw
i1XGw1QO9Ysr9IhB8wLJCs1VE8JpShOjngOwlwQTgIXdr4EmbgAeCHXFcaATDP9prMNuo42HMSgJ
htyaMd5/luTsdn6JhVD13h8d8XyyLhKTh6gMel7LMlsRS3lT8sbfuZsCJcny0mzJAQq9XgRtEG4e
0bJO5/M9UMNYVMwfSqX7GZh8rLeS60bfnLogFelMC46rCJwEX0oH/HUZo+3nWSG1o1W4WBhrnuNM
8taFoS7IemdTlbqJD+RpvZe7kEupCbJlaS8SaXrZmyXL5Cbx3zaVRgW47/7Qxx29tvo7S4b1BB7R
nCCglJF70m2Q1btWjtkl+WhFeVE4c9DFJsFx39fm8l9ycQMBvpzQ8/nOSKxTvpMMykHdocC1cFa0
ri6UWyqRb8hTvuhtX5i79TwuEeR4n5igxo96Vt8kAdNI7EFofQThEtaOaiUKQ46kRQp5Gj2Vo7Co
WRdu1mcDqimdObxyqgKv7k241W8ix5qoL9LGswqYwE/m+higGrv5QXXfcwv0FvZWVdN/SygO1Pe5
pxb/oeerg4xTHXC9n9ywkNRrY2Cf6EMoNaK7zEFNc98eTa9HR1g+CwLIIAywp+xCdDbZHdyIzFyq
SGqHnwMKFytcgRBvJfCgfrhJR1CcXUkDZh+YknztTw4LiYfso5b9Kugif1YiUxQhgOaaXrxMwSlg
5cqDq44hm+DecXfcdamNPv2xVjFWWHyk757ezpN1189mPIyaNRMdmuQ1GG8zViFcJ65MMFQ97qW2
MdtT/Oc/75krT2ldvywb8EjP3dkfDgm1Q/duyYEk7BF31kuxxLpcWiS/Hz4OsbEDG08GHY83/2Ek
nb7DCqpJYG7bOQR6UDbxnBke7AHDsMN46GMpjueEO6cghXSX6bn3KjMglSUVD6sW3Se763E/tRsb
RfWimLry2ZYmr4RcWsgiSqB00rFmQscbSRdoyj9fLvLZuAo0otTOgQwFe78TRtD8jBAH4TPTtzGF
4jOSemoSR/SpDR7bjUjnF4/WrO93PB2UOxC1FGVIWxpWhuzlFT7+t026QdbBiSEDyH1dRfcvAOpB
+YYpBD5nNDFPT4a2e69shtgvMxB3UZJmvUAXwJrj7rfRzE/LsowTdeUTtDCK3c7M+/m4463VUQF8
loKf2SaAGuygfHC4E2Vg/f6ued/C4QkdYdVrUutYJxjVSt2savaozrpcJ13hmz3uA4mUWLLva7dD
eYNnvGum525mFyDaxJI8arYsJgNXgo8GCuNSDa4msnJKnJ/R/QkTpsi/QjZ+WhpbWneKZ8JVuwfO
x+b5xpShIZg5hCQkuabNvAK1kBOHMmIrE292k8ePUU6JbuJ6SKDILVg7Y1uCo2EI90iK93zJHTIq
2mPQEWqZ0/3oROyYPPQAPF98eY2kDvCiFY/9oC+ZG9s32Hmg+T8Jxa4u/tybbnX5Jd1hl4IRRmxl
FRnwQJbpEwYXNVB8MUku2ng3b5kKr2A8oT+sqnH0GkN8OIjSljKXlXMRkiMXuascCzWqvf+zkgJU
Beu5/7EojGECNCz8SaiezzFV5zhNNhXN474XBl8D13NLHLzFR7i3HLaqmxhh8ZdajZGJt0zuh6ea
SXpYvrKK+eatMIa7wISfzgu20AAhQS8UX/dA7jIxJd/ZdqXGeYzG4SVvT8CrVZIDoE2+rGXJYEst
hkEDKxDmyiPBLn5shYRJNoS/9qkmSmipiD57sF0rDEPHZ9eu6i8bOuXj8khCX1njFTEDHZJKvf/w
7Td7l6PBQiWBJGkJVPE4LvJeSA6wl3V5bLYnxV1pPYMLLjQMdWiwxbvpQbRMVVHAcdW//Wym/ofX
R0nQif27vi46tsL+cxI6Nv2OVFUwhQ+gMTK0SkRpwNB/XRgrBOd6Nxe4F73wGAi249wWbjpq5zxD
FHsWPirXSHsJi3N104UVjgZYhytLENmkLR/WxIeIJ7FUFAPk8rurOxG7yDwNvZPYFAzltVr3dm1T
k/PhXGdDmxflDku/jTn+rS6/qIp0Fz+4PHkmdY6Y3dc/QGcou7GxmFdkVBaGnBKXsoSH3OVvqQJM
SNMeR/xMG48lIUmbO0sppjcygLEQA1vsDDMAL9GHPq66R1QgGxtU+uBadYWx6oLQcgeI1H9Y7uGw
n9zcsQPxRYHBw8SWbxm8hQrqwlE88dT+V5QbBtBx6TbVh2CWvbGH1fiLESdl9o+HEQU/AMHZZS6+
wO/GcBu+6PGmashmGqp3qAwDdhdYfmviZx7+1HpdmFl6VWp0y1N+ZhfF3O9D4PpTMjwN+PVX84e7
7HwjQb/VotMKqm4jSfGmyr5saau34daGGfuKNbOqj1R6idESJrJ2dTFJU9Q0pjB18eHINHxKvMcK
MrJdLG42olzdk54xOZZg19V+qUMYYbH8V74wlKBt5Y8w16sz9+obTecGYmS4CuHq8zwjF04UgX8e
fMgBOSZMG8oaffGQ/bjs6xLXD2kDTnT2btNaixvIVJ1kvS4d5DpXS1JGs9vR6Vyf8YLstec2eDXl
XiXbZD70r1qBY8xkJzGbGmyVtyl5vfKvfy2gRI7rc6ZtZ5+XF6UYtFeFx2LucRRSq/PqeJ13rdzp
2dZMCciAMF78q7Q7vOPfeZJGIsyzG+fDsLP16guXBKgc7Mzmu0B2h8VDXGiz+LbGFtTLARkhceUq
7TNVQzSGKdQL72n/JV16HXRkwhgAYC3Yxi+BX/u2I5XgXsjNUSHFSB2UihGCY4fnkG6BoLNFOBwi
m6x5QaX3cwaHMfsjNkAabot94vNWqZ3yj4Cr0v5k7uVnpdBRWu9zE6oAQ7yWJ+w1NISGpuZdeIuJ
WuTc+dpCB7/sQqoWXNZ7qZvqBX64VxZRTDsZRtxWxAbYOqG8IgvtN/BDHtd1sxAnw0GDJjCj4P2Y
FsjvxBCr7iyOwfKtssFt3b+DKVaRtK8bkkvp0CB1IuysBWKXmdDWQnkuv4zJFmyClUGkNs7H2KlK
IqjVvtiSTGP93yt/sKda9tzoF4Vt5o8eiz48Iybbw5/mXYTQi9EhiFQgPhT5iiskcmKtj/qFCayN
tzUk9t8r5oEdJsbclgsIScUGJUoK7XYr3L5rd3UWMQHEDRql/k9l9oFATkhTKReTPgMWjKZVvKJe
cg11U630hePsegtkm/QvZT4on3rXySYqxBubPkxs1wfD+8ju6e1iHKH4XQnDr6z8R0SHe9gM1k4k
7bJIZ6F5I44J5IJ46df7p5DT6wGdUsWvsfylrRKIAtDJzp3LXMfES+NqIGthOtf/ni++yEf8jVYb
z+F4UZW8QkK9oyuOOMHegKayBWesAn1FZOsAD5ghpNhau8RnLx7SrmBQmkUA+DnjTw7l9AujP3iO
Xi459nJVxic9bdQnhGrYlPFb2TczMk4uI/g2+AtYwLtveUrSR6hB86SVSJMU0F43Is5iMKXwPXLn
qxbtAR4qvyoAlgRlyqMOob7wNse2UIHWDRRioe6Del+jboWD5N1bD/FAzYcTVuIy1rQWgFeKNsY+
BMjop1ckJ8vcu2xD7ZKJam9cjFb6SccK6MElVJQqrI81gsvbfNzmsu0vOYGbnP1O6po1z9ptOE4C
XhlvqAbYmb79cfVhHGa96fs0bsIfl41ObKtUvQYI685pGIpdMvqqGdH6kghF9EiMyfgoQai5FSk5
ybdt3uII4r9tMowHIpP63YVCOLUQvluQJhW4K7kc+h4/OwPVURbApgezfAP14GDziuWd+JlCa5/q
LAf5uhSfWiaADuoBLYnXz+p2UDGKRvpxv5gc6b4Nj7rz4z8HU3t/+sq9m+ad+SdKUgnv9sQu9l+S
QoDJtLbwJxuRaRKtQ7tUCbHolxRDHUB3KispY/E5cT+gQ+j3f6nIQc87qTmoy65rpgMvN9zr1oHv
v31dSZNrKpVnLYWQ0ekjgCMF6BsJwVEOD0YjNN0AFbQKPaEfoyzuh2MuTQBeZWTchbF7PsHbY4yY
v06JLnaAFK64+G8jvGZLv5ZvATOe/dm/a+WDy0/c3E/bsB83Mfbz70Mu8PTGjSPFXTPw3fMz9XfF
ZgNnnAL0hPkzw94cor83ezmQIIWWTncYgv2p2+svUYuAv1pH/PMm6Ng3CHXqOSeIsvfYfSg+cZho
ZIlI6kNlRW0ZJgMt9KQv16a0GoJ9Sif51jL17cwkdVjwNN9hrHQVwPU2S5vCHp7kfWeysrjD/s9d
YSkETdyq0iz/cLUAqy34kofFsaaOu5NVwZ4N/qAktXi7sN6JpA8JU226f3EAgvmKOgRS0II+CGaN
I6iwsrVseghEaKtHjAX43sPDKn6Go5SF+eNKkJ5sRLHxygMwISRNIS7V9AEz/98NB5rOTTZcUw9D
fK2xhbMvIdaSZhbXAcEpCF+oZh0ZeS9lFuPOc9Is1udjGvIxTWcc8X4UK2GI7pYp8trZxGkSLiux
JqZzgCRMUd39m24S3o9cGikHt6WwPNwly3DKKug+MxB7BOTncHpa9s9S+15l+qZ9mOY6MILpP91t
kay5bdDpvkJInVjJEuViQ+TfYmXlBC031oZ9/R48OJCsOxfvEpMXN+Y4buM2LDkpfMPCGmPsl499
aa5B3I9vIQemrTaHd0fX5yUvlHbjT7YsDLL6Cstv+3yjBDAy3vqgkqnZmDmFemq8pMZecfHGQFDJ
qWoV+TF4fzRde44yRCtaRbqlz5nNmwUiFexgDP1fun/IG3gWRHilUaffX/MagxqKrg5fGtqFBMCs
Bw62IsyI756pA5X3EBc0wD3BJskBy229wcOXd96gy3bzab/2bHocvt+dKyskAZe4x3OF18WM7kN2
7M4Tf9xWcNMMO3MbPtxXJ/sd5fOJdB3wThalZdMj54eg5EXujPAaM9cGYjsS/+VfVHrmn1W2PKyW
1s4zl4xdg6Xtx9RStabQB7pBzJR9Ikz/2tRXTKsLSFa8rEHuABcVKq+pYnRz/CTZ84g3ZRxPGbOv
hNahlWI17PRVJiel2vkov9Eb/XOZglxU1mOpVP75XFjzWAN1hTHD/R9ryhYii5zQescJLhKuo672
4xHV7Zsxmw6/LKIY4fghzCY4bGdrHW0bhYGk+Dy/qCm4G78cr1eIisRzjzPok1ZHOylxDD+PG8vw
gvPAfhhweYIUnKEK2ovb+khNkSH+a/R83WIkFCDpOt/5d2xmqGF1wcihIcEJ3nKMWr8Ticu0GQvg
0lJWgGgoUrP08C4ngMDdJKNQYHVrsFysZUhADqIEIamisLVp43UYB0ivGFVL1MtiwGA7jQkaM/Vo
1Rl7XVjQ0cO1SAjds0rvYmKzJdahq9ic87wxFSqXnfbWHVfCbSsv003tOex7gCdPZt8uNz2CQ7JQ
WLGXsTk/PgJl8h8r2L/tRIb1Ey/s+M/1GcfOeOo7stBm86fn04eMCd21Ttvu6q+UU+Bnoa4Mlq+F
5tNQvyYMw9CK6Oq76J3MlVQ7qo9f9bIzrJpdktse7luVtrRVjrPlVLDEwLIhPZQciz3kdhdv22zb
/BPNYpGVrX6VXlMb/joRmjR3jYfmDIeBEBxMG6bF9csxC/X3bkvmTgIopRq47r4ogrKN9hPWpsYT
SBRhmyE/jnoVabJrObQgR6nszIi9b3ccAe7e7BrDNSatiUcuLtxWjq8ComS5s9JLEcs1Runw41No
2fnNiE972nCMhLDwlUA3htiIQRqd94myi3/XxC4PHL8rp3t9RtqXhhqD8RDv3QEmo2kk88egd7P5
ys2TahXpY3hsgVpXTaZojMSAgRz/QgHG6DCWqaxEVP6xGPiMXuIbtw8gl5Xpg6w4DUnPBR7oJjx5
qAbn+/H/kSA0lSDP30j/UbW9D5GxCPEnRYfmXgfryYAIWGOraDAzdo95aVBqzxLO8lK3n3v2AkKR
Mv9ZbLFa696D1ctfo53fmnBsr/JpG3YxAsKhdFe1uhyBp8DSN4s/bTKsqSbI7xLqkNSSPO+wMFLn
aCpDzCzbzTZmOCIc6QANLRoVS2jkmg1f6SNSdPJyEM/cT8o7zZGc9FHpieJQ+0vwNxt/6HpNXg5n
DAqlBDD9CdxFESvoF/PbJrAuH8AE/nC542dHDNhRyaB9uduO/yJuhV0nDcVPDCMOF5q8Q5+ObT4i
8N1m086vgfnFXEiuQ2q2l4NNtaaNIyrXHPoSTzRagfkYcvddfG8Lq8m2tqDjYeseiFmCJk4+DfdA
fUirFVDDww/CGsiz9Rj6E8yHFD9zVKV9kOvhf5vkDvf1Rh/FxS3N6XUiaTGcWvCUvaHk2oo7Lurg
qA8SoqeOp0XNICV47bLPeEnWtFKqeks/282/ouclRmcVNPQ9YJhk2gTSQOeWqEpBa535m3kt6xrp
dJlo7aLRRE51YcLS9E7Q3CIBWcAY1S1IV+GDxoD/BUTE4DukkDHVkJaS4tEtBGSsppvXTZlTdKA7
VlGiuCKGWAshS725DBsudSwvVcbfzFFDDnz+OC/22pk+zbyH+Uh1NsDcWE5J0+sgNMjH7wpn1Udu
SvdEHLyCrByqRuORW3YBMSkoLoyxl/n88BEjgrHLXpVuQ4YtLqF987Qc75kMxTalkkDerbKHJkmS
HWIKwxDeT6nR7BXFnu6LYMwN0lDzr/IAgYHcbRlQTSr+MytZzk0FiJNnRmEuRKZDJ06DbNJgAQPf
6nkyZC5uF5FAvr6KeJrUvVfLTinNyNC8rGw78Ogpk3H4qw+/MJe5yF2G0UuIo+Ln5DbdIz6NtNwf
Ypg15XL78d3k3pCgh5GJ343j67RXlNqcwmAbjMpEq0010BMrPGa01Ta8j3W+TpJjcEMljPCmx/c4
vRtRsv9hJzjq5QCy62gOThlvnPXbrugI0ZZjpLPUxxFqPZeu5yK+tWSLm73hVIZCluZW1KcJVwLG
PvXLo/exH2ykcOmLAAM+4KBBQlRJ7y+1jW3LqvnfzyM0Q0JzJJSRFTLVC2x+uJRO/SoSyuyXj/OZ
rtcWOI+O3EW0EDLB5fu4VaGxLqSpEMcowKMQz9v+GRR7wBesuI4AlUvZ63hFVz7d7QnAo4gBwsaR
xezyGHL1U/jmwsIbWwb/UM+xqWayhmU5RtCF8SrgHRpzyYSl/bRzYUMZ9yfPqQoLs6HZIqOLMqzb
OREV+kHi/d9r21pk9vS4pgnYsPS3jD1ks0aoVCq3L5a8uPdOsFalhy8xVmDzFB1+xsE9/EqPMD81
PHa4jwE5mlYqAt7P72JZrf5fU8Ymt5SVX5DcO4SKbBEQ+9i4pubF+u7DkNe71hs5y+dmwiyO4qIO
kzn3CRXnqXaYDhVZNX88mmlg/o8UJAFyOWO0N4Uz2ceuOa+4EZEN4EonGi6DdWW6QwLqxnUiIA2A
dUlelHOLS+skI1/Y64AHDB74rXFrWEPgsYsfQVKq7X/v5/sF4+J6LErHJ0UBir3V9lXjvTvYBhEk
bhw+nP3WdawpZmZ6LuwkdMLKoWxop/nRmPkENB70e/UBU6GRzvyn55X8uipzYI1HGw687RUUHqB8
+qtZWS3zcYP6HxgbzJvrejvFywyy2ryq4W4rcuK3mmvMSx5oYDKg4rq3Ok03Z7Jr2XBn5qFm6J3o
VKFsqQZsmzOpvtBBz6Ih4xikc2Mtcl2FjXJWntK+iesuKgHwlOF/UklsaX6T9WRH/MifLv11tvdr
KnjDP7cVFTRYMi1QG02TwcSgzkqkK/p6ZsG12wE1guLzF/Ze+fhS6P2qdELTrDGYSOEL189/Nz4E
dbFbXbTfKAHgGJ3NQ5YGRyroXjbcP6K9izzQr72jCodDvypgGVRAPuY2m2u66nuH0n4AmLTi2zkA
ZcW+x4pN64wWfZm0oWLGSudkHy54H32FLY++vlF5dIhMyhzF1DIUOgv6iA7v7dT+eUrtpBj7xntW
9R5N23vKSzWuumUyer5BMqyZi0HOopAsmaGYzQ+S0uRmp4+C5QEZHxXSCrXL5FsyauOtrtt5wsUk
awjMdWn/LOJnfhamA96wlOzNSZKPV+P8sPvlLfngaz7QoCo8VOVDnaXd8OfaT6ZD4vWGAF5nGPFw
+rBkV/Lbr2jFX7yLnDwhYoFWgAMjgBCSWF+hfCJ2G3LRV23E6aNVT4zMNMKAy92cFJwXgL4WqQD9
Lu/9Aps7i7oHyzMHwhnkW2DlWFSx7+TDmocpm9mssHgXfDYVczXZAdwXabdhi+h7g1fdC9lSu7sU
kIC51znEGITCuHlH0Qil6n22+b9fnqpWP5bRQPyPpb3Mn5Q6+ebPAldKes1tMKYxUu1yCtIplzI1
2YHbYEdBIbuADWJyeM6EwN6+AzctBurQOKT0K0KFJMYQoG95w0QhrH3hKiGxlGgqHfcu0GBbNDwe
Q7S1lU4x+AjAfAZbbhWKiUF3LhfW3dy/LSGoHbeLrL36VY9Zm3nhVgMeet//BYSIKWZZb2EaJIU1
5/oApyopD0ejaJ5bybHDwVTNK8TpbTi3xPbi8UxY3p079pFckJz0NgMZP5KbElQymngf11/UNLpk
iZjrISubh5ymi+Fo6ba0JbdkI8y4AvHi8pnOrNNTOKs+pLrPeiU4ssQUu0BU1+sbUKEDA+pLFcJv
Qmkiuc/QNxRe+Zxb7UkhfL4yshtwwqwsJlyqECU+4ykSgpxy2D+26OByaesBQQNIvTo5Bg4msg02
pHmsiqTla8R1aUpY/QTYyJZLwjK5xogzcz5d3udIs5r8VIE4hBZt+6lBJT65N3noD93GYtlMH9Z/
wlTjjAfhySWklY1zW3I1yMA2dp7qDxUmfeE0B4LVcxTj19g4D4DM2lOsmGLSCUamni+7RGh0VzQn
ABpBfNBSyx+BnhUEJJdfiN4kFnecs1tC1Nj1D4iOGuQXbfEki1t86o4tYOQBT8zU85bAvuaHzyOJ
Og9pPtv4d5Pgitrleip9y/4VGgNOJNL3sD/bWhVKdh1tiPlRqMqi9d5BYg0UFnhSLe3lUrg4Jzvb
E0sxTmhw1+l7AXKDKDvuPYwQ+ILE2kynw+sLQ8lzdxUerleLeQegmTGCaefImaqpyA7dSTQa2e6i
MzZYQdzb6D5sIh6fN0yvrSeyY2LVpMkoz6uouKC0eO8QIU9cUBEXqDEJ+osI39Fx8Q+mN0oWMYq/
9G7Guj2vrJCiw28QdU8qr9TQnotM7U0iuTAb298mxMdrtokG9LJfLwF6fMHSXYRGdXGMnlYrPZ5V
Htynk0J7/jmearSKA38zVjaPtLrY982/tqYS1FWedo2W7jKmwIsoS3mXaX2fj8CGtxfdPSK7E1nU
cJiEvDa3u/+XN3KX2GJL//wqYD67ayDvNVa3VloAEWMGY8Ck4S+xSDKsJZvdmcmLHfztgU60QvFx
CpF3bXRF6QpEKbz+HZXL12ll6ZvqdS4kiLyalzBcKN0Kueeu//lSCSIbk/6PuhrECRtP4agXALHI
aOsES28cKEhbP0hWdbC5bRAW9X1FKPXxQza/kv1bauoGPUww2yTWwK62laaW2lYxZW2ouP929wTL
lXn1mry821Hes5/NjcoXjAmhVzGZWePBkgYT5wFcpokxoAFKNO9zkYEIfssPZyY1QPlhUd7mcgAW
EcT9CBXrvCyKHovxMoEissN4aVz7scOjZBAwkfd8YzMH+tlh02EVirsPe1ogcd4MhTnVrZYMfB7k
sAzXo+aaHd+cZhal0KGomW4sDS/LjxkgAXEJwoVBi9c3m4EzHwrac6eTJRYwdh90e9IBj7xx+Tks
14t2+DorCU3nHDzRJqUz46d2mbYp5T75e3ILh6EV449nzfdowZHJbmFlTKrtuTwCTNiEojE6IZId
oXjYOmCrjAXNlNueR+wmtazlaw7hDoHomlqNDXTmwcY9y2dXBRtd/XLdNiW5+GrfJKjT7iMMpar3
OYIhD4LkMsTxw1IVixrWUqDGnbhWbZPLQY3YfNtuW6EpBESlN8yR+dGv6UaVeEL3VMH3T4y2uc4o
JD2ko2TdyKXfLFcR6FzwCZZzx8zqxtWyot0rrzgqP+kO8xz+EXVI/w1qVoE0eCWOVmw9cpq0yct3
//pGP2VgCEL0ksjTtWMX2jGRQxNsKAxkjGhkgoa8Dbnl+PgSfHKmoAL9yNM/kM9VSkRHfExpxBzP
dSqhxssdCtjOHPZJTPQ3L1furD1o02iaGQ3kyZpF6+uSGgUPFgN6yJoMYRvZ1wMOtTrATlEfVq/7
OEyda/er3layo9sEc+SQ8QDEkJBbAimewd1U8S61y18WrRH/VmUO+AJdFq1WvreVqGMnHMcp7T+I
b9J2YT4gYXNAzVuGTpAgCwlFo20W2SGAzGalrlFBPktrkaywLBStvtuSiqfMUMI2bePM3VAXkn3x
okUn9akKNGHaftCR+prey5QQyy92pw7ux+b45gtdZL7k6BH49ir15uNFNFm9VMUBvqbODq+RA00s
6GMx6NMCf1BMnkEgU2rZSON+raXgeNutDRDkTjmrrJI0iy2giS+YP1exxgtqd3oAUvmN3CQu1W34
eHL7yfhi0Sm7Be5KxTDufcGconsSMLt7Q8Qy+EGaW84YC9GBKwg0cUAYJos51P0RVZ3gPYVooEO7
Cu6q+l6fuYeKaGZvBRnD6cq8AMQgw7SGHMEeRPesuG5n1/h8EUW1YizdajLPQdmuo6B0oSTx7Pi/
38RwJsyfVSRE1TUb/2bN3qCLYGl/tHSo7HSq23NekGp7hLP50UDZ22Gxfk/cqrD2erwtR7m0A8/C
cZauIVLfKhqQ5eAFvEup9rFAil3WhB/d/5AS/WkhJY1PLN8zWOhllO6LNv+dOZTji0hpUFMvxxPm
mQ/PZ4p6gFn2+kcCISWAZ0MyNKLZgo2kEapgWkCRpCprn4eEc3J7ysSdSfzD2p4O47OghjLPWonE
1TmJALR6OPXO+VKZ57mzyutHgbU+deRQ47k4xRTwI/VgsddN9Qy5XlRfIXdCOADTH4/p8SxFH86l
Gtghbmc0cLDB63J0GdF6ZrRzKI6IN1vPIoFM9yrxAIvik344zyrZjN8cL8xiHYt2IASbKkeDuWqp
oJxPUIJc9C+rg+KMmhVIWtLZjBZtfZmtCIuWHOuNTaPYDtlWPZwoHJs1yUtyHemEo4l+5K8k4KTA
PaWVoYHTIkEPXn1cq8gZ8OeBGabcLw4heoC6/ydx3FtVBLbNQlNyy7P6VIarfGNtgOMKiJmsxXsE
2HGtRB7nn41DZ357fvaa1NFVMqEdNuKSUOKBuJS9tQSnYHGrVl9jojLZxF5FzypxXxcL+lkh/vQ0
o3vnq3wi24M7AD6ZtOV/3Oj1b5sFC8fviWpabZKInW7Y2xLhxraKGxip/qvh12lXqqmZnkqDjABX
+RReEQTMkAj6MEjUSOq+Ai+MoOmt8PhMn7T6MDNKiKZxXatY03tF627VKV/jk1+jSM80IoBT1avj
XDDYKMSU8PFMLJ5SZjhK2yzfySgNzPAxfAZIVz5pnlNOM6/sAugJdjysgWA1TW4c7nPlpQod2ZWI
HZylUKzkjP3mP6HlmcR0bCl+8tPS5HZM5lSRfjY9XonFZXMpd2GWqrm4BFzRjkAX7hj/yACfry5o
BwlJK2udU+R5LUJ4ENE1rd9zDsAJxSL+8Drm3yjBkrPttVWTMnBQa2q3mfKXwoE4wMUuZdejh3FT
p7zy049J30FnQ7pQrIwF/faMTKKAUBkUyGVgncOul9AtqyPVWIAJf4FIjckmaQJDebc7y9bmnedh
PORSvKqtZvVBiJBX6SJdqTXT9xOkD1q8EKedFnh9GhiTrwMctKjGlLpmwjkYm0AjsEopq295sKK1
HBg61VV9RlmNx2V19X+4BR40Zs/HawzFXFnK6yP2+NAkeE4F3e098UfV2aYPiUL3FIljbmlZXeXp
CzGtJF0sh81fEeR3pee2itC0egQNh8a709j8daKAWZ9brZO+jaUstmv532Vo4ER02O058h7d+DTS
ttmCprgpDz0DHngJTM/ebhXTALYyQwwRuyRhBC3tqmlHIX6lxexDvPP1CTx7F8SemW+so8HgTMtg
fGHZqoK0elnLyIvIfuFtvwGq92uJ2zI7Q8t6vcDkFm3Oc97WYqpESnyXXTjNKllkHF2YJJiQEGYI
4O0BY3BkXSi1x3FWcUSW4tA7uN1niBPpEBLu1ohvRGKdklpXT4sokDylsqWR8JGmAiN/T/h5EHXm
YUXEly7ogtF3nLhpaXp8nRIn5cPIoIR54GskCObk8PSOB59dN/cdmxv+2ZqS+SyUX4yvvgfhYaRy
lWXIm0YB757k04cbMQWeVf3zFnT+nHlETEoB3DHqeQeaVTmQvTkKVpZOyYSSLyrx+Z+kLxZM5/Ty
y439rfw0Gol7aMFsS9eTr9AY1H5W0f/+oXqliS6RyjforlVqyR7lxWr3ZjrOXZSwcUnyCoGrrBM1
BVbdSrgaUb315VE9QYPwvJgdxZZ7P6yVNlSVZJlW61sitvSMu7taiTRyS0daJge5g0sol+jQu0BG
kNagqdi2fhr7qFomQ47lv/6Hep1XVUmWedodUPrxaXppLQvRGAP/NK2/+2HTHg2IKNl70ghy9na1
jCrNaGQNHsGFV8M3WbtzdqZbtKRnI0LuMWIiaDchutl0kVZYnYK+4z8wCChnk3FR42FM4Xhea1L3
wvf11U8C0eLsZrTYb6Enb9Ohkv0dDiQtUYLCQ4xipHNeO/futPizYyzO+4+Ly1bec8IfKXT6sZyB
3k6EdYzawY+9xsywau7xa4bNZaoTY4KYjFH9EguPla0lKcxf7rfA3ybDk6swm85JT0B27PQqd56b
jfvtrLuCvIZ6+Pmb8S7RD5+HnMKD531TUIanHDZN9oD2CqsUtKZ1tA75UTSc4HAqPcXXzbYia/qL
WQU4oVLUNi8Q1gzuTFEADfRrVfSZ5ZiPeb2//TYRCdZ0XCdeJYz8yb92xPTAguCx9oF/mBsEKsH0
pTXKL8lC1VbHXoY/k5X8x7iQd7IEgzsXnlyq63zfidAX4io58N2pG3aNTBqvQU+DONXU/8/oureY
7cIww/dY9VtiBDT2O7r5kW2zOfgpt3kS0qSOrmFW263RXjNPPW4tJ+vE1H/XVD9MDtxjtGzN3OFw
SUecicYPEkF6yoAiG2A6iJWsx7Slw8TiT+xQHOt+H+LSe73HPGbT0Ht9w5YC0KJ2OFGnYkz2yxFk
a3WJFeuIsg2OAMlTUw2dIX0aa0eLINz+Tmgwr9CWU8GmFjyBkedet8bKVU0JV1KBWmWMm8yQzUnW
R/KCRW7C9RRKdLQUEugCGRASR9SS4OoKL0SRGliyWpp9O9zSREBsHJEnsai2OMMTUfg3I2ZbZGyn
4EFhTZqsjvKgQKwtiRfkCaNcnrp+BLxpxlD8CjF7Uny9fnCMWqBBG77hc7ljjX3cXaPCnyIOnDFR
pSwuehtRfyM2C6PcYlxI2c5lV8Kilzw1vkfzwuQDJpPc/aqj+aQeIx3BI9u8qvjn84NgLxJC/H9i
FLa5iDe4CkUHHcurQj/fWEHVyIxzoO9BBNdF04jnQXqyrUF21P7CfEV7ZZ9UlTMAEycp7o84Jc+4
VTqfsnFtnlTrbYCWf1OdSVsI0UKRBMv1Hd2CRJW2sPa+Hq0y3XuZV2cYhp7oDf8sjJfi12RP/3QY
aLB00U5EHBjptLyQhLgCLycNriLzZND4e5hilPWnuLwQ2lSKsr/MwB9xSWUcMG6ST3VnK2Oy4bbv
+1aR/+x/s8ufRcyfnVYwHu+uU42INTbbcmOK681OJySvYV7MeZUQLO8Z+lyLvpmoFbdicVkYxipY
TS2VfH6pvTWwVE1tFdIVbxGyyVOH00SAwc4xQ/e0r5CHHvoED3afOOIr42paoy0S/YiliqXNh95R
Qu74Vu5v4sbh42xmaY3f5w9ugOPkaMGPHONV3PufVF5ZEm0VgMltFHrJ+u+Dbh4s53UtJgT/MQua
fJZbizXCNlOz12dSemlfKmg+ZPyeh91ccxAK5jyC+QQlARn9uUm7hjXl7YWEQpYvaG9IJzGOH+R/
9Y4cA3uFIJSUbfOwi0ArDJH6kO7QYU9b0PGOxui7S2sdJIGDJGyTQ9QCJfnEkFwyMEm80nPJoO6M
UDlpRR0cImTC0bN9qAYC67AhLRm17WADpnfgQgJonmbrL2DnrPNBYKXca81d4gDxi2E44IaUFk2v
nNxExX1eiKw8COsgXFrt68Tze43EpWY9Ow6ImnAJ/2nDI9qTz5OCLE5jfywmJZBzEtsqp/yTTAKE
fcAXQ3oMe+vrT2H9QJShCSW6bLWPSOxki08kgOAMbGznCZr4z2gd6FQDK0iySmhgDQCq5USiHSEr
VCJWWdb3eY1POAS6Lvc5qPURy+c4y/1h+jJfo8hIVcnW0Pb1QTOuKH5kBySTlPgF1MfgkdaCcRNm
lG3I4ZZ5QBMypc2BMLDAC3M1nKngAxW+ul08LzVRSTYGeZ59962AbCIvNLnbXn2MAC2l3IxOnsFy
DLFZI7cOap5+r7MBmy2s/KW+u430I6YuIozL3PGO5Rn9EXYzIxj/rFUt5KnmsV2d9tBF5vCBH+De
ajsE80iJiJjKWqJiGQaRNSYOxB5Vk8RP6QTxn8k8gVx2Hn/9/YGBfFfz590bflTzeaUyRBdoZwyN
SArKY0ffmokVqhbzo60foSr1l3N0oEjzFaXKYo5fgEuxNCDPhR3J6X3A9uHIMET6adkR/1IcyLJm
oJiUkracmp9u+ZRQ8BzCnzDDJUZUhNSlyH3Ixoq4DgGQ8VeU3MHdnDOKiF101koHF+RcnII8kHd0
Y2cloiGcMYG293PMkKdXs0RFnE5o5JBYmbcI5ToXw/Ow8c/xRNFCflnVwE2W+fltGoApNxDhH7Vz
33btzJp+lRAATEmbfuHS72ZiXsBqSzkqYK3rPqvuihCeQHGeDPqFYVQCU1bmlSSh/i8tsjo1ajNH
ziAeBfbHq3dbHxMNAUPCi5yjFbdp8EkqP6OT+bHBXxSGl5BudKcW1mzuCcZJcmJrM8nj8AryCOAP
i7EQkz9ZtHXBTRKS2c6S9jq0S2VrRl6Q8CCEF+t1SHsANzR3sCfl7a8tgo8jjdadC0RZ/6aVnFNP
sD0yY+ygrY5G4aZvcPr1yXWbQDNIkrguVagq1/keljOXRkZNFdpUbe0xLEqdubYRoupkj71VBsox
Jyj3PgvtCLqAxEzuZhLYgAnwxeX5n6TaRxslF+RcNoAj5oKA6t9lVaHcld825KZVhJdSKZ/odEW0
deTTedsYu69XMRwKdVBhPF3HHxX49M0vg6frN70JX7iOLAvRtFus43lwiAR2azTC745Brr70qGIN
bNGU10D6GLy9im9NvaeIYypOpud4GzvzibocvoGXLFOrDwuungoTxV9veyTOvXP7m6vmixayvYIh
AWYDSZ1Y5k6n40EvleEMI44czyhYS1W6QmUzXE8xioPvB396vuFYnh2PLNqfoaNRq49Yo6LJqjiy
0lDPSNLs/yAbJbtJqFFmrjyi1y0NTRodrk6/i5Vh/e5fDHeDMVRzbMkAQjveBvWGhdLhuLUcK7YW
pkCYvr5VfvxsGLxb2+icc1LcNm/zpH59T1KDuo4ANNhetFfbUCRKtUMNrfmKErNjV4GT6joUXvmS
Bm03d2WbSSmFLtJBmdrw3InylTDYF4/1v9DCx+q4qBnY3aFdNBIRMJyFhtqRpM1xQE/JdKRVe9mt
L/hw4WYs0yVKGKkWTn60UsSbAhQ1Ho1I/+bimBI0O4ibxesyWQiRm9/kNZ1ffjr+xqPPsQsXmCkS
+O/OHgLVw/X4/2fhEZxKcDxVW3ycV2iWGOHCRNm7+t28/UrLplUA9Koz01Z7uc9r1aUAz6ShQ7bn
n3sSpBfKoRAzltsHrHfYTd/m8NgfVdjelbPMNh/eJuTCR49/uN2EBBZSwT2W2cd9zaPGFrtn6F89
cJmgzP5LTmuLVdfq+h29qa/5Lmpa3KOJkdQvkuqt2QQbB7CDaflteLg8sgpbtUGwKAse6h/EqSH/
Ht/krq1G+2hlgWz4s3xKaDcF/sk2p9D4sYwQOWu/4+IWTA0NYoTtipc7iXtfNjlbkW8lM95WBkjr
l7bOMO8ErQGMyrrpiuH0mgmKDWrdW6aJajT5LoECBt8k5qNbNsKx3XjNNsu9DNxvIG8l3tDb7XAz
Wi9HY2CwvkG1iDw4lE1YvtWD8tGg+jh8a/jFgpaIKLpC/75xwsY6Hs0aw776edztcOa183m895FW
pG99W/E7rr4QjTWiXHcT2NWDCL5MWL+oRo0kitdn4jicA8QV+U/YFCZUHM/FsS3TTXqYw9l7FpUZ
yiukG//7APdJbpInw9Vvsqs+vW9fcLH+C5lb7a9UeAVK/tW/nxmeCEO2lRdS/YGNQkZGIuqwPK5K
nKUBg66rkOuYLFv7895lJh+1CDV1/K89Gxix4w1GSBJD/E9jW+ccofXvlP3BrilYCvg3Y3dzWixD
dokpmJ87Q8aq+ayI+XJziedxyrT/6l/Y13Ur+P2zXLqyoCu0ER2KUIERTde0GOmo0553Kfa6Q7fm
AS3+JD3jBZjqA0492hEI0T7xp4e44Ugi+xm41N47OTw+qCvw8ikgl8Jv3gwlnSXhWQLNXjYRHf7F
ucAS6BwmjKxo6tJe94Lf+Sj+guk+yOnDKxMHmZQXNP3NrsiiVnun87YbH1PBuimOTSXP2BnQS7+i
jhqjXipA85f9wlRdnrdBqHzrLQ+q+ZtUw8SYnX7I7OgKu4AeiGlL97ljeEZWBsghGFr1mU/JFeky
7NaoCmqCNfybFEpPv/fPMAX1EvoP8DY9NOzLo9bF8saSgatLRCp8Ga/icA2QEekk7OhdJyhSNDXs
e+Umo5V/vYUUvHJ7Q6WfYeeaQ1diQgAffEOvru2Ho2jer7I1jgiEbaoDmS4YFBvalW4XEfbTBtv5
27IhQWde7Cy2P1DC3UAXJCvneE4TGX1QUiSK33TF08XQ2cpM6qXIERb9tJUKIwmsYkSSXvpNiGa+
b+0UjwxwBk8O91HuT3+wbwkDtvGzrbDvIr+LDSHM72im89mIS4DrwltbtFd8Z5cM2UR9eAV3UEA+
AEf7koajEfyn+PO/u8ofPlpUk+y0uuqI4d5TSzhBOnNz5vG5DfH3i1YEk5XYsjj4BmFjaLNho79S
Os6EJPyrUQRsd2DWGfnGUyk1S3AWaRGr3I8xYoKMMELYjRUqUjr2ty1Dm9eyxR/uRGNsvP9IHxrX
bO/io4fNwv7GwcnYvvw3uf5pdRP5Ng+1CBORY8nLlHfar9H44VzMi+bHKJQbZn8+pRHxtVRGpY4c
Lvj1X1yQnlmen4xQTp7u3eve7YBIBOtZ6hGmMFHrjnUYMsk/I0j4za3hZgWSt6liIY5tUmrIUTBv
CGfYq3q4/sRxUQDjFeNM5EH75Zf+/8zc1GESG5u95qRk4Piz61QFl5oRo1neu1wu8Ux2KxjirigH
SKVFXaz0q/As1UdOMD2aWQNvwPDrdguQpLM7YFBEq1Ia84fFsP6VgduAQEr5J36fk5/kObpjcOfX
S42QqJqlRGsyPc9j3juAwE40WfdX6OvhyzH00ElgeB+6rEFaV8i1L3tFxnjJ0euHW4g2r+h2POTt
5b1MyUK7Qp7FU3Ynwq2DZTMd4EpQZ0pKTF1XP2vJo7/bJPKUkTZLFBo4TQScV3Z911rpSQvQUFbH
H1orqZIc5Awe0bnuCoIJ743DaOehRLlmO0NgsbZf8qHei9oco7D+rFnJ26yDEJ8at1ZPp1M5URQh
q5rOAb9zTFTCKoGG1sSAYqZwpcsZYKK/roI2VDC4xAnIkgNr5txNDPqj8/5wAdzMMg2WnDZjwHVL
JQRbxOCTdNsXuR4gMGzr7UQQjd6U4MHgpKm/R0DZ41dbckk7V29OCp3AS3NkxaD+OkORV2rluDFO
gIiQ2Hj5xRnkggczDYiI+ScqFy77PuCrHDaY67wsNw+clemTgmWiXQgXVcpeRdu5FVU74k7+yFFz
+GFqVLzG7Fyp6SxvRHq63aGcjEf18YP95CphFgLWukrOtqZ2aksqQWvi0MAr9/wMHnBgyAIEUfPS
uT8r2pdDxW4pLRC12MQ5aIrdRrmfu/1KFalr1EzqRFY0MKEYAcphadfwTkPlPgZHZdEXjoLZqZZJ
h2jHrM28n5FLxFOa0vcODevq/dWFR4lQT08Bjc3WWgQ9VqjhVNp8R8k5bdNacb71+nrU5b95WgTm
nWnurPK2v2NOUagKvRuOY6e5jgyuArQ7fRc/1K8cnGR16ZfdIJ5SauwhfWrULOjpXGVp32Wrj3X7
pDz3rqhyorpCEG17U0AVMb8fV6QSJL1jUUO8rlYEBthov20uxnaunkWMC3oItkuHOQ7+zs2eKEL9
KbW6CtaLy3Q62nwNls+Qb9XSF945VGvZ5S0HJ9ysU6ECxEG+rGpkFrT5WFoBVGpCQOgUPQiZp2UY
fueIr/GqtMccHy2RQ7FIB0qHMfUzF3HW1OnpNGZ9SFz/qf51WaTo04K0Y2gdzlxx7PSWOlYsp6gj
sVS7bErrVzPIMFu0uThIjZEbtxWuDk4bPDHBJUbS2eysFplm1opREJusFuCLyPskzEISCuxQTBlh
sRYGonqdmlPxF02/wH59YeWHQda2YpaABBqRfFYsTpXgWeQHoxVM7siUvZeAy41cgdjEal1ap3BY
h6J48thSEEIyxXYjy9s0/jn4NzwGJiiDh9k0OeV6uFU1StXOgWqla8QmfVrr0IKilAYXFIV+DGDN
sKVjX6Y1FHEANqcTGf4wJDPIIDf6bFdSbuOXrChfhmUc/io9lotPXhbGTRjO22cCtJuZzzPbmrkV
STQgKYkqIp6aiaCUwdUt5vHiNRML2Dn+Lmjt/JK/pK/xEbouLupXQDoUsb9ue5YxaIyzWTmfXRsG
K7xkYOK5ACc+G0oyReum6334/zYscQwiBQRKABj/jTfrfRWCqyTj0kcBb9NBuc1Q/XKBcMJG8PTx
bRCqufY8heOus0/rS/OB8pZM9ce0xe7VjESIislBgUaRApb7azJK5Okx2afdUc5BG08f2+GcWYLz
7x5m/MERAi20lkeSIo6Nae2W0PqqRnRXRYQqq5PTvslD/4gnbd+JSTIMrZK/vM2sNoQyUm9kXiXf
RkDo4vijyndf/+YW0kUYAqCKwVkZgjfPVhnYkA5xvD0VPovLjCFffgPhApuNQ6Oc5MiwAvPsWobO
d4bltwYH4ii4NuH6Q8Wa0XdmQYPobg2H0l9N1tFi7RxBi5K6YRVg1zCHRI/NAY3C6ws54LOnrhl0
y+HRbkRN8h3RtyZ39CvV7G5irm3LMzqAI5u+LpI5zJ4jPnwaq5E+qDSZgmUVfM9UwxYEeXavxGJG
vJlfWtLKAhtBpnRE8PNHuw51/D6dMnz4+6svRC8fW9Jp0ilfLS2aiS7xjD8q0yzE+DhYBR+TWE5f
+71rEX/OWxhETQuSrh0keFahR0abHMsrhcwzRRnMiZBjkpwbPYCrGfZHD+RLILTv5j8wYvWyvI/o
l46i1o9BFxjOgyJ3HzNHw0DQs/mZE1wThk2IlT+Jm7wP0xh2Qvm487+/NHkHc0Z0ASDvQl2EAnLq
476auE8VjL+mifUiG8yPFXqT1V6tTE5UL8HMkkpAnXZunL3FTc2iw5s+B7+J5BxsTL1QVySQmziI
tIJV6wTKROWNhL8xTcnZRMMywjMmJ6Q0C645/uxRTE2RI2QzORq0Pab6arh83A5BkZ6VFAgeih0O
5kQHlGiSBhd8W8RSadD6U4I7Fr3gRqyZVhBAYulQw/SqMpd58SMOjXZ9bXdXYpHVzE4qWV8/+0L4
1z1816s7IFcKJELX3Y3cIoEb7nzqSsXfe7C6J/LovV+sQ9lXzayT9C7XNcMeaSCijizLHCIlFXK3
0dyIzfnuE+eotEbsBpGwWhTeoPjyp/T+17aGJlISXhIXaKe5KDZIrPnPnfXM9YyhTnOJKoLIFo81
QF0qSnr8YG+qCgTQy4oSYJXff9MR6a7yawUPzid4B1NgUn6wnpHX9Nz1pKiGZz3jQ7u/FZM6EPqg
BrZLMyTSr2QKJfSLqvxX0lcSOd18OEfR9lyI5tITOy84hVh7OvAt0N5CUykORuYB5r+tSEZhSKR2
NXuf91lZSpdOOsvtNCYvHC6P6r/Z51WC0C5m6aff/GcCV4FC5C8B8eHEGMta8x6qDT3AgdfRap6h
UKTMTGedTwLFFsUNZgPlalZSJzGrYtUyudn8iLsrOYMtGStNXylCsukqkbkqneCfD6m+oD5u73PH
ki+mGOL6yxo9qz9m08alWobpcP1UuhKxvGhR3CUd+We2UK0c8Z+wjWD91AaZd6Iw0qMLR897Xtrm
ztJctLTwHBhdw8mex3n6zbAbFdobSzTtkwCmFnDbbDDp1/IU238m9gCHshlCNAypQk9lO3uDlZOe
BGMInGbYWjcjblKeZCB2U0C7IbWjHIJ/0jQAbRXoGA3kVJGH1dFdTZIWv2PKdQOmvj9li7wcszdy
LSL2HB0DyUgJ2Cz08hdT+31Am5bSQG+hdX41yoI7uGUp8G2rH89RZ4WV5hAv1LrjLktVSzX66cvI
Fd+UAdrD+N2WPTIEgEQ4lhFd2YXAGVqiZux7jHvy9mfzK8CA9eRn5vhBYrqAKc23rfuMohX9VE3e
YwuM1VEkELrxQS9aGYnI2cBhSz2YCNH4xaEBq9CfZFV9rSqVVzSXX8XSR/M+12uYzskZFJ+Z+HQ2
Vv4qnW1GMsTeRaRB7o1CENl2cx4LcaqeY4qP8ixDSMM2xU7SBK0RXVxdrJ+Kv4Gj+bI5xAuTUN7Z
P71BB6qG2wRdcNd5LnIgqBh5dRvPR38nEKaL6JInGAuS2sLcTw4A8+VjDyF23P0dstySIw9CrNsH
A/nlOwIePwXjIT7wv+H/p+cC6aCH3K1mu8SnRBK/cZoRXN3sYZrwHg1w/0UZvM1G7NJ+JrwdTHoZ
l23IUIvj02hMKqojp3GpK3mzkSzeK6dSWxfmtmyIYvB361ibOSgRS3hHI6nMzUkFGyCawx/9T/RJ
xa2evxhmPZnCSFkCnJpe/9U+B6ZJE5HF54GvQJn7lH4kQnlU1fKaynmAs5FTi52NyN3Na6qggkBC
k+zr9Tg1yNaHVtnZ/owEHvkpKziTpvGbv38E3vbswzZHIIHXy9Fd587hXSoGAk8JDpeVowXufEyV
0uhlEMfUu3a7aRTfSW9JZQW2tGcp/uJYBPdkYOE7StnuC2qzz9gwCWDYx/FLsZ2EKeJ1vbPKeYhl
1PG44yxsb16YszYw1JaCTZ4qDnavXbOKPfnjBj6isNE0388kWG6hknv2gm5lBoRHqsabmElTDc2U
oHgcsRgXpoT7aFyZ+YMoKJrUx/jB5zEcaK8Xycuaj5RYXQCALUVFlAdVxrRg0O320HmLhQzPAFXm
XffyDeO7yxc/3tSJmqbukQUKtGuUyDEUtiDGRGJbnUNGlUigvlmMH9a+lim8+w2AdfNlooMe8OPW
UVDEQVGN9+st4U7OmggDRJmOTmO/uG4JmvQ7LTHRX7f+0+vurut3Zv05E39YtQnv48oeSgE1v31/
IXjGWkvGzRR/1j2vL4gs85uDfe5qIb9Ieui1jzX0SkoXpfO5d1cPRQzzcqYUn5M06Ac46dxGgeBI
IwpUnNAyr16hIu33yjcupdv+nrsZUFD/Eq5UjO1c0y7nPKeKbAjLmlnz0t9RmlBcXb3bg4APF5zA
bI7N9+/URtv3dVtq2NwP1UY2Tx1kVIuS8pJ5fNP1DPWeuC3eMq9EE9QpW1uYHYwu9DPyQMENN7Jj
izUKPhWXwZYnEzkL2uwbpyYqw6+sX29P6JwOH+/EpwSEGvIN/gfko/su+ZkFXpEBTthS3eyAjwPe
/Q4inUJiHHVLU/Viiznep/IAhRGBRKjJfJI+dsmTwTctALI3ihAvgSjgpC1jkFGnumVD5kjjLkos
XCDvCsOOaqbQUtglZldaK7cKtJwJC0dLLbX8XWMPQC8G8BeW/hWfmU/bctAasp1dtjazf//6ch0r
CYVl44oLcDXTxBN3phZAzj9e09SavD025/2grST2RjzJm0Vo+FwhcZnBWQu4hDiuqVRlrxWBHCk0
KSygzNGoc/r9MGNsTbQbfnV8tEMUsCzbiWnjymii3GyFXaEZ4kaj6hdlC14aEfhITGSxlRq/AOWU
DWod0O4bPIJEnAuSfnrJCr0Z3niPJjkD6Wt2j3wHyQc1uMeuxp9ybvGyPD+1C58SuuC38fTnQnQk
iJDKlJFd0WxA+AXxb8XX0Vj1IR6qhFDcr4vizlt3rNH/mNRtyDH1gRYl1QRZY14bpBjO5eSuBaIy
hr0fyXgJO1rptsftX9VIEAW+UpRPXoPR/ye85g1rOCtzY67UEsvoNdZ/Nmxg/KO9uxfZ3QI9R0/G
mGegviFd5ij5a2artsCexp1/Rr9Ln+BQ5gZYEb/03sm5hNrQEg0/aozyN6n7CBI5m4rrUh3Ag84Z
DGpjFKacxz2qS01+YtpQCAJwdRT2mLGZVKWa2E6lkfzMXXm6mQ4RNIxEBQWBjfjFq8JfuKOnMm9p
QbE9lqHQzP48CdO0bDxmUe3s+inSP4WPQqDm73+P3qpW/VfnJ2XFd4GTVPNPjBxz1I2/wMVEDyVH
m5zYoNpPDS2Q4TM0cScEItnV0pyRGaUNEwHTnQCCCE6YnGDC1sZiajF3IEk00UN1yJ68I8YhxJm2
FPjIJktVMJqvNMIrnJkDhcyllAOzip2VGPzTXb6rpoBqZ0eVLOQ4MfmxIeHozpjDBGLz/DItLnvY
RhHOwfljPbllE54dTzaCH5p/6IG5kvGykpCj7a3Y8TSKGzeMdyNnFraOWatDH/cr8odCDxt8iBvo
iODipL0sDJ9QihrBa4uZZjg+6Y6dwPYygAxRQBLYEjnPiXTP3AsqAlPZf1kyN7384418mkC3fvcN
vcyDjAMHRCtejQ1MaEQIPstK8QYQC8Xiw61zf7SX4GzLm4sN2wre5N67AxpXuDCYrM+DawoX54kX
Nbj2VYsMxq8fuv6ariz1UbSSjkeSaYWBzwKUJtYuBFaQlVCBMQPlVY0TPzI6MV6qMJt6aHzRwO4o
bUJ+rItJhHNXjqDF7m9Pr2VYV0xDl63IVMTTJmXlGhxnlZIv5NjUctRDGifmLq6qD2wh3OyBzEMI
Ow44OFsCzuYSRlpLUrVMdj6g7VGxaW/2Rs/TZIJJTD0nLrKNfOW9kpGPIXb6CxAcxWEPuGJlcrPs
dLvvnEGxP0DlWN3HHGmaYQbHEzIW8jZwyhUdzcOvrmkcuxaysJBImxH7NVwp00c1D2ojusgK4sk3
5zqhMtmhjPZ6V1IQ9dLe26IoG1nuJ0TgFYesSPrAfuMd+NgFvhq2rV1hSBl8qhSgEL8qzJeTHOid
q5Y6CQMkCaX2F/7yViBZbR9viwfJQ5LWfmYhVo5QRo5AuYIhFUNHfTd12mT24BY9CJU8lhptlj0G
RBCg6o2xVxH812y3zfzoEQ6EiubaW64lERxk0O8P8wH0yOxEY1dQOLB7wnl8I7Y3S18lmRZknhWT
fdFXE0LGkgRFuAu63trk9nAmiWXl2AAy2DeXZ17PsdctNvmcZP75/2RYMdlADvm9A3NH79o0FcA1
iN8s3di9MHK/cnhcwxYKVl33TYOk/+BlyxOZPmHKOLTmzib+r8cdCpMXmVLlpE5XDALaVfEC+XfQ
DWPWWIDmu1j8kSMgcxC4H4k7h4d/kS66Znd4vdN83zg6TFfT5D53C3lSTRyE3XtJZ0s7MLUjllSK
o/XXCIypnv41K1pWLb0+zLB5+Nj7qLGOf7tVAmLSE0GzjaF1/anAg68DKl7HoOeFxVZHW1ZLC1ww
Vpgl3oxFYqkL3QM6TrLSoBKD89vlvXi+cexow4DkY4OKG0iTe2ZDuGCwa/KWYgnv1/REG0ITAD01
CzNexoeXUEsIupDUAlxC8+8eGzaMuRQmPN0DCVc4zlgPINatF7L5d2vjkMN9ORxwrNNYXOKi7GNS
okp1AI2+HLidHJqN45FV0joLpKQrf6/7EF7VJ1mPK44WREL+YR/h8F7XGacLr3OA75w3hyd2ZEe6
UI+Iy4vDJ8cGjzcweSA2I1Fp+VVZiEdRSrXqOBjod7//jkZieZ6hA4kX0mUTqM/rggaqjEzT1gbf
W5WAuG7PNHFt8wxputecj2GtVWDZ1OAaHtW3iKli5uh3zY0iUUL/eEYDaTwAee41aAW1kUIHNFmv
JlzmqkJRyUfo5nqEZ8dMWNG6dhD0uhzKpaPUU/nkv+m5EaAI55z4IS377RAvH+RtVDDB89ltsp1K
rjjHp1QhFgDk1ofFGcLhO0YKxY25slObqrFZU//Jx3dTOFC85gGwUgHZRA3N4SzNm8Zm8zZKt1C6
VlK9ljalp7L/5Ks0PfwUgRu7zk3YCvmoBpaTM3k5jOICgaGeBE0LtGLVaFovtY1LujNQRH2UW0Rn
BlVlRrNVJR2KCP+ZQxKfljpq2Z46iSK1j5PlpKQqwW2X7EWN2ciPhX5kSE2wcR9VzFknnFlxId/g
GZY307ihVxlwRg9ZwS0+9Q8SIaVdPMBpC7tGGxgEYDmuCbK7kHLfXNNGLa+uwIsZ2h+VGBFsgN+1
RRhmE4uqsUvxivETIeRegoZQP1Cqp+8c9zE1zTFtmT/c4GA7WCd4bAUXOelaqnzAenRLYT7uO8vk
7Q7pKU/cEMWKsVoLGKVUHMUdQnQfGP2EsBvn+uYiwlToD5an5u2oOxfuZkjRyOQ81s5/SCAsRWJk
EWpthl3ouqMLTS3Zq+2wna3PTAe9z34D2eowTIKuxNhCmzBDZn3enB6BVIR+DM1Nu6862ilmEn2t
ncgPxNSrdHcfEbGD1/c25CdSpCc1uSqu4EREZizC+by5QiHML6gl5jNGso5m9JdhqTLV90HLgZ/N
O33vb7dCbfivny/UCo9cC9XVYl9AGfdHeaWz39Y05bXuOwzFgUiI2cFuTRVGtYKoE050R+SZo7Yj
2jl/tYslqHZMTanNyo0KB86yfNyYVkDD4yW17RjNNqxcQElZMM6Z8xIMVB7cbQlbxUJpIlz/cU8O
k6Da1qcIHPJ2y6+k2cQLQ9YMFxrMyHQGLUajXyGNpEmZHYnbLdyWgQOqk7CyPSksX/WzFgMXiGYx
mOSytA+vlOlu1b+QdSB7sgaZRXWJzvbn5G0s7dS9kUaqf0Fukt9YNZ0+eLhi43RZeJ2/8KAHLD/c
VGnXke6pGRDEVQY8LMKhK4TqpciKvNfnP/qzQvnm+06f+u6jh9MGaJQwizHntDLKYDo7Mo+rGUzu
Xm9dWlN/cpR8ArMwWuj8fFU8Tn8iUyXR1WznULj2eN0TOPbQS5EEmky7pgZVURtENPerSUeQrzZj
wVe3l1OZFimFXk9LeRXNBNbvfc9YFz/afdG9dyS9W99N1wY44j0QArih8S7ndlI1eRq6fIrum3H1
Pedh5olqoPpSRFlJSht6uER/BGcZqgCz3ip74f6HgWeDjPB3TYU55ltC0cdt9L0AcM4cia+nn/H4
VTogWiwH6V9EnDKwi0JZFqaZO6MNXr4dY8G1TeVFgXbYD8kwYD6+aI9j25b8HksBj51WoAuaDXRO
jpovJbDGX2fpupIKaTZd+6kf678o1wJfiy7bzuyKxe+aZlF8zKS2o0whJV39IlQ3SQVFUYB8YUJN
HkrzVWxDzAXwmavCOA4IxiW/S1ybOyPB3ChiGtilldTs2+D/LQPrh4OTjMovyvdMSZ0Er8pyIt/x
YF317jEjTyGPMz0ZmeH5GekDLUpvmDeb7CNWobDLSDtAHKxq9BEcJoZLmZP8wVcXyOjixvj6gQqH
jucRPF6ft/YY5GVA7NhaBFehiS/t0u2snluIa1G3XjYAdskC9p3UYldiYPsl6n1L/siqzi7D4z9Y
b/OjinPegHeW8YpPEyFUj1WK0vtE4zJRRI/ZEDpSiQ9OYzRFHmPn9kV70miPKwKwKFc7tCZrVJI7
oyZakDAfC+StDhTxkNNgxUY+CozZ1OqTVvtgB+eeQI9yZBVVCQYMkiWOnJ2Wp07eUWyxnRJsaK1k
qqNG5aKFiIA4/iaS4xz6kx90b6L9xKLpjXZZJe6S5FqHBQao7i27Y2UlUujov6E9+Dc2/zZ+CZYI
p54mkbR26jbPQKRSnJyzIGUTVGZRkoHNCBdW0J6dNC/zObGW0wov+WN0RxAgSeMBLKJTOO2TXET4
vIToK4l0xPXm2V/anTSnO7Jl+KzZ5Q8X0zIfvUE/x9TMx83z7hsv1fSsE66WGvqi1XsCmSiaC+yO
mpi2pOxviAaP1XZqEIZ63o2+Ma1KIZiyi5lloZTmAA59HHu5LJ5eC07E18S0YiJdHAuBYdYK0aHK
Aftbnhf5WWAQLVhUjwB0+lIngdX2DerULCbbwm0UzdtG7g0aJMXVq4CgGM0o4Z5NFpAV05QhtfYW
O1lEx7dBX4SiEkcmDmqFTYpBGMkPKoPR7TRWF+yB5coPQcBr8WI16fGNZKtY/OGigy7Z9zADBRC+
kqwwZUR3JIx8aKMx7R+3HXmFrdOQkr/aRLvIIJW0FEvmNj09CospKJzUvAdIWJ7ykMNfiuIcgsQk
J//veSGT2AOMHe2lCjmR0C6tnwxEddJ25/5SkZE+jl8/JuQuHALuthi5sxTBEXu9qEYMIUzKLPlQ
ngC/6VPBIXZfk/xBO0oJNN4aNU6O08jvMgmUAcyyGGUR70xRIBdlWPUnJKhNLndBogn520Ynkf4M
SQ3fvkdtMH16NdUFcB9DWhkViJyLfZCcYFJ8rM5Gal0eWfaL8x5yqEpt20NglsUzjCC0R02mwqdf
YgM3xYj5L2Dkf74d3BiCXyDlCvd24bPTn4chmcZYogLJfe4ySegFgjrQmpmi8Xra2i5ze/2caEG9
nlPvnyM4H3qmjZvkmrOFChsAsbk7wx9jF9Z13ih2y/KQUOwFARnomHh8sf+giN3AVYESe7YF8tCH
jk3mYklc/D3c9QMecoLz1GiOh7Lj2IE+20Y5daOVxtcUgpo/ke0fO5xJhOwAZdXTmxgkRNTvGwh3
ROBo2JpcbhoNjpCW7xcwHW30oOITjS0+ps0ygFDsjnsYeeYdlwAeDAVwgc5enapnFsMAtoic3TZX
ktXUGJCwCa1ZpZ205OWLoC9dnqImZP5OYQdIkyaSJ9jqQTX8ryEbja/8YGx7Tjl71N6cDiaP2QAX
hu1xRIrxXWBsF133PYNgEmolKGBi/ydyNrJNlWZ8pCaEj5PGD9aWGgII8HuP/zWuK+oRAdmqSDxH
crN/nBw5sc0N+DxZFBSPboiSV7l4HKyxmk16TbwJmu/UgQ+lvNNDQjdJcRMGnt3q3xNKyzgdfAk0
jQNpwF90cKdm89NlhBdxAhvvXppIr8lT+OgMXvo1pvMykvTjkXhTVJwOHJrAemzuKZDf8FCqxFjF
iBncQogsmuegQigVXmbGH6o5IfNq0gRKKVwlzkwsXDvD6Vo5iJ3KfZ7w2i7e/vqd1Z4WXJmvJSa7
UmkZIBZLLW3l++06H94ddu2bVuBN23PweGkeJ5GYj4GyG8P5zN3AGKzJcUOwLl80DuuLL3irHO61
cV9O3vTsqp6vy9ZoGJ9xPKenlfNajPDt6EIPVZwgN3FJD7+AwzR5MgMYODsmjoQUsKKGivQ1mu/j
+mMmN2AjtOKRMm8IWSrM090eB4eRLKU+eNEsEug9idAoHDjnTL5OvVmPo5qOsfiBUaJCxMDMmWaJ
NR72Sr4jPP65UoL62C1diiWwIeZSv2nAnGp7r3NE7ifCV4ELrlpZP3woSYm3Bv6U6xQIYMN0oqGK
sg5dlo/sYg3LUR7ljyqdFh6JjhXkUa3xsVMZI7u7nlzHVHKciDu/Nmx74bDdnU8HwQHbiXHLeuM6
JCPYt9GXBa2zbiEZGqTbbAc53f8YWKUVnzlgLEQHl9SoMeTGC9lBtnf/wL2GVj7doOCI7aHk7oqs
Mhc2rULWY9S9azSdiuIdNaQsWF0wlIpApZYMK+j9HpAifxL6bdS+iz+Gi0an26tsS5B/69I/2/2L
iKOaBYUr1vXHaV/Qryjuz1n+rN99LRVc5QD4HtksKKSKdOh44Wiq0h5zSfpCVrvpLfTqH6+Qb8HW
KWd2xSxzW1z2cG6k0n3f6ikcpD1MKG0ENqb1f8o/thaV+gA8xu3fDZUsqZCE58fDFCzEmLyTfB5j
Cb+qcELOPKQRgAB1cGq6QMkAy27OzGBcI3MARAvXJIK2rqHyRXBSlJ91reaV2IhQAnuoOj00bcVo
MF+XvrwnzNtQk6yVzQM4Jw1y7aelcIgaBg2mDeCcSV3QA4UE21taoXTQzPAyoLM2j18NaJNM1fcZ
B32K9nIMkTNw39EYejByoYvSnsPgzj+eZhF9QLqO1Z7wNKBYkfSl+xDFv0Ry34g0MpTasyK8iIhv
1emHd8ai4zQ/4qBCjzQoWMicVEl6ZAF3jzwWhkysDupkASAmgaELiP6YCVnflLewRqKelhwj5Q9N
jmv09TrvMh1ABY04zSTsf8T6isFkc+z2Yuae4AAz8JR7tTQ1AUd38g4DXJE0F/j++XS6DZVpMhKM
gxWxUDq4QHkgQmxGC0tiYosP1363ijKVf6nyc2c+y3/hBUGHMb+2TRVtbyekxbG9g+wCrw2GlWcs
RWgy9SLLriY4WrMZQPN4eQGHwC56yKJD/gEzy1A0xECuMliCWz4I6oIbcvwmfGnqan22h4HwR9vx
bx+y+Xc5Jd8SJEImeCU5rr4M5FMcRkK/LfY0c+0MDFrE7bLjtdjcN/thDs6tvoxpoOtWNLBFQvwP
UJ+JYsNcX77oOjsTZtbYGiP7gw7keRzSwenTPU2vUKR9V6mO+3G5BdsKX8UW/1IfvkjU2D8tQZE6
pjRoAGHzNCLBA36YNlGbyF6UjXUMeKQrBldRowbCv+QO22aHoQ5Xt5eGOrri2enIQdshWo7mtOI2
UE3Zdsq+n2Ik7d8ziNVDBuIHYjdsJJgdA57fXUukZ2NMvHriZ2ifA6I9JA4jc0HBcCa4XGABNQPh
XssZDxrWM+pRQ+eEvhmU87hI502NQvVUCiPpMsvZPYz/J81GaH6HMd9umxXYjHjB28qE4Ts2gU4g
KMXgcNYvFRpkSRyJNmXkPuc6B/MRdB1ZupEHuHhJyEKhVuP49v2AF7ed+kOiTrn7dFuqO6F5RPda
lzeGqEuuFTfqjJUMfyn5SGhYKSpjLUxmbjGdUcJU5fQ7aWhLEDZXRUz/vQT1m5e9h+avXRjOb39p
3stFm5NAzWkuVzSepjvuwvSd3VeFAII1RJ6xN5iic4ZJ63nR63UnVDh0E/EJwWLvuT62ncB0H6Zi
PCiSGBO8TiiDZTBQRNT44Gme6Lju4fF/M4VQN0Cero9Gd6XczdmGNV5kjRIGNnVNQplfDDx02p4L
6g+jLv9MXaBRvD7UmfYirrjRqKDPy64bpfdpMmCaX0lQF31Y5tS71D5dRoU2Z+dMV3gvRyBv540A
+0G8RcF35U6Q/jvVfzhZKjf9/PcGMmrM4bgRz0Jzy/miMZVk8PbROnSeUcPePBvarl5L8LEXE+8k
K6L757nfeTJP0D03lAFPkQaI1uwnu8QkYT893Mi2lVKXemXZ0L4xfHZlUbpffO10tRBGoBFL1o/H
+XDwZW8XFyocgminiPxJf9umY7JTX8cyYygMgWH3VNG6xFZfqGmtmCyIK2tHYrakd4dq4SJ19G4f
oSxjaXSZnX+2giQFn5jM0vdOOP2DLN9Cn3oPruqICe0YBygPbsqv9NwYvZYYo2Tlrs1gEq7XFbfY
Qebwn/+nhzIdqst8+8YrlcTTDafHwNXFg6EjNxg0YasjrRrUMsxGV6HyQKkTnwwAjjN0A0HUHe/P
LG9D6gytgkzyfpKtAzGmKuLqDeDOrtiTA5X+DL4Eua1bOCqtpTDRAqD3VwJ3FGBuEWM74Ekkileg
xBDQWKcKTeIDdowiwBQvNziadtCdP89oGSKKuCIGlKHqlOflukcUtxMbm9RBw98sXSantSXTJKSF
Ab3XGpW1m0AAzamHQS8On5YSPnap2KPDCMhbiCDu50tHYkmDzD85kRmUoAGFcsuOShd2xnmAYpr4
A1/9JPPSkJICC46OkCqCdE69HoIq/47IJT6BnLI0x3wISE/Skjk9ndc11fMYM2I/hY2UZXiWXKgW
uCknyeQ5tE7EICVC9ufbn4IeRHzsI/iasSj0kr8KaBfLH2rAywbvCHSoLbHOut8+3rnXGRYr9zrQ
IplD1X0Jwiivuwr4Dlq0CIusXq8YkHikxqBsBUaGKy34f8RJEuezodraJVAgPDDwod0PGiWKcAGp
3lMAds91vJppustmUdmyJ2ffjQYe4prqdvmNkW+Crc/9SoB2npO8vaihghWH0yURBE/7sHZNxy6B
YV94tS2M7lV5VgWRZujP55+aJ+aGlqJTdK3UC3GbaHXxbYBPlJP3NF3Ogq8DzT1pQVhqZCU2zo6I
LyqgcbTMCuOVrS5OpV9sECInPmRlSSPjTPe+G7wrejpYAbkvU3EKobelgj3A8BoG9xa8EECTq3NP
Rb0TvpC17znm4iZPEUPcLT+++DOZbzNFRAsRQSXOp1ipC0km7HaVtUxmE6eeuFgJ96S2h/Efl1Pm
ZRr46GPda2lxC5LhpFoqD9WTjpvrbTo8ywpgX2nuIUFZnPnDt+upkmFW1MRIM9pNOKcUpUcN1Ieu
5pPGY7y4LdmsmLNSTIFh6LQUq6Sx6Zw2hVWRpdxzEpExoVdhxaWVJ9ixM92pI/acjxNBFGTVQjmr
kAOZRJDVwPzkNrPElYXXUezqF9Qt3K93CvcvSBcSngzowdlxI2C9kNkQp0tpm7eBtEA+AMu37QTO
XVdy9SzhHjO9sYDoBUvtWAR9K5+J9F8iwu+kX6WX9WedLLY4Wt/UpD5h4WFKmaQH5GPywdFbYXPM
/FVE2asYLdha9PwRqcj+NvbnW1vLxFOwCBEXHx44DCLU+FqfKlAnQqcYZC8Jzmo4MF+tORTq+2tl
ElmQD8VIu6w3KrVdqDEIyKC8+m67OE4xft+1J2Swp38m9HFLo/hilOlPRz8cS6wTVbOn8cGItDAD
5qM098hhUyQCzOnEtUi3Q5aU7pVhI8HRsENn5DymfjGQRlRKVjLnAh6fvDNVzPQt7m3c0KI6q89R
zycDmOLxOZtqY8e/+7EEjDGXyPyIm1sMpyoJNb5aMvDaVcFHSCqDiJ1RBkmZ1rAChybWSkJbhQCr
MpfoJkyQ1Dsg/YXT3UfD0DvHbXxXJy3f1PqGtniv4ByGzjizeMLoMKig6Hung40SYooZSsqg0+D2
RaVX1JKjL2664pxdEzMkQ0QNqpsm05oPKG2Tqaggt9yeM2RaxVpfGO5xQbJygc3JehLjoc7ur+t6
LPKHbXWiahNZImejWt+NIiRSyNcy/oRLs3nEHEzc+BTGLp1yh6yPGtVP1n7dIFsJfBKTxmRhEUOP
Z0yPyz0h8YVatjOkC4VVxl+a7Vh0uj/He2nmnrI34rEI2W89ozXBQy6FiYs2ysDvDBeJxXaMcm9N
av1c2OWcJmpDqwH9olYa0YD0ImQ4lW/3a0MTeDfvt7G6gpS68KsbXHszCPKz0P5XW3LqnKS1gI9k
Nod2TIX2OkTbpuUrR8y78zuKi/98i5ANEgi+4izjEaCaCpJQfJtaw07Lka8YQgM1fZCNKv2z1KkB
iAWAv0MQE/qQ+CF9jzfGFXlGhPMQS8OP8n+j8JQhR8PzJb3nJR5G065hO/tny7aeOUmzyevjr3ws
3zn6SI/DXV/ftmUMd8w9yXBeNwnID0PaFRdFgv9GG6LIWodtCFyueBgxYqaY/1E/zuxMHg+FlkgX
kYDKxTraqik1WnWAvsr1sDiF5+T23DHr0fo2cp1UtDtJ/ClI+no+LwFbrpPXOWSxleQRN1YkH/L+
Tk2xHJbcV3qfbTm542o2LNphslkrQtlPLMxcQxUPUd8JW2EhP5Wsv/3r8wWWEY1iCE7V3AohsueT
22mSq0qdGHMlS+IY7zNuPqcscNjRQSlDyvhP54TPYz9BiqZWf8tiNeb87Moh1WgpDnJGH/ja0VWw
Ktx6Ui/+tZwUTbPBguKaLxj8cMqMMe5THLHUG+i/Vq9Fwmd0IAd9SL25hikOvf2ZBPlugWHZLzqb
IyZRjqrcoUEveIopaZRT01TKIdCWJSrWp1E84d5VbhSLHJnt98nIPjncaj9W4AZS7sTjZjTfabf6
Aa12yvXIOoY7fOmOefrYkS6gw2BdfFm0avI8XruDN5g5a+NG6875fXO8dkdKmbgGKtPgiMTheKGW
zTsfpe9LtzO0itpIFIt/DvVcQI2yaMKGDmF/HD20cFjJUqchV1yAQe3jkOWJmjNh08s9aLM9fjbM
pFqoI/6Izf7sEIXTjmqvSYiQEicaZVAFTuxrs1O8DswG3ojfHB3ZKp+dQuRaCiYaRA4gBH22Ioy2
Tdx116/lLfpygFQSPRFRWDv9OpQGv2lwb+fPs5azED4z2SnKdwhaxrNxtCJSeKi7GiPmSvo4sBPr
GsdjJkJu/WOrkgSmfrRhVp6YskR/h7UZ+0Pu7l052k3Qlb5OifeBuBBlgbACnFU8FKeMCHr+NS/f
E4jYZCrzsn5LEN+fm4XBRZ9S0Suec2dAJWQmF+/JYCD0mOPA3qj2qfnVIamNV7h2MsrtqZnDOaIN
p5865dKLBWw/PzH0h8TB5+alodCJ4dwCmbXl/gvNMihPfocQanf1uv68oDU0l71xAP08kdYA0Vww
zK5g8betq8PYYoWiaWQgTjqCBjHqe1z7kV9fdUMOxIwi5f61dw8Hgji0xeALLo9cWDWiDSVfiwFN
eKaBrMRGZLG9zSxDMOYeO9nS/YkLLvpE95g6qqIa9EeP2Sugvsgf/Wbn8LhCfTEOyrd6KLAxruiB
B4/FZvvOisX2gdjqfjBdfBVeevbjctvk70xtepe5NOitV6zWAmbQfRRsrLqWO2Rw5ozw6KKH3ALE
s/eAn8wZhRkgvhafBxhIG9OclyrfGGeCb629hR4WBQ+9Kgkswr6ZaZq4qMxcCUuQtKLRJbEUv0nX
F8xoJt996vFMfjen7wNK+/A2YJW56KxLeWY9sUVCA5fXlxv9O0takp+aVmVteKO53Eeli1YmtcNI
HaW7YZ25jEPDpQXlp2BjGjoSNMvMb8QR6xqS861AGfK4KGvAtBrIMCsNuWn68pkWAsrJH3LCyPO+
tK8Y3GUhPI1Rq3EF8H/28+V7cxvoaj8DFUIQjfmLw7t78uDQu58+xVaJhBlN2ebm9U6nTC9CeVXM
mzerjYa57RWRDHqsTiGMxwellYLjzIHTNA8S60/oQOVAFs/depUujlAxhkKR/NSulKGt1y+ufIb+
i/qujzZMTUK3Islik0uPl34Hw8G1BX6qJRQdo2uNLKLZhSUAEds2590B2SmL6HA/H74FVW64RJtW
6khuPfV2J38gfibyzNhEaZny9sahmIhCT1HtHoNZgucmG9hRUIXPtEq1efyis5SHd5P4F2bHbIR1
0iVjhbpubmb08AJsck56Cxh5eFTcOEX3NSpVWbgUS75bdNHpzsQbp+XKpWHfc0qej3PAC/5QE9AF
btL/XM03sYaKAG2N46aDE1fc7DZJCDikRCCUOINqw2RQW4IgP6eYq5kpW/TuCwyy82rPhlceADsq
B8QEskWjOSGXFVZdq70vQN5PDm4Wv9leW7eY3pUWfhhE+7KJGDV10kQjMk+rEkzophyRNWwN4bUv
vY9T0Zf4sDeertJAQU26pHZ+j26G20n36BMv953+wUkijNpegPWOC10N1CSFj48MWERL+7a5Bs5g
sDm9ANXfqkOINUtiR+REnoAWOUF1tIPFWNvvD0UsOC2OyY/gZ2FrEymOTSPHqUMwJNCsV61AAUTh
uWmbUn27YUpwJiC3e+OLotVtZPwnud0bKP4PJIn3cO+yw2QXvkmoU5LP7YlCvQ42CT1SG6HToKHt
SNYcqDuNgfFQxmwWckI22lYd7gnXbAx1BfiarwjYv4dycaiEJ5uOKyd6ae/uHQUDldW6OYoO4pH5
7RfIGjVAxKIagU+F0gVH6pX3jARS1YPlxPDHRdPZIVBn2dH7f/xORIw9CQUnVGdwNm6gUMB/dBEM
VKgErbMMnSHjyspHVkazp9xRVG58MHdfKlOODPQr7NguvqGB7YkUhrG7v15SvX7ugI+OwBriWWnl
k/ZPEHskorx4zWV3nUmYLlNnfkmKqf5oeT7bJj6pMenFMrdAxTqHzGwI9KEdD3VWhwQzJUL5fFio
RJg1jpsytGab2e8eDUjqIo/abFOgoGfJIFe+4kQMIDEfaz/T2rmDS+hzlXEhXDmuCVoLnVf2Jbqc
Ey9LfDHJDBUVuHSQDAjt/23pj7heS1F7w8iHHJvtqFW4K3GfEhCtHO1dkEt+zEkXGfcKx3PoNu2C
2ogQa9geV6MGt1tt1BDj1ztKpSuzI/HFqT6XUVJrtKvZCTc1VjBQ6BTwLh5mwid4Tj+zcPFx82yc
wrHulzUAGLNtJyV/7cI8oqYHNeFuOzKVEUI722sXeM6o9TH2jBDfuOTFUb/iHZ90XsmnzkhkxI4J
j5kQqwrYNAkze4UB7CLODBqmTCkaVEFxdRiOtaS0NEzNErUKZzPmhHaUiayH45ihXdpRNiAtGffW
1cX+nHTPEhx6ISLkHiM6VOGv0ZDcfT/RVlfkxsozzqbGBYWSx1VW4cxhCKPiP2DE2FsWoxSoRX6h
WbnhezUdltmaovxOay/c8criuN9kBDhScJZOVBwJxacipX82QLgxImZYHFaT/cjQLx+Dv6IroNEy
VWfHG9/hRjWwWi8+sGV1qZYTfHqnoCDIDugsyQnZ7X6TtOIFkK5d0FHn5lPkq4JmVYRGSZghgr+W
Yb28+cV78SGeFLXQwG04if2L0ing0b4Z26uIxrSLrAOnc9DHfFbucrokR7iM8k0fddOQFcJEXSU2
TYu7izzmYzRT6SoAvsIXlNEaBwWV4PfAgORCp/8rJIHisgSB2tCMxaKdwkW/A9l77E5ZJmPghsVu
UXHEXEb9FK6uX+pOuMLZ96zHuXavpY3hUEZUdM9QMHXPuOgxRQQmCEXuPEQQyott6ZvBGZR/G17v
uu18XuesrufKKrjExN+J6uQwbjSH8u/xR27a6Rbkc3TW8AomVn0JMk1eRhljZwh4Tf8p8DMrbk27
gyawVrqZ9upGlZtNcweJsHuwg2QGF/5poWDJX7LkaWeBwJ7P79z+p/5rXQvmtijLeAC31e3cMHei
8DIQIG/s35045UBwFGmZhCfXma96VLxheoZBWQCMvjUZfdTFaIbI5YE4D44VNM/tw4DePubd1r9B
p4pdMmmcxMlk9cWMlggLJfS7QuhffH3Cb2SKfatB+ZPa8DeXRqqAy3S0t6F8nU0tuNplRl7+nI0+
092st+GPvvFGYY8ZEZPUDvHJObhAjh2p99ECQqeDaVDyEe2mGURXFo0ea9iwNcrc4MYHYecHEjvT
ZqCB/TbDDhfxneldSfW8KRzrRCgEKk8SOSWFKA0sbqPzqCkyEBBGzLkG1X0hrKfxLjs7Nui5n3q/
VIqfoyOP9LPFwWjnRX8/YOprstIXAcELIrSBSDAypNoH2KzKcA2eha8SwwW0RRE7+KJ8Vq8ngDo1
EqFZSyp6eUwotzndTjG+VoNbwz1RwqvJ16fHbxEfcNV154UcaGnyv6NwVrqIA8j8hessX8DFEfz1
iZDltYCNNlpWKL6YUCjot4G884W0wqjpbNgPpPRdcllxP0w1IUuGy/LH8Sd54cXBh43bhusRfV50
n/p3yaXN/piI0Z3uK2tGPNfLhN+Eh6Llsk7Z4In42ggFtbAouwailcgGouyCdvvrc72Wiiivu4C0
iiYSIyW5UBr7HPRErh8QZRoeyErMQ68EHu11dnEW8wUtAt3DT4Zp6xL/HcBdb1GNroCmnxM3NygX
zpHupV706x3CO1lHnQ1WaSM0mRO7fxUN6dMEQef6UDfWfPiMdBZdgycFwp1Y8SIlnfRwZSfzNSHk
MueW1AKN5kc+1i3sxXvTU/TheRztb1K3zW2Xu6sCO/PohMnQU8cKy5iy/YzOx+LRl/SsoMgM1xTd
yIyZYc489rrZR7fDoMpV0l4z0+W6viUI/kUjtd3nMSdk+ho11WjW7beWdgOh1aYnDZThvsx95Qtb
OCMaS2HmqMoUTvGHBISsofjP9Il4eCTo8HUV8uezdIzg5Qno/8TUfSQcbUZEJC9QObA6jClhKYF7
d1WicCF9SqZecdpYlQHcxmhTzitQSFTMjNmw3fvOzQWkSeJyoRZt7LLk25wSYdaf2FhUNFw0yej/
siyKNGrORCFrQX79czgGie+YHn+LUHA1T0oj5zHapu/TOCQr+3RC2MwCdfoy4UqcjOq2qCns4h7s
j8uutsBBr7TeLguC+Rf+azajIrJ7AKd6jDxwmgFKwIL2g2vGLH9psubRZ7v9WyAbk0+08IGCWA0N
IjUTGhv5Tf8BEwoXbOw36F+HJZMxRW7Wpk+igMCedD5m2iStIiLkEo7nXeZP+olPyrgJtmriTccU
PCQdgdqFRpI5iCs+Aw8xUmFhjoFzLnXzd3tW0G8FslrQHE14M5UjW3tV/PHBdUFkGC0HxljTedgU
Yrlx1TlEXlobZj8js+vZeHK065pv4gRWCbDgSxr+qu8+2LbykbkQLrrij+QBc3+jDggrXgwt5w96
nZUP2rV1LVzBYR1Pjv6Wo641oOuskscNhtATclCQZCm6V0XeLpQ6MocyfST/uMDeEw/HRnYQDlyc
/WPOMJNBQ29SIUEIct7Pl7iYnMI2qHHOpBqIUiGSU7SF2ymEaprp/RhiisiD/Sy3u/ExzBEYZdmS
0GPtIiczn5Wl+iF0KIBWYnVdRwrudntklybu8t92zwMLHfBZ9XIxnt1PP85ghkMifv6ODwIo3llQ
I/X6WlFpaOGA1oZ15npp5j9PRFK4KDAtPnozpFMC26UJdOQm6j62J071gsMO6b3m1GdU8LOMV1n+
HByz9Tm3Fcplue0KPEM4NkKXsGE7jyMuHQPGraE3UT0tssIs1T40Ws4xkjoDCUEQAJA1+Rz59Gsl
m+CR9qvD2151BFDs1gNXZxb3QGaQYQmWobrOf5+zl6fyPabe9jw4GH49rxXkOvPoGoLWzdVMS31e
Eu6Rjp0IYMY6Evuxm4dRHq/DwSqkJ4k+9iy2AwpksEHtvks1lk20TPOM/sLlX9ezBeWkQYe3nNSG
5dElJxwPcK2S7R/qBfVIcJK+3kXaQDdA9thdO0Nj6mifLJq6QLTGsyUFmyvaS1HqC4eal/9KoTYY
FmLeJx073Z2YAFqPPXc7Xc7ZWUH+sulXKpnoF8gzzGJZHlFQxbV4XAKHxT4AuZYGP+r2DcbYUDO+
vxV2C+Bo9qYAvoc0vlwQrPPIGfsTF2Rtu2PbrZ9rEU9A8Fdv8v35CDAHb+6L4CKZCRII8xWI853u
UxtM7hmVzq0e91FqPDUr2wLW0qcwNUeTn491ggoyNINA4LmTY3UmOiqkr0+rWODb57PLSZfh3+JH
CjPMU4+pLECRz1dV3iCg2BMyaBEEa+aN469ydBiG0E3t2nF0MvlMYFvrA9rMCU7AORtp6OZz5iZ+
mK/TP7aVxxfDFuk5O1A+VO7cfZIC5vAtqiq5RWu48P5u0gGEF1OVibDQwN+/y9PIzB5QWgPkaueJ
FgafI/ycNIzAd1bQ7/TOzSuAlUlm7VSB7QGdSgduUqVomhg+riBsrWsP7zvje0Q5sxxxi1SSpsVo
FBaZ50DnVkVa3TMx0F+BcW+r5rXPI0J7a3i/zbm7ZQKb1j0sMygFCSmcTjBFcZYi6J3qWygZ6nSf
E5SZrrBtoRQOFoGcifJX+GrktZ19zB28+ASCOM1LsrxK3GZtR8r4k5X97yADex4dDtMbjRVljsAT
YnYSqY5CBYsVYedqcJdU7B856AdxL7BXDW5k35JSCkd81n1s0GmpVMm33QkIzzXXHWNSu+3WwrsJ
HYPTcG5SGpwDCk+RFaW01tnb9BSD4tbqi20SzIbSe/n3GzrSjifapKRcqJ2D3nW3QbcbIOuYodVR
q7ljtPdMFjA10ud2QV9ph1v/EctzoZgthTW6TU/igm4OavJzawK3kwAIP6gIpKrQMBp1ZmTfQdwI
wtwn2BBwcfewjxPyX96OqwPqfYXO8kUs1UFegYJ664uAVlnmeG0ftlAFRcBxyUHbAlpz4tKSw7gM
o4vhNwdh78skqyVh++3JG5DRrDIAVUsbdpKuHu7Hud5L/L9Ucx4PNWLvcWqGjaMHCFGA9MnusFcz
ZJiX6BKRgVhlqXNyLZcnhJ1DfDLFPY7BPQXSKrmoO+C2xkU0h/V5/ZYek/kQCj9qEOosyhPqGUaU
XHWDm7FJPwjl+e1Fm03ppBgW/6xw9hsSjmf7yyf0EYAkaGi7PKIrp8fWN3LcMuHN30tGDiM5mic3
PBm854JQWCyAlL9UAS5jWZG+JHQEc6UDs+jGBwaYhm8PXqTdBSIvEnizURglWJTO/z0gruRQ0cPk
TcHgUKuAGmef6qRSYoupUJxeg28SJ0SHJ+1NwNd5Rr5cImianJi+TdETu3fW5zMs9eoGCQmImEUH
nOj+/qFlD8TfyWsY8dakz4C6meHp9X+VPQ2MKQHFh5c1obiyATP6LRTPiL6gnqmpK0LL2icWVdtn
FFSzDPQn4VrKNID3bkDLTTTkRcZuQxDERjQRgXNQw0xrjgbNs2//gZo3xIlABddyBPplGzzDCztD
jnesrLMSZ58SxJJyqSF1g5vjoqzrgyM6qjnMPMPDGPbuMiGxh+R364/m4/9cOzbRoiSNKAe0Et0N
tOjBt52p0v8FAKjXu+H9WtOq497ITfot2CevlEhOkCaT4ennVEhsr24yTQskwNQhxaUQd5q2gZ0d
GHpuF4UMk48nvfld4F4bKsbbVSzAhi9WPluPEBYG6VmZSentxba2HmER92mnrvhWNdnK4kPoWhcu
n/2sG/aW4WE8GG/vWsMECKBA4a+v0teT0XutU3shQKShNAvQ+TCdvDkl9dzYt8OKGluYcyz9Gvwj
yUPscZ0k8lxDmF/NtYvS3ae0kJZnpEF5O+c8FAilH8iwoTneA3dN0uRkYlhum8Mzg56esX+DxB7P
ahGniatNgBFoJNPnRrtO2xNGv5ZmrqNS1gskAdVBfw3WNywPqSteGOCa3jQnvYvqm3DzWg4KEMQk
RSGO6Q40t8iW7xwuSS/BRsLlQb6/SUV5cgd1ensWHupu9cIJ2rJMe9wJICQ1gOnJG14rZa1s0wRw
63HGdKvZPDB1yGrcp9W3Gf2VlVtAGn4/yxWCcNZnDEkgXWv0uyYxkuLfi3mLNkKL2sJzXEsXCnOu
Q36FZgQfgsduCfRGOAqo41gUSaLxG8zoXlhyX+Vfzmky35Uer7ICpFcXbXzBC65ThK/6E6WDKhO7
zgehX6k6alcI9moqBn3keJ/7vNoLgWlSXXwT4ts89gH010M6FcuQL23bG8s5Hj355zS3qToPwvmW
bVwcvTKGO/NgI56rn/edxjfPrstQ6nxv5cQ8/hw9EbWdwZttAmt2dPd7pfHYmp2WUrRop1r8g5tr
hl6MpQQ+iczzXaBG2uem48qWtIw4gWSeM0KWxEPlV9ykxDgkKX4ybbroR9M9nJw/OF/m5rT5mZVZ
0w/hFhuWQm4VyAjBOMO6Z0liA0EmARCIo9wBuBh0crVZjyXLW+L0MTBWt6TEo/Pa93cMx6pl+Nd1
zRIPzDzOJDlaHGHx1Lytr1wtsiE/Ln4HM62mDt/JQWGZlLaqN34Ud7GvrrdQV/up+qz7aICUPr7X
h6AughqDLITNyZAM7Y/Pen5UCCxlANPU9Osti9DhWT7WgOA/jgOGEwNi1x3y2jrIFHl766EWCb3T
VHTgYhyH+1xLhPuU99BPXvB9yrjYeeoCTtgUdiklZ/Qx5R1VAnMIdLZLiRk2gVgPbaAIFMvIpesM
OMtlug4i54xlP+DHI0+m6BGvTBxNmwfDzmAeH1/4hEnREdBeVFc2UTEVLhq3EjGLmMP0Gzc7eSac
JYEsI85c3Ld8keA/dBRTPIc5195E0lPTb50rCukiPP1CCTWxbiFKi3XWiIJSyRLGMV+Lz5jxqe3O
XuxKDtPKwAS8B2eMItbi9do1gCa8w3EYI8LcaTlFICto7zP/1pXgNnllfMiOEDwWAvnFpgT0wnoB
HOBYgcKUyZ7oHflvPY75X6Qph9lUozSR+lF88BwgQsXnKj/lrRViKvHVk9gneow4IuPTF0dcGgoN
hvsnsxy0k6WXv2GU8P7ev/ssxGHr2HK1ARTjwFsW8EZxKLD1W9RZPF2xMBrDav1UHdGWoEa6qT0A
ypZj9L/y+RpKEfh57x/ji/v7MY1CaxoMFM0aOh7dfE+/+bs5jY7kQGiuhled+vGRaZTysR4A2PQh
s+EaeLQv/3nC9JAI8rS8KfXkJc/Jc2nlDIFVu7mnQ5H1nkHxZuMMOQOkYt7Aaivr6jigRq5nmv25
/nOYKZs8RqjMNQFJt3FjU75E2JYEYIbElREHFS0xyYeaWRa8aepRFErLfM9aj3QIGp4mAlVEcnxl
//OuevOsarRJwgFdGrKWLPIFQPY91I1fqy2YkOezIccmBMUo0STtNkXjts2/BCXL+lwk1k3oKEYX
8g8gukZ++nOiFVmD0H+nQkn4pGCC1H1RDNIQ6a8jk9T41Y7Oq6K7g/OrRbPTuo2d1xynviiGlvAG
jYi8GsU9FUjoEJwLwQU93OfSS9ZMaIt8d38bqufQv1aHbNXReRM9NF4tS18lGKHVejgP2nqYqnzU
YTsEehxq5gPXFw5udfAG4cQXgh+yTcKzsg4i+8r29bwdqpbZQh6S7kUpUOubwGGjJDqjkHWr7CyS
Ol0HQ/pbUOkKRraSw7ZfKLzlLgF+77KTq/gO9BSOcaTvAS5i+Bj1QFj1p9rzGIetjsJDSCau325o
bBhrI0ezHgt5eCWfqH1ReiiBxW25II2WwjnLCVWeAXMA+PJ7OM3eUsaQ/ud7KwZlZTpjWE9qQUFG
RAp2k92264joaJhn62ohBzDLEVZ1r8b6ObYm50mERpczj01TjlE0S+1x37EqH0ew6wvLf9hG/PXH
OeDR0ZWT9cWdCS9HTHi70qtoJCT6o2ZSBcsn8apKQ+vdIoxjcw2liHnHE1OwwNdCVFugW9wiLgbZ
jdd9VpL9S2au9kevazbW8fDKHxlQrShW2dWp9E7Sla7ngeD2fvaiA+WcTpLeQlNhQkUkte3mQV/b
B4ibCkzIgLlBxUXuuI5PbesJTNPZdtvzJCaGSOuB30/AhNZr1sbVJyTVSVYamueQr80PlPNsK2ZM
OrdSLCGbp1P/h4FcOx8IFcKgArbKH9X0IyvzpBz83H+6E9lsnZvG9+bCgB0CaEe8S7juaTbIzaYT
RuK81Zr45Ay5fMDxzKC67ghO4Yc8eoZchUvH2NkWceKTtOsd+GZUusfvkGTpn2TlCKHCVm+lqM44
NpyNllJ71xsl+sNt79h/prDt0AYDeKHrLtGBDy7YU0BuFgry9hG7bHkfB+Kfaj6YZpWQ/WFXLbbO
SdDKGkDlC7/94x9UwpKh5Y1Rm2f+xNxb72Jz6gYul9gHMaX7vH4d3ZqBI9Y9DTKX9WmtYC6flZmB
Bcv2Ly5k7mDaCnoSh6StDNwyE0n7pz+9N/ZSbRS/zqrvfAo1dgWx31TKd4Mw21kAj8qArBy1sZK+
zR2C93tjfXle/6RJ9wag1PsbN5i1BGTNxq/LUg82somoPZvHjvh3TZMql/VKrqVZku1XOJdHLPCv
PLfPnecvThlHEUVXmYsrhLeCOiJYr6mtf2HFmSOdwLSBRx1JkgLWTUjpKBrcbKkPsV7+aCvtZ+fq
opfT4GzhewR1Mu2uGeQPCNGdco9oeAYvVP+2IVeLsPUVIGd4iJGXnivfZwYYzW7vJKLWE4gFX3jN
CkKbJD1QUsmIW7W2XzBPyNEGnjzwFi4Gs5fGIaysa9bpiW5wE6dnA8Bo5BNOykPkzldICYUK9vR5
37JEAlJuBmsYFXzT1OkLC2x+VhemULE7S4bnwbsMi0BugnuulbMZ0LkHJODcAj7GfPz/lq+mQWcI
1K8yosYPUC3msuSEIV2f6BbJfTz5dj5fG/ut2jUwwk+eF/zluiS/qytS4BACL5UWKwMkuWJv6kYc
pQPR4E8e4OGRbe96yL2K0pi/dMTOQbmWv5iwk5xfZsTmjAQ7eHNv/lBf5Axv7rxUmOWCy912EOOv
1pbiHWatmhEE3ZeBJBITUQLw4K/XbNuCgC8Zsf0zxmdodVuBpAsvN2ud6mhPoMkX9+HaI7yFHfjx
ddQ3LcaN2we85+MJjJZp9Dlj3JsWZf6mmYgUyJoxGY7Ws+SHzyeVqWFbg4TvyUGrboGKugQiayPG
j0k+SNn90tKxYw62+AOY3XChznd6ZYogHk7VcX+qZJDta4M1b1ed2NEkteUv5nus5N6sPLwMr47O
MgbjDPqriUmDMxaarnjjU7FCr6FhBLcQShy/gKYnLaTUTl3gnNAd4m5HSdonKBfUSbGrJhZPnnnr
wYc4POdzdwspC2JitvlIUcKeDaOTI6bSoIuM8+cVhe7EufZ6aI46780RPzyheuMEpDNNeN9RtUq0
meozDKff0DiDoE2Iu8WHbhP2MX7vpcAxbejmhv35gjHVTQDB4PBDaNTji8XzaJGDifM0nAQG39DI
Ah7jf4Kt22lXqFmGJIGmZHhvGPIJ5nPaa/v1lb9F+KFBQDXCY2LiUxgCc9Yx64z3WyJ/07s/XGDx
CibqUqiuhjpxWNNGeuvTZ1fdcEYd6O7Hgp/j3BMNCr7xlU2orgYEUIOGp/DiyKlAogeRQspZA60a
k+3XSuY32uXZGBJvs2jzuOujdQlgCxgPA+TOboFSvk/rFndO6cjLCzA0iLr9GUCONfIvD0mBM5Fs
s4lzabOIHsLgUITWWjFULLNig9c0CSPM9nDXX4Eim0fQHhZmtvt2cdhILUd4KiddOUu6fKG8LZnr
bdLF+4Lt2Tt9daBNjGX+U94r43gSB1kBkQWHBDGxQJbCtyDVKIBQiqlyaiKOf2p8NmtXJu1oWYCU
vK/dJ4/seiC8aOQxWHPaSpG8AtkB3GJmqonJLTwIabJ1R2fgSPADzkwAcAXxkdlSnwlokBe0b5TV
jHjGjzuW0YB3tCQQu9J2l39NYqcibxHnjQ6alrgpXL4kiUB+rX/jk6ollH1hft2FKdB/9FVAMIWu
jG1mUKvR4PSy7hsI8RrmijKXfLVTFm2fr3u+osH6G5EUG/sC0S5ryUrPXfN4BO0OxFfl3VKHCKoC
p13mlK7rrP6txYktSz1GEfwn5AFGyravCHJ6B585Y5BkhTrOlah2CxJBkRTmccPKW3xB4G1sqxRQ
e2QAAqAPZeOT/9/XB0hIDSxgKG7tLeRxWI6Ii3qJmJVuEWaXwyPfbctY1ufllXtNsXrv/OWH2FxP
0VFUstkHbPUDMdiRSQ16x9cFMweHzaq1xINcmKoI8lBB3IF3W3ft8qpzUbP2OB8VeH7AxLu4jjbT
BNJ4aC+Xz+FMoRNPebAGT2nygm889wgBwkRjSUCBAaHUpnaP2CY1HV4ZnaVm1V5DVqud1aNwdh0w
x/VpOyRXiZIdT5H7Rro5CCGEZEaswFN5n/PPHCYzcKmDfh9uoROq4MnWyB9xg40ZAkZAT9zlwQ8G
hLjQyVXoNopm0YCQq1cW3m699RilfKpQp9Xg3oPqVfKcs+gESs/CQbN8UYoZ3Ch095/035U7IOBo
pSfglJVlvQ9qJD+pnHCrMjXnOjYgffU+Ll7ZDxlPZ4Gv03p2XVW5liDXY76KBrgAzFwjPxzd2qeE
r+J76Hv9HhuF4ZLd3hQRDve39eiwbOg+7NYF3hAkNZZ7r3xvQHeheANFxZawgoHF7k+mcjTzNomn
BYfcVKYDMYu+ucHtEzJAhdgEQfCnBJ7VAuqJ5MPXopQUsH0mG4PX+Gam7tWPFqD9wViXZS84SCUX
83utZQrvvNgNtmdX5+SJK9hiAGP+kDAEhLcAlAT2jH8NWT+NNi5PLu5X+TUY5OMKnFUbTOr5DjSc
R3dPH/lWvQRB3tOr9advj18U9ezf1TMH1qgxpfEvyiQR58ZMokS59ST89PPbW0DmKkr5XLntVxHs
/FFAj68iSRTyKDUn7ll2LNfkuIDssaN0sGmy7kW3xjV/wpQYc55zDzNkHAuwLIaoL4ksiAiMa2j1
VZFYY61GfLMouxLr1lehqmSapJ8kA2zfazqvQPn8sTyC8Cz2eHYrbkRB5P/q2jcXSOZQBaTTqVAa
+ppx93r+aQeJ+n55uBGdqkjj8mHcJMnjm3/lq3RVHJIuG5vQp6pQcJIHDTntk7JRrPioBWEmL9Kz
pOgfMwShtAxc9WcuqVAXN/4X7/8jAda0J/BZY0muJ/zDVxrWi2ye/Pju94Q0pYq+s4ipGHOVmjL0
MF7knhf7fK8SVz5v11PTxxa+I6vksCjdlwkJTQFfh4XI/ckRJOuLVYfplNcbaWN27EIHYBPCfgT7
nq1byCghfwCw3tDWEqc1kwsj/Z7sFD5DNky2BDlSZnGYWx3hLpePRtIVhEiXAYkAqnkuCMcaer/L
L3ifKlXABP51vY3Lgc93oqxHukEaEsqOnKvdL71i3yRhTjbYtuLsLTfp4j//vGhndDvJR7T5RcCg
7BUQQvmQVBbsK4Tg+Nu4M3s1l+xDHimxvxJZLiP+r9TnxxEgsoYKdrKCL9RhlbeU9KHSvHs+Z8OH
331LiawxA4vGK3xuftD5wrGN/W55fso5fTlkef7cTG7LcoKPwhu/7BcQN+/j7WzRdusm56Q2m/QS
CJqw+7Zah1PKJhZupfGAkWscmuNRRAdvzZju0qeCtTu+abUndAV+tzECih9JMP95T6xWsgq1Z8Dx
D1et3LlN4j+cwZl7u2loBsllJCXFhoKpKrR0OT08vEfFxTKxfXPjmH/Hq9TwzLgjgGgR0Pd7MgQC
OgvUPS1naWHQF8RN4XlBVMWD0TVITxwkR7omSAE6MVXflh+M+0pwdJ0U0tBpVDYdxEcU9brv875a
tPDST4B3127yAaEq6k6byeaeYFkspgXAy/lzS8TnFD9e2j9TFVEzzYIn5cmTCZ33J8CUPoReNWii
0pasY/PUBDhj2kmMotEtSmLGr1MqXNvPyN6sFbLb6DJY1wmJ5PQINXgHzz4Z5PnqeUSnQIev7Bhp
O1GTymEaub7nrmQ1EaBg+YtnH3cdiNzVWH7pzwKu1oBeu44WjXDsZ/+Mu2bUiWG8GG1xlEeqTI3F
+8RwarukScd7gZRCcfwdh3mD+QGbO+oR6aWQXxsQnv+TkrZcP0E6hZtt/o0q3Ms4SQV7zANHuqU2
Oz3qvO7BqrohojF8okAuSxIiGs7FjTtQSdgMwX74qTZs51EIhmpbAZ3gM1LTdenDZGIl+b0+ldoi
0QLSMWWWQGaueu6vG52co6oApSMQeV2sRsUaoKw7QP6y9uEjgHl5dNzl1DducB93yCRFptu7b6VF
jIciNOuEghTqfSE9oKfBNoq7TEM56O9JpwPJ0MEq3rsiJ4QL6UPaq7yjKhniGI6Tj6BBLCqglvA0
9OloOikSvG7m0HGn5jqY8lz+CndVbrRmgXXmb8RiQ7kdnGVXkZTv3WnBKGZLGk8CAtSFli3+cduo
/97kqllaPGucqx5LQperIxzKbEmlm8XZNt89D09m9ITi6qMAGiZNr7qzB0LG3LFwYHvicilxIDAS
dPvtUswjPo/Dpx7fD32XY6Thz3GYprzshOTuTC/2zL6t7QK7cOX+ftI+Oa53plg8fFPOt9ZRC4es
ExLQ0gMt3WhNikc3HYJ2GZDbs6jWzaJtU+kqepPMWdD+pclCSOC6VA4Q4XarUz8wJ1TXipc/hC2t
g/lQm0x8pnPh+DLU0su/ouGQdPO359OMi54ZG5kaO7XecJekkuTv6p3X2FF3Iy1jHVfPiC8M2nHt
4RQF2HMAdnlMFtiwD0sMoAoNVvzJbYouTfgHLk2KyU9uU76mjvSraT8rZJRpetb64KC5faApxqr4
iDxWhGbtnv5iKnEpZT0Ed+CA55KxqNkN0uh5gk+bVp6lJ38tX1TxHp5CxjSyoLUFPdMptxoisDmE
hu+uw4N0WUS3OApo9GrE6rojK69BT1i/+VJ1pDv5Co2/njWMM21VpLAE1zygQDcAGWeOYoNEZi3u
0xBzvQZIGHMW2/T39HR4EsoC5Rgn9LVc9oleJlLMOLvq/BQN3pPKY+cBbhQQ0y02A4VNbZDYLkk3
K71lUlbuKEXT9yDld3fRKyeDpsYAjQ1BA5SAlbtzgYdrQKthUgW5xXEKAjszHPoolRgOH+GsZxSk
fc06ff0l06UmMMoSaqzuf1dK68USeLQIzxHbM0wvmkTPxPQ71CMd1Ppuw6vATT2F73CnlWNk6tPy
kWg9VRCifpF20QrFmy2geMGKf9Vr8q570amKHXcXxKZwqru78oTpb/dSyar4Xp4Lz/8AKyNzLqoY
vrkKEdinRyelu0VAp3cOtV3X+O2D/HCVU4YEIzZHI4NQZTB+tBG7dMBdmi909CjEYXo9/8qOl37W
P2SRAGVw91i+uWELz5IelrAwF6d0XGAy/rYOX3QKlAYnbnei6rx7vUiLk4l6Cr+ut0bCMhgL5gC8
ZPBzzcZHchan+ZWrIf/yfweVFnoGMX7+soRg1vGJR1l6TttTejaPu11i9SQNvLsya9k1+h/vc0YT
pGfudn0+q6vBJFbJ33kHZiHkyfAGRslngASm0ED6ZDI8xlLHsC6v+G5rO/tKXA/vAJPvRor+ApFb
Fil5+Wc283ddqW/ypqH2yQ0tTe5rdTl/liZpWjfaLRAMJv/qpcln4iRhBZno6r4Z/p/K0LwKpTka
2GsoI7lTWpe8yhohxaJbkSzhQVAaG3ylpNzF1GAqeVZRz/6PK52g56kuQP/omCRuCd4C7t2PD5tO
eCl+5o7CZ4s7F8JE6hFmwc/hDTJp6pU3jW0yHbdP65ikbrX6qNaLh/3qYUE09KqMCBayOC4pCP3a
ihdqiBbcsGglUiZL56xKUWqqTvwwJlngJme3LAYsaa17PaqWBkhevrxerH8R9pFyh64xCkjD19Ac
nfnh8vM6wFDv3r6AsNByttQi1yx7/nhEXusDR01dRy86dRxO32aKfHHYgFlVLqhSqCVTR4pd4y+2
b2x87alr89YWBrGUgq8kNjY0k7ODkOKRShEDROLJTQmEfI4EQaI/jdDLVnY/DcH6RntKPRNOXyoo
d07EgoKk5HnZXAD9pEZZ+AF8/NAr2x91Fb3ZizW0G2rrRC5t8557Pmm27iX3NddjXqcu+HtOaWxR
yaxNRnbYfNJ0rM1N6z4jd3IHxDsDQPq2dqd7uHbUHJopWyFXJ+80YQKPJEXHIYuWE86beWqqUG9z
U8jojC3I2uglTzSx5oc2gsm80SxD061/1ldKa6o9ZIDJy3LEvySHJ1Jt91K8LU3l17Wr1YYfyDab
tGRQm7/JsSMcqs/oTBF7AjwHEUYpFTq6owGRnC84keYfBs/qxebzEeYZMJM+u7q51zHer8neiz7r
EYdbtelj0rZk7PFv/Z5lXroJmANIrVBHCpOuMFNKHGwYuwkmxgE5hvLIwSjGBs7Q8ApBqwB/DgbK
nKuisSrBJMffHqq9lQJAtOeyvVGvp43HVtJsVzfNU8JjNmE55erAykEu5Rc8wG9Fy1aA0h2HWnJ+
G0mAaruWV43H9tVfUd41SRHvE7mYD6IlnBnCRSVs6iFKssN4QowI+FTKYFVLWvLdyxNm8SCoOTwu
+ioRKKqC3rhua2gDZTc4+XkUw2hAJSgMu9/mUJMVnBZjliRxl4FGHMdKFf7kGtpVf8VUtZjzGJIN
x1HQHCy7GbvizJ6NhkRPAW7TdterkMzHvfm5ZB/BUy8Qrrnbc7zmT+q4f708yb1rasjZKnGt+des
f8cEj7Jyv0gcfiBM0kfXE8m8Z3Jcm1fmmvb6UrpME9qw7fM8Pfiuemjnj90PIKfC4hsbLQpYxcra
y9SIQgRB71UvdCr/Eji0BO8vCUcoYYE4zO6gmJwnPK3jlJ59+HClmRAB3s5faKyi04tC1HF72oRK
6ZyRt09G1DTKdnT5q1+4wdZKcnml0DSqNlLDrYRssAg9B/DxSQAGYumOW6F+acnlXK7NE4/cNThD
T9+CAomOtvIwBP05y33H3JaQ2JJRzjkH9Y6VGVpiID7rqBvaDwJPKzwCB7UMF/FLG8rFdK9MoATV
9MZ0MHPl9HAHdjANrLTQnwrILOK9wjrF9CHvNJalSVgw5oOG8rkaq7dytjgrhtgZOfD0KDJf79p5
++HRt1/9PSWwVL51TR2QhNpF/fxd/hYB+Ga93pfNBAhWZUKn/38N88kSED8dYOgsDl3ZKcz1Z/zw
p3D2ZQdhdWSYQaWSqBxqEIWEZTDQ055qzsceKX5i1yhjZla5i2Ka4UjoBCVU1tnjRiWRZVqboyxD
HPKwYtZEva1oZosR0HnVGMhIdOgviuA2ptZToMhEYCZ6+xy35v0PXSPCGFKdGHfs1hYtallrgwUI
DFrNaX6cIllylcnavshBXBK8ulbrWkcTkdQpCVEEPK6HjdXfABAp7JQFOs6bbPGangnCKmkKQyvX
K+L20NVO/do9ixYIei+yCLYGagygyqrt+9bwVsb338/shxkZFqdd9xeveYbB6s6SRt93W5bTrDTJ
A/d4/lsvGQZRYnaJb93vqdJetXZchLm6jlIWpUsGwGs3XNCbbe6wfxE+aG2C2lNyMdLhRNya9B8M
JDl/en6GLB+3IGQ+mH9Ar0NvngmtMxytAVKyk/0PiW9apWi5VrO5HQX0l4MYXfLHGo6rDSnX3rZI
YuVc7F9qb+ZSPBovMDkOvEL6etDqNmgjg7lBBp7EVmXSf12oQ3i3mQFo23N0nbK6OrE5kTzqIYnr
3qMmC7kAXJr/83ykYS2GQnC9ySqFKsGcR/IMES/ZMRaAuYuXWRm6i5qKhLmL+kkozZGGcvOI2Wmu
mENAaTALLjJaxWNUIfBlcn9FUn12Gzbn9w/GNqfG/RxYjWN79uK+LJVMW1p1CqNSgIP7LHC+TWkd
qi3ouZp+6SfL14uW9L5ICsTxb5VsfVRbxgYozgWptUXNahJupdXjOFLv7LJfUPo1kS3kPOg3KZXl
9FS6wfieNFO+I/ifM9DmYyeLSvE9NXkO0+87R5ggKKEpbyKarD3hDB2gEg021pyJJvrm3Y5K/vmz
nsLfP7c+1ec3E02czh78JSC11dCJgCCsSFFce2IEYcyCTCkPIdTULEEQ7cYwJn8ZHY7HJ1+/UZJ+
gng1t2KMR2hWG60VGhd8SE+CMarHqR1n0pltP8lr58qYU3b81vEExQ/e26kHk9w4WwwmXDuEnKXa
YC1uIAr/OaDxGdBt3dd+R144jfV0z/lan3BDS5Uo19AdWQQ+cUFhv520D8chubOtisdVpNNIR+7i
lG0h4OjmHSJdSG4RfGGUqoF25kELhYkuRyxSJIJhDiqXhw4PgwduSSH2bM19LHOvYL4vPFD+Pin2
rI3IliDE82VzSyhlzun56NOULrM6gklTHFLvVS3Ak/WtKBz9aPZCIo9l2UmGxFf05AeR8e8igh7v
HgMBrc4ROcbbYx1zT9qvmK0rz4OWUC8Fme3auE6rgqswy4Qr0Ea6sO/a3eSsPsrWlVgYjyaq/sFT
8oIuQkwESUcqlY+fikHmNiceMdrxjwpyslvM0x1tD5J+d9cVttEf/zu34Xs9kTWCP5L3q8ZL+NEu
JmcPnyl3KZMVumaHBWxFl4Iu/1r2yq/k7Xta51uLfsf7y0sh9Jp0VA43XUTwq6WKiiK7GcLZNycI
mDll4Z/pidBC2CZQmn0h2A9dOpIS1JSBtz0nj0UE7dWReSfffjGsaL+KVatRlPKvEMJkr9QAxnq3
krAI2gb+HkV4TxwH7BKYaASzWYT0r0TYD2IH/SdmIX2/1BoQoYv4rGRAO9kMDuOswTM6YWKZ0bi3
DNQaF91EagnqMkodup5MfqV4cJzYzIGE3qExaAQANvVfGtHstG+0ZnBMnpWrKk9PBaXYkjj/5QzU
PVyX/FZHjZxkbpKaUcIL2JghUUWRgoEkyEP8YjdNf8yx7BsPR8+4vm4DipOlRZ0IGm1Rba95bBua
BxqA/HTTmNaKFFfGH0pH393gQ0ScDZ6BBpiay1wYrcYVtKHKn+1s8GZZ6hf4b5Md6OBYEktN96Kr
lMBeUhSq7Pr6fNpKaayVhRmzt657QA2huubOjBEHmPWxU3kuWO3pbFr2gGbwPrL7LC/6IKJXGMPn
0Y5cFLMrYZ9DWVyVWhBpfQZPG1e715qfGfD1N6vEm4UbzLgH/PcEVErrptWAJN8aAr4ksdHYODbu
tWkkEajviiGZQPVH1Q2w/11jG1x4BC326JcNK3hu0OVJjmo/TgCBURyURHbXuQx8k4TALbPBzqnl
OlS8EIKmrM9WrQWbUrTuL8yBd9cG30M5fxe2f62UTgrdrk3x3UJO97fzA19yZ9X7Yj/Nqz7ZCHW9
fqGtmc22UBUIwAuV+B+GjCACkav72cEbkAxtsROX0mLi8RbZ3m3+EVpvPvehrm51damfJlELsCsv
FjWFey39r24pWW4GWIWig9/aKJc/WyH6WktQUE4cJ4jrmlTvkblDYTszBdXvg7TibIo2Eglf8CEM
9UAL5ABkUVcwTIqID12YrO+idFdbIfw9K/MPY4nEJ99jak2bReTKL2qVKWcAt/PABdNztOZFFBlh
tLRAQQXR9rSANZGMgfuqkB3/BCc6zBSt+86LgD37FRWPuZ0rGQzbfR98QPCBWnoNL3ZuRaj5r23q
cd4/eyfMgdubXmXDufGyaRe8YuJeuBYKVh31uY2WAsKe9JL2lEUhpXahyYVRHAlbV4kTYivNbSBQ
H49VyA75CPn3s+hm9zn0rYpWVqGEunmLW8g1WsVxHCo+0NW18l2NdIW2nWzuCf9Yysk5jcJPEOcK
PAzoVRGD1aQNDWDEXPzebD7nE+chJjpPFQYH90m1Asy4Hegc+I4c/+RiYFvWHtQHE78K14ZKSueB
P2uK4Xc85Vnm/LZJR/gZyKt1ujy0TEP8XD31XAAl/Uk6q9h75u3q7pyqXVaeHqp67b5o0PWH82AF
9heOojX8iwEX+ODuDQHYRp8SaIa+xqyUYlfbgbCHkImwYyU9+0OVKdgRQAsoc0+yqXq2wrH8RJWe
TXxBWof3LBe0mJl+M0ns/WyNPW88JdwpodEnI8czbrjf1yxmDYcINSZ9Zg4TsFTa/YDdb12QqYx0
XPEMjAhH/pyhoLOO/cLbUCUNs+jNRycIdWc58acEqNzRT38HmCxHmcUqWF1wybxmS6G0HgyDR9Jp
GkoX84U2DGRtwUwdzAHw/80NNDi/8fmCz+HKSRhyCaJP3RgQoLS5PCRpI6lcop83XSZiAYsZdVrW
SY7y2IJkHQC0bs/zGk27qbajHR3Rv52Iu7ygUw07HlqhZNRBYgWq+D4BkKSOpKwlVNtpRgGZ/bxI
AVXq+NenziJwz3iZIJG20AfKvXmng2CGt9vfsPynz87+wpHOuUI3ESjUzPYmLCyfZPjPOJr3/X5J
/Z71dbXvHbzxNX8wM2bztO4Pz4pLiZRHWSpQLiKM8PwT8pZUEO75oTCYwpSntLv9nMNJ5aKj+fWv
NG50fJ1HY1kBaBJRoVynZW8zgKQOoJM3tdBa8az7fkFb4txBnFVdr3CyWdXpuaR15YS67vRf1O+a
MrO3sBCKfXJvJKgPNzHXumvea28N4m9ODgIhc08BFrK9/+xLOwUC8OFEIonHKmM4BOwEB4uxFfpt
K6UrJpuRS8texhPewBmdbtD2Ie3LWnTJJXa1eUfxijNRaUBuBUjPF2OTlH3KEgfbpFO3V9djQ82U
9J6MAdkCSn+75LDFNSAHmVFMO7OLcBFC5gClFI5gEiqcUCgxokm2ywL5dPe1ZduiILR5RLJnq99i
fplu39QPGiaV6poCqA4KzDKL+pw4j0VnbiyG9qYHhkG6I37pFlzEyKtf1JqwGx0EMPpBZgBvnY9f
8DjSWwMbsXzfu3YSm5MRPnmkzmF5FBxaRiBPP5VAuzRIi1GQlWePSg0t3/5TqTok8aiATqWhkiTL
eyq7GC7sP9Xytc5u/8apKRMS+GwcIJqzUdriuGCBGydGDwjC7AE7HUWabtitpKPxu/aP/+mzEo7F
aZr1WH37byBztK45N8FSbj2aJp8H1Vv+pu9unYutAThszbGhr7nIlH/BmW9LSio+h/9wEX5fQX1/
Htjrn7FAokdHir94KqaGM7adR8NOsUPHsfI7S/UNOrkjELLoNeU2jCr5JQNlA95gSg3XOrYOUmvu
GvXDdQmFb5KgOV99Ao8NUOBPCT0ZYYJmr6UsoHamu69J/+f6BbnDVBvh4RyeiBvx/BF50OhzRKcS
27MzmYx1EjUR1BVOt6I3nM2nQx/L+MNhVMHatMrGWfni2CXCI02Jjfg5jKCzMYOuuubCdAXVm1Ly
gl8LjHDASX7nWLoP9mHDZNwMdr1k+MxV5XCO4gUKWDOq/UdvjJ3HX6H5FI+0wPboLgz8zV6bdt73
psr0IMPmHU0wnQsSvFYDkexLKc2IYUSJflVqO68Q9QzWPqULBKL2GqiH3/1dyDCroB+IB5qmVs18
JODjSnxDlD2iMN4VG38jHTt12/+3euXSCqGQt9GoDMehjW1RuvvCMT2GB4WEq57GW8YqPwW/mj4Q
PrFiq7h3TjIkS9AFDOtSF190NjXYvLeQtNSYr3jaUhPw9qTnyNoRONx1YWDIeWfk9zmQldHjlTGS
lvT5c7TcQ80hO/VdcnHEgXIC6/ugY6yq27lbatpANo2wuFeZqglTe44VAeYzNM0DLEL4uBJWp1ap
Oc6YddML/k4CH0/YJGOKzT9893vssbptNSa9HvpYwuGzjFKOAuVvl8JVRqYC2owyjJGu3pIAV/sZ
SoG+yxrBfb9wIxhO/6XKFbBT+Kpn7fQ77EUTejx2QQDQiyMIdKhgIVkSlxRA7wyP8NXtAx8cZEk9
Kt9+dHRRRuKUmPkYEXQOxjhY5902eQcXTalgEDxHRFD/LmmZeuCxBymx7+i6bzU2byZgTU98jEd8
NopLAUfpyMgbVWUgMOsrpit8C7kgWbr9XyVS5lMs0gMJ7ZR+h50phGTE6gH3OY9tmd5OiuaHimkb
0lvK1rfQ/LWNKSuI6HylxZZGe/m8AY2Ad+f29ZMQl6MevDEu3U8rWbauZzffduT+gQ/rvk00y2gS
FNOCt3xCQobXzNy5pzVvs/ezPCFDWipKJ5HAWnuyw1IQA2lqnJO874ppvB9aYe6GVuCLVajYAYgi
DXyMN/h8lW1kCzkPbuJDvYzsTggWx570IkfJFFmDzl8hvebOmcHcVsqi8tc3reUjnpsOvw9vHmAF
gfmO43NsplgkjxOyfSdMi/07C1zNJFmKgoV8+JwdqDe3iQ8chWzdGZVmWDJkmCiGR9Tl61RPREfz
gnQ9PD8TOe1L5/zKzlairSsD2O+fldN7RiCWo3cdpYEbMJwCVgHuszjb9+c6jiZs0xGQVJ53xwDu
+yX7/L3LRa1R28ujJDAShuSAGWZWEWjgvF6bON1xaROka/KPU49tukfbJiBqQ8MqN4fTYLd+5deq
0fMZQzbpWu/gmnp10i8t8zKS6HpX38qfLY7H6JMKhZZL+v9jnxpCNztxPLoMMwh7krBHB07gIOws
cxMIINDwN+Bc+i/MCKbfpKCKecod5ZIfE1rEr4TDOVjOBAHsRV5FpOXrA9NndoVxQmfvAq8U6X1f
Sty0wfdv2/fRouG+wKZsgZW7nbCdmsE/x0/wkXdZDx5vijILVWnnAbEzrRD3BatQfdbaJtxQEtEI
E03CDlfmueEjioRlkQoWh0GB9Vs/kLDei+YZFqLDdcZRFSDV6CJ6EWEGmshXb/TDdMpy7PKQfLlZ
MaFzCVR/rHXgkvEmtadkJt/36nAKDjgGiXjOVxg3adJs4SKkLR2kui8jpVpqMifuj0SA4nIRE/Ea
6KhQe+LpdfaGG070XOP/V+lKG0ykX3e7AOO5VKWKFpJmpES8jA3oAhH8FvB95m3Fpyv0YvDuOkm8
QWk2WEDF+9Bmt9tQtXBpNfI4jEiHAanUlMrpiZx4RMteNBMb4mE6IFNohpuNX/mt+Cc+6hfF6tEm
H2iVay+erLdzpKezKnZHGnoK2I2Cu/216jn8htqcnANiH2xbrqpVIFtUtmh5d3gup5sX1tI3KyTX
7bBhGSvhB5idDQ2h4chGSwTLjpST/jpO8mefehKC5mHBUukBgzV1whNuV7DiSOEFADLM3WT+x31d
QLWFKldWzYYBnM7qwIcTX7c1/Dn99NzwFcwBPWX+38o4D0EShtfoM7TLMNowOSOH3j6MsVuv3u/0
3yV60T4cHxn0NEisjtuBLRD0RFnqbiZ3LLfHPKUPkA1pAHFF3nPiTteEHVsmHSM8apa3k027j9dU
Y/70Hg7Q3bQGhWWAAkX8SeIGx3Foa4zc9Z4mU6oCusuWTN2KWFkTzmfDcsXX+G/9xp10SQ5KMYnf
rTeozfWnaA23FmWg3nvXXwj+z61Y4KlZYar6B9BCWd4PJ/GgDjT3/jhMais3N87vpBPyWj5/qJhe
7r28oFbK6opWGRO3CN4GiTEamafc2QiuZsSJRpo3WpyZoYFkOyLDWM3HlmFdfRuJyywtFRmrKHFl
kBeKhyJiEpVq4+ET7+DJptgPurWUte5zSO8vUnZtaePOQKGKv/4HcxHfu7CzMGSqPdq7aRvNa7Au
vl0nxXYCOI4VW9Q17ySow1X3vH9tuGxxijv222OyA5D8e9L8fLV7+7Yl/3ysCfaWR0+a+xKmAH2m
bTK6sYkri1fEFhg8snTXOQYw3D5parw2YgAI4UPwe+BIaPX7mzXLznWkAIaBSSErbO5KNExnNqtU
yaV0VHa6SEDBK8avuErcfBUfx5z3vLwR1+Jrk1yT6vlBhrdEffVJAKUqqu+0+MwayI5FTuGBU2e4
jAObXesAiw9jYAkXQxVZj0rxApB2wpW67+sIjEZF4ryKeQ0P4itK+Atrqt/wNxJ9qTnxGUz00fuP
qouZrCjD1jL0g/yBgFE0GEK8jKVauNxqJLCBcrNARaAmtVE0w6wi7+dh6em79N/gzVRh/OQ0qTTb
PTewe9ZRa05feL0bliGHhpbDq9N2n18whDLq5ekBcUubFMFQl9SFearrQcSSvEz6yhx9FBKP3Oho
efoY6W8OL4w9ZTWIcpAafSIVjdHWQMRJXOFypCENrh7U3JlVEAOAeTgUupGBVU2sSJVX9YN/4fdm
VGHtSMmbm+MLLo9QjwEyiJpjcfC4D7kRuCCXIsMxTMhvTWl+9R6viN/CrC5/oO9K/Q1f4AXIwnyt
KF8UYryzoMwPwyj9CX29dqx7pr5AMTSeVXJPalB0KAYL7mT1d7IbTRPgBSy4bbx1yBgdZvstSPkR
BDCz1mUOA/38OskFTGbrrrwL0NXcQBxhxDUR/L9+/b0THB7ghrpA4Rb9X8XSuSBHQwm2FGYvperI
JT6VHPdMxPndbBQl3v58din20pjcSMwednblOiw2tfrncPdItvs18Q7dZ/aIlRuefP8jaW76io91
LJO8+a1nRrWdF1YOX9mORS8TUX6z5sXruCoK7OSL4QWl02SZlGw7xNW9E3B4TFyrliTu8nTqCO+5
KqJD/gnMEQF+7QnUu12c6O4V7VLpPNJNW2GkVdETFQzqEx5VT801zvY3DUKtjVuPAyWkFJIDdhJM
MPr/u8JYJQtNrBNWPZ/2QiHhIX3vwA7FcBMpI4zXVjAEt5eqp34nm689LY7ieFrUvtEcKBdQqI3W
zWb1EZ6oIkU3CGEirtXvduCJaP5/6cdAuyYXh0rXYvNqx1nFTtPrrjmdepIxSlrgozHzvXDebS+v
YqY1tJzEM4H3eX69lZjqr+kZzMl8gCU0L1dv+EHje/qgIsrQ18iV6fNGPaO1leDh7dDEXP5K2EtF
62me5E3Gn4crCnZvTgqHLddBlw91Gvl8xH3QB7mSWw1xq+wAi9x0ay/gO8OHYGZop0IGBmGqX8kk
gy69NV4z0cqKhr+Ej0kp6UGYvDWJmQmAYLs5IX+pY2P5BBjD03rEVrwlQJB5Z94BIj5ZmRk/hr2M
YffmjiBwzYPNMWpNgxhJfqN54dN8jMgILWk3Wn2tdbKc/vSrj3PKznFfu9BHW7/bkXITyOymNP+c
Mxec9M0D9zZgwfW80Sq4q1LSP3SueKel6JTdrbHWXdj9XoxkgQApID7JzWHdsPZxQU+CYaB5Y1Gb
4vkbFqZp6nZ32d/4dviy+ME2nhNELTs6hQ5MKMeuqdgYSF4989na2q5XW8G1eBDaRuSWilZPGEJ0
0DnkTenxh4Vh0H/CC85s2lWBgx+KfaSl40pR95wXWtZYtRy/bu6z7uKggaR2Xk7QuXk84A/UyZWE
dq00sat8gFx7jDTumlrxW6kBmEzOVnFUxsKLivA/RuVP27d6r1KrEbSzg2mzYvcKqyXsbkdhprzP
p8++yRmjTtbCfFM19Nc3W4yY+WFEsyava2jiMCT7DXA7J9uyrc3NjrCN+FtIQJ/o6XGtVHqEm3r3
Ebf1138EBFueXsBRUxiVjENnFJa1OFX0TWfKAGb+cQBYFCQMPI6cbzDGIvnwupmfl6v4qf5YmLtI
zbt/RhkpjbBIGRtbUDr0Zzmfk7wR1Nowa4fNHh1gVqxOy25HkQqSqC342mIjvr0qxJvKPbZmE5bf
tm0WyygIovKu6m5Gn/Hcv4yLPO/r0Nf3JPyaw4inAR5Jo9cEKlLAYgRdOs/isJFdXxYkRhmASDs3
BjInqHXpM67aBrNSCBMPjDPtdgV6CTK9LvGyMLj0UgVj4OqUGK/HiuE7wmZuxHDlamdDbB01R5bC
muH9QhbMZMdWj+kyBYLsWgGBGjdwtyHyeAm4Y929VYbqTuWmDnxLqKjOssuBeqxuMcclBjBSUKPH
tvPA92IqNE1joPmIu1X7CDuGE7Mx1DFUyelQJFCd3ANAbbuDARRl7cET7IXE5u/t1bH0oAAvFxIw
Aj+ykWg54ZssMn+Ex+RMAaGG8tlUvl6mur3M44XBa8F5kcoV7X7lCqzsxZ4niWNOEngxDDVHbA2f
4tNC995RQOehITTJPi0jKfesILhn2TTlOOOlbranRIfNZldlcEwv2CrpYvspBbSj/d903SmQ7mDj
DE2BOPvnHugmlelMwLNJDrc953KEDESAiEmxTSJRV2Qo/Bb/eRMQC+lhlI6HEop7QanlYXLDMDBo
99R7KvjWXipS1WWK1rvySmZbJ5knLnFzl5WR215CDudhU42+sQQN+Av521yiEdN/rZrpCHRHnBjc
10hTjxKcAY/dXr/i5qR10Mv7/fvd+Fi9QFVMVjFQDTDSx34xbFUqEn7ypCLrpQc0WALPotXwQQws
ok8tsWZdhm4ddDbvjrpDzGBqFsP/wMkmL7lfZLGd4r55JUROeO0+mY+fca9ai+oVmRrcz/vd+W9E
cQg9/5eMz6HBWcsLkoZSs9oUnN0xesQOScpBINVa2n56FaTilwo8wz8gqSQqwAYU0t3XaPQ08+A5
+8nZR0WuVc5rzDzsyKgQJADwmZ1BRzcEgzv0KuhrsUWVx68JlvfUtx2WibQImnIcVzOVf2fSkBd4
flK4Bu9BFzCg1XCyuHxrqNiU6vw+YqmoL1yfzaxGDSEDHjN3z9NIt1Dhd/bKsfqfYiBeEp0ERYQg
OY3Uicq2A86pfFaywPoxfJO6tRcRV4Z2aHcr+3IVsiWqOtgaTgVQRvNQLIqzRacqSG+QjBpUf6sa
Wy5mCdCeMmfxeDqPxBqnX2Fqu7BZDO6XcRv6vFEmWIgxjvlPn0b8RLnhrSgO0lyCrnXkRI3cXqtg
DKALQt+nXYmNC1QQVWpwsbUPeEZg85NV4ylv9KKQ1RvXiQS9p/jjiFCI5TH0DQLxZjGYN0xRn5uz
1slMsPHoXgvA2JbUHUG5MlLVWOn/DRTrYD4LUFJ+jdQ/xpxcAffkKNbAVu0qbRk5gfFO/gfFVsEK
3KSsP9Nsd72xlqOAXGs6Wu8/+xLHkbr1EH1BrjvBCTsD35mqGgo1WKg1kP3EMc8qu1EiqEugTP/D
qS8Az+wTx887zuFrg+pz8THCi3K8feDN+6l3RWftcgIhWDmGeRbDBpvuuCKB8/hV50Cxbf6d2Jbo
QZs+DJabwvvpLPuxPHHx4//DfI6fOd3ZT2Sq3v17wjmQ80PSjV6CU2xxgzuEQenCHizZ9Z7LkDc9
/cXKSIKXQk7f9J4MEnTnbL4HjlpgprEYt86wJK3QHwSDCNZdr8FIwg82fL0HoYwHSNlkRbTfHkpN
Y9jiMtRYZkL3Gx1Rh+7UG53wHbj6USbo9IP2YokS9xfpGSy0XZDSnDRmOgPZW5HPQ7alg2tN1RGI
CKx8Wv6rijkmJG8fMxeuMTawCexERBCyWKCy5wkicQsHRVVB56guu2jmmwNYdkKb2FpHZ9vvHDSY
/HEbV69dIpWrS8OPqVshBM45CFcf9VU+9LYmOTIZs00bNk0iAYa1tM3FLMJgMxxTB0OFfsojjTBh
0xawwqyGPrWNHBITpaQjORf4fefHlHXNkzYCppzWRDa3FjysquVEPWVGOXki2Db9WK/D1elZ/64z
FMM5kdNC512hVuz+XvsZRUPBwQ9ZzxMMG9zEIsd5lbdNRL2jeithyn0WEt9xGLrCFctSWCqW/2Tk
AdFgDZnQPnD5C/nhBbeIKi5rO8fW0PxjW2xvR1EqcXsko8b/GbnLNOkASXrHfc95oT2rjw6nW3u8
wvQkC7BnFabdQ69qcNmYg3rA766vaDagvqRBqh780I9ZCKfle9JsU2G5uQLwE9bVwVOfAOaftZAY
jjxQ3rxJmYZYp7FzuEKV9xZtvWeT1NXuHKqBZvvg5xoMEfbbWFwBfJPU8crMcoBQVmSIHOumGUi9
SjNB2VnL0B+ssJUcYwIVwCwJSEaqAIyiXHID///7MFTy7wsmb03tovK8pg2mYBJrF6uPDv8r9G3n
/0lhZsdpArK18q1iKE6F5/R/fBGgwsEPXbCrjqy/qed99UQ588vwDO3TgDzQlxF7xM/Z7GNM1KpO
dIKZeTXCgNlteoRUV5xk6p0H6fK4+iuTT0/wCQP7iiA7SUKFZd3BmkxTBxABWpEeKVHQZ/1DB2F2
GKGS2ElryhHGc1tZdFqoxioXXi+gZp2geSCpOyZuapojeqQIUr1d7npvHpGi2JI/U7jERKUqNq4o
Kevs0O6fmSHyuJTuKMCfEIIFG1NgyISCTbCbPyOFk/GWoBQ2jkBHSusG/FlVsiLpT/ARLbuo+gKE
z3HzoFx5zNIYGHHpZbgIxhsP2psUmAVmy2pxdyQAiQt77a1TIjax0R/236Yxb5mGHyD7vt8ox4Cw
bk9xtK/ZBy1JOAJrJ3J++3eiZira0XccM1xzAfUO1BlYiSKMeXuRBgAuouElpr3+dtttpLcoAr7j
b8CKWGRLBj5t3a08H0wjQ0Pe8A9uFQ13cmT8w/tDySsMgjGjPWcI2XoCYJivHqq8N8kasuRO6vy7
UBzFtkmrnOqj9MqE4jEm5CIZBoQH4kEq7YwlVGpBJfQVpJtPk/flhmyySHDh7Z3ZaFpwsco42sWh
lC5gC9Z+MjTOSjVbkCThCNW7vlDRok0+uTfIsASWXoDEPojkgj7xVOLhood3f+h9uoTttv3RSwGZ
hN76bnRB0ktkAkx0+agp6DEOA/GKjIqS8oL7aerNE1/RNah6yI6gpp+/rH32yZcCSTjaYCLsPeZg
kSHg1UE2ZzuRXglzP2IOMkBKhQE4iOP9YSBJh871W3HMLGZAqI6T/V9vaRVtg0p1FOkVKUH2UvJT
zeUdm5pgoIgtd4PybFBP9U991E+9AgBx799GG/fJk+pY+70ktDNNaCElGIV+yCM2uSxOGw8O/1H9
DIUgXE27AJhtFudUTc3JhvtY67OlRf32IQo4oJGcXwq38564VoqG4X5FENmvPh+PB16h/SHm9krT
AlxPADe5O6yUzFJ3CNPJG96Q48v8RmWNkFfixa7OQ4XgnpmL7gmwj0wa1mqH9rAKDiHieqYqlieY
VqQudev+5jB36mHJvWNglxk9GNJdzXzmRLH12a+i+3wVcQgHpySen7BNx3dpVPMs7aVuIG5qrd7P
3tNokVZTp9RUxBLxAyJrCkQlPwT9of1M2VmTWBEWXMeLNxwc+ZEEreUo0CVGj3/sjUlG0Huc8Tkx
w8G/EKKquHsqIT4MwiAlFkUjz6mGeYG5I8s2DjLhZjUMdcTB2y5efcJdqyUdQd98m+OE2lR3orwm
6FjGSVcUGv7mG2QUGULyQG4VIaYIoPqnWOwzlZnGjyJp3p2Bl417KoFQgBOE7TEfXUQMU/XTvQwp
5qufkitr97cWsVUP/A55w69KPpO8pWJbLKKPMZ/UgZ55jxrQgkM5mY6d28IFb2K8X/Y9/NV35rkF
vLh0kKuvcTDflspGH1L8iylPwgvMBzueIicNdKmnrebQPbTVMaFMyYtfiCPCZsTyVV2PNAh7EoG0
UW5p0xXn19D/xHskck9JDVdDn519ArbzZAqszY+ib4h8+6d3Fk3zSHR67nctDaXqv35i0/v8PvLC
uVH/obF/ny9SfbbahQC5luAxT2reHucG0B7xffbZzE/jZ8t8E3jYI4VhbdCCTyP19xNFf0SOwHVs
Df8lOyYT1wNaEnXeYljI5PZ1H2mkcpdL/b0h5Lg+M0lkdTl74mgktBXbq4xOnyUuopeCmZh1aCaf
JhvPHNFHhoyH6DohtdbsMrVZhN8A/N2rkE/Hdd9YKwXkta39brhhv6smuVip4lsVhg3x1WSqalxs
7Iv8sIuJeIjMfPj1TG/66IAraglVG3SK6Nm0dxVxDR/HIHLcIYjYrGPzTHxyqZcglQKDAvFSYvVF
JnA3g66SPbcrQLB2d4WxYpkIzznEif0oKfbIwpVkLbwkLQpgFvXKi8eiXSPU45asXso+RNcnFci6
n6s10ejKJ7SnaR6A0h+L5IwZLP4Eb/KcBkNVbHTDGU13X8f4Hxc/ack4/Y4L7DHB+KRLJF9JQVgA
H9q3Kn5qsBLzR23kyTUuWD4ME5e6Eor8JVQdZoR2tExXNlKxethmHL6waVNoUcanLfoCz/9TvrVx
pWJ+R8bqYj3BxSW2BUWCrOqKYApbV+eFz1wVNjlbWv3JJxfdoM8c/XkkdhDFeraAUz1Ya9FO31bG
vyRhGZEktsKBT/pXjZ4Hv04vA/sBT6fbp0fT2+iXFt2I19T6k37r6jPxoMVTBx3cPldCoByqGspi
U4vGuxxFNZHJyldWKflNi+7fEZtud8w+DIhfNh+xvu0/EBPMeif8BavJ0XEGxd5VJ4wAveP9y7PI
LTOkXY/9MRyoWfhE7omrdtZRMM07RqbWxD5mkEoxJCDiS0BFxlS2hQNJLXT4Rzghobb5a/rbLhXB
DU0qj5yU4nLv1BObHG1xJHH+Qh+prMv2WsHQTAa44m6S0rfaLsp7IjC5oKt59lmHDcujxZgIly2O
dCeDuc9UON7RHkWwQo2er0+3S7GgycAEjGu418/hRVJKdynRgfV2PH1XE53uEJqYixlJxYwGMOYv
fXSdRW4Py87w1/udR0N+MJio0nJL9iuzoIShyRUm14sUSIh0vCEk4seL0KBoPeCPj6ATXWcSN/3C
WI6z6lOrAF4nxBWVH2xWHam1pmk+SiLTo+B27nKLmwLLS3ZlWgj/2T0lbGHwdR/uFPLT9s8NT3kd
b/K7GDl/xErWo1VmiGInXMxRqbjMs4rSb8F1gJYSpQzfuOb7EX5009IBaI0tkkw+gotjTqvOBLTw
UHR0cu7hy0i4GeaGZKuxH6tRLo1Hg5BKi780RYJstzTZxnqJoInsZqkmLmvdjkMN0pc3ljng0xgs
6/nm3s4Hceq3hoTZFpPfiGX+L5zKid9j4KZfNs0QoXATTdzj6QP1s4p5pFnkr53TMhA/UK+iKWqo
iPupNQrisq2/KBvW+cIKR6l59Uq/n9bnOC4m6jtiM1ND7iEkM/19tidpUoPsi3cgTfz8EzPwpekd
Cc4cGSwh902SHJdErcLA1nZrFm83z5paHj68RKlpexp4bCsG8AYSaEK4p9cZ/GXvETgblxEEJeh5
7Vcq1a0XNEE952X6JeOf63dzq/WQjKRGdx+LrmQFFYW5JoYt6k3nd5CJB2fCozKe4o9cxggYqavN
iTWZ2IhfYNLhg7Jxh/djLhoC/+e8LpxaAs8uNDS+DPVHTtO1vWiFZr39lzKo4kb+dk6JJoOInvo+
IHIp6yS2Zgon8sc7vmjp/lEFqkJu4o4ZeZjSjHJFF2zJMbazmnnYKEgKvSZown4LTCwmANWN2Fxk
VHGln4mLZkzWbU0f0YRsp5bcMJYKCrf4gjUYQHa5hPOV7ns43RsKFytuWcvACClZGAUpwey23NoA
etn+/UfwGERrghHOvadlXS7ajJG2y1cCeZPl/QYF0GlmmFeXr+4syrnFdFM+l/C4qeAw6QeVyWz0
2K8QWxOz0wPr7Bb1eyyo1cghMzcBhorxWKJssHo2DvRh4loiTA26Yiqw0lz63jVxFfRNIt+/j/lz
WralMw514ot5zMBCxTvw0/lSo15hLJ6eEOVpW4SPPlcRBDW+6RyiRpK0TUR+8aNa9RbCZ1oaMgvc
2wluDM9zNxKPKaOV/HtYfqS6pauVmH215sipUug65UEJ/iFVExobbn4CmcqBXaZY8wzMtWsQyMvD
6zsLk+Yod1j6vfXEbyZViB1Usg6bO+4K3MqR3hQPhgHzhv9Fx5Dg6D69wsqEY8TVl+uNk30oWjq+
Iz14YKcyXBBakbEulKoZhSXHQY+vEcagujoUgpzPIVkatNfkF1/YunIQHeld2Nz9BHbYlDoqRo1A
a7B1W9gbok9gPSvDd0l5Gqjhp+vBRSJ4mRwiPjdDmbBAJOg8wkNRWmypNH/DkrgFbI3KC2jSG4LT
ifud8cuupR+h5cifdllYAnncqIO3mqGDcmKwZjYRUacdjvMa8z1y+8QMplMnGV3mxSis2FyCoDcl
N7JyXUBrUsMRye2K4zkl+AswAa5ZEvcKCPm9pEvub0r1EnozASWooC2UW6v9EEjyBJ7EHRVvfyjA
Zo/gNH1maU23lE1mGM2YFx4RNjr19J2QQKo7u1MSZ9ck/T6Q7XzPpupYAjlRkvh//E4OVXFZlaO8
BCc3i35kNS63KX5c/QqwFYJsXBNWrdXxJIazYc97ixyQETuQQLuPlyHMG2TTO30xO1CafNknXQjw
tQsxVB8+gcC4uGen79iQaBX22lwxDaR+BIRx0+tM0bSehUjGFIHU1sz4KUPd//at51mPdVzYnKy4
WmdzVuZ8IVQqAK1TxzlXxXDxL2KK04nJ8cOZigWCYspXBmoPr/rn4Epb9JZP/uuh7h0Mjj+CwDKU
bK5RVivAtU5zkFnO0IXxAPvz8TaBDSkhGS8716Z8OcDaS+JA3qF1f+LENYxJFlD6UDX8Tj1ss2lS
8Bxdk0BhzEU3wr5GdFP5+bv6IW07+PglfhcaKkFC/OeSK1+GlOJqbKD5qdi8/VhymfcROCjj7rAf
5GvzSFkk2xwp4518vgB3ETAZwK42ubTbDPHp4WGQt9EOhMyXcuPzA8a5UWZZy4uffP20Jwmq87G2
0pHYoujZzCQD1Jt+XhCemMqpzw7RNp7ZqQB9IIm3xCXipuqE3QiCw5ZmboWzp8YX3VYjtpE+xzN+
wwuhivzc2GbDRQazaFUHr2/OspYDwSRmVaUzg27CBQaBUtFMEL8GVCGJk4dKi12bFUgiaizdL+8/
o01hsqxz5gmCfzORKUXoMUxnBbJTR0BNNinfwTyzT2Niww5cA+79v1thoolKD4aI1uS+tXEUPkGu
b2wZ/Xue7gZckFmHZxBIkPJpv3V7LfjIDK5eJomB8H2f0SWVUjBqKGgmyxBo/cu5RvphR+naIa75
lRGrdUobRkuS17kUvplU6ts9r574KWkI27gx/sWz/AxOS9IaFQIJVBrp07qAvt/xVKe0dV10Y9Pa
OG7ZMMC/bWg7wyyhVnt8/f29ICO/Ul7zut5FCbG92sEek15sOkQHjEdvuL0cUJBH4paR4oYgRpK6
6cw1EA+NBJ5U4eWJDUhVSmoMVgjvudTXOJ6WdL9JxMdwiu3Bi6v+taVJgvfBGLUMQ2OAMPBDBMTS
+hMO7yEl+AGz677fY7ZKgcIdmoIsTIvTFLBkaq+Vf177dpAmuD9C5E44gXYvYUfY+P/NsS7zRCw1
05bMVc/7NH/mn0PBJn6Sq7Wfh+dEPXq7gbmym9QHyw30yBoAYUjmoQyl83cSXDcUbbi4heuTGB2p
oQVPkywCGV8hhdc3ZRtTTcxYArShzy0ax0ccUQ/09osAKIKV2O9gY+7RLEcIsOYVWXs4s6oNYwga
FeeFpmcfGg5GKCJjMnM7NPpHyViIH7AqWTv4wLIWrM4nbD3ZnsWvD2la4t8+iDAVx2yHifQANKlU
3oOqF9m+CixisxYRGXPgok18zLO5qAlNS+qXYAeqwQMClKOdf8+SLlas4h3aPCqMquO90T/qmBGk
a+ZMgDN0f0Sl9kE0l/gClDZXzG/lu1isSWgW+adazM0hJ6bSvAstRwDNq0BClWrnXfGqx3hR4ODt
81PyKGVFYS4QVAHSaB17OkYmsAOmVvrr/OHx0xvqa3YZonc+jsfbmohkKqqMtsJqlC3/6+sbKvB2
8CEEh2Ta0+lq13UYcF9d9YimgNW6RIIONb60wcW3k+OMwcqnIUAywTcbGd8qV0ZqeQwD1aOZaGYX
JgsBn5rSQhtBUXWH7DEj6TFIN//t10nuKhKtFT4YuRbL26xftHqeZNQ3+8x64Q/rqT/tqKsAnR8V
V8hynk3DBuCHxo2/S2pwdlgOq1/PxW2J80yOJ9Pykpal+bcNbeF6V+H1Jy17mdQIqsHO/zUO/vnu
eHFzpyYz2PnCW8Q11nDvAifADozqgzynTukxxBsw/pj0qXP0Ufo1WqhwKcadmVOkX8qd2T9Skr+0
dt3BxcrbGPlH9MkpxU2mY4cUhYkkY0yVR9XIFCC0VL0shzTYtlaM/jUL/DZP8fhC2x1BSkriews1
Yxp8Ma/cFIwFVJyjfVRp0jEeqHrXfAdCPklHqK2gxkGGudHLoWtIKWOe0faHEOsB9CAlEUk5a8F3
cn70RTthyW0jZSs3jcvYggdqOcgI+/kSth5W9G130xGIMWpQcFyfNqCEBejoRyXd4eRpD8Te0jG6
T/FXf4355MXjOdgOAyfOj+CORp92B3Md/MvRWt9sFxGAUd9CQfVkkob3gud4pJ5uKJb8JqiotRDr
qwTwGrBAHD05lsnw6mNzPB2rwD6/YpjN6al1u+7PZ5RW4viInmTJWJmNMIKm8OTaOV4f/lvJcQr4
6xNtsluBRono0KAT1xgk08K7HfaV/Uq5CUXmpcTnyq8+bc1djP79yYd07ZzMMXziv8xvzL9HffqE
Q7dEeFmjkxhy1TnNlyicd1qTsepdkycYS3Ymf+kg1BjMWMhtCREPAH/BixW8Q7M3c1wT/dlmQ9VV
BHN9KOIUH07Wg5iqaqAj+s00McUG4g5cJMr4vDT4+nBn18mkZ+jLZYLBcf1YMHiUk9t+TXAoEfvW
zJ2F6NxAlkjDYptcxy1f7+t+sKUeVs2HnsurKB9ZjRxxjLqEAZYvCvJne91yIswFsuvwrD0P+IBO
BUd9T6anx7sIv8GvmUKwRguzG2TBVdllm4gRZ7yjcyPfjJaltKXNYhTHx0ad37UZvkesbzF/o6+R
F/4YxkvXWviCkbgOkaLHl9MaNZ2AzR4JyUS6u4tCP0JNk97yqRgbPebCXh7a5oTlqR1lg4BcQmWh
11gDDAjs0srGXAhAMSt0dw9IYpwoRhlemdE2+HhyGoGqdPt/zop/Gj/X+t7TwzFV18XqvT0Lx4m0
CAODXYuylNUldrdbpHoFPwwVBvDUt9op6PS7bd2uF0082loTwnGojV9jxE0I5XefFmle2SUBy5vH
ujM9H8tOizaB3Y5A/DqMN4gHSDU9c1SXRKtc2HlMG6q7u/UuDJF/asUpN9+BcwOzrfy/dRNiPF8g
WDQUCZjXJ/j1PVFO/IaKfjv+87dtvvg7d5276m3cJ4euq4ZfWLSUF51iJL0hLIrBY0dTkkT9dr2G
RhnNmvUwBAQ7Gd6WNj2bXJMnh3FT7s7X3HRG+Vgt+pOIngZKe6gBu/3rB/qqMCedkbLoNpIRZDsC
4P9po1PtNG8vUYQGmUcqfpPiUWR2CYvcHewMJYo1Yi02Pxc5hfkGyYBUsAmHtLtP91HCJSz5g4mS
+9Lwu1rjoz8c23ryahhXerAe8jaYPXxqvEsdg1hxb7WcUjoKnwE4fPPPcY2UD54bzKBLKyrs7Nuo
7XsqUnUy/vXcZjlUlBgvi4DsqdcA4su3gRsHWcyuLRc4AGxevo47HEeenZAZ7c2mRuT4wRUkh0Pb
eCe27IAJurncAwZh5cuN9/2xS/uVvTMGZn9n1PZIcH2xN+hfZO0DgI+dRwBGshGX9dN9wPcy99/0
+y51+zma2S7JU24TIQDUV+vTrpMtDawQChcO9EqXSMgqFuAmMwWyfrD6qhkVM3HS6kPI5iyRCF4M
pzpc1L5tt6hW3j9KqAywAmKd/HLltI7erhJtXdhvNO77DWautRCyrWv/j6f3Y7W8QKhKaTE6wk+N
8k8ZgF7nmNZizXmLtv2Y3LC0H5KWl+eYeYItcdIYkxCaFVSAQlgNBV1z41nFLXGMh/7Be9yi30Fv
uokvDnyHtXsiKY/y5J9agHh5Diwz5TiI2JRKOOEcJNfOsToljjI/G6pRWrFagXaecO4V4jXy5R5B
8j8X66pZizd3TbBuCHlWtI7DrqSuqLwLWVf4LGP7v9I65ZQAoKBvsXyFckT1T/8r/KtZrrTiy1VC
1B1VNpzA3fM2V6Wo7p/T9psPvfTjXIWkpOjIgCZEOQXIjoaAPZWnd90EcDDxGaBoS1lPOtO3nH8u
dOx2qAvhB4v5rWNzr8P1vImbAHn07t74OdfsdofCVhfXVuvtZMpvh9v4ciLDbMuH2ktfg6p/5e6o
2eGbpoYc/vmBmBcDQEU5VuBMHN4wsNEbtcxxlgR2Bqls6DpSzGi1gZb/9PIEDG9mXfkWa8O6Nyk7
7Rcu2Bh0pvZZzCteb9Xx7fTDEpm5lsqfliEbhurLdxv99BYQsdT+Ij2qulVRI5sSrvdFTiyLnBvy
lhoW6VIhxqRgW3ZlBiyA+VsJTIJTC91MUPIRvgqp1n8To86X1OJnoNHjhPNn+7xfdds21kWXMOuI
L50upqPGpFeSOe/mOk57yFEKwn2ZQwwdHdgr2C3wwMBTnC/PM6t4pHVRsiGVq+qKWyuvysYyqgjs
5Sv+P5Fna+6JcuzaVNfxfQPIO1inEqtMFPjfbhf7j7Nnn1rkBSKDfDvsbweZJp9CKbcTooRdZ39C
32H0iRl5kY6iO1FHU2OG6d4k625s33B/AgMBsSCplSYPlvNQfjR6k3kR95jprFJ4nmmpez/rSxqX
3JU8zL7n0Ak/rncJ4QxC4zQ4ARkvL/joVoHuxjXJwhVw1sAifnpzU/L/vsBXHA2YSvHRVsdr52A0
QaY+6oCocs9xcCuprbx+zUqExGA7Im0u05Aq1imFVkg1BYopJ0fQpm1XHBM4ruPqGdZEK/nmPng4
Ln09JmUdJI6ZdRn/FC8HkmkkdOeD7WM16WnEuQC0ADbKoljDr7oZHan8jMuplthPrl06j+4p5OzR
rInnrZvYgeHf4GEh5d7KAuHlULkC12giqBylsJfIq7WcJmi8/hPtPO2XaP7wMvClJepzIUe/x31U
7oUn+Pf18681sw3iWr1Yx7vG1WTKTnMIwkAYg/9H0OPur6BedJ8TFWOX6KFYVAj0bEf2HxfLqenC
DSTe04DIuCr0+1vOBq2mpFxud4qCPSPpZlgtoHH0NzjoK3ZgqMcDB36G1vhg5V0A856ZJJ6e91eF
OoGujfUMQRxy1hM0H96NLg0ZWvoUU47VmxXPhgVY4a8bZCKcrvMgEmWKD50cwnCExPJfEkFF7Lfm
/m+8Q4giTP5be/7krXXKOunOBSYM611dOi/7dGBZqA2R+8Mjjvqi1kEXVxev7b+UhF0re7o98qDk
VgJuGpC17FcRiMWmgt+oZ6KyAAOXP/MGieqIK2CWjrbxFiIOWKbsBblhjHcTGX+n+6HDk0B0oSmp
ilX47pRj/ZAwv53xjoaCkDby0uV/t07sxv10MXwyDtT+tjCefZXT6W018p7nwFP4lvcu3qvh3uXW
vJ4dy9Hz5T3SYnQ6lECg6BO5casz7AvKdWaDNnQ6P2xR1FrquVl39FnRCfHcvNVN4Uyrg3SPKcvm
xzCJ2lIpdV9nfU8MfHy57jD7K9qFpxj/1c5wUNuNwTaJKS+CkSUYjDphNbHkPw48iF/GkD0PGN4e
6F+YGBp1/8WzObbQZJwgO449QWdYYE03ExxwVWRfI/PvmjJh1j2A2y3HXn3fkteUdJJeRUPzTHHX
jdtMhz1oylkshWD4+KrPKfTax3D3HEYewSHBH9axaaIfnhC93UIi+shVKOHZE3i7W27Thg5B1LK1
k6wbEIpaQmSwJNaoE81n6Q3RSagSCFSzT2NYZBkqKOORaPB9srY5hSYjeSjFflEL1eZdcxuj3aJu
xX6aRac4XB1E6eb8e9LwVC5Saiudsug0hYs5zaNM8cNJwy2m0hiOYharraUDb/y/BbD2WsiV5Exa
eQwDDfky/4tjR2xYpVaVBI/fT8Or3wHjXiZQatlCuWkuxLqb61aFlcE1sM5opZLg/DeX1mX/I60q
9U7d2tmWt4hx5vOoQwCeOMb0s9Vor0Roi/YXWiIH7zybCK5IlpOhiXVgbo3esz5JUFW7Drvtld4t
AhMPR2jYZvmR0GgAteyEQV01AK/X7tsIzftleoW72lNFPbLrh2347xnyNLRMKok36YpbdWgJ+8zs
lt89oqWBTDDKaZnglnhUC65Dzuw7lENTVO9BC/2jhzu+7ZKje4N4ECkVse8gJedKd/Gtue7Nd+RL
ZMWgdSTotpyGeo89vpF6WN36Gs5epe5gOVF04l33ZwjTFdUABYHnBuNHbM8PJCNu32rMZ+F+SDYe
22BzaajHm2Dfe2YgrkqjTyrOQcjhL0mZwwzOtGGX6b0R7F0zwTkyrH66bgU/H7PYXZQC0QgT36Ax
RATwS+M1FV7rbq83pcNPkr7ELz4oC8NbU2GTv5L1dgzFSGhFWi1pMln0LwQWoJAhqR6BNcWBuJji
/ELvPM5O2yedVgDcjOzlTK5Abl/fYDmiinJUDqgpUYvT7U7QUHPMxHw4a1FVh/YbbmuFWAdeqLIp
0IkIAcW4zTfHYeignXrdhlZoll6nN+6NFYWvW5Xo4M4AOTK1/t4lA+ZHwANenukmPRWJZMiG4T39
4xlzu5mmXOvfsB+uzU2jmgs6c1HVS1P5F5VadgN28Y8k5FN547qKsV5q2g01TaVEEeuXUdidUm7P
fLzf56e4SOjq/S2tQskMK98q6ZdZ/2r69p0tsEv2YVPR0odLWb5U1AzPXi6VUr8DL5sUGZXDRUaE
xs8Z06/PDrlDfgPqtYvdqYDR0m9Cr4rlWHgJbtTXXQjKnYgHA5nM21VDo+H4phqRzkR+NbMLHPKM
AjTjyQ/bGklzFAInFOeeFIKY/J81qocsUP75Tvixlx9sR/5wGfA0d1alTILWrxK3eSNlxwYuDS2X
p663MnEqFvmsGS0F8tBmuIFlGBl2r+EZ8OUP0oH03nbG3kdZ84jC0RNKKGVEaUXbGTdn7TaZ2FbL
I1ylucRW/DY/EIrBAdXNeyq0Ou79U4zRPYJoEMc9H9ol7k+chs+dVp3PyN1olwHnFWmtFRRzRUX6
PD4ym3X28Ke0IK/Nl7i+U+n47aXtmk7lq77yNffGRO3w5514dn1T/6JJW/l6d1ZoxBZ11nhPl6yP
wgTLor7/fRT7tvIs0kffk9Iyy2eyXO/GNNEJR70cCWwgqtxKyanW363AIJ2hJxs0BFR8oA7dMwu+
S+rEoVpEtWWKulNd5eWHWe/SVIKNGAhD3fTyHAmIDd4TWPA/dlJJ11z+muI0fO1gXPpC4uyRw+QV
W7ZVXq1IOFfo/qLNer35v7oaeVuYYkmKqMwY7Cl7ejq+luvaVqWO1cJCgtkaIQnl7fi8kcAEep4+
V73IP4nqi8EsGC/1XpDLRSMeRI0iD+hQkT/5FtTIh2hC/0fU/HkBsC+x8qRgbzCJy7Odp9kwRNo6
efgB+rGrWjdyEqOGmOXiDB0rXWIah3x8YNYumlpmg6qHtGSQrMII8wMy0PUR5DPh4R6GBHdAtovr
A3NJfWseWMqU8qgClkRGb6rcQ4RMR3p0jMvn2BWSjfmDEMKMHz9rrdNgZWqbcE/3bGp6FwG5yXCT
Qh6Kn0A5+s5+QOBoyhPxU8FRhXxiM5yeD1ywpgP8nfbxei8Ru3rgnlzZPCG4p5R81jHZYHfJ0ly2
Lk56o9OBR+2YjTsrhTHe8PoVKLWLxEseBZqR21d0zY5MMcJwYM1Dp9KmzeN9C34KPtGOUb0DBRo6
t3syaDDHsMpWKtGDq61IWr2YPP/syAq8zBn2gqxqxNGDlE06Zi2o+X6R341KreIOV2nCbqEnmDA9
40ZpI4tP5AcoQVQjW6gdbQXVNmQ8RqRB52t63ndafibRIbuvubzgegVFbiY0XARX0DmRLzEDg0SD
+QCYbU9Pyk9HiQ2wbmeJ4BRFA6cis8QPeQpgGjnAwIabdsHyR4/xQWKduB1iqI59Tgmq1u/QFW1t
8s4Ar6+kuRA69HAua6k6eBbXiz2X104r84RZMoEbHcXnX9oMtgTKXpE1vP6np204bJdDH1k6Af8s
aHzB4XqWGQEV3bN1K436zRhYXIg8itRhJEX4HGJzzWz7Q0pY1i8NyQ2oFm8GmswjMCmqKCP+HVhR
xnAyL/Ix5j4MCGwNZ1Hzl6KFGV5F7mElCcwKGc+Ze7jrs3Bsw359xiIAObWU7yiRKhC32atHvJmK
ac+neiGf7aRlSows6pN9g1M5KP3NCMqrEn4Gw5EnhWdAhGCJqfvE2tr/3W6bpPSY7zZqBkP6sHij
Y9s/Rn6Ps4zFUADuZmLkIjrRRykbVwJ3j9HNo3mJBQm9y9XiSWUQGvYZSXoWE6oHJT5lk+FQF5M5
fVJoCyo4ZBVXlvL54NTWMBLniYPqqxeF5lyzBgTbMDflNcj5PUcrnyci75/I0OpKBAUXu8hAu9fI
xbRgOhk8u0BK2r8U5rjpmQR2tXcUgxkllEN9mwFejbyplIGAm9rdH+N5IzHd+ECoLxWGWVhySvPj
ysHCxjRPh9EfHbrb/mnSmuBIJeTySqT9NjW7bHQTUwH5DxJ34JWEa0aAlCW7OJSoTtOkgVnDrsf/
BdF6Crm02eHeR0MU19OdwRDvUZM/oWnWxrqh7zA19mOxIVGTxiNDe5yziU4ktGiB8d7MdbUafp4G
/QT4SG5VX70CHEuKoqYMwBfdBktC2xNgeEHjIZS9AU+aPZFQ7ocp8CZayULLZ83HUfo1YjqqlKrj
OPLsrnlJskZuEat8HL6iFm7jpPhLhnz6vS7nYBlylWFB290tVTFy5jnSuCaF2rqPjCGhIG4gkpdQ
qgaQCbtgP2AfFTJ9/QPuyp6L1tLRa0rZVklIANjFgKX+N5dP1HMSx6YMc/08lwQ6v6nYffBv/lIl
B1vyWbHmBg5hrvwDwvP4tJaL5DSoVbQVUwMEWXgQrBBnQd3Z+hcdbTT2+uaAL+j0aE2U2HXIGasQ
EHibEs7mNbIg90lH9huAXNtSuZgjwO7ZyLtOh4pX3hCzgUck79+lOnuHEHkG1cKF7WDKW9Z16PX1
oAhks5ACbmaohRuyjQ0KQwhLHEupDsfxKap7+ZdJVajaU9fQqvf46vz1bQQgxrJcwajjPpR2e4wW
rGVYMh/0p2tq5tlA3OOd53NwJ2ovARqPzbEBonl2Edm+xVFHj+hGgK/0Xeh0ji93Dj2wXiJ9bfUx
6OKIaEXHiw7AWHel9wFPN0PsW1vPt9GFkt2oRGtix65BcyaBYj/0FqyBp24iDI60s5Pm5zmBPnu5
5tyPn9PZIbP1xRfpx41+aVamt5gB/k4oBkT/d2oZo5MZwOA3Yd3rFkIdzHYV0uRUrGu9IGJBQ4uW
oVlYtzrsOKu7GqpRuE6qiHS/ozXGgiVtvPy9ZfocZIzmgxb/qWvTn5unv+WSM75EzgUm7HM72KHQ
LAphtfZpFAhMIK0zleSwfiSyTNSDM9NldfpMHjiBQxen5kWpRQdQmfDBMXFWPt5jebkLuzAxxCxu
mDqpKeAbjdbCSfkb4WdV/9S0HJ4E01GxwzYlWbHEn0KAKnJQLE2qbW0/BfeDdVx85VFf77w/sA86
Bk+UBDf7Mm1O2Gl7cx0BCCKbqlNoioXkIRk5idXe85q087Zz6SwRrrK3gPVIabCkpVTZWtdeNsvz
xVogeE24ayVzlP2484zK6HkSje9P/fJhrdDbLyLPh7ViRRFNWWCYEFtG1r3jyFkZdjZ+uPNI+Om1
/Lx9dSjXr8hk72u4NLmWcC8dXhwypjiMd73eS/bntcjY7Kxx9gR/XqZzjkkbepJ6x5HXyygBeUVC
E5qDtHQtKwL/fBFOxSSP9c+jzMTsggXU43uchs9m5OHDGIpWHHpZwiTuvXp/AAhlwukHjhvmvAiJ
+bZjeEqxnUJpKTCJrJHba+PzIERDo5HWM4PvssvWm4QJyY7vD25BD1C6bowwMZH3mM06inhq68Bm
M/CrbD+AFc0NYOhmNWyApkPracj6mpkpng5PoXNXD5EQFOrD3pE0GHNKPQoAVIUiB/DQGq4wpNnP
fhl2XVaXM5ymvfin48ljToT69WBHO+duMadUgf51CXewDlRaTua3G0DblYe//84+kBdpmhl/ZeoC
dTgNorTkyoOigRpoK2h4xRQRipGqepoDQwltXBJr6jFZ1npWO9RfNFGFdzbT5xvXanf9XuKxuaBQ
M7+ieKBYiLGeql5fHXZ1P2EY2Z8MntsE24Y/nmcoil5PZi2dDQW4txcF9oFzlxxe82vFMhGvYf9T
v6KOKkYyCaGxy8xuPnzgvlgxnDlGZA9ZSMiH2OVozg9QRukdyKzNOAoOQr33infsNknqydZTMa83
YdXzqgJAOJDcgkR3OW3e+q2Ek9mR6gcQc/1cuOTqwEMN9tMRKQ6Al0Jtoy4BEqsrwboc6vtp/+VN
OIN7ikrY20JZLGAdfZyuavo15fK/1TpluQ63BXmmqvXvKk+CXD70qVXkjecHLsLbKlR2AYifISOQ
StWD3yfcqouXWtw7ciU4FZFNie0ZZAuuznxmGjxrUIlu00TK5NCJaG+jA6KZGsZy8W3Uge4OQdDQ
+paLZ2htYriwyX1Ryut1A3UWSTNiUiF3ymE2PfdS4xszApztpjIQchetWejl1hPNIQSM0327HXAX
8m5IJnnVSAqovgojMk/mEMB3kPl8d63gRalx9LHxz8MZpe3JNWPpJbwZ+6drBjSBlTstFwLgFwFt
ec2KDv3yC+UR/2MvCiXFcdxkuysvbgsBwotCqwLzl7W86WeEv2CVt6Zl8iu20yYEZBvCphS4ydTY
/1ygFlzvdEIcVcChVBWefEhi94N2ekbsD3BCgMzZ/H5I0ZFcaUF+swa1iYo1O0Ev1fXNO+fqpkmW
2+VJilhXPoeMsbZeOfNWAVP5qlKRBpwLKdcuc8ygnLttse6hoeqWtfZDvO+PpNObJIm/glwHa618
1gUuc1qPyN29zOq6VoF7kesI+G7lLrqFre84/yiiWXGxR35ql+P1gspC1S4stuwKmFCoklN+VXng
SLVaRNJ2jnc/FtYP3LRUUpujtbwHIKX8MDE0TDHTKgW7EL3PCOsYiSKZo0fGt8QC9yoTQf8HCk1C
bysS/Iyl9cGtk7IX6L+dtZ6Ihwam//ClwgSSTS+3wiy6E62vRo933u6XAQeqgrLd7Dsu4Ne3JPRf
oHAcWV7eNXymIu5BAbY7uWmoHp5dJLVFiZeHAZHBLenJXWLMZ8lUYRk6JD8X9iq+vxgx8fKWs8Kj
jR3Dnw1K9xMkdZrUrMKsQVd2SnMjTKNT95SalBTmv4u7cS4xLJpHYUjeD6QAXpalytERwFawO29u
aE0r2K/sj5Hjv4kCXrYAjg5sjIY5th4lPTLcByHym9fbr4xrEM/aWXZYMnWcnBFQ22jpnZBQL531
MTOWHRJMojC1Z1Jd5bKtu3EewGq2ubAJql1yP+FIPU1qG/D1TrYoay+hZG2NC7J6rpNW44in1f+U
vy63vy3KL09l1S7X1HsszCaqTSINBafSfTKYumNQsgTKpk2Nj1xSAMPA0jWUSmQdEH4mD2Sk4/E7
YhEl/2rIvsGXteKrNnjTA+P+7G6BmG9js9Vlsx/TQYizq8N56jENFC3nHJ2QzCfvdVWYJk/HTJuO
hx9TafethXnV1ADfzubkLnPk3cnXrrMglMYAPXgqw8vTIhToqCeEpgF5nlTp/Vty5qSTEJR0Qa05
r7t4ZE81X9OfEmwAlBpRBQHOUnE9I6jgVykwYBHkqeFvWKxEYoR5EbmIE5jQNshsC1gNHuiIqV/H
XMZxDnwjS7JhifwL/le6sF49WIyX11TU6RLQGZadbVm2Cky4A7hKyN3vRH2UhVstOUmWkOa8E9xJ
OOam7niU8r/2KPC/gV4J1bNfFdvniT+eOZtsR5XeRNJILNWbxOcJhmNOpGGTcGJsQuKGxJRvKZon
G702CjAMu9USpcpjQC02uj9QthAq3XErlKGV2ubEbsJGOcF87tHevNRBlOHW+zWVMwLTK2CHZZhU
nwHh+1S8ECZD5Ue/KyQp+VUEw+bcwZECqPcG9lZ1Adgue3DwsezFw72uvMjLzDfC+ak2Hs478ZUu
zaP7GXT42SttNFas+R8QU3K9LeRjHHUQzrC8z85EiEAwj6Yxvg99krWxM2AqUzHk1Bs1P85MLPEc
8J/vacBIDmRITAhWq2yLXrQIDlyjAXf72LnB7XK2dKHmu9B1gAzJlmX2l4XYBUdbW9b0nVe/bDNc
6hnzaxBZ9segSIBZ7yfeGG5ouEU7pzDeAGhQRfqKsuV1/SVjgtHidBy8tVVI0870E4PA7nZgUr3q
qsJy6B5JwobJMKKuMPrpYgCniyff0TTfow0M5c0726noEv06kF3i/49zh2Aj+wNIl+OafoOCcL24
53Aaq2hLqHIinI25EqyiR9aGogekZFbDiDgLTvjZOheK4nt6oVvoKjpSyvwHsxhn2+gh5QxE66XX
ehDuo+ik5K1RNdfI1TzoWZ9wSINCUPpI6ogt8Rgk8FzUtL5CzGsIYqHnK04YjI+21EOHL6rORWwf
Ajf3KPoh+jMkD9gZQxBOMawBBcw8mVc0gAr5OwX0xcfMYIZKW2Uw/Fy1cSP9sKR9cOsRwy5Xj2DH
kxXoJ7NIr/mlXruiTwX6zl/zkuSmw/Q0fXL2F9EP3BBeGIcy1jVXU+u/BYuVtCe99Xp6BykrAKLm
YEs/fLJFqFiUFXwuR63nR4Y/PkFHYNqK12kYZnmfMn4cF1UI+m8k4l4AMWkIKEBo521GZ5CFDGVj
zNvD2bk706tRXwy2/j7K7Shnh8+IuAqx7uPezR6z68Yj0NtOFuXt2NSGFUX0PfUo7bQqFl6dpLKD
S2gPP6k7oRgwHd7TI2r7gkyp0Lzt5y2LR43tUATIxEuUgDbBuH4nncuxjM0/dkWhXZRzqEMclYYP
xrU1o9Y6HTfv10noaGrW+9WSaw4Sg1xCiXu5cq0h68l4kNtt2bpgXDe+bFgg93Y11zdR1vrawG0a
OByjPdxGSprqRakTtziKeQXzcZTrO1Z67LyqmuC0LX94Ft2vP1ZclSZfKwbgNF5TNlK1f8Go8+g1
8XfoD59gECzYmrA+EaMWGVTEZsVfLRvQiV7FbC5yo2iFd8iS6ipmjCCjIprEFY2teon5z2SomCFa
JIbRsbxZ+Jj7aPivCZ4yMCf/OLeT8Utv+WUYuDq2BZwiK7mglUrdQKZ3wQKrKubQJK1TXjP9O433
Eenl7I6Vw8UX2lcJFPBHvZaC06fgQq5xGrKaS08tbWAJZ7SqeuhDXJcJLJZ34PvxAVljSdoaqNhC
iV910y4uwjNyYEIPtJcQs3HWk87KvkUnpeUBj/iaaWfFjDvuaQSR8H+eCfb4T5C6d9RpXxEjiLET
nZ14R4f83LKIsH1Jbsr70bkrpO4Q3KccHX/4nTsdceEXTPtz/2IPM/23jhbpQRtv4IfeSs6/pp/J
FCavml8czSOL8ctAVo38n3dMGCpPnXl7XVAuzvgkE+p7v/bmwVbjuWkwsTm/OetdHET68HAyJItN
YfgNxKe33ENGtOw2DtQ/Gb9can6XTqU2EAr/e91PB3lm/Zv94IPbtW5RIYkfVtK5VmRpYIi37iBF
VAGQ0byeTVtb7JoLYDbg8IZznU/NLIag6rnl4V4X/iU3sl10PITFAJ7zQLKyaAMK96Nq64Td9b6t
yiML+bXSLbNkW1zZrdn1OlFbnfheU6vaW/s8usjpXtHqZ1oRWX57YeYX+jcKhLI4We0EAgufNZrq
Hq4Lb4VMeOk7ShvM+HFSdrY7Q8+09Z6JEkXPXjC/qcgo7mL866IbcXFE+wLK/IvfQnpmboZwKhgA
1x9/nXNN9HFhvGV5yeV1BLbaIKKDZCIbnyGS/5boBXI2/wtk8WQTGs03sC/scnPDOjq0AvRy+9v3
zUeYljPHF2KK3byPzuaSQNwY66tugVL4ZIwFoXxG+x6GWM6aeN9WygIhWpWfBBshVYRIrHSgZs6n
cyDuPOd7wblUij+1erAk4tsL79B6J0RkBjpty2LgGnkE5wPz+tcrw3SA5NKCE3N0ehxGnMVMQggz
ohMM10+hwtn9FcwIhacx98k9bVlWiBJrjS20GFG4GvQBkQYSALrFTrYdTaEfuMo6mvgW8YLRgZGa
6eL3gkaGKHxQEVj8YIqdXeVEIemX7dezU++F/2Lp8PsiTsigz4eFQxj4qIDqTWTQSj5bf4otSfZe
A6qkKZpO4o5Hnnv9GNsIKLbcHltPqPoiTLwpHMikV2MjvAmtzqlS8Yx+uM7pAaurUhOdmU7/gPVk
j/j52F7+pb/PBpgDvvq9fGF8sSNlhl9bbHsSMuiVjvJMJ4vMX8gkRFQOKqv5eoUfG5F8snBM+Ha4
1oGwaPJ2j1bcjJjsh9iY3NK1dRaReRppcrEflml67bG8dDecGVjLh2TNZbyzU3PxGrTWW9eUR2H3
UXu64W/un5lJnrSCfn5d2eKWJNH5VuXmAENBTUzw/Y5hn44ySwQTEHvuFf0crqZJGR8yyC0t/tmn
HXA67fuHC/MFnRtD9IdWHuT3oeHOx0muW29a4tqvxGtveTtdWgYOYnUGg3DBDmlzHVapenYc3igy
jadL/gm6QYccGhudMiy1IwKIHgIeS+2EWqGAMZ32dGaCW4cQm5441xdHahnWQx+z/boeLlkDaDvF
xcGqU7Vx7plMG6gFhLJeefKWTy2K619fx3GrTEDX6zDpj/vyghfCY9YBHIMhK+59oTje6YIOUbnQ
CJgp8T1CutDttnjLaEiJA9o7du6FV8kw8arnuSZ29pw6p6EyUIriLGCIt8gwyAvc3FBBXK9K6KgD
5nMIK639zcZoz2/gs3Mwe5Grfq3BNjS6ZW40Wu9oImQ9z2sGXcQSRUmavXtzho2dSU8N5LH5U9K5
gkaL/vmx/tBA4yzS7mUhh+8srfi5xi+87HqeOnpW49y1pTwUXSF6RdrPYXyPJr8QK9Jbcq9ZEzte
BJ1jEaYkWm7m4edJKWuKVjPZmXCttOaj8knqU20pzfL+rgOHwu5meMEte5jqkszZmza4zjmeVFcf
o9VRcl3eQpKxJTck/hy3h/NeaUMiBy3UhqF/T1uCi8rdWSXAPHvfTnrPTjsW6ehPlqQ3kqEuBXnY
CfDbBSRwUwjT6y1tjCRMsxu/SMqyUG+GRaZwhWiGN7MI+stpF2m3wN4yppAtKqm8phUVIYYXFm10
zVc2H63VP+nNmGFNsdTuhlAvHaeXuls8IzZOSWZbH2D5MXS8w17LCxLCtYr32bjpNf+fW6xJ/80o
Bk+4hiUVo3hHETPOzWw3qFSqRkNEYmsL0b8D730Wh/FwImss2P+fn4Yd5oQr0MwzPXttocPXCba5
Rfnt1iPQfUnmgxOlzapkM5i/+5hkvm1NU7LPOgEmoGMiaWsS/OVpyeXcFX0ZXJpBFVaSJ2zkNiP8
TFpNWA8znKLxSwuwMMzROVegyv8EybnrXP5vEUWF4pnx1wjCji3pTey6AEToF4pNYS/iSAttnXcj
6VFK3CaQCVhjcg4fPL0lwVHdMtzMYUeTm+71fY0hcQzh93Q/mekBbSbXrT8nXzStWnuO0xfGqZgT
C2WjKydCulhGYvJjN5mOqmSDXgECjtw9LTObtaz87b94jyCv1vKdV+kqHiRs0oNeI8j3xLfxQ1do
6wXk5ef4i5r+qK9CuTXiy/shsrB3aNSY4sk4K3BfZ/Gm51Zzn9+ek6abInvkWH5/4ZPvbrWR3adK
bPsJpuXnk6JWSZTGBePdRSYm4Sn2c1RMWp3LGy2LREqhYakgLXAfkkUoAgiD6oLqQA5xwNro2Ny9
sNecOrE2xA2Z4cWAkQYPgFDKoeYxV6hq7szIXR7kz0/oBdNxcbgUX53Ie1vMmxomyb5CEJ7ZQjjr
0YyE6zLP+DMiDQRBCvTCsE/lUf6itAkFXDCqSJWUiijfHFCe8Up+y9GmeOFbK2qIXmyc2jLK9Y49
CogTzTTHe44ODrvUcBMfYSihwCBsxiUPZYckA9srXXTP3j5Dis/fl7C4RD+0dPm17jyj8cvvLtJ1
rXB4i00LBGhmCNBeeQuAmufEGWiqABeYYGDNF8fNqC7rp5uhXwwaxBAWFvnF9XlLAQvnaSud8hTD
REPBNwb3ejMeZ0FXfi9noIB0022gNjtltoAqWTv5J2T6nXaD3U1v+fzrh1xxipKzJg0Vi1RWdaPe
naHohxpS2JIMVoPsl/bSPOwjKpDk++vuuNdhS0r2wgHLrLcOqzpfsKR8DXkiEujw9t/ItOlWtkAZ
DFQerfAZ7ug9JRABGBIj1ycOWhmtxJHD9NVXgQhKmzj+a94CsY3SbtHwDRQw2hUDe9XVkAZudqac
typ82TsRwljDokqF2yHGIkr+HjDWSbatmQJ0dGUUJ32B3wfP1ZCfaMSf060y1gUKeCYkEl2zfcvC
Q/Zx1NgobmTKjWsdnq+04Zqqh+sLpySaVlEMv+sVIQZ3LnsFftlipQ0DBTMk9+KVIUpOnypeUUi6
zt2MeGBGGoVIcGk/2ToqanI7kDB8mEsi9ly0s7ba35Yai70tK/yiCVUYtmHy/2NJfbGjcNGgF5EM
RIMXPYhocSGApstZktUnwET8Y3ZOpZw0zMciI63J+n5gTPPdLuh1T19gaUKQQsMzQetKyU3iBQzA
/lbSBDhA/H/cEIvoxMduy9aFNhxqZ2FzNps0XDYYjOGd0BtB5g21/MQoPH+zKHL2cJtpdZdrbRyf
hQhfuDvSwUQ5LQbGiBdC8yJbZvVxs+LCtB3Z2VG628/ibJ5q8eDXmWxKWJKi51DhCnSbWD/Sr0KI
VngLIuK+j1j+Xscbcx9jaAQ6r8kmdxYFa8NDCtZBUbHkPJMhHtuCWb6H7lzShQzATYTp9sCiBHRz
FEHYJi7wjKqV+2pRimIqz/uTBcXdqUqJ5xikvjFgn7naSevs2oXhF+CzpHi1rqWlSmD7aGaGhpry
IyetmUAePETXBtE7ohp1Qr6aMT6RsWqJbFtbNNxliLsiGBTGx9JJFXnBLJ88pvG7pKS4NUZrul81
Quqq21IAI0PDD2d3BZjUqKSLRLberNibq3/m0e/1ftPtARXiJ+jHjtofOa4npbxve6R//JTA72W5
Umytj2rx8Bi9lY72nZLIKgD16dtlFIRNl2Sw1vOXQoAqEEnces7oIal5ZzR8AMtbZx5QGp1CYUm6
J/sXBHP4TIkdz7sPlp2WTtD0An0BwQRo0B/NYaM2r+p8PeZh4r+zN58xGye2rcnHTLMcQqH+twIi
n15mkQ+Xm6wcMooSIJHxQgU1j5uXhHhh7Xt4CkuoZ0YZGuldjhXSP9kFmZlpyxIwWpGgJDOo7GsS
c7ZAxDtcSjzdQg4QgmdAH2ks1s0h9nz/DnP4w3nZmYDUdSmA2k8GSALdVIpHYV1718erDXRySwpG
A7ifVH9VKVExvx5dT5dihCVV4FDkr+lZ+MZOcwYURXySbxk0Wmn8B1W4GDMM1Qtth2IdQNVaQGe2
epSStkHuCpYaluC2MD17u7kmEcjFkxEB8n/5xxVXd8FcXO7GVF+j2nP81ZGXbvYn/OkDGiJcz/oR
sjXidYSHHwVWIz8Z7AHYqLrCrE/i90Ds7TlFMFILFttx2L3zjEWZQuRTOeYMdq3QVMyE4AvknhXv
hkLR5lnnYPXIMBKwZvwCxUBoT5yvrFzUcITxnK3+Ci/GhTEv3hh1GbsFZfuwSBu+b39DsGNc4DGM
crJiqfz2chkhsWnCp76jwp0JKB0oB6glZ9obsJMPs1Yta1YiUq0Bd9nrdVO9gWURS0hm1DG0cJBE
/omjqaKSCSR88Uz+jFDW2RufMNJSAMQc9+Krbuhkv3KZPkvrjEvT6BdFHkanQ6obRHRAZpuAM6tT
rS7kDGrCLvHHn9Kp+AJg+sXXhC6yYsY080Jmy3tnBAXyIc1qqMprlfchGEe7tG/JBF9o+Zzrajac
3tVHjBMpQIFYXpaLtKfQAC47fl/xP5tHncG5Z0mgHOUYefGLnr9fId726oGJqD0XfbuJFOACnVfk
iFHYtqfmXwh7624ceKWG1Kvqjw/bhUeEgLGT0zDFd8/7NRIw0jg27j8TDN05278iGa3lgMW1HjSN
2QGm8Zie5IPYO8qLoeCESCZpN5NbL0EDAMrZLK2DX9iPVMNiqhp8fIHt5yJU66KeHkYZmV0axD6H
7RDubIDiKkjSwJBr+zUAnnnWI1zkvGB8HhY8mBBj93hJ+eFISdHKceyUaGpN11/MUMvzB3T30wVd
qDJzImYXBXfZ0jUcq2HRUmzfOAcqCXFpI/u5gFM0CXi3SXJb6P5RnPbqwxUEETT8ZAi9GX/YeRWz
1MzD9t31DNlCr3XBXJpY0X8bJyoyAh8Vg08LaIGhKI0xKQx25GXVTQ5Y/Wu//GwiMmr5S8XiEGdO
wmtvQ87QAIjreAC3RY8U04qd0V4sNnTZHOSBaf6ZzYxqOAFGTHE/5q9BLceMC5bV5WFGHgvj5m0O
GpXIOexZrvYxCr5bPKzJS5KLK0tOj4KMtqMPgkMafYfEgmCq0aNTJJyCvwdaJSHAfKSMNJOsj7y4
OgNOArBQUs71izPDAAP8KatqFSAU626TmSUCoZPlN4+JvJcY7TTeFdX7s5T9zpKupt4640CvHuEJ
KCTMNX4h3yqZvkgYP+tjJ1cbO+Fhusa7XrXww9wUtl5dfAdnqqpl+x8QX3/81WV0FnTA4uA5aoiF
UeoTgqU/lvmj3EzcE8YCB5xzkqlefwgaCOXfYBvzjxO0ioeVr5o59T7u9F4f1O+cj6c8NNz3T7+w
Z204OfPJyJLALvbTLxtaj4kLjavPefRz0mXRL7gHhckiAhU0GlqhTAhxIbZmOupzrlg1BQbOoybl
Z1lJCt7DQMDpti/Vm/Yn29r/26x7g4Ea+/k4brI5Nde//Olh129COVFX6FqW7vZ9wsbrMuHexBeU
yEdZsv/n5gIMddyFoTq2Rvi7jENvo8PkzXOruBBn9ki/uiRH4hd2q+wl/yt7euvkuBmI1QA/GoKR
2QnqoPus35tIiJLjqym2Sp+5E9aHAqPxXbmcMyxbHRBTiCGUtb/CE+hBAl5aP8vSXw2S03wpyU0P
8CdKxLAd5POtQajwESW5jrY04q6ce0yzFKf1J2VaFOpqESexRlvh2fBEcKW6MwojLckIsl6Bj9OY
Rbaounp/mF1a/I5TEMOOQziQWgsTnc7/vr+5fi6cCMHYxaTQsCHnFbwGR+Up8VnyWzqTsxa+TqsG
beU0dgw5OD0pCIcRxKFJxKM0KmY3vsszrZitTNpver0jcPTFeY5ky+w5h3LR8vierhlduGix8tJN
CqiKrvi2tj86IhkwK1WfNJl5bruqWCmIRF/hHOmdRbOplACCv/vQdfH061z/o3sTVs1TT0NT53P7
rJM1vHz65WJ2+dxkjT5vQ6DtP752aDKZTiDSQu4qZq9UBXryuX23mBozBTThN9hqAmHqcxlU2kQJ
BLO3AMP2+KJ3aGiuKA/PeySz5BRLrULp6KLhPy8R3+jCdPem9woFpDERNDPbJRoR9/koXU73+/vc
VrWUlddAmju/k75wdTLkrCcaMgk/lLPl4kqQl/15skfXlVdMK2k3o9rpuy2Z8n+M0gLz9V++gLmk
6RznWhpeEKQGSN8qa32bSdSM76y0C8Nf5zkmAiTbhscrmgo3jWZAKteCULlJTe30LNAWwPnRvHkH
e7xMEFqDvmsiEQe/k7zkWE1BWfYgzN+JqXKbf/AfdtfZBqIMd6euMLwih30Me3/rBiPKIxmw2oiF
QD9AXXqQ6EfGp1B6PKwS2PQG2quLtlpdK8vXD4WZLAlrauFSJuJJ4q7Vg6r03xno1WPb2eB/x6CR
CNBLYguFaQVav+KFfRkWIKAzIGpA3ukjzW7BWHPBc+4cG8zMAPuxbkAZoO4MVB6X6MKLZhnZ7hH5
SgHtosnX6MDtFGbH5bpdAfXuWqoLw1BKv/k5C+AMfEDI/32fVzvacpTsV5AZOSU9sr7Lc0vPNmos
ssrZinyFJyeeXWsmus6MFAZMBDnC6ovC2RgRTF5BKQu4VpREbjtrPyefqd+azHamaEENbDGYFQag
KpL/OzoRfCKKX77raHhzjE4BFPoaLDgT/3yUYRiPsDedg2uvEADQ3EC+v31sMz1yX/Waa8uSdh8/
pYKF81dAsDbG6YmcrvhaPkSPem60aZu+PNADxcbcwon8iSoNvJTRPekg9xlafjoXZ4YIo9Vn2SDs
OEIJHZ3OuwUMZ0KQf8kO678ZcOMh+OQZYVyOuowRmcJYaMuDjUurxahxJdXyYKEjdxoC3HbxnNFE
OphHZ4v6Kb8onI6+/YlENhMX2sr++yYZ6nSB0uC/A6Jp+JC+FtnBWqoZWEzP7Ze2l2mQ4+sdM9zA
/fduZJ7kG908HBZpMRgW2nIWTYfJDpHO5fMq+hQPR6RWntOAFMFAx6+uI1h82NF7gbWzEF1cPi7Z
yKqOTuA04gQ+pBMNG15rM3OITM9O77joP8NZZb0dyxfE9zY29a8BvScuROygagc6wiwX/Y/9mz5V
pz+PtyLXLmZurWiFH9kevfersjx4q+gew87azHVdPFqPvapiWrwdsdVgbzGTSj1sMSFfZgCPSIwp
4mPGMUkGSLFZVIcoz2f88dff3tkiC/qISahPvxLnhI9z1ZI6Wta06hPoBelcUK9wwWXT6kuTfIFt
n7wdIXYc0241sKw2ZfcpMFPUvUgVfd+sLXi4XUaY6dfaSDOqLxlRqGsqOtan5iAVRQ9INyoVSHbC
Sw0ebsXHh3Dl4aVCt40qoIq/CGn2lpdtHh1v/SHPwmkaNbG8bEI6X5ti0RVnhqkk8GBbXI7/BCnd
HnmIYTpEc/T88uPPHpwyoeSB/jzDSzrgkm708Y6fIq5wpUAboYtk9DU9H54vDDnv7qsZMEn1k8z0
LmGN8Q1GKKvQvBljLX3YSthrDe9wut/LEM3fCHI2HAFVoQoAfjXRfb89LzMlXO1DHnVji7xkKuC/
bG0hgglUwfY5BCO/D5Sd30g9V1XokLN56IlKmfzUZA8kohZpJskhapPsYjHYFUIa/woYlmf/hHbR
SSdwTLBuvypkkIEIubpQuIF5pPy4d88Oqh29wnuxWl9jFGdGCcA+IBPXcPjBhm+PApOMcGx0IAk9
PgaZOa33ZJsGD22eO7OOOrWYMHToQir7ellZR1IjV0CymKoskWn1Ewa/TpYhJdnrcT/tM8MO7uav
qIXfaBVVrb7e2I4X1rtHPPCa1MSgEwtdgZCbvMLcMlP8n4Zz6jELStscc/O4g5PdKO0CJ7HGmMrt
r9mhQ6XV4iJ5pZT+jWeJhE9fHfWDTL+Pxg5FXUTRUiODhDvFhX16KhEDxcsi2rTnB/eHtASZYAOl
SsKZFxCnUjc2AmUCpDz0grVTNR2rmlcDsmFL4V6bDD7M5VmKfG7nl3iIQvvyeHqQOBmRHbXlOXKT
+oVsAgziU2rDEytL2xcPdFRVVopvPugLW06PE273zCR3L2UzchHZjFHn1A5KzzKFsneXTgusmjHj
mBqfumjaK0W98KSVDNHhhz+K83qfHA5TE7MFAdkEU76urujW6EqTOCacKr7QG3l+zRMMZRxn+6+V
MSKsDLvF1oQ5lXZMHhCV++fZw/h6Reya0Sbu1Px17VjIsziPWrINEQaPXWMg3YC2bqJF+FYtJB4R
Vhh9WQMmdkkh+Dlhtx4utfxpcchvV//jnK5GquUzUBbrU+Qw4CoTh/UnllOq0957hRPNdsgEMKhU
odFPTlZem1sjJNvUcGzddqr6/XYuuwGldfmZYxLy8BCy85cfo4EnkWUI5wRpajumttOZA0eQwJzG
gScCHYubKWcPBTjoanrSc1t6vJtKZJWwdsSXGpNas4+sYbn17ZY8MX6RWwZS3CUU6PejL99b6uOe
n0XVYJ85CwGy3tmXpPPG9z8fUtLJy5W2xx2lyszxMCtoiVLeYA/P4FJPmOp2Fqic8A33oP3JV7LI
Kj+2wNH2pzE6gAROaWdgZPpZTAUHwFdL+/sT2j8TTMZt1Uf/uIr+itLFZyb4QlrcKqL4AEd75xgu
2bx2Vor9xgjkcN1uU2AjYmst1c4L8BCcMpLFc6ZOm6Dvn2wTHyu3lGbEqThahWdymM21+mz99HsH
yy+c83bwKhuf3ekVVBoPijEkifkCFYhEA+MoEh4XTAPZkfsj/BHQShpfrdYfiD8yBkBF5jby0tW3
g+lqj6EY6vjDV9SzeWexpJkJ5NM0EJH1/hr5Q020knsAARbfgRG/tLbwBc8PWXfH/QQT0yLJvZw+
z9BYW3/cNVTRXBuNwBI6ubisndS123FQhMzRW8fK08jzTCudna/uHvJyNGLtSqS5dIKe9CeAg0vL
0OqEBXZ55QwdPncLaMem5MYIgm386ksFwPhzDn8yH7hix+QepE2krmAh92Ws3ZDp67/d9TYfPpDP
aehmd8mOa1AfUiH8CMKEaLluoeqUUMBtW9myBTISrWyxf7bFGteppTpoKR1LU4TuXGqOhq/JiH25
9P5BUhKjaP3PLvTy7XDSBpgiw67svkOITP6qksQMenphCvkd2y5fqdzwNoy3TPjkb3a7laOPg1mk
CN0HoyH/sBFD/QI27haXX/J3DYr1PHBNTi2z4MZwMJzz2zEwEs4uS0h87u7qmaDbBCaxJSC+gx+K
G75cJAUjM31csI7mzQ7tZca/AOXZIMbH9V74fXYtz5umjU7z81s3y4PSiYqwtiO3jP7m3EZIIPLs
gsyUQThIfniSPyDMiyKLF60BUHmhv7FvKeu8HRaxdeguYXvAIpg8W+L+mFg1u3nqDOEpWIfK6ISj
yF6lzgTo0sxaBnCu7IlsCtjkEdtw++UH185Ag6ib0NElAXEwcs74Md3fpDDwRkT+CyJuVTuynbDV
NNgZy2MVcjrDYsKdyedfTvNo2u4atFPyUnP+7YsX0aKm+Jwo1hzvjH0XNq3Q9gkMfj1+DIVMeWbG
7qpoByEcrtQpl6yHY9VFcXYofeRTgjxnng/LNwQ9v70IRRjwAf3f6eW648LKWTjUTQCL8dhojPvu
eZ8ap7l0yASvCUm/Q8xqY7SklBnIl0IeD61whSCQc039V+8dDsbe/zmR1xF44gD6Nxt9QV7SPRai
eY9U0e+qPSmYJ+/cDy/o+PbAv2CJh2lruYVYBPkkURrSi/X9iwY3Ttw1X+lRC0+xGdimy6+bZN6f
YjAS8hL3dVHFZG2uCwXee212LAmhiubCtcGoh0/ycJjI0p/6n8BmK0nL2cBYYdI0vP9woJ2ab+S4
8j3XRyvkq1IODIBhp0YGcYQUdI3FhuWi1LN7GAP+5v0Wcu3eF6CbAvtKOlN80zEK06ocCftLeKbA
iSZnG+qz/CRXBwrk1KHgXx6tDfXl/Hb/uqnyuccp9o9qpFimT+r/OYQCs5J4XUafKlMTohAgINMv
Jq6lG1ttYPK49Q2ecg74HOB+SInjrebvEbk+yX//XAbNVH3YASCtcQR14Od8m7voy0ITcAjLM9Lu
K/wLirxAbb4N4RJKxtSGlU4KAyUT6MNCN6UIgKh034LxlhDuoLRrsFAkkNXb0aXugHSha9LyauyO
++J/ok8+G6lZZ84hBTW826dPc5vBBepYb5UUpGo+KOgayAGVPdNhe3UCmC/KQBuD26CVLf3rRmsJ
fHuQ4ut209/j4dDuf/AzDt4uoxhr9W9OVTG2btrXsm9iTiJQY+tnsRukpRiZmGCKv2n/a+zbf3Jb
dDQcuV+4YSfpO93LGeOUrYl8n0KdB1j4dYIX2kxyNbemGuRdLj0DuJ3EAP4QTzB7cUC3cN0/x0RA
ErNEFFB6yZXAnhPagbwGCXYKYB6HfP2QTdZZ1gIYExiYfVbbz8lqrVjijGF1WEtAeWxco6xs0Lxk
rZ5R8M+LZvtojnvrpzGgCC+i9aF1mSCyAIFOOgAV5pgrdlGLkRMTFtSNFO7WxgE/Axqpr/eSxQkM
5z+zO8BxMw7q1Ppaw+0Zu1Nc2cxR7X/4zkqD0MT0UyEw32V6a83KuvMbe5QPREoZEFXPq2uxcmiW
/b7yu2pu5Fv734AYU7MBc1axUi6Zyklq9KG+9CQDJoaENBjxtVzTWPw8XrSgAUlbghP2lncZ4KxV
FKGiNqmX1T+7xJtezj+XpnhlWHe+2FvV1mCB4O2xF/pTXmyNOoGQB0kIF5oMDWKKn76UQWxTV+HG
BVyMAWkPgb+VTg8WzwSY3faLm+QRqzGUwUd+3DXi25zomih5LkTNoEjmhcCiGWFXPlcGXURQ0NcL
q0DR70zHrTGNuzbxJLF+q4dW+fyuAcVLpK3ik6h+99EvDv5EcW6OXjsTN1Xn25bzJ/VCD847bYgB
m2pxUjGcwBbMD/roZuNLZZCd4vwof/fhmntq3kOBBVwMEuqbCc52dC4RkMZp+R1BZv96KCSBzT9U
TAGqZ1ZIxJyJVNL2fESCG8y5SfWcyTyKsFky+pL2t8dH9cXsbDB25g9IDaxw45qMAnrtnKE5K7qL
7ndEjs8DIlNvTSGA2PZkwA0BQjrBSQmDZMpOVyVd8LMNFC8HMqSQ0m4OVdsd/65JsHcTWZFbmByL
jnpJoDK0o5+AC/W7B4HjdJQrxGVXyX3HkcdWCOeW973dSiWkWdjsFF63R9hyAqVCD/uSzrYfKtBn
+L9P7EW7+PSP5jOWiH17ZBkYWWcL/ibNaVcmug4dL+zx89zY8rxYXYtjq1GMojeahIlJe4uQxFue
l3WHgASdOLR+EJRJPEqMTh28za7SQJv+OUM4F0UFlOJWX0Tzk1JDE8cHo5VryLagCjwKsVRKIWoi
dNFPX5t40LQ2VDgvu8Wu0+TXfGxz7Tubm+ML49RGV+u8JHjMrQ3RkpvPCD7EoJ1S500guZAq3Tyq
BPyFXPfccNV83wx7ZVSCFy4AZRacKD4iJauxigJHhHPe7j3S8j3uBHSF52ofwqGMb2g6tuo+lGxN
HdcnxgQvXnIQxntAClaRV/aGzKfxrOA93NmPBiPNsruC6PIIupasd5OZ94B84FjBheqQce1I4CSN
6wyt04tJzCfHcMkNyeVqhXGnccccUMuv0Z2WG1LEkCwJApyrka2VhqhCABmQnly6pTn+SyzJxyK1
C7VBsFXvIWvOeFtYh8pZFiKpmh4OUOTgwaCAX6sg/4v35J6hinQTMAHooWDYK/WhCHS0UCGfls1A
d03JjYDI12kIAxN00Qer/7f7PEeH/MeHkx0lYSThacEUFoz8fYueeG9c4PMDAZVvjQiv1fhCkS1e
7pUdtNYfvBALoJnDf794CGSWSkqaIBq1M7hcco7TOKlVE8wMRjt355UIWiqztBJQfLN8k8zz4/q2
f0QYAAdM7qXwzUdKDYTbDZ4jIfPdzN7eHL7sfv3UqEWYHuG9Z7PpGswp46JPBwhMI5vuIVIq9NN0
5CoF345Ke4vOWrvCm4Hl3/zLZnD5zMe9sQqNJf04RFIcKyfnTS+984P4P6+P2OqaX7TFZ6qVUgeB
qdOWy2s2IsK5OXLH7LzDva0gycS5pyE4SVmMQahjsxFc8kLPLOfUcozrgzcEDb8OgrDgL8goKAcK
SjpB6B3x3JcbLq22Oy/PsTf7kBM9xyupjh9i9YhIkb9UG6jIDGXNYk9CRA2vpyKFI78/35QWZKpV
U6JoQS2PegflvB0uoFgpR7oN53vVkTwwQBfs2HINFh6Z8SlZZMXDXj2vR160emPbaLIuZ1b+Dh/O
w1RJNF3Ki+ixwDv0Ii0Om8U1rY51TFUDBs+O1V9B6yqa4tFH1F06sQ7idjv+yuUXxdmVhd3QNAKC
gkKjNqvQIe4uygYxBqT+tBBKr/LOcSvJ4MSmTQFGuAGN1dDQyEr5s1wt4MANNILsz0SCsCnCvQGS
Ca/vv4SPul1kkgDGEVOjsYNYMK+ckJM9TOTVltE8rQniu5bFFiGYblhU3FVfKRdTdvkYo0Svl02B
DZXqKbJeDxV1PoHD/6XwCYd3ZqZyHoFSG++OFADiThgQj7mKrWiBSf+Sv+oE7J+XVdJ/OWico1uj
XWSs2Z38JagOdBAZ/qsWEmIJIot52NS8E3eDQsLCjFlj6kLKOAFbjOghsu2tE62ipv7aFRwH1T+T
FW9lFpwNQmADMZiN2+l83Uxu6pg3oNK/TNfyfMxyABMaED115EfWuDRHAUjtAT1kYZ4ADHAVRUpR
9IzAC2L8c95mlAmtM0/7pVcCQPXInBpi9mCtdAuy2FsvqdoFkomYrqmyIxtk65InBLvotBwjdZ7C
HCbK4QcMWA19FR9Skdc41m03sdfYqcDnChDQI4TyTe5/uZMF1cuIJWR3wCbfyOCGOjzQZr3xdeUx
GwU1pqvJAnUwucV3UPQqIwNAYgDU/ZITAVhnymtbN3XTNJfkW8cN5eXn+BChzwoR2drK+hDP8bjD
0o32VOGjNDs6XxYAt/39R5l5h2giPLPY0FrY8amIxEmgOYVnT+BwgE1+qWUipfUVQvxzreWKFc3q
ZNmkCPaiQNx8O4Yhv8eNPFhFWWDMdVgopSuKWbr8eNUJlpDlWgg3iJ56E3o0m/PJil9eeSTZnx+S
jgrKp7kI0Dg6POd6B4ZMtAhxqiKT5uqsC8wGTzMhD+/LhHMD76RLOUfjDfS7zTQ7Uq35R+FpgphT
+NyeUX/+EdmhvYz49lkr1+mzRYLMnpcvefcPF8jXmn4ChYqR2DA6W/QJ7xWhWEv3FItqKLZjl6WK
35ML8zKQqfywh3qhldQ33tB9gLt/dDPFnpR7kAs8F5YeCVj2RRkMHcr0FgnyM8Jz/TNwxpp0OGFp
Prxp+4qUmmGev3qCsKju4PkE5frZokrMjLypBiIMaZNOgKXBb+ErgxvIgKzVlWXzSBn8xhNG7WhC
u1K08q247a+Dpd1NjQj7C85uAIM26GoY4X/qiElD/a1itoJhUp/mGoS0yYAfBsaUBZ2I0V6/OBbk
kQwzfoewTMme/NXcN5Adk0pWMLSoq7ntNcGctSL1CElLcz+x9Z6gEPQoJcPWYGsJDW9asRixLDgh
v6Xka9zo7Gj9+1SUpjZl+2iI1Z+WuHC+RsXNU9vSvz96QUOC0c+YPrbzu+g63r5cttigbwO7vvEU
GvQxfBjUmRvDeFK3qY0Hoscey1a47My/CaP589Y1aWRviW7peHBQl+jSbyh+NxAJE41o7bgURpfT
i5tt+K4Zjcf9got404kWH/sNZSPO8xpozN4AHwbNWqkfAf8u6kP0jDTbCI+8XAqkLvs1tattn4eI
GNL1YIIOWT9OjCrOiffj2vLRyZoqBH8fahFeWyAYHiqMyWgi3M03DN6TsfqE7j7HX5qNrtGgfsSE
xHDJeGlE00kce9I6ul9z79HKIQ4lD4/xgbONp13xgWcOfk/aEqWQ+TcLdiTtIgO5poZUz03yrwX+
91tMzi4XkFKf4S9TopTN2bCXZoibhBKhXTQtenmDF+izUPAXTUY5TcIOmtWODOMHEcCbHa5eaq7N
Qc0iYfLU6crl5fDkB/QS/UeChTg6iyrqBll9XwrcrgbTqp9IqAxp/Y8EO4BYb8UkHUzAP2zrDOCD
BxT0wRGx3/GciiA3xo61y3o2xmsnxsG1K9HzefbbaTE/omDE3lKGvZYxukABLY4LPg10mVtokeIz
3nngGPaoL4BdRUf/D2IGPMYQVIoxpzzDORETIM31z+TAgURUZ62NnJMOYqLbhWq08smxN5IxuMYE
ahv/E+6t6wMgSbcsVL/Ib2NZlwK3x2ritR9VjNar036DHJ/ULODRjC6el527/NeZBkv05Z3Cx3fV
yyredNISABj1Rul3To8Qcbuyw7VeRLE93ArCnR80aIxdLRJ5U1O+m28HOgJ2yXpmwz49rpqLQ63l
8IGB5j5RP2hgA3zvq8buBnOOfuaW1xQZBIEG38iIrIylNP6lJ5yqiBlzy4Wie31hqiwXGbOYJDE5
gcmeVIhBOvKWd63Sv7Lr6B8aRXl381zwhdyHHStn/Qchuj+AvmfUCpYg4E606XWQCxqPvUSx0pwx
ocu6caWiUCIHJCX8gMZLchGPJem/58YmLEgnetmVGTFaTobyTUFim3mhZV/aG8/xtAtkig+wFUGT
KlwSuzFAI3vRZ0iQXhO3F9bTrsk/qdpCGBfy38gi9Na7dHVvUsbNPpwC1AqPyeDPqMn75VLxEIb2
271x/gP0UsJzFfia7CHWvRhLzmtvJOhLpJyYE5COcKcEkdjK+KiZ/3zdOpuM90VKwB5782t7vQlH
C2KSw56ynZ3NIEOte97tiDW9bSVzkkXLKmMZptKexXef8/ftR5n8YJqq9eZuD5SaC43pB7QRxSF6
ywCGQlbU6iWgBgeMqepJXPF4QjwGIysMShnblk9IpyzUhj+tC4njDqsrzHx+hVxia1uTF6NC46mY
+ineMsR1CsyZJpbTW1kyYNPJ0Yy8mhOK1Iv3alhyd8GzczclVvd8JZUM7UgecOiEHhv3QuoT6dyk
/SQ7aD/SL2AXgYq1ZdOVIH3uN/o5vc2/KW1zZHNT4WXB8KB0FcpaSzGUlGKDQqdCz0kyZXEYIDQk
gwzGRvweFtVpqDOrEU7M8uFzHw65B2Fbor0EW/6p2agCEhIz9jnbiiXHHOLD2GseaHiOYagKBG3y
siD/ihKqAHTebeYIlZC3ONmyPz6SuwbYUaxnk52jZjfKDvMwMr2nr7b5nN9ZkeKcy1xbi9MLN4aq
37oq2TthXLq7ZoUE9A+BtBwEcAU+i5UR0GWjWEF2tfDvZFPc7L6iJLVpNF1DG9/bWkq4Ss31CDMy
lESwyUGTC2OB+28oFaD5fychRPrVxUJOr9y+0wYvay6gGJKCd8vFu2vkZxorijAjTy9YEnaq39k6
bsMjnsNCp+r9ygV+BsnJJ2kU1Jkj3amNbg0guhjxmaOXgkYcPlIvuH/Az3JMd1ZtaxJJNJPFe21l
vJ+176k809gm7/ySQgPV8ND2iBY8NscOP4TDe8NnPo4QBu/BkT/BZiNo/MT9mlZz5uC2gzDa0mtU
zoYOj6sVwgDOCXdZziqoREvCUsEHY85Jqzp/sWIvCck9Y8+m/4sXAX1Kq2+rpbJBdSrSCIsNqIn8
3mqSpiJRWXJeULSEvGW/0kqJLn4nGQm43vJBFukeu8CyRH2BQgSWmrFttjkuhpCFJPESCTLv93Mi
oJvLULxR6tmq2ho528uRIN6R1TyMNH9iwATG1WoSPgzne86MQm5TRbASbgoiwQvPyFcTnQA+3W4H
n4TgeeePRqA2zOJRdHXmn6evt61Foa/OCgb9WdIhfajMzAdJxJjv73Ts2ECqBiEHHhiJ+RFbaEEu
7vODVbNt4raaSCRtO2opYC+l8U25sDvb9PJHrVhiFDPjrZX5l7Kll3cXEEKQ3JuUWphjlOnRaFP8
ORUIKB/uW+1PSDfi4IESa0H0mAeeWOftsnjFJCHjOX6Tc7ipRC9oeMJ4bNIHmeAl7fH4Pr5cYMJ+
jN2RoVSrG4a7wZoD0clGRbUybRWqLq/jT3vefBgROkgHInj3uhZw06yoivi6kMJf+QrjXAeOdO58
EXp9JML9B/Hy4E93lIkQh4PRIkrqm/LMo8NMb6/Bgvxjn11P5wi/V3sgIiy5GBJd6tvBmAI2j6ZI
SN/sk1M75dr8j2Xh8aMrFITPeLS6uKGup9MyWZvWmMfLVrFvS5rhd8aSUy5aFIyyyfPpX4ZiT7Sn
WMnEtFDdH/2mVNYR9tnFjkotQ9ext0FHbEP5CQJ09VpSsOHYq7G1MywV8dXjRVo+PtZnBfRiCn6y
vGPm43zw+RniHEAHAmAV1EjAAHa4XdJb3aP7Okz0hK1KfUH4VZm4Rr/E5DyPQH/mkWfseX2a2UnI
LcAJVIwmlVs80BQt5vgz7sQs95d2X7l63eSKi5Fw8YZ9LKc6uPmcRGlPho5LarEI/3uxnp5omUxB
z/XAfIiyiMGAOYgHu9+8JWxBhfJfzspZh77nMIqUEkxpf2c65wi9KS1SIUk7VjSKe0XX7hAFQqTT
CPZOdJVcOV9RVnT6K6z5Zk+FTTpBQ2nQoLOayK+6UBZvZ4SFIgmXD6EolwGraJx5ZaLyKy4q8FO4
X9lS1N/hJEkM5nutJ9kxizep7CS/TU8CLumnFpWc47SQe3216UIiVcAdEDAX+/QfuBlQHd/+Sqk6
3SjRlhUqhLVOwudz3suUfuaYRE0CFCqdkSTz3rnW+zi8+6VB2Vj2bAu1vhVsJiRHoHklUT42TYJl
AdUuuLW23J0P4He5Y+dVEP4Us1r3D/n66BJWnqMxnK4tMRs/lBNcRKc9ybz6uWC23LR+3A/vcp5j
6Vp8ofohJmXmzIDo3Vb/Ev3mqybRD8FHM4uOfi3sK0H1CHkctJDSag9ztaAB2YxIWAwM0lbDcdat
7GedSseuOn2tqRBODftE9WmS72OnmNC1tjuvc0Oc5251V1vWWfcivS08lM7nTjsx9oBjjrXpOZSz
KUUhf9hf6LaKGFu8xaUhAd3qMrhB2l151qEerLnYusYs37IdnLyZLGP86G2pOXtyMTJnRiIu0kCb
eKOIfnBqEfylcHJDzfbLfHzNMFckUkKOMX8a8uNRJtOhSARoU4ln3Ixg38Zr5hAVzLRWkAfCqKqG
CzqPElhz3I8aLBCAZ+JQ8iYMqdFzxDDq4apU8ffbSbcANzqzBTOy/N+J4juvxdLK1DzqW3PXK1eC
dKY6pvTRlAflVbns4GRXthkOv56B8RhRTwebtYqV0wJBRH6fA6ccC+tk1QK86/eq7Vc73Db7ubHr
z5qXZrc0VEM/g10yQfr6naX2xk4/REn1TJEYr9IkwpkFixrzXh/Zl/liaQo7QHug+NoSQIwmmzGW
wLiEggUlgXCRImjNOGbFy6/f3eW5waQ6EmPJBbLTkHumM4aff6X3hzV8Rqw6m9er5y17dFDooI/M
POP2PSuNhlX269lgmVClINGs2+85UCdHfMJbN7gmPNQEVahEclGgdlRgrwOeiRRSE7jQKmgrbBVo
csUs0EOAkARnyShB7eOAeDnhm5yasU0xwb4fvc4u0+wZF8uWhwI5nOHTf1VSH7KcrfFWKV2NzdWc
+LAzZ1X48gVGyNNM5uZHN21iFXUjmrCrbEhsKGCHJxvWQ5R/NSRSDc4zdbaAyklt5ofYRg9+PyhK
9JfNmGjMlADtL3z1aWaQzedgny8YtsOYf5NllgqmGT4LM08aTCYB2GVKv4dXZk8aHmHjljRrboOn
mPOfXPwyYBYjeIJbBkvE8VSZEv/IIQP9PviuCZNJM2wgYPiNj5z0HX1xOYsarCklZ5MB7eGz1Jph
Ijuu5YAhIB397uwpTYDBhJchms02T89fdU9yQSQ/D6PVTpIUNQvd0y8aLfiUXvoReSJxXKSmCB62
xcxMMXrey8pIYrYRymID4fLG6eX5GrgAp70iCVoaSqex4qOEIPAJDCzRi+69qHAgkOSyP6mNUrAr
GS1xBVJMNQCEzW7mo095q3ysS/Ho3Z0uUKaFJV+R4KrkgcNpfgDC9C22x+KWJ0oc9twxrvZGr+fP
UQZdit96oB+u5h21lT79HVRATUgXhaFZd98vkLR3WNoWKobkz899T5v+RmmMjJhd0HY6u5WcdMVe
paWdXJRC+H/vykW1wXzCmy1h5yqatB1nSX6dSL4/DXSTU0dH8L2H/ol6ZApEricH0KzztmAs24kS
MOsj0NjmMx4bWzZuMnWEFqcyRGEq/nICFTgGk5h5HpMSeE3d1PB9WFU41Zbuz4Xc+WQTRNvt6dMe
wl/1x0KEzwSxsqzADzNC8aY/ED8jjTaTLMjQdm5q4Jw5k4qCRgnsp9mMhE9qYWoSTjo2fZb2JK8z
KcURH4QIl5JRgPHfK+rZ+vGVar5aTbTX8cjyDwo4AjcHcUWY5r4UkfKYfHq5aolWc4YVTAyymuKV
SEtmb7f+ND9JgbLhWbUbGFskUam8q55HuL2SIGwQZtiFmHC+/sT6XtpSAo1i9QVbfbvnI0v6LGHI
O4H0fro0GUJLZ3o6f2sCJMGlcGgPdq3k7PTLAYcSG8pZfIKtlEIi76rlP6qSTNibVDasrMbUY64n
E44IIEHq+1f3w8jn6MbJmqpmBzsMKm2Yjqq5dTyKQ8a+gpzs//pn0XNrmVPORQGXoV0a8u7QW+3F
88VDe6d2LYF69HA/AMqLeEqWzSZEmlH+O8Q2qjdI1qkQU+4WNeEAx5bx+WzgmopnWaPGk6chgj8J
lmROmSfNsrV2mrRFLhcxjEDpjJnRqLtYQmjkPorTkE4Kyv22A7bjThC1R8LiDfNaHt8h6ao2Pjf2
Qe5/0hu+dU43z0UW0tfPufNlk1mYWHwXmZCWuPlj3J2eaXSX36/khQAwvfMbzdPPTI1J+Qdhurqp
uf9ayQ6JhLAnhuMB9L538bh2bfjTCBNc0rUrfK+xpxfxDitmp9N9ZUgtrd5+kPcdQeR6MciWelq6
+4z+8dlDBXI0j102mOkcYR6YCzuFys/ljjOPFuItl9AEXBo7Jh2Xe5RQRIGpaFpsxdepZNmCSls6
zFIzwtAAA3uQpGaOZo6JSCpGCuwv2uofOZCHry//4OTw5KQL4EAzKxwOuNNJFwiYM4VAEGsNg0qB
aqqCux976OniMSpKo5Tib0i1gYYJWGtggwMUb/7/NXELcprRjislmeKuYhl2TqD6EH/mHZdQX2I+
bIU8Ga27DkNW/0/xbkWpcT4D0h2VcxJ+v0o+1F0toHEjsC9meMD1xfz4JhIxRZTwsaJLrw10AtlW
UJri3wg4CPJglNjSciqVpzA5eXLQ6WHUEDO9IcgXBwY/mbQeQEsQHmy264aLIacAYvZWFfW1ZX8m
eS6Kcg3JE3FC/sO05XGRIJFXldhQD+zPSdNwiOqYyih/aiudgbVmYngexplt8uSMd4KkZgQNdP5e
+1kcuBOl+gIuUfDp+c1oqcmBxbzCo+EtNL21mUhh7MKuOXWycAs36uBL1AOllbndezbxGAOFodcg
FmbFZBJGOeN2/moTU6W2pJZIMEVs2VUNF2hrhLCF0Qag9w8M4vlqDEGypzYVNOHE46QCXh6Q0jCv
Euru1EkNlnUFrOoI5pdtPfOAuvnYbBLnVIRKCORUfr5zO5PftvoAHi7eZSO0hAzrga+uiPA6SAyV
kRnDo28H9sAvyndZHHuY5PoL2VKgo3XV3mL0O9oaiubiO74hGjzFd5B8Ga0HSVc0C+/6rpIwNFhH
dwj6eMDyu9abQhdVmmd+iflZcr/vqZ1NvvpO3xGvJVA7L1XWLVNoJ7rZDT0jL14Z3bqIyrwP5sUm
O8OvWOr3Ds1XUP7R2pdZFQGoajcHjFYNkTrYZov7L5sBHZmhwZh3BL6PL6WFDt1EGJ2OU8yEZEM4
VQtUEf5SLbOE3uYt8v8PzHX9aUUx+Fv+gROtts8N3LZlvg+TDvjhbSfUhURLs7nEov+EQNgmPhKN
XR/pO/4o7ekeVzZ96EyIk2hk2BLhhJycXUU9MHy4vy0UnEnSXPrdtk2lzoxToL0ANvfKz02zCJkA
0inOh49tgxnJwD7ZzEQPJ9Sxfxpc3BMKn0EGVi28wWbb+ICOvskXqc1DTGJss2ey7kS9369+aqC6
oeuQtSj2+ReUam+1UG5FS8v1ZQWvRsWVQkwhmU+CDM8P3NJ4sMNimJ7D7XChpuxr2SxCGSD94xbp
0NU9FmARxCEKj0TVE1vmK6/SQihNIkOEUelEp+Q+l/NfLWQvZzfPmuwskLLrjyWOsA6M26i1cp1A
4r/Awf65/MPgut+AGb6vElXBbN/XgLYqXvv9ktOfV7B1aNqEGsFZd7Vk1Ko551EVbJnyJ9gFainm
6L78UcMhkgxUhOpyK65po87elTpt++QqxFuvHoHN/mOH6Y8T6tKVcuizRXTlTZZ54QNXSnjPengg
oVU/QhKzKrF4KFbvgVe/ByZ/caIkHkGhIURvdfzCSvQiREkFogiYMj3xqH3CuVKXxamyMYDRwn1u
IXcKVRo0hHD4rGbm3DG9FdM8yP+f43j2zYcGARRLqGZMMqvaszSeULltdcCMjzzxvP0BossWu578
a23akMCCheVJJ4pP0aO9Z5lS2GE2ctCeZgnOI3p8q779iyBEtG4ggxyQqQl56ZH3Q5REORF4b+J/
i5rxJeJhBayTaaddYrTAVUQ4iZnsg38bB3LwxCazBwVn9yfyj2H//szc3jTTTVMnRWletWAaWN0D
O3dv0EwrA2cs/qQXAJWtfwG4OFd/a9kTssh/jxe8ZWR0asmpQQUvHPytM0D87xMhoOiMxZk3sscH
6GH1t+/qVc4bO8d83e4no3PjOqTHykhAbGb7jY1AakU9ce6zlKNkl6oBbdOcKvqmION+i6VNpGS4
lFVnud4Ylyg+4ADNa6TeC4GK5OdK+yRQtEOXWaP+TnpEl60W9qj5fqBXcWWdMlaBLmHRQfjGaXmY
QmIQfzs/0DdwvmA6p+6RH05Axeeaviaftf/g9baXGVH6o63jVRkZGfWDC5uOjnqKavDAAB8Ujx0g
GHWJCYsGwgyosds/rfP+akk2NnxER2/hD554Ry5ozSsjT2ioS3+jVlO7CG8C16DBV25ehVHBksSk
P1+SRHYNz9SL5g4JpfYRQWxmEXy3p1LFmpBQ3heDt53loTXUt9hxK57cwU+aXluD/66cT7ICxqtg
2KclP2e+hHZSMWUIkX8SYW0yqWUsSpz/LSdB9qYs1E/3FmPL9So6PraRgCWgzkRQobhDkwJA+e9j
R5A49ZhHgWYRMH4mpDnEXqBiSgYrQUw7FsN2WkMrTnWDagn7LKTyiQKyUQMA6S6WHP7m5u2DSc+8
i282syj8bxTZZqZsvGELSYDH+c+s+OOp7dxZCUFEY0FIcZayLb3DdDdCVtMswtRi93vQg5WuH3YQ
8xoctgmKk+TXdfUOQwrM/rLrpOZKAhAeqgv8auHKoiMcYoTikCh3C9I2ALdpW4RKHNtTBGDv851N
p5tHgu9/frGKaqrTUMgaaHNIbEJMirpCXEInJNmrfgoePv1CHuta9KRJrs8T6sRPJQKfwTtPrOE9
yKX85CxIADlKeTEBV6sSITQGBWRxk5BtXcNVaM3g/4dGUcSqTFolqYiK51STih7cMb+hhL3iYd7B
mFHIevlanYIpW4JQYLpe0ziJ1pw0uP8bSNfuJXygPBwn5xkIN9bwNAfjcvTuCbWXPOokqOVrHq4J
+kjKqzYwLhQHmtgihT22BbwNdl67HQurtGqzbFOi9qEJ0HK40hlalFYvTXZwB5rkNnMFUCyP+wGu
wwoVTTenbL5gkM+FEYq/ntJGC4wcb1NutwEmn9Hc2I1Azd9SXfLPIcpVN0NTNyi7Qxewyq1/v+Ux
FRyXqasvRD/54IExK5ph9fqBF7C1/xapSoovNtCqYIiaeF9HWK/r5oncwSG/O3HZCmKYeSiOovb1
Vo77+8M6De6WYUe87YGLjXHjxAOqhxCymd74XLkGV49SPtM6Nhy7p8aWzhTbiZTAXhZFE30jaX4A
k180sVMveF9anTKJzDNNsrnTblNRU8W9A35NJsrVg41wxSJvOMVp2NUJL6DVmCc6E+QNmRP/bxzI
1SXer3EsdYcxjxC9jZhr1gioC/SawUZt6YoPV8xjMruvIY55BUAUQWmi2cC+FcbZhp8rfpqzosrV
No2ob9LhY1eUSesCRBIkOJjuBmFOM0VMpF6bbdHgX5B15zw6QdKpxQSfccuylEnSr077XgvFiVsa
vvxXedRePeps0ZTsQo0PYhaTcrTCGOGEetVHvWN0KFoOy7EJY/YrBOuBo5lTZ1oholQBFm8SGhVQ
FcJpc93xvAaDn2fpqzTp6813O6UVqC7Fv1Cb64bTgaxxPk9ql47QfeG4voN1Oc8SwAa5ZsDG1Tqb
kU07enNqhuMXWN1gt2K9YJva6t1JQFVlH3pZJKNo0R787uey8dBzQN6bZWnNOV/WzhiD2GQjNljr
dpvvZITv7kNbx25gGLQnUvsMsqIpHgUszab9ZGykhyFwCZbTW6krdPMkkS4qXKq47VsOrnBL/vm5
eOMm+qM2WaTDvofJgnLEcvOgTj4Tj0HdDPR+ANJScFhjDe/yPVI8hFB7mfvOGMdVzEwwph39KriO
eMwwtqhOBffAQwbUG/im3MIzBdpj2NGzZuies00RvLdeCROX77Rm0/a6sbzA4phNr17IOvb0T6SW
lgiCLoeB0T9r2Sa4BPWBjr6uKRzusBmXVI04lhX0DtTU3QDffQRfbxxxFyAoDpDoQh/N0A1xeoiK
fFtxfy4bSM4STrFiUl1W4mvRz6Cmu5d6eqBoFrIjZRJl8jkPD4Rrp0Oj8pqb6eG+/l8ZTnc31qCQ
kSO0Ik3mL62ycHLA8iu1L87GDW0fyJIlsgdBZu9RM0VZJmqzzofN1PnZl9r97gt3WSAfNlical/h
Zdfvpc3eeYl5O39L1HmRZmGPJSgjbjvwTNTnevWgqHk/V2Rn8FoCP0O2lzrhuyeoAdEYtsDmh6hE
wmKp3DIVsmjyxz4hlJy7wMrOuRT4TgoP4ta97C8eob+n/lXaQdlkcSednF7dKU66tmGRFnyzsGD+
AWRd9vK7bG8TZfwqAm75O1Lwcpd9Sneh2pyWACuNLbcoDHwcneoRWaOv62lq48oRHWkPKzPlpMg+
aDGuGXYVRdD2FYUnB3OLRDKz0fmAHwOLp/TV55pkdtgtg6eJO3IC26I+IUJsSfNC2wRXEzTVYdXr
Sv/9CNNQqsbjvtF/ejpd9baWd60uJHNNN3g4rNnu2tPirdLmhDX5/MIVM0coyz0d6fMCguiqLEbc
jMDVCV02zn6C2xzJNulYV7iCg2Ufl5yullWb/xpNBcBvPxTBReESvjHipbgcn1wKhf8+X9LxzF11
qXhA5QkVXqwbQ0NvbCuw7Dbh/WDoXYwOJKaBezSjOAEk+kEl8hr0EHVL06YoeTFin/MZjvywBHAw
k6hd1hQRsbx23h+lYbXQLGxnqnOTH9s3PsZw8Z+lBcgZyugzx8VVPUGUmnyRnjvFyo0IkV1r1lES
izyLDQckdrRpG/23ovoedfScfnTSDUkxS9O2SMmfJiQjqR8c0CFfkXz9o94BFkXpojQAjEcgaujg
9LdX+soYmIvIjrZSRjM7vGKvegehFDYATVa0azlwIqRTk2p24ddMZpw6c8siG97K/fcO+EFmD76X
hkUJrIzYAkyPGd6VHJDYkDZVL+haHRDNzLmA8Is2Xob39vSRfY253/USOV52z9/myIwk2VB8H6SR
gSYBSdko1rosTOikqfaK1ksEzb/+oxj+XBy2pbdpZHw2Pko67ggAHX6/OAXyGfbJ552Aax6vrWFU
Vk21xWMHysfCX0dj+uNJppGHxD2lSxCWgENlF/IB03AhoCjTcr2928OQH2Vx/8CNRtDbO0jQWxof
4rTwn7dwdgU3j9+bjpbj21oUCUH/Nfz2m0h6fiyCxPyqjhTKYUXYQUgs/6LbeB+VFgqVNQtPdU7A
PysdqQWX+ham3ED69ZgT4Col7gve/bAT1VUBztMf02Tgd57sO/ed5e1n/c3lAWLMPkVAVkeuIiEy
Y8PVS2capgnN38JJQaPNnDJkp39/rCbmqe4FEuIFzOIQR4F/xlAPoJDYnuwMc++xUdI3YNufJ2nG
/UdIiwCt5gtceNafQm8SbBzLfCM/UXd9+eN3kYBAcVdTialWqVHqzsNuboNEoFyWVGRNQulWttG1
VGKP9Sh4KdAgDPb0JqLWCirk836NbHXG7bMc0xZAznCyjAi2Ch8iknlZtvqHacQrKHSBmpAZBLvs
pkWmBxty40XRdxZimzjxn1V68NTlMh7Y3GLAZj6C6bdmCkEm6CDJGxELsUADYfQOdnWSjhPcWNnV
l2pJLhgEw7mK8YUaNymMIFYhn/GV529gpWiCszvvou8YS5v/Zr+16zjKtuXJs7kKDw0r0p/3yPqx
BT+dNjCX25UP16OsK4uJu8VW1vRvsSp15dL3E3shrVRH3i+sA1Kns9E1unOcxSZ5mX9COZ2jNVGs
kwcOYcCcAwqOly6WEuMZ9GU/xXnPyAMVYA+9fUGOc4pVaV8Bur43kgazRJp7uHLNovlAY2EH6JbL
r/Xb8lkqjZRKo3gXhpl29gkUl3WtbSX1Ya5eVv9FFNqHZYfr4ppPGS03NNNnvUj4m43I+W7D7Fl/
ccVEH2QkSSMS75v78Z/YuFVXhGLeHtm7V342TtA4ve6R8qLMru+uIA+xYvNkaDRCZd6YCRkO310y
BKNv/4MZb2PIVX+9mi5s2DSs7SN3vGCTjKIaq70OOGzcmLp1FJjTqoyZYkjcHQIP88ZSN/MCVAfR
oBz9TNbY8WJhWoycwcsXdSH1S4hXu3JVbiCrmghxBwklqa5jNIHFMmS3wrBj03nLCYUl5bWS3vQp
y7XdEq4qBSrvSv/Qm8PIHempec97zoHXGcn+CdnjiG24freei8gdwkzGqOxnWWU+4eIB6PijRfob
L1uYhJo1YvNPC7my9CNRaNbfuJMZir1p/40b4/LihLORMijbMtN4X/qsrlU01Wn6cmNJB2Zbfj1s
JpCVfidcEgfk3CL6VHP0sPcRJAdfjftYac7NpjNtE8rCf+xEuM2ERb3jIQKgMH6FoJhCIhZ1bkmz
HhdmPsU2dXUWHQeN8/86RcwPyIaJTpVgfuK2KhISemPmGtSUAbdW5evVxPwZBqjMylNwioeLL2pG
ChvGm/TrDiri2WYN6MoYi20/tVsSwdMGiggGiEY1mfJFCzPV1+dBv1CeUeAg99OdOekGFy8Ajn/N
dTcuJekSNofShJRf7Ww3BcsMjZep/elUmOcrSo4uSbSBQNN83XnI9bFScHggI/FWYognlTFBgbsS
Vx9pqhqpXS9sXjsVE7k6j6TyRzlN8c2eY2MRBgHqyF408bJ1lgm28PNEM6FndCvW31jb5x395SP/
bDJ1IclnQnRDRxcE/y6unGFihuYBGg4eCFUG4QgRDn2GLy8VGG4uxPOxTIkmXYXptrWu3ZGfq90Y
P4gse01HEqorqV448BGLSpGF7l9jeToLxq92jqhgwxrorcWOp9wLyih4JIU04Vl5sA0e7SkGKdhB
PZyBWqzw9VD0PRC9a9ughu0r5gLrStRj5ZVZOMe442G8FJIxgdBPZnUxnvJVfalk0EwNKTtaqM1A
Lhz/kvXaUk0q7ZN/+RVAO9PH4Xm8gXfs5L0ai7GvxZQ7iFzugQ0w/Bfh28K5IsczZx/mSE+ILYBp
9mLbW76fMXTRVBXo/BVbBte+EB4hlIcuBYs0Jpv0iuR6TcQ4sErK6dNL2L2pQN04qfxghKbqk+G1
B4kVmDRSsHzF9cxn0uuyNR0TRumSbpA3/LYQsKUtrOkL9MPS2J/EWTUFMx3vNZbcjXPOZfywTZW0
pLdtH7375OLeFkWMm+ZmLwoP7SHFdeopvu0QYEiQ6ei6qDFGtjThOBb+OgDLX5Gk/h6S907gXrnt
965Z585+ukkcJeA5nrGxWTT/lzMCyZ2pVMv8wNqzAkiJ3aumGuNrDxUi5U+PSwMBwEFky/8ZTybu
hI7//v7ntjbFjz2Aqu9Fx3MPM3CnICSt67RFZ1kSaXMrwbwq9kzfqPQUqSongG2CD653RHAcdpzx
kQJNw80MGNQ+7EyTlrag4GlF4cH5SSq8KiM0LNCP6L0kNXuAUY3Ljp8lqo7uRG0TcddG/ig8/u1g
/xpW1f+G2abGxXGYZ/Pz9pK2VcrTgWx1m4W7B+dIN5sDbKXtTcXdq725v9FNCP8fZkC7mMcylj65
mtkGtK9MSmiidpR5UAamms+sRkxNt6x4JeGYH6u1rsjqz7PAHSfoulgMNyXHxffU3vWmZnAM0E4A
FWCD8vp6fCWlcFFO1q+QxW02QGJlDXsU7WBqUhR4xWLD5Cf8B3WYxYY3h9/W/o9M4UK9KOTXodtX
+vWCWSG1NpiWI9+vbFzR5vdmWROXvUYFYP5BnTRU3IAiKwJ+kv7JzVAvCpd841YpRKmKrvjJEA+N
3mc/NwGKC0IIDVkzDC8koE2SQJ9ZAwtf0p18jlnyHZ5n98VhYqNsVFOLfKWDNoGYX6f48fTx/FRx
a6rXzisVczn+b+cdyH7XwubdizgGxOgDUsNeOJQ4Pa+igOPSspVDWCbha8KjLyf797BmuZ4OapZ1
0kyolL0B0alUMnKSa+EGRI+lRqUxquqoZx/LIdnG3Dx0ahwhdas5swww27gZP8cEG6wwVYN56QKH
/ZxypwanTj1L+LnvGnUKahm1PV4KpnZK+GS8kvQ4HjBWz0BoGD/ltZCjsI04H2G9wftY2cIjZ4Vt
MGwZ9v7QwgOTE5zqIFU3Wwv7u1hOZax9ZVkcPIc5T2BdYwy9e6XWDDV/PPS8O1VJYm9MbHxz7KkL
5eY9iQK9m7n+D3A8IPxgr23NKnTWM6yXgieZbpNh7QiKKp56i1zCo7mpqq4h+Q4FI5J/Ok2s0vkK
WfeCc7lagA9hysy90e8qyMtgWCvU7WBEiov1FiSzbPzU6hgDH4SgEpexrC/mvfoitkVqu2KGYTYP
DW8KRns8OiDvgyeppTOATXo03oBfJvCSFYDkJ9emZ5CfcAMhWsfERAGWdKbXVkeNUX7G4Z/4Tvus
4QnP4i75GzGNN1IyPCvYiJSpbl395nW1YEr68bDeoX4YRo9ICwjPTyy9TuDw/dtFhP7YL95cnWu9
Wg+snOxL68nW3KScYWQby3aR//1u0BUIZkGQV5FRj2xonT4kpwbd5OCrKTs6Q3KjFgTotmZLi0wq
S5MwTI+loCHe0UQ4hSucYGOlo77Zg1gNG1ryKMsJri9ImV8FIoY+xAoSsWztUlMVWL8s0p9SZhlv
HWXTJzW6vWCxFHC8gslvnuq7IKchEtbi4SEF5euKmcVaLL48XSNDWRTEgMgndEtvHbT/scJvSIA/
Yplmsjj2ImaClwbsjRdz6/OnIMprEfJLS2L1AjV83VRLyJ287Ia8pjAHyeO2nvSdVwVmj+03L4jj
N0DwfQVGYD1F9/Xq+pBxlc3BoLXfnny+COyM1RZWmpG/umIMNbrh34aACd3nc6MJsUQXo37GpZbt
Fzg8ySCvzM/75gGZ/qPeLyjrPOQrBSUYf7lcU4Z2b8pbiZ2TFbj/HHPvx00D+F8yDQjnPGnDC8r/
9d5gDtdVcgpSZLUqwsaDa3uP98GSQxpUAaCbEA9R8wwogy6IVbnulYQ7OSFUVdJGMzt2SyMhTQkK
oycneRkKxlttgAcFAYYSo1EeEEdXg+czxBAOHyHByQNZwf1HEpCiI5NQ+Jy919GWmEakqNm2gR9e
26hGR8l0hkW6zIC775Qw5IcSDQEnzaMmj4TItaVqwIXTLOWpVB+gN6F2/vWM/jnxGQeHaaT++3ny
jmDoZkZXrcRp69tW9nP+p1SAHusKDCUqOc0oRziLfmBquRJv8k+sWqTTumWwC6iQIYhpEu4KuKvd
Thmfb38wTBOFfj1WGPK+V4eyTWYY0GH6jJJgogKDRqg7R2QsXG1c3CpeqOk0HVFibBuNKRK+QVru
WJ4fAhi7Og9XYK6r5f4mvvzSaLr6mUEfYeG2wE/icM9Swj1VNzILgaD3cZ48LkwbWJEC/JQ0tDSD
S4En25iqNaIvZNIShY3G5MHYP6uKMn0rX0a/B5O4mH+nQBOh0+n4RvupXtqzIolffdAqoL9hGRKq
P+DGqjRNJiMkCgtLhNMWrZ7h8OcKic15r4uXtj6eLgFU9tCJJtHBv/Wt+h9NB69ZPI9Dokc6FmTl
yKIv6+xRuvCXsJPog534LNLLNHhqe47vIomXom8R7VgduWDWg3SEtzqGKUxPZpqciZRvnvbKEkOC
wC042gYKVCQzba6WpBLY73SUXTA4c5J373BR9HH+dwbJcW+e0p7KHwZc4ht2oMefwk8ewzVq1xas
IBySpGELRkCAfwJhX1UdU/dmyfi6n3izlEm5rNBWqvy6Cohk5Ca8nZqVnGJZPL5CwTSrDHR4OCbO
ELqlK9FOhQ19J84Y7UXadrNZVVEhmJ1pal+2FFyMF1UGfw5+LZI5keR2rG3ca0wSuMQhAZGUdCTY
+R8MWBTpOpbijMgaLRMctFmDJR3d6n76o+U+5DtWIBNhivoqtEEqaTjj7eLGkiCLW8qbm3DG27Fb
FBHePF6/1PnV2pgYDT2+rDjvi1RMsr6pxHnZHrp3nfaFro68Z31pcargAOW7meyw6zdEZQXoBZjZ
rgDcfwu/xmGtmjDFNK07ZIYZaAJahiM/1aRJtzY1/cwC8EaMBh+uRfjDSm0n8ujJuQwi130zz5d5
RpB29TuG7+f+JJVGgUCngWwwgYK8I2VnXWUWXDhGs1J9adsyXEuMc1sZtTZjVrPvNnS72X+lReBz
6NIgH7br2Mj3jXejiSZBbgB1uPKSs3yL5k3jvYTpUa18gecIWOcSVLkpKjehA1+ipWhbNbS3iNKR
cs/cdItmE/J4lBnSc4StQoKD2mYTR9TozDaLQcpzQ0kW3s1WwyyB/kFfThPk0QCH4f0ArpVC2pUA
jjN4BrNxSd0j1TO4/21S9lQG9Zj43NwhG6hacr3W/AXo6NzFAv6YZRqUJzjZo7O3IBftxLoEAiiv
LA3Kst+ixD59laPMFwTr5aozxWj8hTafZ9q0xSV0yYgRQ6N2mysKcExfx2fjaxGIkAXwIipkb6n4
hLcotH7lKBuBd8iEOSQ6++rS8Oh4VWi+jBCEiJ4LWlXZfbyq5pMgX7tvIXbrE9c+K2hq7D3b8nzg
68Kk0QHt8d/LAFlqZ7ShLZm+1PvhqlL99tVN+5kF+noNO5KYXx3Gdrzp/WOoti/ZtVUG42QEDPii
reRUkPpvBKx3m/Ek/UlqAYPB2gHp4Tn4TAMkx08d63Wl3+Yl5NlBKyy4Obhmx0Vvy2kdjFwWZLfH
qgIVBbu1DCV3iVbgeI1KpXX9qcJYLsVG7r7VN+r6uyLuMZtg6aeTbpwmaKworBInzL2hbr0w5uhH
AlnpSeyw1It/vM58+z/cmMSuysU/LU5GDu7ZdoC4uO2vyuVtUQsbI1nnMiGokqDdvmt4Vnu28BQS
WUfbzTqvmd/A6ovjUptSJ5AWRzqGYvYlJNCfdEGSe0AcXhdZRXJPN5kRpXBYMFICpNBl/jviA4Nf
/YKqUc7ELWemFz7XaL4RhoR/haerPGhe5aNTzk//pUCC6nDmZ2RMJKOBqHDTr0DDKolEFvFyA9xU
tPtzH2bum7glqWnP94YWhKhT3gwOACscqmvXUqQr4j328CMjCWYDBC8jtfRJcKhoLcTi3nIJOFtj
pJTO20aozfgoxXCdNhH3DOZ89P4h4rw0XPojZQ0LLrF3Q/b713KSXf/yytQ28gLtbV87zSvTUS/9
YvQ/kZoMqSBY5IERvZNQb6GDD+s/iLd6fCfmLrgCma8pfoQXaXiveJMdc3wlTdMIeZ4jRb2VwSKT
qYk3c5FHa+zalCSIc69L3Jf36bkUp4KvOG0h/oHVW34OTVpqUgkjIvbJ30JC4zgBOkCoIw/KAZwj
mXYY+YquwBoqt+8MpiCjweuMMukvuWh5x0DhYDfWEv1bqUKqNwDZ1/v30TX/6Lemqm+AZnAW1xwV
KKzkg8reSvKWA1ZtHX1yFIhPSNFPYqS/TDP8D+Ub9oYNvFjWEt97nAKSfdGDDLaHumC7b1JLbFnO
c+AYHy9OxhrF8TFCmkEOQj486W5Y7u4s10KGOP0g4zO0nmoQxjaMSdODvpzwsFGgt2Fqg/8YAa9m
z+4kycAED9wbJWDnGk2FxadmUzw+PwhhzpkzT2b1sNfSYYksxMjNZf8OByXwY2xcMRab5KRxPTr8
4zRUYUDv/0Pfmy7YrGqLmH0nfpBiTSdvH9oNG5SxVfqdTohGVi1WkM99jnJeqlPJzOAh+Mcg53QD
ybZC3aGPM/rHKNu9lmSENqos3/M/xjQTRy34pxdN0FoDqYJ0QSpJyEDX/O5yiFKSVCDBdcAXJmgg
r2lm4v6eXBVQJTlXyBFNJi7GXVKZ8ZEmAms7Ozuh05XjJR11Ea5X9adP7KaLBc1WSFYH8wl1kCqK
G54LMLbKKgGyA4vKnSd8jHFayFzwg0Q+tgWuyeKpE1ySiKkYPJn9Zl0JuL8XQVLh7xa/0a8EA/BO
QU3L5AQAL1u19L30NtjtDnoMsVH3o4H6OZcQFmF0pG2qGgVaqwUwrqXoKnKzLQLmTOzorQxpLuRG
GyLtmpeNcNduewLwi6Yto1jzUqMGs7FSh90NM0s638T2y/wqXnMgo/4wPEXnfREBRvflpSCQ/Mkh
d8JgRfTMahk+0sytmZwJAmFh3n5NEY1FxHhf8DE6BfCa9PLsFgSaf4lidhnFQjvmB6kfR8Rfgj3P
hJhBUVbIfTdOYcHHXOybKLZPgjgCVUm84Afm5YBVg2AX5avIQ3Fs3jTLmfLp8s1AUqwqdlRM5lo/
2C9L+heoi4MHcmnhRlHP8ZOET/7/EXuYRMrd33Hp3KvqCfra1Aozu+/ngF49vIABAb9riYUCISl/
jMO8u9Cr9yQWBMVQ113gjaqDAUwSH11qgiK69G8xw/VEOQ+IGzvkzOVQ4kGjDP/zc90C3OEpBAnr
5MSwxETJqrA1BxakL4/W23z2I+/fBQVzxc5cioWNM7B4QxyZDpLW6EnEiWX6PcOgoS4029fxz6GX
tQVqVBBEV6pHqI91VUcGR4CF1LQR6QNjzAftSk1ERUCImlsFQ4Du+Y0BjTFTb7OgfxR05fJq1tnd
th3GDgWwfQaDyKo33Nk4tbfBF4+fP614aDeKSajSG5xO3LjS4MlC4gkNSjyFyVwqzlc5KQxdN+jQ
Jh+9S1IoWZ9VoIPNQD/lGQjpSW3A6Mz3yRGwbMunASG4HimsA9uzd6OHOrZjcepeCYZj4DXfwQHs
hMF/X+g8ExCTM2D0XZuK0jpYvw4fcRkJFfkiLCLbg7hs/lGeTQn0RNiU+Hg0yanfUbPhmO7T8Hk2
RN/oQLEVBOy1GYCjiVD2wOjXyq4TPLsPTu8C73fKsLCyCFovUKB+LJhQuBJkjnNkpXRRt/LjkxyN
A5Zo3tA3Ex/kOF82sa7TcK88Le3sHuFJcJdZPrnBv5uTaYjIWTlCT/rozen4fbyaWaIcgGT0EFA5
e6ocW+ZcEf7eTbTzyuA46nP08O6UwXxT4VwQNDz7inwtFCUIA4hfsWgPv00lrZADRe7yIJhr0GVb
j8L2H27vcSNwql2/wZ8p8G4qAcN9csLA5DVrsHBSLbk8bFw9Pq33lNZbr+L9W070cv7h/zNYlwn2
K9OcGrFon7Zn8cajyh/wDPp2kDrjQ1sIRNxEiDvNEYhbYaZyoq6PoPQiNImvWfNUcpNW/55L7Kgf
AGyeZU5Y8V/DHtXlGHDpV4DZf1FbnNiee624lOQE2RrlghDJ5xPKAJgpNtk+4yYF6xgQ+hNaBMPN
JZoQTZWMrMckwqcjWxQbtalIszghDVtRf3pM5WxHSF5V8jb0+qDqRpuW7RxL0MtfK0YZaEWGDOMe
zj+pKYQBVreV2mVARPOvWE5xbZphGb79LGdSAJ8YQAWlg9XZOo6jDHBts0uUPHLSj6qWl6KptyNX
FNKhorDwhJhPRXI7V4SXWELAKmJfidKOflizft3GAnfo05Q5lEV+0DgJYukPohex1S/U50hHgK//
aqaPX+KBvmnr8cf8S6WZa3d6ke3XA01QTAOgzPzbyaUClKCAGm9WPRq3hq232w6jVyvk9LR1FZFT
aeJ2X1PIR78ZDR2XTR8IjJEZG4qBGPIHhqEYurMvZ2Dyev5DuBFuwFyiNNxkcLaNXrlLuLg38nEj
ikDfL/yNjDeQJB9X5yLMhPFExbtL7rnk2VXW5vVDBjR4ZxjNCNtKXfyqu9jdYqRUXc8Inw1J0WMy
cmzLfI6IcLSCm97R/VVjN0rBxnGNiwdZY8D2xdnDz91qjNBkpgExG4r32Qj/ucbkFJcYYI+DzXv3
/tIMAwU+arfp+biXneolkxta2vksYl+uT6Hi1CY18eS6dRQQCrrv6qVfuVoPfY5CwrUoGyEcKq1H
/JBKYzv/WpsANuvwV1a1Abp+RgPKW1heX5VxRNLdIlqAO04KIcC7zkOL5qXenePTU/tyGKrgT0+r
S8TK6PCMlDMq14g/WxfOuVSBPYD5kXQS+r7bHbjvtA0NQOTCvDyOvaVVhqwW5PxQ0M1ELAdaxCVm
LY37xr/QEs35Wo9wueWDlJkfoxWuLbD64yNPrDMs9TyXcw0wpDAEL4hNsu5SpGcYHnXUcPGcpaaB
sSYW2/0PfWvj9Z/mhROnLtvtXO1qrVIAf13BrsbhBw60Dub12ptkbp7k7LyVBzKSVyzDBAB/LrsI
P/8MeJfuimcpA231unJbHdwNul9AK6fBg91AIYJ4jlboKB7LjCnkdCJ8/BMvxIoqigIU2HvX9oP7
2CtSTcMB23qK+RgI3LkeuSkx9Zx/NeZulazUpdWCvev6E5XLrJX62ax9bZIkdmIliapYhjaaXumB
bJxerHojJbIeLSP/DRCL/aYxjZt5RPhvNcE0zRWcbOhklmZADDcAdQ9sFLtUur/NRms/WJiwOwAk
C5SObU9KaCAgdmKLQxRHSCxntZsI9RurpthRSBxIHYKfrV88YKZdCMDzn+yIYbO6+vURzYbwv4Gp
sZPhHL0MQ9L8y9sT5gmy78MyfuCXwHAiYTKOHeNap2OybzzfNJVgCjZI7Bc1S553+q4w099pQbv1
ZoBrkOvvH3+VqpEKA8DyZ1Qam0qBzGIXwB33oW0mvEi5lTz8Dt3GUzD3bomtYOjRHc6nLPmLHGXd
1up6iw0KHovwiGVEA54dESsTlv+JLnBlZ6FJLWt/kba1WxKhO5BeIkx2hM8APpiy3rVUq6zjuPOe
2MQZB2NRhhX1S7Jz0ORPnlxAeDA3711ZXBMlmyPDaReW3aI5DiBOz1C7eGqOsMpdsT1UDqbCLP3a
K+zjwByJBxaithnc/vD0wxz5PvZ6ulZDZi8oDdkXhJI58XaRQbLofkNhdWp7lBPzpFrHonRSH5HU
VSfCj3P6VgPXHz7GxTaUkn/gUUVm1Vxh5Jlhm9scnVC+4D00eF8lBhbOBkn+dFGN3nmDt7lT4GgB
Nh9hR4/R1dSLSG01FDyzN4tTk6NC3fmoDojFzVGjbGkMLPPUftVxZg1/gv13gf6F/eM+TlExWsfZ
pgMaTdKjj4YkGQQUkH2rNippb8sWCpenZVQK/W2jrYSVQX7GptpU9MDEK8hqQnXqkEW6j7vNLrYe
u/sUsXAZW78Pbj+MxW+KtOvCGFbxVKjxKwDlxaeD5RcPk3Wnir9ONU18726HMOIsuZecohhDeYw4
4OdsKCB/0vad1wvFn9+CIYoqmF8m8qS0Zuuwr/+W1FKq2u68E7ip2xhR9XvQJ3hruvUwKaUCA6VD
Ot8ZIDLeAck9PwhiPG0L7+TSazSNjo3Ta4/PRv100jTVPO/y2+CHE5gUnmwVawpbkk8YOorTt3J+
8AobEpe7isnDhOZocggiTOLRncvqavDkKq5vuNQ6OVJJaDD9zKhK9G+kHqHQHOJRul06W0Ul3dvl
7X5hPDVB7Tr3VhJmo0TBzzxJu9kKvTcUf2McucCsIanNsisyaYwF71l93aNc1OCV9dB/HUmopouW
NIb0Oi58jDMlufROwDlWEFP9eLJeTg+OQcIy5mZP6h+fPa+qSsZd1T+IL7KUSp3Gy7YT3peb62Ex
cdaT4GWN97En2Dc3V4f1wBLADS4tUH8HKpPpuV3kWGZ836qtaERqeMYr1dYGGnvPAUYyGn4gfOBM
dgbtt1SYG2yqPGJhD9dTDe7bkoYhNDY6gkn2Orgq+IzNiAPpmVGNra7fqu6y+1sZLo2Moww87LGg
+YH5eJlEfAsnYWH8ZD2CM3XaOHkCkfSzBh97vehDHvJ4dY6MF0G8BMLGFYSCm016kXjm1ZBIVKsY
Op85aSZvR8+picjKM4rAvDR5FGvXe28b4QyBij6obQ+Vr5knr24v+BOrynx9cyGbnApFX8j51JRL
tgLwALCsTPzpFUM6cSmsZ5RswzLQmNgmwEvqxtLNnSzqHvTIuncEnvubu8cqoKyVAJagyI17YB8a
EXHKaZuM/aPdJGZSNjXbpPZb0lX6guL8dzJpOhJefV/esplwRmSnRaP0O8xBsbPMIriY5R5Z/gyq
1WuiJgOu63lf1Z8ahyWKStNfbsvCnZ+C+dpQ0uiMK0soh5kfj2HUnJxKhWZkrLBiC69QaM4wigaE
oM+p1yvv28Y4Vi937rXWMzs4H2R9RS5d/pOIYvVg9WZQj8QHtrrfLEw5s9ph8uLUSvMlEsLQP9Sj
S82g7wN6HMOEVIZEpqXe9te8yhoAhX71QhKirhJ58+mKU71720rIlrsKy7WFk+0ftdm7iZF7Pgt9
WDpQZ7YKrOPseXogszVfQUIOp/at+ulkoKCEOk4LoAkTM8JBKHCJkpl3lqTZNkYnSmLCrDBSd2Oc
5dpERmKtup44HCyubAe5HTCXjYn36Tw5nQXR07V7d+CRKPKvgFw65se03uEawtP0bwOH6ZKULmka
S9StwnisGgSjvRp5yGgxw55mFIrG4/HhHnvmWARMbVnjvwCrovWynVy62GTstGn7GVVeVsrhinCc
s7+auooC68Ftt6jWqPnBqUkyOydcldQ6vKzNoqBNvVJEi0UtbhMMXE/bTuSGD/XiZdce2IiB+b1b
uFBfC3wSt1M+0YTk0JTXfOvTfT5ZZWq7ZtrcABcRfjbYiPhSQv/TopjMDmasMvD6W9PSgW8glv6T
FkUyfyhFWbzJpeBL/Odl8Amxi6fFsnKzVEbQajozA+g2JEPw0bIinn1vB5HlmAUeUEB7bav3Rrp4
JZf01TcWgTc9Uw6MEytmcTXs3I2yfbDzBUTPQR2L2IhjyoF/e9RcztxwSDUfEryNla0FwIgSkypo
W7gITWJOkYA3TML49gspniluyVuXM1EPQtdTgYUbmFoCbxcurNRj6U4Um0GtY7iTaEjyKDc8mdlW
pdECvXvB2txlqTx3FnRXhVm95u1/xrSqtK2B44qyPFE4YwmyYXZwG78tul9oyKC/HgVaqLqF7dO+
Vx/1wUDmJ5bJfpeB3YB2DRcp7MRkgpfgGVa1xKKg8+43mzkgSxHVahIBdYF2nTrJoZOlbNoXk7SO
AmSUHNUNHo/JhuwiyNvcxfOkGwhLPh5h4yFKYLOcNZIs0mNZ9n4ISIZv0uQ6YNjN3TAPFC20HoJn
2gUDQRKQvXvdfXpbDOphh/DlF8k1MoVZgpg967jzJob8K9LxIvUs2Qtuiu0C3EJH7d/EW17xmcP2
PzqTs0FJLMCe3yK6wVta9jXlvLAMH7yf71MLj20o1mFAHWM360RR/HHCUP6ozx2lniLbA0He3KJc
68nHnwoA3l81Wgf2UbZOzUDim0zfp6JTe3WSV9JvfJPyKXTqnJmY216dazkb5kEoiEtVd1/zb6G4
LYLhamEbrqapK1Iye4udXWgiwFPiziShtgHRPrrjgSycunSH/sWTtaaHXoGNwghEVlHV8fjfKan4
nM6IrEQqMSaz25Nac0a8GsilYEs2Xxtn2cuLXr5OzKPUmFjAp9Qf+JCv7vAQcCPSTNr61u7rYRDG
xT9qGmwvcP6/ushmIzQfkPCmVGEOUmUtGCBraeoS96wwaG2Au95kEfCXXxxl3bxqnKYy2SHsyDoo
H9aK/WWG9FBMZICkzo5HZ5YeScweA5fxCStFUUhIgMkD97V1+tVtD+dUbevHe8l7GijlapqP3IPO
qABmmSuoT/rEQmXiqZ+y07UtViRLVWz9Lxl90qyh7Pfvem2VdwnRRIQKyPj2PApacqH8N5YrFvaC
vMzSgE3NjZVeO4sK+cvaLSRKXazkLSAjcwd0iTAotYUd78e8vqkzFxaLGO52DerFmXJhOdpfv2yF
oRtKYTejjin0BWQInyHDHsYZy1MA2z83uXvhGPXNKVrrSy8iBZQwhp9sttPGD5Rso/i1mM6+409e
pKSlvRLgvR6UivqRrpJfFVFc3IFDFXwXGxyK3NXaQR+NZDm8XX9fzXSqfdrvvBPAgvc9f66f/jqu
C4mw5a1xG/OtiFjp6y3cq6kjp3JvJbWAJeCjEKO9VdYiEpovSWst8J0teJdxwIXrS1IOtEUulos6
LrdbH8ZW3FGWw4RH2odv2oqnAOSdj0iGBlIXtdzRiN2CdJn/rebDnA0b8JrDMRlB6mexxgzFu/VQ
w3OC1ei/4U379sXna1r+PPflYrblYEZOF9yGOBpoOI+5KnhS/Nj3xVf2Cv+KxkRtTw02TevhZ2nv
hCzGLYhEv6DRlu/FzeijoIHU/wG2i6WkKWuGTm9tuB4BRe7rh0fd0sDvDZQu61uPCD5VgAE1g7eZ
6STeeqgQGZ8cgsPl0hFCpq5kpeiyq3Oz2pYn6Bs0rmylqc7i5CnBqorlPasWrP/hOJRvPXJA9WAj
b2jmoGyiwv/cxko6uZXPWtkaSHBVME6dbneKmSMEd6HtY63K9VMhOq3ykHQU77iwfwVW2dqBWKHG
DvfCCtykOOhbkfT53SdWnNafUDbLlmKGgtzbr3VlhQvCIDFX3S2CPbrPKl8eyWcHLcT6dCMlbqvP
5RjVPAjXj4oo9DnTzL12pPInT0uLqaXkD6yWNa3rGuSh1/+A34F73JGj0qDlJz2qx1SoHb8oFF2u
/D1WsXWXLHWegOEsufTV7dGdZJzk1tXXOyHrbnXmVUZgpseIQiExr2Yb76HiO7r+bJ5vp/aRAJAm
x0wKfzkrrH2t8wm75zBxUWwu4FqRs8bxhh1umg9LX37l6qR74E63jg6GGwNI+2DgT7X0uExXilPU
GIGf3MQ4Vd5/s5CTfBL/mqrJqkhOdV5WQyVBnzcSWaBEWs26TeIfDpQAK5OHGhEHhmty2iXV7Tst
udj+0iRbfkulc32FsBdATHLXO9l1+OW7TPO9QCD4xSn43sFrIAU6TUbLFa9BErWrijAqIZuv3Y/u
2a+V3u7gdw90Sd4dbSTADiyB4U/RMq6GjWi28JrGxIiQdjXalWY6y8mrs5+x/az0qX+c6sTC/dqV
VKr00u5X9vVnZVKtQ4dhhd7sYPj4CILIYwIJ0kKaLJ3tEulSpNdN8FMxg+0Evf784ytsY/yagoZ/
jFlVUlIP02FPMY1SzoCtoczyfqO5GHvSdM4fXBS5dBqWlpbbyKatd9AyNeQbWmxc1/pGHJ0gfL9y
hAmuDz3FR/oMloh6Zd4oQudXRcecB55vfv9QE/8eGGZ4AHU85zB91Xgx1Q8ikb02O49p+vO7JYdo
F4njUYXdW3bW4syWQeAlY9wKb5NzvdznYrhA/T7N6IpaevIrQZfmzKkejk0xlHCYXK5ItdYSZbrW
xTQo2bnh+a5FQbVEPk99JMROmmuvq/zfLQrO4BQppn3Wzsm6FQIZyX3tlVxJjdYL/W7FR9ay2eOA
jzkmrUXBEfBa5CG7x6+x30mavqS/fmhU3KFEO013B0FYZYpZ+LfaOAZ4Lx2tJvJcJ8c0W13swvYC
IqgUm+N49U1HfRRxL1YL7NWp/il2/ofYpRR6jVY++nXA33hx12Ckc/um0pQYUJmY39eiwD9PvO6P
fNMKhDkwdrfBrehSx17j4KWVYguIszbX9CUt24okwWCtIhnd9e5L4PS52U5b4g13GcPnyxv0Zh7P
85sPWdoa3oFfY2hMBroh8PIRqBQamvoxQ0GB8eNjblt7roaHmbF5YnUbgtCN6GXe4g8o89Mw8FmC
pcG3BV7hKHmuKDpcg0/OrtV0uy6j4orZ1G+SsWFqm+Tz2V4PDiY+jGllDbPSGqEtji4lfC2nUobp
xife/hdhmgC/heoQrdXWYSZfqXP3HBlAOuOG4/xqxhv0RzOAbb6DhmkVa6uJzYUDmxyIGkNK8EgL
Lkp21HPtFU2D8Bo5tgUxzJ58kExwV/S35v1wSbmbT/eYfip51dUe6lAz4RpC9vq+9U0+Nxu95yZs
7HkqdFsqWddYWqIVaFGpablQa1w95+DVl72TioDMiErxfCAnMC55BNCMm7irauB75kCQCjN/1LDV
NqbGvtoenDVaEhsRRi6tYtEcLbPRgDkbwsB/nHhqXE0pInzR3FPI2C53zDWgkXoYXGiuL3+Oc3Ew
QACx73646NVyJ7GtWsSM/SFRr2axZkMJiST8DYQpPx01ppN5SI7zIE83mPn1fwClwyAO2sHc4rg0
+9l937FmVqd0IaRdWwmtB43o/WMbUpKUhyjdmTsjuewEcL8mbSAbozFCH9R+LWLB0tXCyA9CUrvN
1ISIiGkutVAyCQU26SsQwmH0i9Pd0KvVus6rvg5s/u3LoI7NxarXPTkso8aSrO+3qOqTRzGdYu77
rN309JRQz1Sjggc7rMgVw49jb7OF5oukiHriPIVrkL/6w76muw/AiH7lYSG1zdTB12/Epg6tBqQ2
/CESeL9IayOzmTDAqWoUnVpAGjK4NyqVuSfI8zbFfQuvSk0gH5yANNV8hKP1bta7YYWhVqST7Kwo
MXVrAbpY88ev2HO7RHmR5PowfD1mQnpoh/+L9co8jB/FOJRxqQ5iY+RDI1nD9Xcvs9dRfhJczq8x
u8WqUQ1LvuAbHRRkWDDnwvnj70BiEnG0XApFWUAW58ccs9PitaYNahOZkQMId27tYcwxU/X7Jkj/
I7cdfyIcUuwAvmy5xWe40+vIrYl4ehMbCaQp/WdIBxnmuH9n+QMBwlrJJN3B8HvRmXaYl+q6IkKF
A0H8tjZOlx62H5b+aa7WFmWRZrZA6FFvtXrxVN22a6AiqZdoDsAZW9qNSkJOgUDlGZGqbOmjbSQb
wH/0GwmhoxgDQ7/YoXl93lsthcQAEPxDNg8zpsjd1uFNFAkirMOlr5gjHYi2sNxHyfs5c1zoBmHk
l0LDj1R8Mar/taYNZcuYybo0KBsZcYobkUWAHRyhyDsvqc1i28ZeJIBJXZ2LSrQME0++tilpzgzz
2jP9c5+v702/p8bhbeCuR/kM6l4TU2+l/XJbwF1/13FY4NuOimTf3Ci5dV5LGzs4SDlKPT0mA2iZ
k73BkdIvfYDpUJAS7LAfCLP5LoyzOo2ohLa20LGEsqkhHa2nNYLBvw2gjNLsl00E7Qttn61neIGC
ncwVoC2wWMpx76Xfu+WsBBOidQcVpjs8/5oBkmsYT0BaG5AYg6+u/OvdsJkbBGyNVSFxu2TmHnip
jGFMepe3DTr4LSh8KxFKy+Kx8/jSRuHqaPO2oXfMRVNDqLAj6OXQ6MOEFnoHIsN0BDNscIUhjS+P
Cx2hIBJbGqFlM+dyMtrHvjdw2U2E0jCqY9Wq0+DZJSp1nJnp3rioPFqlQ0cPmR7ZfUcc3nB5u5Nl
FDxXbMgJSs40/I5uA2E23o1B5m2oou4W0UlVFPSL3DLYaCUDBGGMAOWpZEtrvBNREjpqtfpvu/1M
4+XnzLuK0k1SUU4itD6n/sNWkKRVAsc2QgJImMWJ2d2Ry17PZlAmH+0qU8+vUlSPawgRqUV9Dyd/
jJoZUIYuCOUFGyNWQ90+J2sFhjZz7Dd+qZ5obJeTxNW3RwrIyUTSyDqvkVVD7wtk7vpot7zNc0+h
0WQ7XzRLB85HrfPqdSliiwNm5K1XDPJdUTPl4lvM9q9OXT3XNcspBl+Cr6TRW2GGu0hQZf4IkpxY
HR/+nu+V0DZcrzloxNxni8a3ZAIUwmNsMZyMXlh7CN9DRyomUm42cumMmY6F6sJv0znB+TpZZPex
rGEbZWhclhxU1HCKDB+eNiE7lb3FXUSrAzM9td+wnY7/gzUAU3h+97zQMcI2imG1flNtOqmntgsl
xyNhg5O9u0I4eWcPPYDYxs0DV/5XcX4IpbLbU2xjJNzn9K4JfmNhpplut+q9o1t0Sa+dvo5fykRx
LUii8PPwPUa+qj2t0uVzWdvwm3raG9Luy5IdQ6HQfVoB4YrXHa4J4uwxE9XCl1mbsO7q62jKHNnc
bbMaAjSM0J3hX/BEGxluwQozYW0PoKJtiaJcQqz9Lnl1xR45UfnhpDfQr++81qN/i4yjP+9oX6Cx
Nl+E+w1UFdGcKReeajliMrM+IzS+Y/xUZKY4+Eq5shx8gcu7WOC6MhLhUgyWi+aAFuxRr+0GB2E7
4hoz21M8nZcf+M1NP9FmPWWqvJTUsXgeXje2EhDLx7587/P/oBO3p/mHraKykmbzzZdlr7CGl4hy
kTm+Cm9F4r/FH/9Kn4GwUrHX6IR03es0LU+k7tr6YrKpYPSyU1v/9e42xtUz1TsoNtWUDvFkEUnU
S9UnVSUs4725BJoAbsXBFD755toSFxIRbIK7mYMyZEpm7rVdsY96+f9GqdFeTM0xPP8TrFMyK+Cs
n9P14ejWwgwSywZCfsuCfIwSLGaeQ0X5RIjvnC/72rL58c4Iqwo+hElFDOsd6uRepXcG1G1FAgkK
dPYRMGb9U5C/1QpfvZd1VC+Wb2URwIllNl7YyFDzaOq6YCGDbyZlf7cQmts1f/ROXxXAwukW8LC/
nKhPERtPJWNnqhzsXjzrt0Pb63E5ieY100wmK2HxcWscwuv1+eKjDmNfhSjSMWOxmAZT9IcJTwwb
+FAd56W7TWWtpPULicpJWgNUebXWx3hKuNbT1EGNeLYMKbMxWD+gHOL6jiyd8ldprnmaPGurLcIr
HPN5MAt1husiMEyDupX8vSdSI4sLVUAFIoPvyVQk/W0shmY+KDFlgpbAnWQ9CcNalEUMAMcW1DUk
ikNS4os3/2H5DhIxKq31YDHVu/jhXbVZSLAooC1f7aLKSqJilRECd491Z4E3FJAfEyuFirsNS6aZ
w18BEFmMVF4uH466P+9dwfwwK9H57TT+Kt5aDffixXKMsRyp737RPzlQEAhF0ys9BuQZ3oQbrfCY
u+0UIuefeOL4XO0xcFJWiJpeatDlynH86EqITP02Ml4ZK7FJMWzQG3c0hxPH1XJuJJQUAimh9r3o
Ld+15GVthUr18Wxm0YNCT28BP3t5FZbo/47gDJxrA572jCq4bWlwYXF3wY3cMinrcoKJIUBLxhHg
93TAdXFrCu7P6BmmKIGB3IGs++QD9p4Iu+ya6Q9PZ6brnZmdGVA1TCqswliVT8L/gSM7pDIBPrE6
8OJ3ISO0nKP0oRbH/uk3msuOHwvKZJjuvMPMyOT78tZDtRD9ut4WZoRF2xYTLKUmZFYLgiAd11LS
naTV+zaiASp6q/gQ+Wyyp0QmHsT/Kqf9UYCMKwQLVlRbmbHjrpbkd6urj9S2rRsKbEozpgzhworA
fImULeUQmzrEAolSonxWuAPdsSbzA6gRDQsDcGXxi8IBGiCSeA3ZoqfB2W0lYY6Vl1OWJyuVkHl1
GyokhfWP39AnSD8csb7SpZcVm6DfYZk7E35yV+nTasJ2uZtqQ6bgwZWmssgj5sp5TINr6mZjAff9
i1teeepHBcmwd3cwqcqJ3GUzG6N9zm5Jc5WnuI9HVbZR0y2P8Ez9APBeaoBwOMJ8bmU0f6thOggt
abNHOwRUaLPMRgRYpey4WTrLVmDU4v6WZ8vMhD75ODyFsWIQKC6i/AnrEXJPV+/yAHB890ok8ViZ
9M4slg3H2YagM3OtAzPmcb+tfTlShdgAD66RCbEpxbbm3DlSRxg/FO87GFv/Bo920i3v3K9k3qSM
hUy3OLtFrgeNFKMJbnFJzKwT+3l2LTMZslaloLh47qioG2kT5rtAL3xmSdqFC7e3vzVv/0t3oHIF
3k2E+Qqdc3f+9kf3FWpQWScRkvk0p4TvT1O/QICOdWKALzOtDXARBRD7IxDbxUSuRkjtt1dA8ILH
5guTW3fMbi4jIqvZ/qUBDKQ3KY5c2W/pgrnyQofn6na+S85IqU3MpGgF1rSMgo5sTUlLYHoFS0Fh
7jkPqw4ZapHN0EjcuiDHNJL98v6sItmZbr55CcWJwfhuMZr7MWRaRZk9PYC1XqV9+So/kjKTdYwc
gzt5pyC+TdFiubXF+VBvnpzpnfqgTjJ8K+yPW44/4FYkEa8YLQHlns3lclWbxqDgKtgaDanj5m9Z
haBk0axrBn8MXcccfw11Df2sGd7ZfjtA2tTPUGkYri19jAe2K4XB3vWFj+KOxyakSpEj3Sgnajaw
lgp1pPUSjezYPnNtZUgZBMOCAg0hkUHWj8ff2YEOK9Yg6GzXlZGYZq4w6Ola2H9DmvH0R3/CZ4k4
M+7Pn3P4okSpa3Qb+UE1h2vARg/y7S0DeD2zg6GILj1N+s+tYnwJ7DdQqBWPK+6uInyAjVhLt+Mz
ofiSWgG/exD6j1T+NT7LQJodsDMQj3RdNYlk6HV8uVNhkNLFvonilvNG9++IY1uFkIOrYFvZbax6
9QI+NTxgPSBnJ8C4I278doi99Qj0xGGFZD7+9S921eL8JuNxET1phpPSVgbxm/uLMYnpX69X+Thc
+mZi7OsRdAJj0dVDen2UB2wnUBa9ZlgZT+MUxMoTUeHno1MjI3/bYouorufcMTnFQXKCIo864DjB
5rsjPNqF360DC+CZIGSTk24iZjJKtOVKzt1dR712AcCq/LIZp04E50L92TOFoKKxUI/XgR7in3jM
5PYGCMmDGjOFzdmdoSY60y707omDSl2S1zG1WvVvpuki4IFyDBQVnCIbecgLXv8VglW0d8t+krph
4D6FZamwUAJjJMl9/1v0xrdw3JXiIM4ArAuBtZ7XAeUdIBgXFnlt/I7awK1DGSTgnHS8SD+5+TkX
bbCXE3xTvkAnu/NznH/hvXmn2GtA2deHJuv9oT1Fhc66Xv5eepbO0WAJ28QWw4EGzcaKAuSyfWi3
YFsWZv2o9AdXBJopdZkOMVvZBPnXuE97LbXzio0shUy7PcpDCetUDEhP+2O9YI89NPbG/UdaAwFW
c2N20mheRP683gx1kXV3bSYhIelXX/gqHTOX8zE4jFfQNAEJaS9Xk9MU7QU0aMEXxrHDypigI5Zf
niEsGZHvMnuzLRGBs4X3W38F08cVJ9ZDzHxZQ4Utt/LZwlITfI/fS5zHsRnhSSD4XUmQnq7uz8U7
iy45Ew1PpvivcYQ2fZhmWgRVCaMzoxgq0uEsisf31wfIJ1FsRhwdGiWF3N+vhAhaua1J/W6jz2zo
D2EhpRqfh/3TeCHAV6YE/lf7EMKf0vnA/pBlRCXBCf0ZJqsGEO0EPPfCdtbjxtgm1nEJ+dhLcuJq
2WLZ2tNdy8kEbXvR42vreqeAmsR35DrMIg0pan7WwrOoN9UztXZcIqGMqwlLxPAcYUgPpv7Sz++m
hN3TRmx0FwWniky2JzxB3/sAFm+f6G30cyo7zA4NUxElYbz/KRo/wAlGLAIbC4hakSh7kKi1L29L
/QYyIcGq3k+0Z4J9gUg1PZUfhpz9TD2eVBZD3fHqCcrK8Yxe0rKB8nmXI7pymT4hREeqF3idl6OL
U3gxicQtT3g7jxeBxrMRtx066CZw3DbzDe/8cud131H6s32D3PxeO6+AtGTearziy8W6g07Sv2OQ
9pMQo3qeayT8VoLsq1Tsi15NBIog+HgEq71s3MBtkgHQ/QyHi/3MGX0qCV67RxKG+asw7xjWHsuQ
6irkyxH+/NVhzEYHhRpLMht8biWTxNhxHPTrCYxXfsld178YliJKjro0uZC4NPTUJfTsxLbjM6+S
kBPS7I/1t7ODqDdyR0IsX2abPTPi70e1hIStyATQjo1Ev1wQMaYaYEFKNwvGePBHTm4wWEryXL3b
7org9US/wLwF4JyqYq56SYzJT3GS8Zsmm1f/Jif0NfpXYrkfdBEns51wzuVB479ZLjGVh4v9rtwB
7C6Xi2gSixs+TwMqJXWlUhHbVqpUlqJJ47ZQAlJtio7d8gb7OeI1B9kzhic4GTsDsOHApJfdN2k+
weXo6xTPXYXEnaf6Y6h+93uTvaGje+K7+tZDMgNXmIKIM5qMR/xsbkAiOeByXQ6ZVHhATvzIIbHm
HvsqK1RoCrGgKk5lmDOUaWkZ9aa0avrbkdwkoswDml4yG95+M1TA2xAQ5kmgOol/LF7PxR+tTL41
9Q7+ykeQR1HQ4o8Gzng2s3f9t/VC7GscSDc0uCMK0fHIOE2q2FlvrWs1rV64+N5S5jF/bF0k4WV3
On095HwpsQWVa8o9kYMHVCjYXq4Wd8jy20YhWvmmXTKgWtbbirtqsvhnXpEquPvf+JACY3zzNmyS
GDQEoKaC2LYDLZ9LV88X5W3ZbP9h43muF/RubmEEYDQn2HPDimTfQjActt4xb9sRs9MsUNTRgA6S
YrCPVxeKcAOWOIrE2+NaB2lsP1jdwODFeKbUedcs+/RjbPJXkjPoLE3X/ZkPgMNlS1+JB64Fuc4G
WCADj7a2i6XIMnfYkM3vVUOLgmu+udFtv8Q+jz2rDiw0JCCATuRIW0IECy6B9FIPWsPLkE5iVLgA
M9uFK+AnugXOmp3GeH24aBuKQxFHML3P8KzT/nwRPYlG+Tn+uCbLWVSyDejp/mKYRT+XxO31CjtD
Mwm7h8FipgX3ZmH5ibHkR75/YQEV6NPD4IuaGO2/l1YjHRMiCgKv9+0DNCH2MI2SEcdjuoTKpxZv
oPwlpBbc8ZvKnyIEZIVROYFBgChDz+tLUMkWNzOQWti5K882AlVruvm0jMgukMpDuxn/lQFQAw8e
ExgWld9Z97LyIxORw36s+hXi0CGpokZw3iVjIrg1lUieYwRiohKE/VjhoH5tE6SP92ts3mlonTC3
nLN65qoX5WgGwdTdouJLbydThjcGgj2fRyujN8uI1zrabUe6Yq+livsvVNro6Mqh9oVXBj0Zv1lL
ods2OT8FuIaY7MAtO6wVuRdI+8kXJhgqLratwLnIckVxmhGWORbV0wWUGan+TmVoM1KeS8BA9B+o
z4T+/iKcyIBZ4Li7LxiF76UYBOzfBaP4yVxD0Of8ODXm0Q65I00j4gvvADbLZxpwWk6rt/iCfsrG
33ShV2aeE/LqQOXN6gprAFKONqpgiSQMzwN+kA+dgofjGwNBRis6O/YCht/B3DaXWCbATyu1R0iE
0ubtoJCPKRUC4oqqFN0Azz68yCxxfVMWjUn60E+NFKzVz39UHaVN6NanFp/Pxq8nGXtMQU7UYuuu
nrbWhtz1uto09YLVOL7q6RXpMaYvOBEJEtnkN7NB4bmquP0nD7QGqYptLgZD3P6Wi4XMGdDAMPFh
12DtmV1KW1IYDHv1W9LDj5mOr8Jz0n9JAjTp3LtHMY7vv/w5G4GZScJGBe1QzmuFYq/oVPVVCRyy
wCQ3uLKd8iq/Q2FsjmIWTLADuhPGB6n1eGUWBpC0KcAmkf7E42UihiS7DbYk4rlknl5F1lntMGeH
LqTZ/QDH2SJkCQUUCcD6A0VSHIppVtmhphzpIfc+rhymwBvjVc37hnk2Zyc1tDP34kgFCMJhqNMI
bbbTI/oyMtLkG9RzQwGZCki0VtgX0Fx7S74+SA+onf91c8AFycPYMg1uvSLW31BUh6g7Am+0tczi
2JGehJ1aR8kKtmdUpuCZj9LoM5MzQzK0pjsOytDZkc8pE0G/+PCIwHNIKHFeuBF2sxbFXUpVvzPI
CMw506okuk1xNaUX3/6TiiAdc+MKYKI5BPaHiySWyuJu/KP2DlVgZGSJ2ZEmCH/WH7cdNXgmk0Ox
zLh8Ds9lCl85ED2UEAqGx2M/KmkSEs6pu2On5lZxL0e+piIodh0zQ8rzTNDaCvVhJh5s84dWGpCz
Dkw5fiSzgkjhzxmUVB4fYPcVDd4YsP+AKGKS+ySN1GUbnpzrYsq0ISS1PbiYrwJKybUBXlU6ThqG
9/8tMmOmZatpAuKO40eUg6SWNrMwySw8ewF1TnZ00aE3nrK0pUJ8IeWDye9GivWk53gMaAluXuVz
xH4rPpGOl38uFghPbTYeGwHRcol1YWlfQA5X16I4Ywh+zL80xFHcbIGZCkJFcDmuycBVnGPUDupq
x/0W8CK/e2QARV88MsEROo/o9cHnmrsjUS3wZajfyWRJdvJaSzqgHu5oyLB5JMVdxEQ6NE49/zZH
BsNU+TLAdFR058oNOpEGbn1D5cdaGKqyHz4BkXxqC/gW9W0sp9LFjQAADEuV1ARZIp/y0JDYUDkL
pCWT22HjXgJVlanzzggpN6szUi6jNmPP6H1xkqcMgOfH5bspOiVr2NEZqgZt7TI4oZN1HUEutpOn
VPJcUvTt47csXfYsLp7Tq0AfECf9Hzvg8swLSqQ32PDz9Dcx3YqYZ0zaPbsFd9IBY+y13oX1tRjv
sps67iHN8co+j24CpihXe+ZY+V9WXGQmcKPs6Hm9ufSNw71KWodEi4FQ9a3EN8WHV0n+zE2pxjyE
mnD/yL88rHAgmRfoQ9o0anbfDC8kY0W9+hWykTaJbdveoGJFAJvaGVgdIDyyUAsL38pu8IsPes6p
H3MuAzCadPlMvR6spklwUbBD+GuT/DS/LDW88mIVRxUbIG1MqaiXJAgFEcM5D5UBVHAjBK2AvpM5
QDcSFHk4wq1xBRrYTFEUFEomDlOhJRdqzwboStGv1VJgdhgqNXTiQz1bAVN8l7Hmf1nB7u7YPz4I
zZ7aoRCyVOesuWe+cvk+4GBz1C1iwJc+yUfIgS3GWPEAaWHrCeV9v8lHlomO7hKab0SAPPciDb2t
HknrquGv4Qb+djsk/wu2UiXz0E+HchpMDBwF2HuqRSz6oUlrGy3OXQeeY7g0IOS4wgYq+zQOCNPu
tfweemY71zJR8DsbJTCVCcYsNKkKbbu2I8RAOssSwfKmzwvqVvWCVdNUvR1VWTqCNMPEfrcNl3Iy
M76cVmV2XquOvWcOXcfxX4kE6vEl4QFXAh8YLKO60U8Tx9qKwei28DCL0tivqMbI6kqsCf3Vd4bG
8uRP1LaTb9cYCteq8QPbJ8f3wo2NCZlhHhdDdSmN362M1vyIntFY9aqXxKKLIL1BRj4gvCXvwSug
t9/WBnQVPvCQ8RcdW16kZa2d0o9qjeCew9PwVYJ267Nmi9DjUTu1ebzp/e23ZQUzD/i6hLGNMdJT
bhxReR48uCHUUKegvM0J8Cx3VQB2nQ+xO6Km/mGuasCOFM4UUsyvVXMXJNrb14CZX9UsuF0u1K2f
fHGMfrU4kRY8rJBs/nCljtjHtTJIV/5FWWlLZwUH/tVywBX412LhDwTNclbrN1ymQXVm3xN+nj9a
+qPFoMrMcSlUYqnKXgx1HLlz6whOnxRRfuYvWq20h9b/JW10PcHVL491+Idj++kU9UOYVQmKdRY7
ip02nguoVJ/Z1Zo/XUej3rQZ3x4kXuMPHrf4RaZRzKhNiDA+NiASJ/pGyaV5tsVB7M/zDSOgsKg+
Bjx5H7vWD4f/r7VrhU22AeRfsvR31h/JvlS50/lQvVtziHjKksZTTeMN4hZuPm8XBjTxbHhPUUT0
gCni+vQEmlSsB8/qtgKHQOXJRzt9hW6O1eXvia1zjVLwugej4o1bdtqyf/QMiuaTPtb7NhQwneXj
K+jDxvdcSeQyYVEIPPFfaR8sZ4QNKrKub3Fk3FiePNTYITD2Ptlo1XpeqDhgkm6MgcJGpEFN9lZu
dgYoI9UCyR+u1mRmQbno4dBpluZj198OCj9+zgXVZ7lZvRHULes+RF2p9BH6EJvjhubT2fSl83qq
9NBmE/rc36UR92DYItXGKUazEu7ZSrqOZmZcW1uFAoKtZYmyi92X4b2azEuQN1E+1b4uuprga359
JWsls2EGVgVP01LDfxipieZhaE/FwbaqRsvmudbX7Cb6W4H+02l7vGtcDMUDMVr7XxUg6AKLT4o3
jFGfBLj6AwesQo42FVUfMt/SgoIB4kossUzOG3oOLsQDBdEA1QoqAHAgUz65gkp/EyTPX0iYS67a
ggOpGfnGB/7PF/ZpzZ29XnZTJWOIC7p4CqKAUrMdoht4kfK8iMnIp8KRh4te+b+lktzcgzb3+XvY
MuO4tNXn5NxCyVXCnZRJjhAuxRJKqPpDmbVSx+pH0ae2TbvsBMlNqdqmlM8QWVv8EQp1OrC9azMm
uUNks/XwZEHFGbeMnwwqtIGhKr9iO3AK65Ea5c3rNR5woPiQtZ0gvN6/dLAnX56leylnaQOJ8F41
+zk9mhvAJg4E58pOYxUV6GDd/chJbJXQ3wZNCjB31h0isxOCqWAERzrMzuMcE3VolESYrZZiPysl
cyBg/ZTR7KhEEYE6/X+7u20tR8DXbnka4OmScffYkmJQ5ID+4mY1v12vVAs/bk3Q9G5FLNSRnH53
T+34n1PCFFXvZYHPYkglwoR2YNa3/9EmN8Jby+COUy3wXuYGvsbIWz54Sb3ddiI48IHS3D8o/NlV
tQUVdQFgZNmutnbtKdd50kHqbacs4H5z3L2di5aGJc5LH1BIVf/edgSzjBn3VGs4dx85qyZ4PLPk
YBj3/cYrFOVMH95wkAkyYSR20fUwnlB8syeuBf4RCTOC18fxUXQ77rNbxJNSIILQ7VOgINFcnKt+
zlrV+sLxhbABPWCv/1Yt1y1j9o+te5hJTvRCq3Jrsvm0eFBHh/DKJlaLlnQu/TB8Cvn7KB/WbXji
ejB0XPmqWYmeMQZ1VI/jBpMNjsvsnmZigXXa7o4LRqQXMyHEeB6S+nJWU4VH3YsBMHUlpK36xE2F
xrNZuuK9pszA/z3H8faz5ik1hSNqFS8UqxivsnrimQBs5Gl5xCbwU5HR3OP9v16ARcrsW/m9YhM7
VedcQgfqmoLPtk/CWttZYgM34t0mh0jGdFrOAm2KSJ+r7gubZXyLwgVbMBtzgZMNEoICL0aV1VFx
L+BZd2n+nHZkfj2pW71kNnnuHDb8XejyChelTeK1wSi6ceVhdgcYZjXbpzX1z9eharWAEdGWfC3a
g2ta/YLcyzkG4+/Rf7jaqgWIjSGZdtLJhv0D6C9oKmNS5N4WpQ6qS8w6z0EkELU80JO7tO8IugLe
2QXoGB/fzeUGjmu07Si1A2YLCeF83QPkw5Oc1Bp2YJpK+o7FhT+Z2Fe2fqL54iKRntZxOFfuYiZk
IRDJza2HrxAaoQ6UQTWGThntIN9dg1La3LTV4xYUE2KrM6079Xb4c6RKQgSdFyGU/P+/9CgVSjxO
c8ZB3zfkXaqE3zstAk/RteICRvDkPBfIfV0DdMlEUzFcQCepj5yeaOuntSRz9Fo3Cow2iKKym8Wj
jco7AOCErn9U6OZeDX5ZdU72QYOH+HRY4nrDTZtpmvaKIiQLPTJjUeVpccX88a4TCW6isLIuViyH
6NFuHCkqsTLd2ZMtnz0hzJpHCWhC/1FADUehMcYGLm7HiJDmlBdUNwgkhvBMznm+Iul+5edBCID/
3H8WoERRPMGWi51pcWdBfVFHMGGJy0jx5mWYGv4Q/dGomqDGL0iP2Sa80dhXkewQsz8WmhkVw3/a
OhjuxrQsXywI2vhA3xmHxED2e8QbNQJA9ZKhTgWpcZw7ukj3CFTRDFJ7l2AJytGBGRLyaUmzbW25
mfMa3pjO3D1WFAtIewTAgXSF68omfh49ACx3Fmuqwjb6c7yjvVmuo9XnUyTIKWuQ/4JEj1yRbvkn
OLlHHvZ048opnpLWMyfRF3AX1G/K0+xgQFUr/r9ddzO3mGxDK0/5gYT5H3VwhNW9FLNuoG8+iDTd
b0Rze93lVZsLgr56vHQ7LlBURg7Dfp9OkW+EIH8LtgTVGSoDrNp+sIAbW5aJbVgvAW+sw3GKCuxP
4zUg1r2R76lGse7/mx7wu8JLkNWJvBcOvQxQPlAkYj2lIQ/0ntv0f10pZbQ1uqKtmfsMvm8B+va1
0MfWIzD03/6WDDzOh7cig3GUw+GJYWxwLXEENCxgQBLuk4Z7zy+uY2pTUbRahBQS7cN173beg/rN
KRbeYtt3qlFQ/R5V7y48qCOpBQK3yF6+B1JWU1yA/CHUhsBG4y2j6xn+hBg2zJr6XwGM0thS4r+B
2otgDw0wbF+i2oqeqhkRmSa8tXsHmonEJ18BmKuTz7X3zwebF7TaWuUufrb4Zzbq/P811neoqOBS
1FMd/z/MojOYxkVk8ebJ92/dRx/8AjROr8/mvLc5fc65CwWzgFrYSrz2ig/he0h56OYx4EzkPNNF
KGIWVKlZafnl1ekt5wFHPe3ab6NPqYQ5NYj93wCTxOxt0xGSKyiX2OZXb5FHpp9Dg4xNq/Fh8qDx
bBIiZWD7YdmHdmiD3V+YcFNe1gT/FoZHb66S6aTjvSsmx3S0XFwklSWUB25/5Vg1Kehk9NGsGlAq
FS4uYdM5ZBz8ScQXe1tQRvee1lO2knYDXD5IlYtK32sGBXjhgntCH8a2mcoBiJ1gL6EiMxIpJ7Js
vg6YevLS+c2/W0OFvl0B+t7SZLRDUQdPk79h5QrtcGFseLUbUMz/nmCGNRCfZ6YrFeMZlxntEc9b
s4kgrEAc6EtKmnn813fXO170+AGnIERtAz5Br69nEtRPMmFbVQfc/9qkVn+NMx0yOdlDvt2dax1O
Dn8VCP+50Cjbm3hoYkBP8zW9j7Yb+XmPnjMhQRHO0R43L8uyqLDHH+CO1X2YJAKpTBopzHnPurra
zUPwaQNojk6rOGhVQU4TzsiNTQL7WTa8IJ7fdzv5/bVDocFnFATU1xE922kl1X4Z5EoIwxDIKOtK
IPxKSfeoys2Cu9ImIH4RjXOts0pf/fpVNEBgGTc22JOkT7Kb7z4hQHzKs6o65f6KoLCLgdDh/cCw
kWfyml6uyQC9gCjau4x4rL09ZRS5x4Ys0O/X36MuPgFzi/x/mc5l3z0RjpNWbDDwT5/KIoSryCEl
iD4bH2Zge2b7ZIBxCrqHYHomG5JD0LaofbcO7yY9LTqfzkd8CWeFhUKWnBNY+yTwHGQcLFz9Masx
hxI81S69FWPZo+7QAlePCBc5BxvbJurJyGYsUZ/XQT4XxENn26wU5iW2s7UDMOaN1XLk2UpTe5Qa
y77Ht7zSmJwa3eR0VA95P8Ov+VpecIT4ms0mFyx/gWh/WcS3X92XmPwPKf0RnaHvy5UOJGyP6iWp
SWKH97CUFPSScCUXCuXaojxjXDCE2mop2qDRSatGTl4ZSS3ZX7mb2cz1EsRsJqMkkTowOOcsR82x
G6RcM56jYmTB4hPKaUe4Flyf39mTYnV1ny7GzGBL+WGF8bUmYsDGm46N/0JwkgIEtmS6TfR0GIen
Hdss7Y6mBzD4JN1Rg2+VD4PZT5nCE0CS+ZgUdR3jzQN0yzXmaCfiQNXGGVI2wuMvub6BRG7lNx1b
XgOW0IiaOGKppeq0PrufxQ7R03FZz5oLaqRJvNxrMCEW/BKK4my0weGBwwbo/20uzqI+ZiXzBQqK
nVrr00lXelWtn45pQsU48BG5l0BBMKwZbsFgPtjKC6/X6uG+t/2mdjyVCRBzV0GOT80xxlym1eWe
KuqShNNovv85yaGh6kC9dpHa2OrCTdzFlsZQy2jEUfIMNQf89mvWMhxtC1MfOGP6+DcOX5fsQKmn
7xstd/tzBtD5hE5IQ8OucDY+hrA1apKJ7AK2bySF80lo2ywmg+3o/QjBXjxi7Ov/hCvH348HmD/Q
sS1pzBH5TnmgUXQe3ShS31VfRgAOB1BmNmrrsHhaXkqWW7znmhqWyIKdHywCkikfm7GkJ38rIVzv
5CZk6oAG+UXxia1QC8VTxvoPVGjpJZ0yTxTSZdNVbmO+8VbRroY9J3xrt9aQ3yHaNplXO9YK+F8z
Oo0eei3J4b+DEpulLEUTft0TG5/ygOeEQ9D15uWsB+cjUOAKbGuifAa3Er69SdjjRH13aqYAoRnX
RDXMHpDXmr+xOs128J0PAeFw95oU49rJ4oGJxPkWUOEY14CptzhQRLzNil49CPuMtn/hZyQkhF/l
6AYqftXIGU06/IjjK3bE3beKGzAe3XQv6oFmlckOjqEq9mt/EjZTXHJg4fyIFSR434r0BUNrIJWq
7AN1mqCFmVxhvyUvl8h8CTyd9ky+nNiut1OHxmvFJYw6BzZH63b/FXuQfh9cMIpLGBAejpKNmL97
720S9FQHM7UI1Wy/5lR48aSScmaz4MCLHWtiqCj+pUxgUubK8SHG73/R9vWpvWQLZF86fPojdfws
IxgtS0bdEFB4/+F3UrYArGWf0ozqdqa6Azbgpjyq4fGBXwiqShjarn1ZXlTMxw+1c38lxHYNj6gP
NyzatkFtAwTkU1q0X/GCQam3GQ54a4mCw5i0j3WT4yCOjgqVk6QguQcj6HpeBwzRZHH1ycUXdNz2
/PL8fv8XV0ZKCye6iflV4a/OOWn2j+EEDtR3OFPQp+tqztrrtoV+i2H5ZPjcmUBcgY+o+4RhPYrM
g5qNZzRpbwcKqyYfzehafmOUyAEwgtzAIM8URT1dOGNeMol6oFCtBD3ecgF0Kqo5gkwklByKGhgy
zLsJco6Hi3HEJZBWZgCSsR+hJuwov67Br6Su0+TCe4XMcNk1mR1dt0RvBaEYwGHMQ4HBLYHiJCLy
RNgfUvJiflmfvNDgn/6OTMT7YY7v0pwkjCZAI0rsXa87gMr/dvg6m5/NMLD2gxfopZQnuMTUjGFm
+5/arujXAf3yXaO2WLGtVFR2OnJOHP2GUnRLwb5d7Ue2p/V/p7EakcW8sjW0VM9NWNRHMm3MuCti
Nycpt8ywOaQjSh9sv1YgnBBt9HhfVfA03xSwuP7R4yv3P9yrQCD2a3qJ0na8pPx70Rvq+leFC+Qw
OgB+9NTe3+zYhexy9vYa3t8CdjhIifh18v2s1M+DxbfxmUg+fCQR7SRmwBLdqmleB2nThaA7GleG
tTX058Gp88OLYGKeR9GKyzZXD2LkSP6Pyxs00EyiRVo0W8AGGV6eMeVbQ0e3HKY1T7NO4oo1b8xN
BO3T6Xamjm+WKQjmUOUWMoTJrUdOpN+0RBiAnBhgo5VipCaKtcJZl9nwa9EshCMMoAOHnX8ACTvu
2SF7W3OquL6t3FF2xTx2blmvuGMFCp0lQDhgubPrxEsVQBeFNremGNh68wgTe4PuVeulpdqKjIvl
SLyiPxVICHj8PkEtapnT0HZ1z51a3ce+Z9+oxJz5/nTLAuk4ypMLgZxiKvFIkJQE1GiGhe56tYJr
rPAMG4gjY6f5OZ+vJeqppP7R8sZm8rmwrBcnwyQf9XZmwiijyOK3YIsp3f1GL+QT5ShcsKDmqwVm
PMsOINDJTAVmeQmcaFmggmGOf0TPPJn5Nj2ObqJOR5vMtISQJJJaUmTbPqdomJfdRjLkZTAwjhIu
Z4RPPrLcuB7E9DciwirXsegfqgcp3rVzkn/kCSeF1Q4RJmn61T4I3XYifOffVJkbAOHwd8aKDCmC
240rWZHHdUVWfr+22cmU4dSDruSReKE4M5+CJmA11uB8ooKUQAhDgaA32jrV4swYD+BN5dtjqHVf
ym3HGzWoEqnQGjCOuQiMB7TqJ41jRxQ6A+gTZdqfI6SNu7hT45XiNmgglfPA0Gvdjvzc4TJlLA+n
mdeq6z8ollnDnvHe2IWnxiLiGkOIFlWf83BBsksgjNEwyDixqn7ytGhHfRmbO0TIl5TUuDw8flvv
TIBHJ0zfhBADJf3RbLxdPVH6QYwIonjdI7CjhbrICaiunxDJbqqkRXVn0TPB1c3+g0ISZwquUe8/
Nas1fb6ihJuht0pfTkALcXK0GVLx1i4IhYM+jSVPJ7eLkCGbpvzddWzZQnnx+PG8ANhCHt3S1WDN
VwDuZ101WuQ6jLOuqMt8Qf/Rq418TghXMbWBSZnCBqRGGzM2oWUZjDoWfYDQAjqGznjl0ele/4Q7
jpA865KRXWurACCn/uDvR5IKdWooMZX42YReZyk9The5Yt1zNjPjnaFGlDX5qWvhOBozmeXa8Rb7
k5EV5EIofGp5unEmvMkPTnuUOwPx02L/wVmQU6Dfs0souXw2WedO8JwIWGD/UcT/wJoijcVz/9FY
AlSRXPJUDYR4wL9GgM+e49CNc31PmVV7sB3a9wCO+aeQTQpNvcit6GurxI7au2UfPeB/86BAuDRG
3w5IWLtf5Oh14tvtoILRNqJsK/J0H0282QGG40FBj3g2OjJ3+oNXzE+Hwn8G8hCu6e/1NC3ea3Lm
XHEdDr2hBYALrbKpsiWypONo+QniWQg8YRnVVe4QzqNzJhaiN3ioWRJQsZNk20LgdgIvJNThdvnu
i0hqRxtiCbgwzL+P1yKqt3V9pMCqGDsd6Sn0uHOyfSIflKuX0EFyC3zJ36B7MXCvXpeqsINlXoqt
OJ2kWXYaKxALxEVTRTvfcxcARHfVYGv9qT+A8vt/0KI9Ebqp096pRX9J51HmKcqOLhGw4A86M73U
90tcw2PZat6d+iv01AT6E6wEYdTgsQk5eQHX6NhC22+n9rsJfbla86OtR+eNBLYaDNrWtwKRH4E0
BEF5crun6au0AKqnsmwvUh58N5ertV3bkvFr6aA7NQySdJLhe2raREJtkW3cSNCElGk96GTQnMiQ
x46BMS+lBB+pq6Y3oxq8yVDN0v+MGFKdzI0ogHXYrp4UxFZZcTwWosxmGMvT/dgVn/JKE8sfJmJK
DCHEXSadu9LaiA1bB1VPi7ZRDvD0Z1VKm5QresyyT7A4Q38PI5udLy7IOcmkhb0EvRM/7qTrNu9a
qaAieGR9PAsfpqYbGoSrc3/vNsp9eDjhVjs6XHkKYsy6fbSmfpI6miWJ7DXec6vuozP/icVHJZxy
PemPhU4EVPw5OWp54RB9Be6F+lQJDA0WvY0CMJAD7nFB7QPzgjP+t+gK3mUVvrZ62Jlph6gUTqeY
cCbLV+T7FgikejpJT1+3o2hGZ8tfhIByxRqN3D9Wvhu5B/ywqk8HfMLeMT6A8D9CMDEpkQCZ8gib
y9qBsx10SLdnyVWhil27NlgS+KfTchqUo6lONXhUyp6MayiZ8cELEIz2JiB4UHPTuDBkE7bEw+xi
7LWZ4+EkE/49UJueqRvrMbJI2o9RqhQnMogwrMaOxRFLlErHclL3u47TxtdpQpsIIPkiSR/Hq8Bv
lsl6vlzURLArlkN8oj/3DED33w3pNam02nHM2zqJznMYAIcjKdJ8+bL0MXP2qO1G9K/kzvEkq9JL
/boaOMCY7y/Yqr7B35YvyLtFZGrP038KXervhgNzQPKbzKQD28pRZrHrq+WQWXbnkdZhWtlZMCsD
c5ARnLDuxbAVIoeidRaVod+CmE/0ivdbBC9BjmHnWJ/6mmNPujKFrGnVZF+yreCfxoqRJLLQpViO
3oCPxd7d4S/VnUG5Eqp/8AVSFz9yM8x3P83krTdapFXf+8Fwlye83nT5pm8fSfOvR4zN72OyHes+
DDcdAL56HbsxWLiE5i6QkMKIL/+UfSGlJcM5R1nZD2S1Cyaa00e6XsVvmHEvBgZ3NGB9HvcCFvp3
IvErW6tYCSsJ5ar8VrWJmjfbfiALIwvaVeNBHnOA3jwTScFi0Godzkrb8FoTCoKKyaAI6CBMFqru
BF4g58Zr6mYZJ2VrpfdmTrEWJF0iSxRcaMdwee7eu4Vqd5tmysur9iDt78jcZBt66y2OSPnRUU6W
YXMeWiRJucRyiRDztG2tfKQUaZCOkBsOJeNDxl6OCV9AJ83Ocp4EBbnNoIjMRQ9yGM/8rxpGX9ky
x3heICSIaEXmhp2pC51iSK8keqVzaxqw4N+LTIh0ONmfkdNKCGe9gO1kGLu8TG5FC+typHHLin3f
ODnIwyZVGMexLqZ+XgcSMbyNt3ptapbag1GRMIjjQTDYn+7blm2bt0GOjejtoESwwxc2tyVHcbCA
DqaBF4oVbhB2KhA5QoBfw9hNaBk2GgWq9wQnfUHAWUwj04Kzv+h/pRn7bB4v55lCjpxe2dL56w6Q
zslD1cKq9Q2M1li6eDPZ2LmaBJqxsBajdow+zoo86NM15Wfwo549+31KtvWCp2DhWMtuFJCDOD5B
GcxtVTDtdVN7XFxaxNahHr/cOGd96ZTrY7qLg6BUnD8kcQrkUoE36cV3/Ykvq3HHjabtp4KE+ytq
OICNJ57JBPKfsQ9rcHio188XkFAEaxA2QAadXcux0d2VwxAFeyL2Q+Cb3RQhUEz/akkOXDtBlfOK
Z03OdmQkrI+I2X2xR6yvGkXWjegQ6OVIEED7QSqLnQZwaW7jYsDlwJpJgtj4DGNLdOvqkkcU9Cpq
K2LxYVje/9K4MEFFMFEOByrT17sByoXF0A29UvXuVcxCwwfOKlTYYBw1tAZePEs7tczgPnXZLXLS
pdoAECKq3fh9SzbewWhAjN5N/Qeo3FS9xFzUqcwdyQ1l1Bwv55QGd3OmvVnZq79lKg9nVHaurQGa
7BkOdMSF7rS4ujtO6PqfxYfEl8eAjUhobGhzSaVVB/hWyem+UJMOI5kVBm1evu1AxlZc4x8bTBra
JcJJ0uzpH4D11EDq+j/mAFSCFB7/3PkZEODy30TFdY+YIG6mtovYWMzhDbFTXIEO4Wqpxb0OZ4uE
2egq4oTjSbI1SWA3HfqjAha7DpkMPTjfwMDM18oC57Gicx2Fgqfg7it2/XdQ+CjGy0qDRRdDvAaw
ks/NRcvjyMPs34dvI9cRAIDrgAUU9zwqIdlNFzS5TIaYvriQekcfAwHQGpIObakDiwWZTPq593ao
WS2NYN5Xt2pxGXk4FYrK/E4PdJHTHRI6GGaidYWVaM/WAkVE08LCjzzDWGBdP1TQaUjoMe3vCS1l
rXjLT+wfXpfheCP9bPdzF8xsnAmFc0OQzswsSfZNYa9xu3HA2jVdoxdN4arZ/RvQhykfhiONuPpD
lP6PslAzGGfpv26v1ujY/HYujnxnkwgmFpRd8lsa50HiKyN74MYsN1Dy6ctCFdjgDCNNnlLv1bx2
L6sf6OgPwuU3lPPuECASckzvQEkMfK0pgTyrxiucpGbg5HfWPa1HzLcdQQflRc+C4VvM/9c5ubhY
fGlYBd3mzkvoP1hzQD+K4KWIzoVuSA4iBiy2thj9bSAz/Gp+sno4/NBY8N7B4UXL3Q+oxMY5TKij
VFWBkAtHn+BkJeVWXjzHNi1XKY0BC8LTLbS6CLsVAhXbkoRlHgeNI3pZEfdTntaCxgOF0nGO8Q/X
QzfthlUoWcRNCgb50DfyfGf2BFGQjof7TFtCgRLfcpVtRCllWpgWeGWu64GRCOee7cNxVL0d5JzJ
3CFRr0stWTk4Opjd92B2+JmJ5FOXzlJy0kg5T74xNu5A12PiDR9oPmFhuPDgmekVH9cWtiSjnAdY
+RFsCpzH94h60dY0GgJNCLTgc0CrAc84td4A+Yl2kOXIoVozzIxkbZf1+8FCvdDW5dMM/E5qMbkC
mp+bxA2OiRQehnKtUTJ0l/KXlkHO39MYFImllmushkA6nri7K8qXJ+X0kZiTO+UIhEOzFkoNJQuc
/F0GmRdT29IZGwB45+dsWmG1/hgKcprBJ7IVkSLuCiaqZbxcehUdjpK3qIaEHPeStkbmu/Mc67DJ
NEnOf7TelCIxEDfpNZxaw2JWVlkFtsgymjeQYEOzr6KFBj69lAWZysvMhteiAzwbHXo65opDtQ5c
dkpybKnZPDK8+ZR/BVk3NRQah5a4nEMhlIQw7rS6+V9MQDUny1twFLPLfv7k/mRq2FJCbq5lqPfE
HeUHXKxfzW5ebJunR6gCN5kCoXZMynL5JU3a6P0QpkBGYJUHDASNFEbBuQkE/YHrMfFQSD4NXTE5
ITQFP685hRvhFP5rYt2esUr1FeEExeaX0htWavNGyouYGFeT08eoyz2TUgMmGbWQsu1UYHj7qwsc
MUmejiQhLzXYp+zSCkcDMcDHUZxYnVWL55rRPfYsnnrq7SXA4hNj+SwXiF73Yq9LY5RmGeik2bnK
7egI2SVw4AGdqD105CbquyU4bHyD4Z8nEG/mSSGvPPXeV6hbRRr0UNr0HMJ5NRu53GeVqKkpdnTZ
oCMZxiXvejzYOPvUE18g+5rbqYXy8UBUhmd8OuzLHa7IyrsFrTawKMUkmceecCcZnM2GqDx7mhfT
2m+o5IJV7axC0mYn8BG4NcBoK4EPYWbdOrnDLS7w5nwu8phcWeht1UkXlV3JGxn653CoLoyAU15l
IjLaptsT34SINWzTvoHA9RS0M4b02d6zSumtvLVhzbQb3GF1HMJNtZ6rf+kZLFHYNrLYgQiLHaDr
fKClmPcHCsxco0zUV+Sq7dyDh0cFmJQEmQIBSSXdZjasHQIcgwZShYZtevhH0E92VklMZxKDpM//
ZT0L5U2lYwXUqAeDo/WLsebL3obbnz/XgqLfry7Bz030TwvfRaYiraFQpeauA2d2oA/FeUDygAiI
FQM99MKeQ2uzs77E/qFCTFtjOvD5bWbs5tewg5nAPtTpWto4Nj+ygbvSQX880yQTXgTcDQciFrRK
WKa61edwktQ5eZ/qe/rO0ceHNs7DJj/KP7jB0D9R829kldZXCBGbaJVMCCZUUsqGnPx7RcaSar4I
55UVpKSbMrXdW1klr7oiRazG+xUYvU4mNDeDhfTr9IbMFgYF5Wd+eQCZMpeQeJ+xrO9CvwysNFFU
ahLGDKcP1DNbtD116PVOftZ44pbAO8asfcAMhbM3Q3Gy6AAb93HN5qchwNB5OxwJVkEmjFWPDOsi
kyr1HUMnxiFeZClogkcZXJ/YUgRL0gBjiigs3LxknK9nuRJ2+nKxuSf00paspSeL0rxWMGO3Xjka
luYFzCL8E+dh4HZ8nDGoxFD9xz2Tc5GyCaOrH18a2DkBhpfs+1V1xdvlqo+bVdRqQcJqezK4aWVB
6k1K3XZUxEmZxb3tRZKbxCS2wJdpD2NnA1d65+nh3A/hs23LukKtEO4ftSNCvffcEJ/+z6FbVWR1
FauE060AoC84hTkhQMXUUHsK2bGIVbJ9J3oX+IzrhT5ow+BLtRqetCS/vrPhFBUT+0n+aflIlUO1
24XQc6W5vP5/f8FcmXj2Df7jBcEvLSLMc8wWS9J5wUjDOIuaJxovZSyjPpnyCHmHoqVdhblVNEnV
t0neGOurwPs4p3V5oQ+My0p6ZwVS70h+RJL1icj/7hPBn3p4XkRNeGTl5cl0uO2+PgScL3tCgt4q
CJTHS+4ujurBjI0z1X4uuM3WWRx8IqYeA972cBUyJg84fh/rsnuM64DuBNBX4Cb9AjuBZysW4BDy
D3xXt+/6BMeMgpNS8FP3zwL0s0w1nkACqhyIL8OweuZ7SFaHiOztRibS+igZZGvVqy73jSTXHBr/
9sgj/zDpx7dBsiuAjXIwmU06kSSTyuBBQzdWvvg+E9jitEURWkGv5ukNUftoTLJ1EyvxRE8UMhO5
8SQ/rjZ/UQotEmOelBgGJAO+EWk+BfPVKAamhf2dvEW3sblPaG+Jj+3Y7M4mkfMNY/SdQKiaxAlK
eKnh5xK0Kz4rosG0cltwlCzYES2zk1kTCVPKZUlBA3NGJgsAU2krb3gaYnEmO5ZBciMEZJP/3KwY
7AghmN+0bWCV1cfwSM+sMyZnIiU7nmhYiKxDO9vbTAdDeITToA5ezSYK/MtihU3+D0R0PZ1nbdsV
riZXnieAwg0SdQM/bK1Q5Kax7N/isYW4s1wCXoenzgpDjBi9Js/0whQ1muPZhyOpuXaurxQLenKh
4GxaqTnblaCbhyeX4qHlmSrafJXZgZ4owAEfQGj37foffsp4JFHPjcB0NuWq7xvIqlp43jJ3Z/sZ
WZkgSqG5p/aL5+yFrXChOUIMPpdwtax39qdjO4NBHPeD7Px61rjoN5Gh2RdMghfhnlcyJoCIKTIN
BFamrbNpDHyfb16tmzm4rH2dO7isNDttirc7ql4k3OYc4ST1eHeSji/3+FDeDCyYqjThPGhW069r
rs6OhkUCBNpgr2WCn4Ixtx3NfUs0MtUqluw7RmHRq4beM+M0jyu6GfIKLfIfzF6hZLG+t0L8xSJo
JVlqJ2C6xDv6dAEQgx9o9FklHZ9zA+JLD4e++/Eez4HZCm8ig/916TnKz6fkbf8qKwbY9/4EFBro
qvAWKO9NMVuq1TSD2HhDn+9RipA1cYYSqu3pJH48W844YvAVtGAz9lZcvjOGOJvm23e8CrSu15/u
hWHbQPeHVCmPx+4mJysIH1dKP71Q6H4bfx/uMtks6yHqbNCnuj/sGoA0phs6QfSafPYW8KH/1ckD
pzeXxzfmtVgyHqfW8+XZ81jOi/9jbFFenuRvTeN+4BNujpeQPtGtCRYlcKhjbo+YNcKqi/ehEj+0
i6Lkh2FubRPbSrqI0744thbwEXS5AsknJtYGbZZccHNrQ1tdoD83ddJUhx9MeEN5utlNfPuKKlVN
Pf8JgjxS1OnRxwGCkUazPkxFbWBqkWbZZg8Dlj/BB135S411ov3h1MxEsibRGZslb4Ipsr5P7zTM
lJeC62aOYc5iCXJabBLQZV2m9ZbkdOxGnAI1dTV9AK+SHIDv+YM/tEuSAf6748aKsAQPKbEwAYiF
fP5UlGwRL2qA14gquY9oWVKhJsg9LIYMD93YWCxGPT84+RaHCYaMeSK+sO2yKMcjFFN0vh7mgQ5S
Q0k23emKMEadpH3h3XM6B3Eh4uJ+yv87FF1yyBshBB4SbWqwwlyQ7AG4985Ebiw8XPtzuczEtNbo
23xxXNQ4qv4Pn4kL3MKunEYDe7/iXUVckWfoQRFlKUAN8bpLHDVXriSZilEMaH6mF/sVjZbXDLOT
nfoIIIFaNQF7bCU1RZc5OkkGCSm+hpgU0mHk8MgglRzyt0GWdNna/kVPQ4/K5aTSrco0BMtk6hOM
WITdUBVyjv7qX7HNENEtEKlo/bl1135u3E/luGeuTiBqFWEHMwyIXj4UpoFDvyP4aMWbJx/aAN0N
nz/A6FHhj9WMK9kBDPApk21e2NGx1qbFuT8QSG5o5rICelrvzNLfWT6fkHxJ58IToKEFSFqUKIdc
saft6J1mV80InGUjgA8Yvd4t4sml/ZgiBVrfzsJ7ygFr71wwpH+8jTfNP16XmODPKX3+pVEwstZG
r64J8UIsANIol99gw15zBnTiivQ52TaN3f+zsF8w3SA5EUOKeYZ9eUdfuN8+TCRxWlxJ+iHtaCtg
RdWFdhfcqf3LdTpopsQSqsfGHCgvgDJXU8R6wHwRRbjARc3P62Aj3X/lzMdCj415era/tetwXERv
CaJwlMU/QF2bmqtc7HN6vWV7ZWHwFWN2rWLCGG2hYSTqcsb6qXYfTss9qYRg25z3U3xAfm3JMMaT
wbu6MfN2CAjSXe34MTk7E3UDhdWJXka1wZPHQzaugHCQ1DdTdTCGsUDRDeKBHAjJuo1zC/WpcDvq
MNXxn+szSQCEevfY6VN7OlP4FPnIE45kI9FkLFnqgoE7KNFA02Ao+2pVFRGG4QBzumzkXl+US9g7
9DsWQiLi71E5bG+TSIekWcQILXk20EnsmJcJdYR47/SiP/w7Guwk5uTWvyyb8bZDI2DYRxbliTJb
mlEy6fzWnNau6ciQdxIJDIZ4Tf8eSsBgnxlIFEH9bz2sA7aCTCGkzBmQCXYQY4I888oG8hxQkauh
Irys3An0g2wL6Z/p34Yz+/JQqMUahRG56RIapmHtCzJeFt2KJZLkfKWIov/tn6D07YNPIQdwVdry
bqVoP4i7VB8wlbvGP5fv+hhCyABKp34DTXR5NB1GCnttD/m5u1Cl2FE52VrXBOLTAmpAsQwQyuZ2
eW3dgRZu7GxhSB3d2/cLIaSLR0NVc5Fs6ipHanVKtJV77F597dNzGDJ5iklJoslPG97iecAUvV4e
WfdCxkwXq2aXrY7VB8mJiiINdc3vNtcwu1LlEryDop/jgKT8TLANGJZG9+yDASP3h7hcqBaycWuk
eh91gmwgvIFgoFS3EvGZpBJF1vyDhwsD2y7w996MFzkngPgJbCHdZYYooafY8UGTDE02y4BsWhMh
21W2wDuJMEumeFLAaKi29q93svJ1wPZIRj/sFOFwylsiNVEUlIwbeD+18o1gJew++BA6iiUmSNua
iaOZEb7i9F3Ti6x/+kIdfakuw/OJ4LlFQ0hEZgP9+R2Aa8yZKA7kGoUS/TZHbGFncuCNbReuUF3k
k4HzsPK8Hog99qzz91lC9dLpldHbv0yuSUhOWvwVOVc12hOtTBVbfFpvfKLqXuojp1Z2dMLsIyRq
7VrARd4R7XW0V2Br0OA+5icLqUewdDM3ujoVvDceujv1YJqptNfe/Y4DWRN71AtpfUS0BJVKrbf7
AHeuVYAi335d/MCrX4OD9lil+iHcofRs1z15INIlbfx35fnKGv8aI1v/Y8BszhF2iQ2S4PW84QgO
W6gIM8uuXOKQ6dZEosLPgPBeBVIjRhLFvsII5lnV5raOc0H6Dg6CUIteGZs7+qe65G4g5xkKliJk
J51Ce7QtoszPDPHsZWOG7wfy1GnloiUVEC5qfQdCoysRED7X8EmxlNyawuMGSULa2cyR7mVE1KvM
a8PXb4keYP3wtYD/ExD7dScwo7D79xpEP2YKNBuT6cj5HbaVlmR1Sm8dVzg7YVBIKwNFDsgoSSju
BTx+5rQcrWiF7aHpjrP5yDbazP9TTzakw6rehgb3+lhuklrfvJfZ5EnMkgc/IDUZ9ouhgKUxS5/W
W/KyM/WY/mu5mwrJWreS7a7iJUG/VSxSYi67l3Xg09YcFDqGSosM2T+hnwgWKKhosyQyKeHyTeOV
BNTkZMlsaF79BsaoAle07o+T4vjw+QTKYx1DfA0HWLASYrr1j+4JV8b0QOCxnvOm0Zb9/zgrtsUn
88mKejzflJJuJZpZUQ2qY5rmoF7blg4BMhh5bcwKWpmYoVsqd/njVVgukiaY6l5CbN0N8YcMJCgl
+/G3ItTlqYjwfiMUbgRpHKC7dyR1UPYepBbwxnXzvpgpYFXzZxRO7SpHFX3nxdyf1k/sDw+j3RYi
dgNSKQkhY/dv8hfUv78xqt05pnAqiFMmoYhYOZj+4Y9CkoXpLjUE7f9x3I3FUG8noidx2JhfIfLG
j+HiMB2crKfU3ATYLLAjQP1vOkyQ6yL8aHvGAr5dEQjn5lMTCAq89e/bshxSSWPTRPtut+aWOd+W
XNvgMIrOtXlgA7IfHj2WiHsg4qr6ZfGgtexUiuKFjdxoV80z/+jMoL+GvZ4S+geCa39Aq3qs0UV4
ezBnojYGK1MIsaTkTgQ8jlFqj0de6p4Js4yGwNZbrYKJClCUo0pICuOcl6BM3xiim1Jcuv/+VBDs
zZoTCDFw90hGSnAppYWizQM+UxHtEkNYtRXLMiIRiVZzzObumScYNhM8ajPaFwR9DAIjucxQPfLh
XFmwKUJtEN4a+CZh/6taXzGZWJ/grXbcLctn4zj5184tDr9wENviV/+3s4tFzv0j3DM0CIwNBYoQ
C3YhHX8yRFoQBVhftbZS8OTGexMsV0q7y/eXngJa3rVgbZEcOx9OaDC+ewephcK7oNu/By8NRqCD
vKETuewsxClJyz7mssXe36TxdJGlna0ZWiEumjCZZqAebi0M8uLEoJ5keteeBXS/JOBU6ksFuG/G
9MDY2A3Au9ri19tw/GfTYks0U5n+JJLm7AVnkziCcUUEiJ517H+lcqYPeHMY54JnX0mzevZBHL9R
vISjkkiATmm07RoZ5uJSWv4QW7JYmEcrtkzi1INySiGIerGIfTleiHCHCJGt2ytDJm1J0gTypaFJ
y0EoErpJ2equmreF5q/xg1r2r+u7bzTB1dCLAiaQNDX5No1nhL1Itl5+nK/nAwQO5BRrddE7JbkB
LnxYuq3mNTZNfcPY1gWzIHJzndilyy4HUhjpRNlj4JBbL3NXTNRaRl4bUY3vU6S7qrE/q8T4UX9Q
GF3hxO8I7rJK3/faM+D2bRmml4weTVIRLiPtDgP0FvRVMVYxK2jCbDtMjHtXUa5vpAY6iUXvuWXk
o69zkF01IfZc1na2Kne3F5Pl/JkIRCPhE2A2kFCCck/I/VWf0iKAI3vJX/y2HBrvrK87th7jPzlj
x7c2T3cbSv47GSb0aFzj6DfSN6clLl5Gb1LzrRgd4TmnjRnXkXpsNXriMiRt0jXbRvh7rgNlNkqm
y/OHgqMrEhKhGrDt6DuhvQX+uF/RFjaKfpOyuwJbUExpX7Jj4cHwTsfGN3Tak5L0IJq4QkAHMLR6
nPuZOEgruxcVkkpy58Sfw+dIHmJtDwF9T9mToMpVz7MIeQIqgwNJZDXQj8d9ECLa/C+Iae6z3940
0Lpj1giRhRxzhnlQNUhyuDxYTGLDEi0ViwCOYxl7PUtT/J7Nf4ZUwExjKFlb44pVLyAlvIpvFE1w
qTgvfsiJJAoC5dHMq2z7HhPjjCFP8MVeC2O5F/JKE61PIA28hcnxd15/goOYhNtEoBKRQuIc1zlf
UdagLngjo0mSzub1rzJ/25QiqZKnlGeK51dp6lciRY7YOV5FhzKLgj8tPO3czDAfi0G9El7YFqE1
zRniGdsL1sACxDvwJrX0ZE5LqsQsbS6465DtrMVtkSks0W4KHp4JnbUuaWv6K4XRB/rP0GFrRh53
lk0BEWAP957LdRgCt4mjnpwOzZXbAJSqglWzcJr7LEISWfvMQJcXZABs7y7pMuZjAZDFphuqr+UD
CMtYkq8fycg0jJKebzBu3FSDOoxl6Sd0L+0e9hS4jeSOrl1+RAD7Hh0uiPXX2HIX/8bAxn2s70Q8
LNiEH1iD13IAEx/RDmRMjymaUfcXfChRNCs4NjkU4CNTPn8IpbpAX579osCN3cwtN52kU5FXLDnk
WjLtJ+6MofkTpIP5Xd9NbzwPSL3VqhIgEl7jsUq+x+mhIGH1m22riN8kC4QpUSDRdhbgvjIZ4H2a
ixFJ0S1+QfpWtxCU42omkhPJ0uGenhZQQVp8mU9swCFK8Mg+/AkkOH3LxjCjaR2LixJtoOiXFRLl
WChwQxQFk8kloFHS0FQEw7YjNmMSxToSIhb9aNExPIMZ+dTKwWaO6P5iV0npkZ152Cnigh8lrhJ/
DYedMtBYzVyDo+A3v+Uba28Jt/ohBIOpvmX+HlCFmoQGCsG9GMh7Es5tbZKS4fjAHUbbBWNE/l/L
LLat6I+rQby2xDA1RsJyBCSrQ9VIQiy0jCbmHr3ClzrzHYbVtMvBrXs94HjyMSe1Is0uV2isrOt5
qkudiHlLwn5jtKi1cemloeD7ZxUlOXl+iayMCK4/14xCcCIXWWfm+vWJGlaYPTWaUN3CyQo7eETl
GfklLyMzs58Lw74/90KHqP0zkSnagcPI8KISZpOpSXrg3HqfBKolk9V4sySyhpKzSpmCHjHqzccc
yyopYifLG2POzZYuDN1ZSjDwzAfZMvoPh0m5CGAAtbWStiuax5fcpLQ3DjEHfb5/G9P+RZMU00ZL
fBL7EyyH0yO5oGJgdq4sU3QORa///g3/GHZKheltTp9FzqwpqnH7u9FJfirKyVAOaWzZeRDbCrAg
eIU5PKgwsAJGyguIKaLlWmVrGLEQHGhxkIAoHVnXwTojc6Z8HeTvh3D5z4eTvPlcFUj5nfqRDKqR
1yJZlLlgz0TQBzqYvi3eUES2Po5Uk2Z2BynChHaAgY8F4+imo/T9GKnOZHZBZMB5DS9d/98kMYuN
oI3CR6bajq6REJrGsMXkXaJYBXJb8S9YLYU530P22pmU+Ly/rJY03J3YcWuFKT/j09Z/D+6WqXPC
/yeMQLH7k0hmbgwfcp01PSOnaAfVQ9I4QRQbrtxfCAbDDRihdHJwcL4vzh6ch7ZjVIEjLCYqUcL/
QZc8hiKAo7/4otIJWWeKZKpFMmnjM1AxIRklZGFN0rvAZKx1biLRAmvNxZAF8S958FGzpF5MJBeR
qoo5hmOF0bs6tN2xgm2a6/htbPplO3Lh3go45e0GTIpOmLPOc4lOXYRWxvGR8xnfUjtKvSQEEINZ
3Wqrp6DpMqdWbhCxogZaefpjXfKGFsF5DwGoiPP9IGeFyGpGwT1nHeaRFCoZtKtD6ggn25hcJ3Qj
z1mgFfnRSgnt//HJiws8L3VzUh6641dF2T8QCTHoQNm+NpyHQ/U6yduixk+wVZQbf90s3iHrtMgF
kSfMAGSozNgEh4dv/sId7UcwLLIdw7gRdZeVQEM4735iafJa4tRH59CWpLgXMU/vutfyk6SP8SZG
CLCRtI85JyL92QuT0BcsIGzhbJ9JOreBZ1hq4ioo9Wu9jJj7M9ZQtIpdrxvnV4aq75ADmjRCMfoM
yfWo4cfmTvIY/kG7tvKCRr9XpgnCIFm0apdwMEIcRM08dgj4z4COAU8vH1FwacQVOo4nKJBZ3zz2
dkMvvP0AxJye0hAciR51VkD4R/rmgAWVGSQfVEOMWVK9cemMmPwPJP754pGBSKIGZLIrrQkrZQ2q
qQ/5P9dgIeL6Ycu4r7064j5yHQVz/SB33VtWIS4GaoJuX8e2w4PULlfjrzIRrOq421aQy6OwxC/7
HBcxVVHkv/imRK/uXOd7xrbJ9P0qjioQdQ6UGgz2eYIQ5t102qS8TTNebeeKJjMDf2BgxsL2g9Uh
pXfms4AWf8UnRCYHcv/YRBljTvpejFWjx7M6t7XZHn710kliAYC3M3PfVH1EHhrN7WMv1pZ5yZHr
sJbSL9qeSIRzOc3GAwGE4lGAxqv5pt3rwWG2OGLc1p5P/uszrJiMPuEjw2SUSbb4gCYhEuEuRiwd
PJhVNdUFB1PizDVoQAKfEHnSP2R7AkknvgJAovhCWEM0OgOUNMsPYfQ2NALKWvzcAeDmWfF10/UL
/nsXAB3WowgQJtW5zUTP4m66cUReGl8VfPO7D8+BVDNmEYfcaE/lKJXKe9/IVydfupW53StC4I/E
4skTc5AdLwTIojGmzMGMWT+H3wI5E8AGPEvTWTYuoicqbngX7Vic6b7wQd8gart06k9PdXz6Nsm6
Q92C8P9GHJqUTNrY63Z6xKtyZieeb69Atcgt8E8aev8hRtliKoxIMYG7+HFMh0jECK93i0j5v4Hw
rXnXDYo9KBhLqzIzy97nMIR3r8QQ4qj5/D07hcBXDDYGyCucY2B66TE5OisUxHr7EskDbwf9ADdZ
l+66g52sMTsLEUWZLjMdwpDE0K3LnJOLCMjVF4nd0+Wg8GA6F3VXE1JwZVGKEjsZ6nqiSizzZNuX
w2Edq5juJz91f1Cz4cu3kyutteOFOBg4iqZwpHne2iU6RUIJjK25xril3VBQ9AeAprZQRhtYFASJ
4uMMJiGIhSsOs2Mmb+OKyVvnv2TcC2pNZNlSpGHkHFH5dZ6HvzG7ct9lKhhfHKigJsRgRu4rdNLv
/UwZRXaEOpaNi8icLINP2KyxW9ZASYOPJqAxCS+Tre3fE+MnU+dqxowvlN5nMnmfPA5Jiol+EgfR
vNps9Wqj15YI9/K9Ax63L4CuNGZkBqbsAzw6qdaHT2QR8bald4U4tgIXeMmrctRa7vVURCCkQAYY
cq3f6F9Qj3WUZmVSMXy4bkiinkWcE0u5pQQIidlJLBRnJNa+FhLI7TbX50VLEFTzMRNlgMW0IX+w
t60wLoYnPSy+l8mB9EY7ZBQM+0YjnjTMqnxuAfWf2h4JiImuRrNze21bSsBtv9aCTfqx5usqOOnx
7CH5tc0LzfTHR+WTyj+jWdOok/oCalvr/QZhNZCEBT4t1O2N8uPL6xWX2fWm8cReiUIiq7HI8KgA
DiaOIV4J91oMVP+w/+27uTx3GlGApfpeNIEA2hmWWvAVNDaeFcgkv1MFHEb2wLQ34e+D+8dS8K+z
iAS7MAm0LZc5dCy/7KQzxl/6a1uZWCBf6xJoGbRt2EB+V8TOq8MXVNNyOR30heqO7t+6aPdtWUwn
A/KHg4LahWtPe/8H++wbusViSzH5zTcBVYlzAtCpelF4rDN8GZFrn0HO4i1eETMY2Tgjz+lkQ2Lb
C8KW5ua3ZBqBswlcq5l0qSwaNiuUSdkHfLA/M+k+zCeZEtKrPd8XSsk+/LE3RjtwJqqSYktvD7mH
YmTLWJRNUnrhs+peBL/iZX6zRvAHREw/BYyCJ/KrDrqX3Vk+a4UIOLbp7nxivj4/ACyxEaIopaRc
anCMke8FdVsHAnBPWDhLl5aQQfy5uaBKiOKrqWzkc7G8Zobez2/cJEZxgvyfpHH68k/Fm69UcWlW
B9VceOqgUOL+JHhHc06VF6RXYnvYmweXFTDjr7/IiV8aQHuSKqUCdEhCgr+G1fnpl78QiJA6IMGm
oLETvPU/GNlLJfh03Oz7GD3uGiBRO6tJLt8RazJgMtXI8lXHH0T1vbd1Eyd2j8dUl4c4+9tBzgkW
mgNTkzM0t2Lilh2ONQnTt+R62Hdi+7fJSoEYFZu499HoNOFMezh3rVquRbIamj0aP+UmzrfS/e7N
qXxY8NCxA75LUKBglFGpqXv1Iw3mig1oZjTCp+rcIEzfTUthEvrTZuxZsuMOlgGVZh6xfKGthlQG
HPiQOiGE0a6SFVhMBs29ex7naVl2foM9b63AcCy9B++agfgfBYDvu0nxqwS6mshqUur0e82A7mbk
mBKz26d+p0XZzOPIdxz1fY2ZX/fYvEyjA22BrduLavkuuacev6S4zHHYrZPEqQBxv5BFf0GHoiIz
JJtmzZ/QEihVeOMig3D9NvQCUoWX7vMlJknpcP0+1JDHAZw8OtLEtJ8/SdICSYvgTaYDOD5ojHNE
qmg3T5zhv6xIMeXSmMvRkHVQkF4U/Br6udUs2uOgRNLiJrWYGnSyOElqpKPm/66HRLQvEIylV/K2
ac4WRdrE24d4GDB/bPpHQe8z3M/hTFyg1pzQ8jWJKUmyxVercM40hmekZc9DxlGEClSIhXJ4gvD8
pJLuCAqYPn3CkAb5OHhXoS3Bj2IrE+Ca8IrgkNCYjhOCUDuuFlv/l1lDsj2qDzGZx6LCZ62dw8eZ
RFj8G2y8yf0YTd/Mw3Prkjt85sIcD3wdwoG9ao9lA3qBCd+tyDQDv6L2Vz1Az88FxxnYJ7nRL61e
UFTZ0QpkNknvPl2F+TegPsHan4o6JMrvcINOL5Jy0xwwm/TzTAWKIW8F/uy1oLz7CPN4BgYBQo4e
FxiHtVTOayw67JbTu3tQ7dDMN8/f3fEw/bGJ0tk+v8EvTAEDB07G0ggZKM8NMf5oVzJr5fq28l8z
JZc4+oa/lXbbkTPUORs70l7q9BDFxWVLDf7m6RWw0H2kk/ofZer4o8SDS2dyITSr+E27pic0CkkD
KYJgIaDYl9+pyZTDktI7OCxyHya/qCSbHlruAb29RgwsEEdTdRk/PWcCTGkmH/cwYZNNIo3SUiNe
vqWb5CLVvQc24dHAfvaGh98ftcyr4xIdgNik2XABwcQVkd5dpJ+6XpSPCywOT6wxgcG1govuiXqT
/tWZWqX+xWfSxJ/+15O3dzsM/hclOW4CkkqhyETjXqnaYgrxDJUKHdhn22UIhS205yw8I/hWX9bA
io+e0WIfRV4+2CTbVR5wmqxSaR3Nq0muZ1JPb1QQ9yAfaV2Zk5Ow6Vm/wjlbYH1uTD36eTzxzJKS
LPZfxNUbkTqQ/HXLoCQ09PaQIlLoQm+jn5i2kMxylzluaAh+ghRqO82CgeDI4wUqQRN37bjyd3kN
KdOUZF8Qpcecd+56c2MJqvBJ/LVGYobS0JWdWcWkzsQDgUmGJhaoz8Uqkc7446JqmSlEEzl86fXn
iOnjNRNebL6H0MpDbOusz4WpfOnUT79DNzcOA4EJOZNzWShPnumCoQ6ey8JIS8VPEQcEywPFes0f
UbVMtDe+jj2u9vK7ehMbjcRU5gCiRRgGnxAiroExY16TYA5FdKe/tVKiR+FWJnQUr6KH2HSqkvdB
YXdDntjg6mv/OMg+wcRkSwZ9YgI9YiQZ8JEq3TvSGrY4yTkgHjAWmOyQSV0Z2lwlt2fTZVyBuX2K
+8SQldJNS3/6FiEKrbi5vOj+VH4n2UlXosgSeP8AwV+eIEzBIoz++l5MlXbAclQ9QSA1bLKKxwGr
DMOnEWbTGFRyOkQyD3zyiD6n24QdrvTSqiiX6GU4pmxVf+5RaZK3bqIXIidIsYlpKLD1XjtB9hGv
h+X7BcAYBWU5ONMGV4v7kTiaY4DxKXxAykXRi5J9KDK7LoDEnLQwzZzc489K+kyDjW7PrkW5WKH5
F13z3MUfwasYb3fpS5o3dJ4eZFN7jBMMqoWASCno4Mf2I3CxRxxWIGIObMsTYjnG28+juhQrDZSo
CYeuL5mJJ+Dv9TXiOWd7ceMikjAxrHieVyf8aly5+9R0c8nyMbjfaL2ieJPOiJ9SKHnS5D7Ojzvk
SjNs9wjxnomNrXeWp1N+z45vx+nnO96stcWKr9Km6SSpkn19ypjkVJyH5chN2/h/kuVix0KBz4AM
QgMvSB6Av96qkA69qaVJiKsY8JQIbWquZrLYzQc23UjeLjo1qEZC1go2HpPoXqcpAc3ZozGOkGqI
x09Qclk+h+oY4cRwoByE0vcfXPHjeuHmC+PH3YcXFfGbpnv5Vi52tUGCegK2SADNfqufDrswfbJ+
NjF+pZKCKMKCPkwq9bRdEfpJkHyAk5cUDwMNIaSEG19IxNAtAh8qlx6H49UYy9FZeKeGmUl9bPMh
1DosKyXEWpVCv0/Jm/gW4x+wUp3k7aeeYP84YoRjc6ERqAe+f55kI5IVCNKVo4ZmrkLVG4W4Jmih
v/YcFG5d/XmHJLp3L2oaUu/T11d3bxpZmLw4kuXk/j9xsNN7qKVfswf2kyUoIVLosT7KrF9M4mC0
LoBkCRNnhW/SnfjiZVVWJ7mS1TfWa/XhhcI2oo2E1IWOMUO6oJviIGtKKfsBW2P0WNjfphw1ZPhx
V8uLPk5fbFELcTO0wSteSdcSQkp6AaAhyPqAWvIHVaXJGONDQEk5oa6B9vznXEFhsbwJaDJbDZjU
3An/V5aKBVcZVrwmRGxkRnzYk8OcKX3P7AqQYYd6LLfjQmHMFcBdyFQABRWc9SZuxIvd7m0NSh2m
X09Zpuz4zGtikSgM4FHPeP/xQAwQbTGTso81dYf/MATT5S481zKtjTmDiNYr0UlqyTIzB8ghxjbo
aKAK4Mg8a+pqn3tl7tNuQXSKC/1PrvJ4Mu1EF0x1huCvbLiAPQtN5Xt6PPTY8gqjkVwwqrmlfsEb
PgosuAYouiMjt80UH/K4KN5KUOx3lIiJ8nOFPb+/tKakjT/+JWvhbJXUZSCh5QEnAMVliEHT5BBI
c3fawXmpo9EcijbewHtpUO1ubKkBD2A5BJ7qMUuImr/jvDfz2ihcd8pkGOAuAEwHIoPqZYB/X6va
sdmwowi4tNc7H3dwVK/uiE1Zcopd2CnSGolU4ggQQmrZACaR8iBmDY4gyNVNnGK7kIyF2GIpdZvI
d6TZDO5GvBAafLlCztTKa+MT8cSMjGAuHgTI9MWPjxPb3yQSe+hxmVj7DQuonEtINOYRvNyfGtCL
+ihPcKkcdCjE2PdzhtrK4JhVVAZ4q8NIvvbm7VHmonS5Hk+lZPojZ5cx4+StdtPGiGNnm+93Mr9y
0PviRQ4oqLuvr9HrP2o0PFeI6HWYk8SPn/Q7ZcW1P/QWfCvSYEO1mMY/xz0XjWl4hPEfn1cyIOyS
QgxfSLrx0ZVzYQ3aqExv6LTiskP0xIvdn4QRKNFWZQAjulCHyV6rv6qtJqosz5up1YaNLX+to28y
fTfmOiz3tZXL6qrbPAhJYnDzwTKDpoKS84nr6JIKsWxzvp3vSLAqX2HcNLpxWmRqBwvc0tAh2xoR
ervtuPyPxwR4ovPAg4XdJ5xIm60RVGlMJYi8bv9VEAXLOE2XEFPirACMPz0C2vBZ4ixHnVjNkMgC
k/ispDILde1FldHmq+GuB2vQEKmVkDkzZ5xlzg2h3vgQnNE9Mt+JRkAxGXGc263NZ5WeuTLwmy4z
uOU4WzTUg8HDFUhpNatHfUMpFTfVscTKGF0ZIiuJ9qwC9YXjs/q/DCvx5r9KnM2lbiixLpcaL1tf
5+0MrvkghJ/4M4yvjbhuhx48BlaZa66rKSXiWSxwE7C9A4DtKVaWFwFd68wf6NM+7+TlETJ4MV4z
Sy5Ou9tpwPTb937CXcWNgDCiYrgJyRfdvv/cpMsipBUUB5UY83FFGWv4UnQu306+t2tcg6DVILYH
QDGuzKGKhOFdHiAYKdR6EdWNgH3TJh0xOAObWq38Bi2fgG2yC36By3NUP4iY34DXY66YSgXKM9oM
tIJwxOAhfx4zfvZhYT5+xX7nDJ45uy3T2ASu56Z0d1/jlBJY8Z2frKbsTwadG1xeOPrb85fju69K
NWDCGAABdsA4MU8ik3cuyH0r8dFQhxhLpCReI2ALbBC9oWyP5TjTqVPkKzwZjYGkun+YMa/GHptS
JJpyAF8k1BWOQR2RC8Hms3L1kIWZaoFgCvaqxUXpEwplgPpgLoOn1xvTNDANjeE/ypaTnQGclxwi
QGw2a6qPvdhAAUSN+MENrF/0Fyrl/m246WhW3EU34fTpjFjX2jUPf8FjI/ejJZXqfk9V7vJFmaOA
wXiHDqksR1EYzREltDoLpQHKEdNVaId/7KzVUPrhX1xouvCL5Q/E/lNqubbkDhHJoxIvifOtJ5xm
wh2u9FLtd23iiISq0NeBsCxD944/tWtpUrJVA4k9BIb9yx0Y6GGTCJa1Kfqym985zJauk4u8AocM
P0fVP1sTTWTabITGHhtTKHchFNgeUUrYL6Lzhv9F/IOngF2H0dwOIKn952208qwz5EM9yhmWX7j3
fE4RQ7orW/wmg1h9PB3LYOGNdgO5s74OmqOJFbvnCLzJlVdbSCugARVKV0i2uwAFFClMpTQ01puA
nifwcAslCiqmsNAOK5tai40oIvyw0hDDuHKg9DhQzQ4dvYeMqPn7LUalJ65UP0yEM20CPuDtWrky
qLcoWRSEwpUU9uEVJT9HTVRGvMpY/s/oa3Z0msYbwNnyMF+nKbhTftz4A8WxKd2sdLfkKFRxNh6v
UsVdj3/Exb7pZJ+cLAgxhtv1hRYlZivsHezupQfMjAObNyCZrgf5avYUBuo8zeTvQMwvcd6ARHjf
n4tf4vT4FuTAs8z4vEWuDm3FDZDmiInekOW/02ry2qByKc2ZUYWqF9YHtxcmkiIU+EoCILTrjk97
huqPYtaIA0Vipbnk267ByT6pGFVaMg6/jFR6uBkrQbWfZO1wZdG37IEm/a9baSWnCOkCZ8b/Jt8K
hLQ1ssSGuXhq24ZhOFD3+biHbypVUEcwoPU2to4mZ2JxXZqVOT8JxF95iSiJxNRto3i/cZCWt/7v
+bWvaEEwNyG/m8yYv2MfkWWdDH1p+zyTdUhl1bHam8pasjgYk7mXU2dQBMDWUavvb7FHnJgMoeT4
hkLj5J3GSpA3gi9iNfv36KEj8Qo4ieAceDMyWuwOGfxPu15O6GlaN+A2D1hwRQvo5panEV/8mo6I
gWj7ijv+YLYApQGdqs/j3+uAFviRsRujKKyUxVNRUQTX/iwymleaJJeV6GXdm7mHoZYiBDrvs8jH
PzM2egGSHDCiOxlNL+UExZep58wm0bB5hLBkxhJ6A9AWKqJT0c80p737GMO7AexE0wnUpiXhP4iT
i5NV/m6da8+F5rrGj8BX3gzr85MugJYIUk06ItfF6yv6NuXg+Q7oZcJGwYWA8hHvf8++puKa0Mw8
9RW8T2Gan5QNvyx3zKDK4xCJ307ujdkMh49jxi9lRf7se7QiL+G5rHtcMTIwX8DDcGHrvGbQOYHd
Aa4PFk6iBGV3ceOGXvFyfehQhecSPogFhH91OVBYzkfqL6V8XfZt3QKcfYcVp4JWDyyVNq3oYJi9
voHTLzR3TCNVEXFNx45ulg3TU8FiNDS67LwglSIq9KvcPc7mNHOEwtAEKG1a0+vuMcYmqIQqNoDS
im/uihbZ/P1wFgv23Z8TW9rS+9H3hXRUjqinuOOnZYIivdqjLTXq+LprTa/CbAUZQxrMaRZVyTuq
IVxKShqKP3UXmaIChc/8H07WpxC3xq7tZpKV7G0v83MfF9SjbO1tmKkWpGO9fxUJfdfm9hnVnaxu
LnUcUr5UKZjReJwZYrpl/H8+m7hb/CfI4T1BTmvVC7x5SkLjlfniCp1qzvtlkJkYVaGra8ZJidiV
Vuk7cm3pkfeeDomIlJeYC/3d49ydYVkwI9grZfistWCAaJIAeBWSOeyJqmkMX/2m4nj1cbxiYSq6
7GLF4LVBH1eeP9Fg9WuzrqzU4sXE2/SKppoyTMyxeJsoHxmR0hAf7CCrvbiGyzTY4tAXptLx4sqX
DdvEQ5R2kI1an0ufJ8UuooR/HXirGccX3/7SoMjgTGhRa/P0FIeX2Y8qQb6DnOlhKIKsAw2fKZa9
mcmkx1qSPpovjfhC/3SVk/c0AXITYTzN6m8GDGQz+dk38Yahq0mqqU1jqHoHnTIV4ZLIPPcB8Eri
hnELk1TMcDhSrvlvgxakCX1PGkGHsyayOJEjCwgtH3fmc9fQ8PHSzPPgwnt+a22AcD+8Q2PIkWvO
bka+SHEv6WJHZCfAS945HVajNQpOb7pavsmPQOQO5XhO400SOccoTNkV/lkKw89J837SQsGqrOw8
T+qf88PVoD5uH8oRuMC4XhEZHngzIvOqkifuB9eal5upAkOcSeYQuh/+KK/6R5xtFdPDnHxIBPgG
rWLtazFQI0+sCMAdRvo9CifoSGITCFFRLyZAwoM4SvVAA8L64ht0P0CuIh/Qe28arRplv+ZGXPaC
hNbDtC5rpMZGUVcTQGIfAC5oj+9SvxDL3iuAGX2omt0sNnBvaLDFYsDddYOl/u/fzkBWN3/+QLwH
W/YlDfMnFX0swtUfJ9s7yNIzdjcwvChitTVgBVR+Q+n/LIzQhjCY4tGCrFfC0pOg4d0GnUvicOph
JSgSEsACBvjfqa7h/GIxuwh9IsfXRVx8qaBz8uKPifSwsseK8YG+IdksuCIkr/dqMQWEhUJT0Bf1
4NyhZCiFc+geTMj6ihqbVdH0qUtP+uSvVTiRDGMiM7v9wvMm+Ad1BG4bXo7n+FahgzV4Swfztnn0
NPqggiYgVk2ycLWReVpagyx9Rv9k/LvWM9vr79yGr2XMdQORnd5MZpCAZHT9xq23vFz0fYELeXE/
Xj2ZsUL647uHPs5FeOC6/AyKx5j1j6rxl3Se2DJbE00tYNrDgfc2XVbPK/XN9C4GQdWFGjcfHdoZ
O79q3g+G29v3i7MTuX9GnMrqi+zVCVbaG9gzcW5xdL+v86kwGPX0Rv804IDSdb0z1br3Uvc2aEb/
U2zYm5vy9xF8hupGwJfH7TJXpc3DxkODmbZP2tRWRIJDVvrUnB1hBpoa78hCOFVlURDWco/k6S0X
G12X68zmYCWLlPxjF1LQXyJGOkuSA7Tnd2+6EefXHHhTqouyScADcKDQ1SUYQcZfdGLNocAE97O2
repD53vy+KxNbCti5CU8r+cqcq1XyrIlpxDfsEDQFcsduecplriMDzBPogbb8tKcpJCKIexCkUiA
+EiWSNILDiZRbeeIWCNjSGzs4JaoJtr/8vH65PmM+R6BoOjQ5PsoRYbS5dpabkqQivCwTsjMEf2j
NaCgYRsoeoN+M3YbeMq0gzPoaJpCmw7J0YeDMjWMTnK2E3pqJC1LDXPYsTTr7p+roH+Wm0G2XBwn
3ASBxDqpVaHeMfjzFR3fPlshFtFL0HFn8KCnGuMWOWPUgX3/YvevuIo5Jo1/FBbO2mfRYZW5y2d/
EVKplc8aPLCRsSIjDpkhZNKfzSX2h3Kd7hEZ+FH09iejOLIxUV6MyBYXQwEN9b/eJnkskfFLAOkL
+Ezygv5Nd/gLHv+fOk3EZdneFk2SxBmq10tLiE3aoTG7LeiYlvM7Pm+lbbqvlos7JV458UxfzuT7
4qQoAF5dPGFl3AmwYPbyZ/NovUykJCvzGXlujh9Rus6lrBMpNLWqARF/fjGFQZ6zuVlkRvo0ccwM
SfVFcjeNVAXXeNbcaVQjcE6BV6/kMgAXd7Ttos8ibaSjs9GU8sgW28vR83dyAbau77hIg5VazQst
YJmrmnVoI0AB6Pt/+Tegmav0v9yNxt0mxgWh7PsWqMqSDKrKqp5RjS/r/N8M1ZOGmSbHF9xsc9I1
ITaCe600xRJmgVhxrYAOPw9a49C5BvgmOGRZL35vLHqaRuG5y2k5Sikahwjlro7Pdwka9Y0wUkrG
PkDTKG/fNr6yYt7vogH+Foae+jMSQcXjWKhVE9MsunYl0PZIj/czhTzMdlB2B0wbLCWaNzafUFjk
32DtkAPtErWIL4caM1fNwbNR+PmKTneDIt36Zht3Al0v7qsAZ8iC8CHVCI4zfUutY70NJug0iW85
tZECpUEkImsugPok33ijyzvTSOAkX1nuWnU/G9iwYF+wo0tb/LsKAm+pA9Sdvd9WnqRCt7s+WUqs
TMiLqUSnsNJMjZ0jzb9AsM4g7jPN9ZTIv8TfFHx3cUkwIIrVSwhGKCJjvTOZQzOaYEaKv/0k5p3r
x1eTTjmEznfFqrf5kjJ6WpJo8uHCzMZui017FEro8QCB27rwcU+DmMQF+MHlupsTXb/7mUQZWYvW
DIP5PKm1fi7nz4175Jzbs6hOl9J0tRP2dz9BR+Yl/VEqgFOzoX68rxnRtVvLaNKfFvbkQU5qxcJJ
xj9Wu+ACUYl/hm0MfM7rYjataOU3FoXq24aLpR8H4qa3Fx9ktkg9SzFkYgrclB6ByQJ+4lyqbLT4
cusfF8GwzoDWsJ7zZoibHttenPf1CpDLq1qD3KXntSdXJf1BzaKD1bbAa1Gwq55sOtEYd0Uda6os
ES8K8rs58wLtcojdROI4syTcP21FTbQrpGsjAruwFlEJYXGonJljHoMr038vFEncKOE8JmCQNH8V
dQOMlqL8t6ecQn2hyP0iQkxyZzVqMd8C1qRRV9PpBx6ct9O12YXrrjD7WD6CWv5ZMMa88GPksNk9
4qE0BckXyqgrG/kjxHGaN84SpnBOl/XallD9vaaQAp7sRsUrL1U9pwVTUnrvqpVr28yE3Egxbm3k
i4vhVGuIsW+8CGsNfN/pplKcFi1oytsToUmMQEhsqZ3lo/lMYVTDJQQYJ/APgV62ykr8rGFBeL4V
iIZm6Sa7ztQXC22r5Up4+2YbhTK8l+JCYPIG6mQqJlGhzzQxrSOqnUYJ05tCJTvMhYUHJx0+OPH4
b3UhCzvOt456r81xX0skPZfVNZDldNAEuUAFCdbEZfsfPRFbzlFX7JdDnME3B6nK4SNzcRfPE1E2
VkCRs/4s5QpCOmeN+tHEzAIGScqx8BAI6PrfTP6t2nOar876cmzZYDheQklUvUi87T09oQHcqZxS
yGcUG/KlNc8SAzvAtb/TelfCZrFMbnFFNbEtENgQCC/hJownVJvA44lk0aazBya5wJ+oOwIIwXcQ
DGxLYmQSX4iuh22BvnbccfOM+XycNjJ1kKx24DINHFLlr5l4qNPzcGykw+Q1p/Nf4ZR0mum01HR9
P4MyNMh7NtnKz0dZ8sBbJzM/+4Uyb119bBwB30BOKCzg7EM8VmOxGtQkFEu3Uitx9QaCFFzNrdq2
vxRUBRZkWFICbPEYSG7zQhNzUGL0zx+YbOLMrrSLaOSo+HvZYxMLDuYe18bkP6Usq43hg5895R7k
wbmvri3KX09M89EpaPtSltE+p5T8gQRUe5V5BNZI17CbK4VfyyVEQxtiJTOTajomL92rypCWnc+3
+QhJWoiMpRK1cFRmNsjt9g7OGaerIYdjxnclSIYfzwbXzWLK1w3PfDjD8w/jJVbG+nFcQ4c/XZ6c
kPx6AY/iKGf+oGzz9tqyUFGZUCwZbaG1UXT6X24Mxxr5pQ2I/pyAQLdpntq+cbXg/B5cKndrW08m
R4BQPNooNs9E2sO2eEEsgSvhD32w1cd9NdbBHo34Kb/aC9QH1MEHTwSXZBZUnk10YMTSOvxRTjJ0
El5PbTVfIlLqce1fiRqlLrndWAlNjLM+m2LJLuAY03aAFUVxlvK/WmStVTJ6H18sBj5GWGGKeY2v
6wx2RxC8Xjr3JrSdXPCWPgYIsfDf02/8l79l+suiV9I2/SGvJ6TN+cZudgETqIPX4jGyRETK763M
QGfiiB9RtYJz/xgLAZyL5+h6L9fkjW9LhH9QJ10yJyvuhafLwOgPKqkI9NMo4xXw9YpYk42u++4E
2/vHdcHo27GECniYr6mDGZH9WJGq062l6W1MczniYPQMYhNeE8uATI/8KcnN7is51lexwnzSFo18
6MYpTDejyafbwJbR3et9QaDeteeQfwmKX7IGnpj+qoK0EsCOCPpyoFru8zicSgH0QDWGRKpeUOUL
3wWkNP85JGi0op6ykmVGnwQ8Ac1SkLWoWVHSyYBg+QvLA6Y9Pv1oyme7Uc8dxnCaXrYWjL3jjc0Q
0LW69l0cxJCIk+8Uk1CDWnMx0rdCecGhh4m0kE+yGCB9LfpwE0vCjH9o916kdkf4AljhlzagNyoY
/A8Aia1EIX7EbrRfeISN47UicQOrymxDnVYPuUlnAWEeLEPPUutgY32t3PMABWvV+ScAORSnYB6A
/HqyegDufHHtOCDjJFoqymNg0L6/A/fJi/fD1BWM9BcXDRAivg57FEJNmjhs+O7xY0uRHucQfQh7
kyp/pn43Kfg5t9xHGZNtiBiT+PWCbbgHFoOzAZlmDdPP2DZlLb/SK68JzQEA/f3IXYPngBjhhHDp
oS+mCCxbv5qkCM1SQdyXrIwmh+4C6xnV2hNBa8eolrAAh/R/JfhICNtod9zChbhB4eCyTrz3UiOi
vNOAF/Chm9gHr4wRBKHMk8KD4VaTh6EG3mw1CEKaE2dk5nIFAU064oE1ixM68G7YfqR5WCGaMjZJ
iAu3Qnxn4d8aT1gYgXx1nJq/zVJ/pw/qRsntiEASVQB0cheBwfPwnkRZfgLA68WbDClDxqYamYBK
HAdb9rK9yJFDglgdSKBdzkIP6tBoyl6aA2QDiOnmYu+JdT9yp7tfhhVz+KHSpImnTnPKn6eDJhfj
ww+gPiKwhk7yfLvkZFskTB87NmiL90dopexjANVAQaTCI5O36skCNjjMO7SgBmNSUC/dpfcPdb/m
A+3Aj2Pup+/CfH5sP7TWvOhW7zhmJ5+g3jVlgMBcKwIA9rvjh/L4ERzoakU3QZf0z1ajj1tfK1qx
RzurhAlJ8bOVdvM9Qdbs8DwHgm0+Z7f1bpjlZb+K5VDY0yx4XH9eJ3cJV5J9qWqf/25np2YWNvg7
QJC515Vq+HyuX9GHQOxKmW7Mr+yyNUnnS2kEt6CMtTqQPRohb5xef3qMpTLV6Jks39d3JY+AFJqM
XDojCTEMyWtf4AgWKbhvXNfw831UvUok2NFBj82Z9KMxA3GfdiPUZH/5WMuNCKTZ8MozDTphk9Z1
gJoR0nPwLVrnlv9WMhc/H4fbeUXsepXvNfpulXsMgqrgkF9/+woHqjaVkzCafGgVyBNUcnuKJ+oN
i7UaJxvNljZKG4lWsm9EJT8h+FyA5jf7UN0XgdiSSl5mt0sF3bNPfsGeQP9v2npl2QZKpGGAbL+W
Xi2OItIuPmmCwb+iRIndLRPX8kmlh8vjxMUpTfKvcpB52fC06V2jvfXZUbAZIlCZMRSbnfwRL/zA
SFNMbr9dyzFvxyZck7/vJDwKxwYPF5jkPbm0TT93te3pgO5rGxvSrlWbazZkDo0gf5spwE+OBTto
pjf4ZMpaMO/DPvD4nhLeXGnEPDabNF7kjXrX4nhe+5X3/JZcuZ9ZyM68JC0wDzuT8LxkOohw896o
cmvYD7MBGLmFytTmcmaab9pg0aE3e0+gI0dJm5VZ3h0UYRtUOueSGRGxHvaoDsdFOHNPrG23mbMS
pRPI4NtSCwhMIAFdcPJzpPlwfti4/KBWmlLaqanIK6sHSPHO/Zb+2zhOOOON+EZuJCF/tSn5pZD2
TgzSHXydtDoU1Kzb78idiedgKlGbL9hk8OyyhSPK24FvSP70g7bCh8jYE0+ACbL3rkt1cz2/u9qI
FTRgo3Cw6UKKhInv2IbXyETtEfkRtZLj5JjKtf8YctCbW1zI5vKQ3cKg38HvqrtIPQReOvZro1zm
QMkNrMcwrxeDTfLX83mticnCpec9K3YKPzLQoXlaDe930oZhQBpPc+1ADxuJvCe9rOAa2N8nN+uj
YJabIR3JSjjsuvkd9oax+qG7IX+XRzWKroYz3KSx8G1gYUS7WtxBeUPTq3tRxA+0kbFGCE7SXHS0
6pgBHY+UsKZViDJz0ebG/Mi0EtAT1ajQrQMWiww+bm6UR2Bnp8KAQZBYUny8Tpxxg7u6WaGybBBd
41r76q/yHA78pYfWZ+W/yk7LUKm+4aQmAxn6jely3/R1cVk24lFtxiyMhWrd6rmv3L+dJe2u07a8
nAgZKDmk05sSdLaE3Os9Dp+YgVL4OFPVJ3MP1nOd491qKwcLVWtrq+MMSXNWgghkH4wUOMOGKxYA
pCUoPiXZPB7gA9uXC7+2YOoBU4K2KBM69GpuzdheIdZeZ3j5TgfbP44Mk9LlUYAehEdORZNZgTHc
JSeMiCdcw1tEzV6bSbaEm8BX211Kwz3lkz9svmqKkf7cIH1mT1pHF96wJYRt1H+TnjoNH2wVkLYu
JAu5/Hby7Y1Xyu/CkAHM605FaKM8v2wghPCBmtMqq4GzVasogKJWZkYWPMfgYmTyk41JLwhrbshj
+RybXsx0DZwiM/sqHveMT1dS4FJaMa1r38Ehu1YZWT27ECMVe3Oi0hxHgq94LMR41GFjNIm0e6Mv
3ZBz/aAIwSMVLvHNL0pXhZDvp1+lLpO6Liih2Ij2jpQr+O99UDCMZp3R13srdJRm9qlUKj2J9UZw
2J6OGiZPTxkkzqZry99cfji/V7xjLe0Lskw7FB4mLC/jyTFjJcjb/Z2xHCi8MnvgL6X1U+wYrMBQ
f1U0144Qg9dv4S+qJjIvmybh0V2jqXQMZzSKppQYTGrXAEh0Br1VxWalLdhwtYQv6GvC12Y9jMTS
40Dpt+AFkfx2dXR+65yfnhuMJSsX7KqD/dju/Vm7aaOSnXWveb+1oBwvkrfflecY2PLGzyYQTa1y
2h9w6m9bEyge2cYb7WfQe9TnsmRuCebQy5N+bqQY7T7kP9IlhIyQgCZyx9m0ylX4ZGHPXlnHVYwS
5Fm6T03rsfDq5vRWFGtmQlC2PfKSaYLErVkV8C2SaoaR5575OQvJR/1udzcm/R/FFlzwWMh4rror
tZ8w8ZaLze367Dmztp87p0pCi5F3DLQXHU/+ec+ITY1Ghv1eSv6+p0FXf4S/Vh4ExZzn4eWeD+7G
YvUxp36HJKd4Dg9ouLcw5lDsme8OPmvDoAOqcz51iLHP2g8ATZCUqAZfN1P556c4Z/+T3Fm1m3Oc
mag81MQjH43J+yOAADIDj5U0ufIc4fH9zp416XDA7GqJXthg8axSxV+sdOGG6rTlTEower3NAtmm
td5s1pQD8d63wBD082lk9D+gFHbRTAzcZ35hNUsNVeSXjI7LjSphczYMlonjhIqsOCqgWKunw4kH
mqmc0B+zj4X48uJjehVr0SdqEjh+/9OdAaKhNB43RWQOBIcCNK3DR2qjvos+aO67cYAh6ijRxj+b
XE7Q0kkX25f5o+xRbg2BnU5G+if46dktyk+k1C0GDj576TU3Rv5Ewri9LfMfm2+vYuAzA89kgQWK
2n1GXjtE34YZr4GvVoPW8qDTDXWpBWtBko2bWchqGdvCxH5cXObT8iTwoPJTmx3GorvhhMQ9J9QR
FUTv33tyoJA625/raSuPJIO72JyErTb/Il9Xr0KrrizzAQwfnTqOUEQKoBHa9j5Cj16mtS4ceotZ
eciOiB1Y9zop0+luxyTKREaL9Lyslhj6VGuTe7x+0vPK0X7QwdZUoiA02FGqaUdoQ5z29guZqVtE
4xkjWMIH5pEJE9WEd5rfHYDhRIEfGbfWG2XEQVoWfziGiUXQyeZ/ZqoclUx+ggXcR8/ZE+OI/a2U
lNIr/RgSop1IXoTbphTVKEN+xNlN0FFJix0XbDiDPmAWNdAE2ncNUS+YKNU9ioGBxyLW0NNWeLZx
OI0e53n6fZd4+yW3DxYGSrzneEOTI0DOQDLueUQgm4KFdvijs9G0zFV4gQWalpMT/mnEh9hYAH/T
rrBsLKhxk+b2Fk6JixL8bY8z4fH1HJhdr1T7Rf0rC+ZwPsWi1fP5nHnUSgxrb11c9piKMJe6ZqpJ
Ma4qpX6MOHD1j2u89eCoybHvSepF72E8MOBXMZ/dEsKPDkcUTrfA1IPRM8TZ24BuHZhLVa+EMidH
Xo/TfufBXO3byq0uGiQVV208yV9tkQFgKWrzWdAXDRGO89CzrMtNLZvtXBaWTK1BRLWATmnZwUEG
m/rXjI7p/cEJNWXfueWObmCagBwTuAwQjHIU2E6xQ5felSIkubyJQtcDhTJ+lMRlN8RmqiIOYLk3
p28cEEfsZK2pNkLbujDyBfEqt9YdQuTHuKWUou4jARCNHAL40QZW64jDXCiInwY9VW9gogPbY6td
DIAtQTv57OECGzVNAgy2q+Bm0CoxMX9ErprDxRES3Hv5CQov0jfgHVaFbi4HirXJ+LHfM7IRn5be
CzkBfd19pt0e7Y6FJ5y4ZQEOBfYY1H//lvmC1MiBEUEHM6bQLLsSr3/QgxsXT1/E2pADxuLWuBQy
aleS8CfzgApTGHfnL3tukx6yzTxtEbP6g2WlJxkPScImrum3yJrKBGcQG7WZpFbihKK6A4XvyBY6
mJ8ec/srBkWFKMtBI+yRkaIGmkDtX6nZyDW6RG15pi+HadqUuI7uf3CqJqAUiNJg6UhbVxF6uD4F
zCGRHdAo52pBZ15DEzxGHZRhTn1JEQA58vhocrGH3B96ge+OLByfn+7Lz6l4nQ0qJtpkTvl800Nz
eIBsSv0ncXsHH7rA7+P4VXClGBOhNuZfdn+qE6Eyf3Aye/PsffPVWRtFKQyPsZg9iz+RxryaJ4f4
6A4G8jtWQ1/YOPhFanaMdsFDh4VKKSfwX3JXNetd17nBNwJWVqu7MDXjpmwO+DdrfL4Y8XULnqwy
eRqn6fDlq1qbJFOu1fBl6wFamijoy8H0MxjpVrbaJ9TxxXlZwgxKMHYVukliBe5Ltu7LoOCpT1uB
norLGfe2RFhUfZRQ0t74B38TLNihVp4OLUG/tHeIvJ/7wj3ZnXqE0rzDiPUOgMFwg/ZjEl5jOVx2
KSJuPUM1C3TQhAUwm/vmWSwWg2WliTk7nEupdOWkjBy0VrwqztPoOk/VNnGdhruOGE6IfhLLhfus
tdz53QV2aF+3AUCPkQVjLT+ao2wXQZCvAlRmZO8qF2GZFjQSdyQC39VidGVS8fqTQNZ3OMxTG697
NNMg0NUVCRnvY4nxxKyjl48n+F5LDF88+oDLV4Hhj3Q5uXlgqOUW79RBgetdiqL8Nlp76EkyAE6d
BUIL4fC/io8eEEfej+8Nry0RaYxNQB/qYXAb72ilRx8J78Nwn4UNe26cTAT93vspAorqFgdovRYo
fqSyps2y8WokWES2CSgyLmORHCaC44eFM7h0mljHkPfj5tohP8C0UC5Lh3lAEW0juDlQOgtbB7oX
fo08Jvumz6/vS+SnSzcbexUhYwZTNf5tGZEv8hga5aCh893mLwGscBDvMi+oirkHuzdZgYE5KjYT
FD0Ro3jdPEYuDWfScKJDRqCsV3kKMyU0PO3LTaeM0Acg823Cc79AHNiSwfQ5kvDMF+ktUhqFkv3d
wM4jzHEKeycbR95nD7jZAy5Mdkeg7BvpmktRoz6orrh9ZNY8GrIz47qGTWtPNoknAbCByNutxyMj
sSPIli4lQPFladxj4UmA9FF8paIogABkCkXWuFPhaNpTn91A2c7OMComrh4rVwEmvJfxwqoLKwZz
brb3HaWlZTbijwco9Gj7KajzXKwGU0qYMMlMgYsNxGUPe7KifEue8a3MJ8QvgUNUQKNIlYw1ruRe
BQufkRpBZLJpnFI1L17AqUrHgXnOqoJEQbZMF3/crLgKdpydEDgx0U1HmD8VTqw0GpkVHUW0hxCq
+ZhWMHvJHk9t/xrQvVqhEgivbL4VibT02JM5RBsaE4FtEIr0PuTcA/8DCqXwMhbXXUr86GBnb12V
JVBcx6IcG+2bk0Vp56S6mpXtAsHMPtHNDUrmaKWELQ9+hHDG+XagkEutIhZ3/AUpTDj9if3GteNi
Xq26az6TPtOLMQq68+PazzIWT3D79x/mxDjPSY9R8rehjk1IblegvaWIDa+hHOr0s2cl5uQvkBnK
7f7YVV08NQGWYLTYXFskWsVzkELdm+woHSxlnrGb3J5uw/lKqqVLWPnzcCAeOvE9z6XEq8DO46bB
mZOcIVEo1Qqdo4VSpG0gb9irlNp8rzFXuNx/z8IZ3i7R8mfcF2WKV7pgtThmQ+xaVtSR3LJJ7wv2
ZpavsGodXfNM2rMiLQDGHqcplqomtuUwY2Gmn0u0ogzuer4/8vdeSQ/PEXDh9yHJ+LVEvc2gHCq3
EBEKc9kO+aIfBsRyA6sRbcQwihtyYUPycQ0mMLxu8REEuUN9ITs8PQZcMSiBLNmkz/u3hOQPVzIr
Gf0WtjlZ9AYkfYWP4noQoJz+Gpu+tqd64d9KLrzdn4m4aWiQM624QavYl6S+xRvjhMGOpwQVk7wd
6LnIZA3AkdmyD3wX0L2GlUs8mE0qY/VBY0QjncHSBVEWf1y0QgfUKedZbjbUZvKom+5W1F0x6VAl
uBquc0gh4qgeFacsJfl1ldjLrUAqFt4YhfXLlX1b2NOkziR2/1iCLyury4S2x5Cnf1/jh7VUEqnb
OsjuiW1Pbufmof4roJLnS7yZA+NIsd0QkWKxSIX3v711Oa3JZNYa9uzECwOQM+o96cpdMO09yrj7
BRNTXhNrixQs6suVesghotWQFJFGHcn7gGoNsiamT1ej/XOIKRO52+9YsSqXpJFCq7qzQJUVxfmR
imCXKHbUiRgJ931aWoycIXVKDF83vRrXQM4qaXuuBTWW662PYtQIIRM+SDZItYJfHAR4AInlp/Gk
ZnFQoST9j3UzDhvKCp5PVAbCu6SwsnaBoOzb4kfrXirLC4fQm3DHGyy1343kEPoAYXLAOHW/8hFJ
NPQRwsj7zrVoTEBKaURzhboatqVf8lB2LSjcGFdwfRcwe79lGQaaIVCLr3xlZN/RsIk9LE87fRJ6
XIugOGbY4/r5ZIHTL1LFEyy+9RTgKtxDwWdIy3iqaHJVK2IJVExq0yLbYJ/ax5yEzwD1jzc640u1
Imkr987oB8PSGVP2qYebVVbVr+FI9XZ7oNbhMQ+DtNng3ipzYwp8UhaWuwNnbgQWiseTAaUznSeb
pLZtjsaCWch7KgZ3+dvovQDOTlahLeqC0c2G+5qlRj+eudWPIUQbvmoZks2k1UDNAVjHweKsk8rr
HP8cwN25PYAjZsIzC06dcbnChO21GaTfTnRvOfQ/iAFyj9OvbmkaDiLkDZIxaTLHjTSBQHReA/83
/uQFAiKse5bk7PxXA58Y4XumLZsJCMpG7Vib3SToYfifnAN6mkd1Cu4cPsapFJQlftCfdW9GF4aX
W6OXFWi+5rYWx1R/J95iS+nyd7LAGSPhLx6mp1sOG/47UdQD9hNPG7VhkyrbP29znKTaXd4rWTl8
U/lfhwsI3WvBU35fzE9Uck25AtH1+ufI5sMu1MJ8dtKV3KWlAWklD0vJorqy4jiVgXLGoiB52nPG
4ywztii8L2zK5r6+eXrBQ0srePuGOUT2i78Um7wdYx2fnLhX90bgzLOUpjUOU5zGEbbgyv4YUy/f
LHVNVyTAP3yDSopJPVirq/VRKiVJ4dcEXy+1Iy665VtzBspvqBLmJCeVq1jGABrn5aiLIeYnbAV5
puYFr1l7GSMCoXWXxK1uPxSJDNzSQOib6xEmSSoeR6Gb3RrWmIrL2jLRpgO/wi8Qj7Y+aBRaZzw2
tBg4ajd5JkDk963wQMjleM2QwamCrbOp/PcwmH363pyTeXM8ICHSg0qr0wwbibjsL9L93/YBbaJ2
wB0ho2MHZ2384625O2u9gCEbZLNEn6mV7ZUMDYewJzuQ/S5bwDz0uTznIo0hzgSWLW/BXgJI3bIt
8EDjs63XA8et5LCu6ieCxwzTI2IuAcqTOAYZ6YLlWndc0YcEuWbhysegyd/zrG6r8I+vNZln86C+
SvWHxIb0mL1QyU67XqpTHYor7w0BVQpEMh9N2AVplh0gdy4JzweyQ1rkVdWOJU26/Cj9+M+d6BH5
XAsKhv4+AtyCMIXvn/WcwYiGPLTWTUmooOQaBU/Yy+twNiSVCWBg1921Vrl5l+Pmwx8Jh3c0ylHJ
3oSCpb9ivp/ovIh0OkxGYZSpcGs/a9qn8VoSwjqAoCmuNbDPtUWOP7/2fDgAaRp+4n65N0XPFHOS
tHmkeQBhNmCKUl/8j4jGnN1Xt8U8StYA3wYxvG4JzDtSHUnVulnefzkeenibH9wBPCc/kSm1a2Go
VKwECyqTOmpwxW2ar1bGnJa44J06wSXxA4LCaunexCP5+mFJe11R6STfmqSwOEBwvZlcVj7wO0Lh
tKQjLNAsOxASWKwbtb5bsmb4Tabqw0v8WMrA/bY9a1sUf6XsXb56dLA8t6esABj1UDlfqCRQhDRO
myx1E1lfuvQBUl/7AnWesvm7VVzUp8d1qHpHDL1d1g5NhtADs76QNjmhMqV9tLlW4onPy77F/S0F
3zf4s44RP2/iPjfNmF7dsQpv/DB1wK0KyqOEKJF8sIXjrMgIM1pj7cQ0y1Ygb00C3HQ4yngWkK5Q
k+lqSs3kivKLDOU2WsbzDXekfmxKYx0po/nPJAmmLErDrxdCJYHa0dOGqi4lSgfrbteBXcKLHXdX
S7vwnCI8cpt501QAQqvJ+72kVRlu1PwaYlfNsoLH6H3AfFcgOrsEx1uZhRgfKWxUMdwol1teQ3kk
i8OvTd9SZbF3KMwirFApmYuF9fCNPUnrBS7Z1nBbXejvbeDqKVCi9yICBLa5sMX1LGHW/n941iDF
RqbFMvxyiWxgNBpWyHfGVhHOaHuakYsgXpW0tQ2L482W6z0qbe6Fqg24K6fwCYUxlYGh/a+WKjFi
guPa296Aj/Q5kljIiGHX3h2VhdXN2b+IQnxeqkeQXCWd7B23QrnrZdeAcyQ/v4G7kqwdGkkPMs78
JlzYCDppRLD1cQOrxkD4SoTa4a1q8vhKVr5RFEngiPOxCHirkA4lK1xH6j4ZGb6Ls0ZfQRPrNcHr
r9Us1SUC+mXpj5sdVfY1WST8ndG4j/dL6WGOkka4wFOP9vcsjCSOGRMWwptUBBIYwHH5PMnaTszh
oRDJo36e3K8s0+u54Wl8hU7TpY1A5jlcDgqKpg6+sW7C88LYYeWW5+5V++I6ZwXwlbqLC1VmPmmB
EX8vKNqsIpGUkL7BYFwa93QeHT+E3R0wdZidb6yKwJB6+2z2cLPH3A4NnnW3TJUlyUuFZ9l8xGWC
55VrP4Jw/I73LQ2j24wgXZEgRSlzhRMHXNecQ/zieB958gPb1xq+QKF3IJYNApuaaTR1QAQ9g5Na
yDJfqG2A1uSnelgPAYGQAq7/zwVZUScZqcHX8mig8lkOuBMYgfFnoyWrp0pI+dy1dcKzHFq6Kv19
J+iKdRxT8+Kw45OKQlMQkq4DnruX1QRy8ycG2vtcNYADr72KVGOl4j9rqlZ02JBAsgVE3ppTrQJq
JffU14NCHFUQuzALccaC/v9Pjq9B+wt55IV1Pho7qZ+rOHBo1+yJIOt9oxxAkf5jyWfAnswKoraL
AI+pqHWPM1mfW8FLDxMj3Rh+A/vJCtjl5yD86SJKNrx2pcMDKDv+/ykCD9K342oKS+yjHKGvVX18
51smTKDxkJv1qdQZ8Ec+M79dFZHyYFP0LZrtmo7u0hhHwfLirLIvlR/MEfPYssycy4PMzxkumHTQ
ic7Aq1+KbRCs9X7ekQrGT/eIEnb8fZfb61bI95Q9PBGApWCO43MkW9TaxqlhTWdz+kx/8+S7Ebt+
sj64ScykUntC8OmyNR7vWC8ViD9/hzIOfSI3GLJt4q49mjDhTwYyo9+9EjIj2dscCtYZn8rQ/0ZH
tClk6lqupkvxziAMl7HW9uD5kSTdoiilCclrRyS3mbUOAS3VF60iuKADgexvb7gd0Dfv5n6EjmIr
8xLLYKUBPqY3gB5XggDddZDmVdtQAfopTbwNEvHKU05Ne9b2M9Ij+t7I11iefVin6tSpI3t3/w7F
UOCq9jcwsBrmLzsMT5KKgAsJL8yN2ClxCzddB3JMUvL+H2VYxlwVdUedNfZOBVdapi6xf1esQDaN
vsnMBiu7Np1Q2QpJSb3CPr+yuFhtDRK/zUHqE/4NW3feFGuxBsiSPYtlu/iacHOiipKgNc+bvGPS
XLHDZmC/3TsUXOhlGL5JI/K96ZPtAyhWBXRGHJw9BFJSj48ycvnC5wRKkV1UyfjnFZSWsQljWTSj
dhZXh+Fq0ySqZCn/KYOLqwgEia6eZcfLKsvP/0U6Ra77MhaR4Uk78sUrqRl2o7o0AqaZs6+8issr
P448FAlzm4L6c91cehQ+9TAsBF/3qO90PmiIFZtYLaP399o9GaXbVYkdQrq0XUnwWUR78FcA7qfd
KiKCBNGu6zZI5Q2nD/xlg9s6iDNXdGdjLI/br493pJyHnfmNDhbItqg4h3LDciC7kYctKxGDNCnD
aPySdC39Xe8261hPh7+MGOa5Ra5U6M81TPnKBw/f6hQ5ihlUKMSjQHV08eQpYIpr2Wc5mZRfh5aD
enM37qnS5N49pJvekcdyvQtenxYP6eqtc8j9C0oCvn2Lq13KdvK2DgB1lnmXGpZYKf1dY9znRjvx
13f3voclVv6t1Do9kBVh2kLHW85rdA7mucJq5yo7zfdm0gdvkwVekyltDVUqOrlj3qlM33s92IoY
AR+SCs8qMaogKl5mbeBOibSQMqyx1UCIG0c2Aw+3xKaTVyoExDoxqEnvKCge9T4GC6OVkkyN60z1
6MMbV3+EAo6+gzeMNuZ7Ajtgi2JLTPzxJeEKm7DlbdAxxlbXIRHVcWHz7xwbo8FyUjBTbOG0wYkw
ZYHSu6l4luW9HG60B828wB13grlcX2FBsAYxsfvhAL6dvgikoY1iaSaLZiuiOL0ONLAtvs+nyBjW
291OFIG9Z+MSOi0dKtMC2F2CsWJtu+n2UxZPktv49NcLtsqnGyyOEzHmlutRrb6UCuQkWxgi+V3a
SH8LWbiYupH1t5vCd9usGigEWSzkkSbD30WInvMJCSGvCRVvey9yp6PKo3uNc02b96IrbjegHuz9
gI53m8QmILhoxF+uWmPA/9qJNHaY6JjXsiDvjOXVIZ2D0s88aQt1jhZuiFQ+J7FuFZ3la4fyB8od
BPfYQuA33RyICUfNJrsDcYSzIDcunvunAZZTaUP0AYmDUEIKHJK0tnaXwmRHbDXGL9An1fcz0S4F
NV3or6+8E2bcaVrYsiEwhdoCpvDEucrygzEQo5wrcV0amgRz4kKSQF23RY8Rih+gCSX6gFq0ajW4
YrkXMcHACzk0Il7RVz4JBWY4xL5wOJy6og3M9OZiFusNj/m3wUCJXpyrSUqAT/s3ZvWqSG0doGjG
7j+ThRKwvjb5HV4Z/aqVzjk/BEC2+ucdYtKWtUx6VC2q5CXYRqxsY4wa7w18jgilIx+bfxJ2rmFT
tJbi4UWtCpt5dD8LjEXHB522SBWy+r4MW7poU/HbBv0vgB51ojzO3eLaspYeAiJPxP0BoGqU2nYx
GYCY2NK8M2Oqtgkq3ZbcAN7FDkdGHQJD8eyPldB3bX4jayBTB8u7Whquwd//XHfpQI7cNwqYB1bq
BK+gWUSarL0uJ1p/btxVhEQ6RYeZsC8y8MHdVpSidP0bwzq5GAo4jnG27I5uyA+mX/CeWyN/HwAd
i8cjz77NtOxNMzoh1fYdC52Tevqi6a2n8EyCQ5NvsXcLjYKEwIKqem/SccuTHS3/XRGHbqGNOx7B
zjwP9Bhm+P885uXMyUE40qnntp2aR+6M5hvLoNYbzc2AGov6s53P2dlnehz+mlmT6wkHmbgAKIZw
EF6G5PdQga/OJiOT4GFEk5ZqugxNBphilGvFgYJ26HpYOQGv8Z1+U/UpK0rYOAeoyK6exFspalwj
HI3Sfl8Za/o9rOs7s8zrCQBSZ9r5LZT7UsnFAkQEYKGfqHMMtAqnoh9lgtdIbhL2hKmIu0GInDwG
X8kkIB915D6G8Vz7SJiIUCHOfIA8m12E6SQjEPPNri+esWW6oXzbLgQvkgrwIFXjSBSchWuGkCE6
l/fudJI1SL+PnOFRIXA0YahL5z7BLK1bQT7lmqfPzG2Mneje2pWbb1F95UptdF33tDo84iNWz046
wx97w+Xuwl1H9S6KGZjYbgH2Uj7VIL1p2ySW/iT/PjOIaiMvoZH3it5C93x1a5/cZ5V/hpodAZQP
3Xbk8+Xvwq5rCEY57vHOG4rlbb2d7p7dDKU2UOCo/P2wDYQ4Z7zpslhcp+OsZ2l/cc889vyAyep7
0Y3h4j9UhWGXBxLiDS58cKvmZPYH+ZbInmXBQIlL2moGD35ykIWA7rP+QdEfqOWt2G22i6+SUbQE
faXPEBQRAe4/Dqv926RlUKIVzxR9aqHvvcSRbhLzv/lCWEveOfgOP5duHH4eNjaU4Bq0rFOkgnJY
HNyuixgz/YXZpvO1jYH+PcgEIzwcmhbsp5QFLqk7e5dZn4kiF80F+sfdCibBhsYvLGwEWw4ocP+5
EwUgzvLADNmWd6GOyKbmR48LmbM0BTrkYTfq/qTiXnA2hU/isGMLcYmQAwYxBWrsAZTHeKt0ATGp
bO+fpAWMc0si69xAb1uIxlS1Clo62WfMhwdNAmdRPOm27b7ZdTKV0PySTtM6jYzm3HtotPS4pOmt
ykx4oyLIIQTd2ub6/3lmuPf2+q1AkRB/FWWoNBRVoHAONbW2DDoQ7aLY8HeCBhyCDrLbbp6wsz2T
OiXrDXxflTHCxvY3c3yF9oPcNIUxaMmHDF+kIpR/N6rRuu7VXf/OvUrOvWOwShi9ZDahD/a6r3br
XwU+EvCAKP4sx7QMc+n0pIfddSJ2CSxSRdOGRpXy3iwPuLjeI8Fpd4QAg2N+HG7NQ9I8AQitWecn
mxLC+DhQesFHsbapAxAVL3Byj6poeRNo1c+SvrcAwf2zENXsBDnfi3sEvjc3/AXnoNGo8gCrxlKC
lbJwLbjmDPt8wt7ggkvlBQ250P+sH06uBZ5LjTqkgHXBhzIqVwkylKWU0rUZ/Og6p8glZikEF5xV
CX8XRCHFzu5OdmUM1+kf4Kk8YSwgM3AeuZO3vlBv2TXDGhCOM1t4zb78iiSkyJu3xbFMphzrRXb9
pw4g4RrtaNyAy/lqAODH/KimOFMz0qrMymULMmxV5TY/0HIaXkmTDRbqbI0PpUnyLzmlxjYpkZzU
8BEC/Rx5bgJcAKFB7Ng+wamDUeAxh0fqWtH92yg+R+3hNEkxcxI4InE3Yh1b1XL3IFD9xOybJqzc
nI24QpYZgClG6r4S62ifPV8Rsy0uv/QPFyt4PQa1uQvHl6lL6wrKyAROlTKiWtSN7HUGH+sAjpsN
FrUhM5ntJwkE6OZ4slBC69h0AG9YVXEbuGBepdiRS87ZjCtiW7YyGJiHlXtW+bHDUw8sd10xw4j7
MkUsAMVlIljRb95jlMIoI0Cml78fVhLAqn/psYzItBKuP3JvNNYpGY9E2LVI4RcBOFSviSkT7nFq
3X/QRPJIrw+sG4BjMrWvvY5LLCmgIhGLwVUZYBHnXM7Ga0mdSmplfDRrmJrsHqQMOXPCDaS8EEes
+DPROKX/B5lJ96qSs2UwDfgESV1yd8zWOjnOR5rSmvp+HtR0Q1f/eaBFglcKsFaD/ANHmMYorsJo
KnnyQDW8ZLErsqksWk74DENBhppwRocVsMkO/LgHjICLEk4niZe6RviVZ8gcFNX/oJC0pecgIYVg
cp276A6QxhtX3ID8mj+bLYCuSVwN4yV36+goj4Y8UzxlnWT/t61FAIF+KvLtGD/IX4CfEkXZGu5n
lRn3CkzYfyghHW3KZm7sfnacpDYE2LsqndNWpU7yLAIHarF0LE8ljXovg55hE6eUKLVTpYQBhwdb
9So0dTZBRmzMD1JlQEEPVrO/lPhjthKl0L8ViBhs3fiRuf0HL5TIeZxN3bHoOuhYC6/85BpfAYPW
G6NiOOWVVYz71Lyu+uh8+ncDxserDQawrAg+HbajTHEe7QSMpiKYN+U/SYko3eFWVSD5rV36HyLl
FlA0NdRUwGOgijoMJPDXSec2tP8czABMMiTdI9NxXmJGxGM2n53DFcQvAMmoOFuu3sk2oROaDBrr
FJSMlAsBEl3XOvcgwpJ4ghBeG8B6CDBsrhO4fVjjx/1ecv5N1Ickf5vn/3iRYZCF837lIWkE3kKb
psvoxi7LR+VQk/LA7L+OlPIrqK9FX4PW96UPlyDyIGjFnnu1kOO+7DtuneoPOjRqea97tS/aXfB8
Ah9IpJI2krcseJgJqaxy641bDnGvFb4EW8Li6enuOgSmNkXQjlh7ZFBL5RToDxX64k9qJjuYYpH8
xpcaFKWQ+1dSwWbDEfI5WHyghSJsmyJwjk3zOSbtU4FUzwZjr4uNMG0DrwMKMCJMG/kWtgqsbWIC
TBtZTk4O1ANUgi0QmKUqqWeS/jYnge4et06coVmlyFvSGOaRYmjlSa9stLu5897H3u5X53AF5G9v
hXtQvKDv4DucAgRHcndXgLbiO0SRgjrD40lqW8fXVwyhBDAANuHrReh8eHbmvprwqqq3CB8S7RfU
1BXUixBsRto8fHH4z7+fR5TZO5hqscB4tx3pFvQ5vWyYZ4Pgr9NIE8VsoWMReH0z49awbbfFyCMA
vnfQ3JWTTFR+ChOqRx5etB79NMmGi/HhRKx9oW0gFT1+OjUnpU2gGLBkPMp2HGVineOX0ab1O2lE
bqr+p+i50M2zZQMHYkl6dEW7Di/zXqQLlbWWVKkLlJNh56qvaDaAZ4TA3aaD0M9J906m0yK/+D7S
fb1OZxwE/Rt5wHKJJnFQCiIJysV779Vq1bkFp8e/Cjl1zJHiqyFXKwgo7qqJxY+CJyR0kFWPmKdr
oY04q/E6f6RY2q8kIHJwmxxSTfctkkp6RK8tT2vJyWQzLJAN6FlJpnfQQMpXK25PMfFAPQq+a/ED
ayRcx6XMcxXnVjoEUT1oPQPUlRTPcoRE5EyD8xRcIOfjHod/fy7IPLvJ4terApxY8kx9d0fsijHr
5vAW+oJNaG2fzQY9rSHY3yB0hByHrIUDiOoF8UnQMbJbkIsxKiycKiDWezfT6m4iw0qPdI+fNQ16
wg3aZClcUFWgXu26bYZ14Em9m0KKDd9EGtn4NqJsoQuT7mdRsks2JRfFBT931qZ+jfZzqDz0LRYw
4dLXK9fu6VwLvQaBNj2B1GexJ/05qsPJ2+Efd8nRkxcDzxR93o8ZGIjLWq6evJ0gcwHpgXnuBuL2
zEEQMVa0VgZNQCVzEgC7kzIdty1q6O32pc6n/WnvSZr8SX3UNMW7FuWylZw8FIn8utTWU/QtbV7l
Dy6K/LmERT/kw1gjH5BjpdgQpqijO19QRumtaK/kfcydRhMvqJpvptp0y5M9n6BGSnbB81jMY5mr
b/5vPERYIAgKpioiPYh6mCnvlwiuwKmBikuX9I0jX3Jtmq143S9rpwXvP+lby/9DU8ROnoN3MUfZ
ItAidDWErEcafIXetmPSU3UbZ3cyyFSX8WggcvpZj7JZTws0W6Qjy9Pgu7SGnkjJbq8K1vSByFXV
c1yBaPVzZMA7iSijHuFdIU89RhnBiYETn7akNIiA9i/7CHUNQ0eZpu6gDCh6Ld0iO8G1BhJzlr6/
23Yul5WFywx4iBQbfQ5N+yg+zZ7ri/RXqmIGZHxaVlcSWeTxANY4nM2WmrLyos10oE4Zqf6YEvrl
E0xWGsxk66VBcE4QoWT3vtWBgtkCdvwXCx4heBE9zqxEUr+pQqQjdRQuCpHgM4uy3glhX40E1YAr
32odcgtEShibVOFnBJh1xnlzT/ErILb7CPMMgJhFUJwqMeAn1aGMG24jLKdwHFEFqzbzn/tYeGD4
UCtCv0hrrLmn1vJbwwIXd9t5X49IZIrX5nyjYcdtEv2Li/5TcaccE21AfakRMIBjtsLj+HBJkKrZ
AoHcVxPdSAEJzo8xjbKDsmUDFqM8fFlA3/r1DIBXt3YXNHPUs3hvCb1xpF4P5lBEF1CFS/p3ZByh
LBLq3TxpOk+xWJ/EbfqcfT6XDqO+Shh0lQwPXnk6SCD0jb0vlQrsTxU8+Ed+Coi7m1MhAiFkXw88
P0rN4aPqEXo2Q9zvyH2NtlktTBVE6D0Hm+GkCqGNyfyUMFRASnKs84JT9MnJWss1l3i+vygwP14K
r0XV0our/0jlq4dqFkRfxH3f+9+O0uSQdODUj8VbTEmcd/V2aPaa5wZaFyNa0FIh1Q3WX/w7fuG0
Ij80SN+a5XLpfC4gsLgZ5mmgJOHvImjcP6J1S7gzP6OBlYlP+rqOo3sAVuJiddoLK4OXPuY3/1c9
tMt9iboWXH0zR284pGGbkPosejNc9wVzKd2Q6EMQPOAGwt2+xcwKzn944jsI0HPEYd0EEp8PF298
+VoOo76dFElt9mMa3Fxl9qP6/glbwoNzXt02+UTPCbEeI1k9CqdII2Or7bK6C+niUSlKqOp4DhN3
CDDWCE0dS9m/g04ryzGF7LIlafJOe2aill/CIAFFxQapMn/y6XfmsIh+zFLaDO3xezSNZb5wcalc
PNxKam56JitKxaV4Z5WiKVr0WGSrUb3/o0sqdYMykyc5fXSLXCIc06pJlyQL5R0czqcntZwAPEgu
OzZIM94w6WnJDewXBpj+AAg3RN4fACfPu8j/SNyGRSXfgN4Fb+qk34oHfRujLc2TOPZYyTfEm1nM
qEGLwcQ6bLP6PTnO2dXdUf8hwI7mOQxSw8vlizcafQQaNZThq3JrCXMGPugMKm4njoNGnxYvrrNc
jbtNCvQqAHRfmHYsS5Fo/FfIYYHOmdFA3u/EaHUBi3aCIzXp1ernpQ6vm+8HNkv53wt9KMo2wSp4
rmBmS+vV8WvzTRHEWHb4snJ0WK7C6WdcM+zktrI+piZx36ZyAUYvywboMVTdWP5THF38gzZQIZUP
+Cwnzz9e29Ip0DPHMh+oaY5VoeQXVWexe0ZORWkteA/Xtg94HXMqX4xqxWeh8IYLtqsbganPpEls
NtBIWvqva21ozj1RZ+KItYv3AG54w35TTuPPsaBv2DquwJtOG7O52JM8Ei8lyyDkbRoIbwH0SJlX
zxItpk1eFKVlaL+GJG9fPW4bjESHAkBi1yZ3OW1PjuLqYf1nW6WqQsWpNpaQ3Xux+EO3A87XDAJC
w95ge4CUIxOKl6GDIRRTMI/GmORwULXkdzMTixyRLqx+zXRFvuqSA/IYIq+WWsoeGXW2C4vOMNJi
JROYmCUJOZtnqss4+YJZ1/f6Y5VSDXzRTS/8i7dA5K5Jt/ouFZetimGhL7veg/dlU1+Wv2VTreeL
QXYyHcJXMna/6iSjp5U0jsAb5Gl9me8rDk5jt4fZ0WgPDnkQTDnlnxYCobtlxA3Kioats/0jn6i6
1XxmJxIFz6wEvLOhW2zU7dit3Zq4uL06fvnoSIEeCcrzMISiRVLT8LCX/edD923Z/nF0/8E41Lv+
Tdim1j5qnrF7Rqn70GzKoTWonGigKxyMSybmq6kSuf/b6ZDv/UkiCBlt/78qRPQrf9A/i1ZZzh6W
EPa3VwWpWwW+uMGowP1cF+I5h3rCa/gypSFd28tLK0ac395ByHUesZis/40HANbsWf0tp2G6hGuz
YfNxqI83FsysKITyZGnvFdS3dDE2dSX0cMARlgUdlZ6CNeWHNt6s1H3ZQHTbOjipjCytwCpXBd6W
g/Oh/PTxS9ak7P963Q0oJfVmR3MpD0OU/atDEzB8YDMcfEwaBO2jS9jTEIqDsrLEM9U35tPl3Hyh
E8uO/ByVQKnCWr/lk8Eubg381en/+BsHapsG0+LXpUtU+vLwyG+7WjcevvDZG/SSTvvbaQC3R3g6
Jn/HxP6ih0mil2IWksQEHx8rJJphkbmtCtDA4tOa9hZqw2WNC3EM4Nsxb7BpuvNKQN/SY+IbIrZy
3g9WUi6CC20RFsOoDLHrm8j8RI3qFdlpCA0V2r9aHC9GvSKBvJmRqL52iaOdLwSrnY3ovk0FRgct
5yG1InTYM4kLUngaKiqYXpslTvKKTBLenDYduAcJzgtj4ESoAznNRbehQKcwMu+nuwFOcxn4S848
vP+7S+kgDU5Sv0ciK8GL8j2WUIEpqDTmWWX85UeBn3WIGwoDHNgyOAa8egnpYYVSPU8v4khKUVhn
G1D0k6y4FS1E4Evb0i7hJxiV+YP5kUn6oAAKghqYD68++n2vsSZY+z6l3AKPAMpSp5fMt9Dx3L3r
dwFoGwfFCNNISGyhQPF+zBvW8ozgBbfF449Rd3xil1BG4uElPMDWgCMZw0ltIqF7sausA1CgjOGf
aMTWyy/9B1zt89buI4kz7gAP4gei2x6zab5N1VTeUuB3ZTWMoLDAIQJtNi2Iu7VpNGk+dgx32sNv
k7bVZdig9DgkGDW3CazpVsrhBexidcoXwfZ4/snkrLk2rq7Mylb5QdBkc//zlXIunpneRthn70Vs
0Ry7u8tn/i8PAN1U/nQLlotHpIstKL3ltIyS6GEkh+6L6xOe5xDTwp7vFJOnn4as5k88wkm8pxso
uNXWJx30HPaU0EmbK9oGOAEvz/dvAws1tHi9kLlC7J6IWaOvO/LbvtLCvfCCViArdyjHXGdDhU9K
IxjNMcjDfjL0sp20MFsgzv31g89faHjBhgii4l+qLB7MC7Ptx3Pq7WxHOQQVLHSb7jEb3ruLdfhR
MD/axrU8RMjXfupStNYIdAqXlf5w73ZgaUh81L14RT3uRprqgziI8fIx1ZNbKbKdRceYKW20KWSM
GiJ9myQuYQX4Dfj2mG2/jYUuuuSOOmOx8AeynH4kTgl3vzAwWlVpEq1ML7DULcsDg93KLiHGWMUf
Z9okCmxDjHv9y0ch0t8/fJY+Gx5O5iHHIujNTfb7BV28/KOGbVAqEvkZLmxArwxAEg0Z76t9vYPm
bxz3Jw0VITjms21tEZk9HNxCQMvkUybljj7WzvfpM1VuaJqmjKh3MQV89npve4hHI1rVNc+gv+BF
xNPy1c4SHkLoBpksx6PZAXKULngy6Sz1vL3EjKTeOQ95Y7uGpkm+k+WsYvluZ0CzwPlfznt3A/60
EiNg9hC2m2JygCfwueGEWQhFiclbl1p8ibBP1dAlU05XGfpIQaEBpbevjLJdfSDKkTbYmrQ2cbH5
1XogUgnKtfyCfD8yJ1gUQ3fSxLoGk0mUm0mLi9bFOvKXisUobvp/5dMS/pAsNk9G6rWKsZlVESb/
JjXZSQuog2JGX/sh0STdTRzkZTAUIgIFOe8NdUS9oMLXeW9fdy9cAka52R9ln09THEK5LqUO8rUF
24af2wq5fylOy5oeXzW3MHrdpytI/gLjExMORIPIiZVP93ZTNA/8MsUIG4GC4NZOOO13MlPM5Eix
o2hw0RfXJJeXdTqf75HY6rTy6ErpOJ+VkWyHB/ja4kB92MCHFbMFLWbhvRQy3FjPafTeoSv6BED+
vNeXGZZhEnRAY7n4DlgH+OHoTtpIReEfSv1v1RnCT0cGnqRI4jw0FF8dIo78PJTIi+yMdcLwnKLm
fKJtB2d40jOUEedVrbhDM3lShhChq80BmHnoJ7vKZkqMdfGPnQ64S/8ceSQIO5t/L1IUk46aviIj
Jle2msSJRJkETr3CGI51e6twsU6aOYhi6Z96Bu+gdTknXRZIMK7uJ0IVs0Cd66FUBQ1E93vZGCPo
n2hV0S5HtC2BN+UWN76sy9StE6LGk6nH/DW4KZ+wAVkQLz+OVs0aRig3QZYPYbFEdX/BW283vY26
MyD0NELe73OnFGqyeuOKTIdXVY0O9OwftISFBgRgoET5vn6Gi+zAfxvihBDXjLnypDu1X29zJ1sJ
plExzDAvvARt0CA80XbNMrd/lENK9hPAZaPRp2YUnJzk5UnNHM29HFhi6OGoxN9W+dO8MKhYGHUt
Ia8XTaG8S1QwvekWRH++/uqcMvl0/2/aBE043auzgzPgI9/ux9IkFstWXr98gC+556eb7gtGMoz7
f7ZTdq/x5SAIbNrX+V6HohGArQvnsPDiusFDJQOi7xrZEn08ujuS+3G+nG9EOxamDN+lQnmM3wjr
xbTB5xOi+cM5dCMCElp+w6+1d2l6JGLv+L7svgEfcM90hmeArjiKfRLLLni4HRvtNx8g5T1tY5SF
iJ09f1K9TRNwclA4lKO1442nmEj5jm73f8TN5aaHzflKZ7c7BF2I+E8zVPrTXPhoLgT5V1APm9ND
2BGHEnFfdGpGCiczu8SKqemwxHp9+J26QRE/ovQFbNNmQ9fcbkrQgtr2i2pV/Uuc9/OkJrRKzM4f
ZF06E2whbXU/Rb8Z0ffjKGiBnqcApofIuOvLrz1Uk8uWa8Tnna2z8CTlLxRFpazB7KjvProN0Zya
LebTP8jA9tBnE7bshh6BrywjdluO2VoGNEshdd/V/c1K2ZDRlPsWBHkE+LliIpdSGdcX61n2+h2p
40O5zdf8gYheyEoVPMal4qevRkv2fLQIue8eeqeGa8UZBP+GwgMR0hr7SNP9sQSUKKeU+Tu1bYGk
lYd5zJCl3D0uEN6iC7eq8PEqnZ9wAzl8D/dhx4g9g7xCxGDgDJR5uRJI6EmV8WpeREzh9L7WNUTe
G0SxDhvrzTEkdZRnEWl4CAN+Wkn+6TAC3sIbnd0Vu7aPqhhJvxa62VVrYyPIRbDMqSW4rF4lUyCf
Q2+x45SepjazUxjkrirJY09pVXQPXSZqTtOXpj5bi88lqBgbCCi4+EiIU7+PV4BVbXSzkY+KFVnC
/DBipXs497l8IhCcDNVdV3REu+nDQesSenGH+xLFmo3YG7L7rMmfJL444cvouvocbVE2qIGXh97j
GHM8TUi3CrQh2Ijiu7ObJ0x8z1L+lOm3uzdvQWuBjEI06B5tR5KW3u/etB03PNuFVWrIa/iHxx1A
TT8ZHYSxV0Yn4IAPCzYPHJWRC1NIFqYO5xJmmIIiwCivyFEIfvUV2FG3OVeoq5VJweZxzAYZJMMV
RD7uf8zUq1X5vqnF7lxSqQuxvi3WCKuLPgn2A7CzjI2xg9G7ZZFeEYaOwi3V1UF1uD5iMIXYxJ++
ZxN/+0cKAyC96EnxOctGpRqjSkg+odLCv5b3yEDuFSDSemcE6MQ9X36e3esH9DGAHZDL2qBOvFn3
ccFUB8xsRRAg7MWmjdO8Gr//FNRscEDfoioQ3YH/Cjku2eRxZzB8rzfzVueN3HkQg+aNiabYMOge
nAKKj04p/YMX79jtwMPvA6mSqpyvWj1KLZBqQpsqjldKzA34x2NbPCZbxGKUxfSsHKTYFXZOpFzS
JttBEBTBP31w565gIkH7qijS5iHVfzdnyVOTxb09k9UrFwlG1/i6lMWs3CqnNgMYNaVINzvy9OOk
1LtXyWGJr4Qx9XjKKXGBzGeE0goSdmGiqwCGyFNdDfW3UYIE2045T4DlIBcA8rX52KhyF4Gz3Hr+
9QXDaSea9488cFPcmTMA/t0XjvdXpd8Sp1vFJ1IFOBZSbHZ/sdg/oidDIpacs07McV76F1yjPS9P
soUpBbsP9DXbvYto+NqrGPajL/zBTsrTMwLfjhU77AERLYU4FbvRfw94T3GXh6QEg8jRBFbPpONP
xADGECiOaOs8qCFAXcuqICigWUJ/3yTPzwbniGF8yxBmgWnqsrFIQBYT0U/ZLxxTNqFy+srToKw6
D+FY+jHJVcPrAjf61PzasBnR9oMR7MKOm27jsN/F4d+Ab0mZOcK0pYvd6ULAWZ8HvGo4fX8lrb6S
MDqh08gMJfBjzJVoYIKC1cZ2b/2awgzmUX2TGJGKRw5U+NLYdjDv5lrxPRP9Q8410r37L/BC7RXI
O9xoGEUvgW92IGtaw1ot9mfZHbpgP1qi/+6E7TKVcOD5e78KKlU4Ai+CFlkW0yy1l3CyB198xU8K
PDqLZq5l8AkMSSS5n56pBMaQofYzKaZ05Zarqq6zs9AuwsNkm09EsDTODJcIEMizWaRG7e/nUaKM
U8L/a5F/4JkWA6eeP/Pawl7t33aMhc0vXedSIt8iWCiU12qBYbMESrncHpt3EEuFEZKzTXagD+gU
cFUO3rveBQnDx6LwR7+ao/5pqXfcAhQ3mRXoU8QENjSrGuyRsOsblvwcUKMn3L39Cbo9/RYJ8DVG
EixKwzSbfjmzuXPe4AE/lQgOuaT+qJQCWs1SMG7e7y5MDlGLhcABx4m32QXfqBHlmB/7VDIrsQiy
eqDySVQbtE2zX63kYR0aQS9Exga0YJRegDe3tNlvrZjKVbD+5V90JPLAXqQECoBPHptf9rj9CQGp
985R8Il3McNEtCrqWUrqiuBQNn98TQhj4zx+tI00sTM7iv7dGuSQIOMg+4S9Q8ZpTVQQE1T0DQPJ
HHbdJU+wOtIpoySeWcAOoE/Y5Pw7WjxUzXTO1ru43aArvip3OMgud1r0mAflgW0RN/Rpl5RYC1Vu
jzkYxs6j4oiz137RCcWNju4Cr1OikPK4N1hRl0UPvncV5gkkXd/GdA8DpcH7xcfc1QnXPmfcILnQ
Qva3+hmAhE94FN4ZGay0a/1uvfGmhKqy8vCxCZPHKWOGnnXGmz+V0ULIaWRIU8t6FEdJtCRLP4bi
ZW9A4Eqw5Im3Q95yYnDGPiOdnCwrmRRz3+QBAHuRVHhoWbZYz+UNrvf91cVAkGDsQKHXqvacaBM4
vHyq9QkVLoBjucAwLPqvYfmEk4J1nBi2V5Opo84wpX6ZUbb959gUBTiZMSIPwsRmb2NNM9vuqj/b
F5y+F42xy3uXLpj6st8uo5sj4K98D4PI+IcG6Wpw8TfeY6pht58Y/s73sREo3KB7X6B38TjJB4Xg
4P0P94eG8Abezf8CBMndjyTSGgZO15an7w4MjFE50cJXysnjIifoxRpr3xNH6I7mX9WbJARKod1G
1UlST5BvkB/HVNnF5mlqmHEFKsjzFCAbllj9Gv3ARb33wm663lIjWldTT3TsGj/LbZAWChY8HzbH
DvG17UtH8B6geozDa2FViLFgSy6H+EJIbap5ZOatxXkaOW5I4i9WYqpNM5SnEH3Nn6kODUACQLzq
u+VYYu4wrT3GDVjpT8MvHzw/SrfVK9GzIc/Q5mgXiYbuEpsQXSjeJ0v6ZA6E8pHOQHQ3OPxkkvna
omgTw+IGglf23mNoEQ5PLfCZe6zp16kX+i5Zabd0ZkdH4LP/6WmKPOqXPKgQXAJCP9/vAMW84QOG
ExGb/34Zo4HxTp9pEtqSHmkK5YobXuEA3LfZ3llZmOgq5w5UzSkLmuYywgJ0JIS4y++CJeqMJaDu
4WbgoI3CkdrdCTqYclTLWpDGV2LU8fNO7kvCHGsYwOe4ICPjP1yPFbWHT7rxAPaXLZm1S0wwQ0BK
8br/XchJ7IYqvyNfKXpze62jW9XPlQJ1ISkyrfO3Jx53+NkHbAux3YSAxsIrwbVFZzyCOblzN3zS
JtVw5Bm9ywMXMKiMstg/RszD+WjphQTFEbk3r3M+8hePzZIK0a50Ow1tJ3SIGUJnekerrTshRqDk
LEguYTgkLIryr5DI9q0u50WVwRx4fqcUdHvBXwB1de+6rAEdXF2TAwA45hARO+INejlBnzR+kwBP
Hx87wOVyWogVzVS6PMWrZkxZ4wH03G78pVF0X4aaLHASekx1YYd9xv5dtCrKH1iIZ4Ce5bvkBTUl
o5cWAnC2K4kNQTmuPDoFZPfYpADcnpuQ5qgEpTbd2tPWY/zX8xiNgOg0cl8w50sQeCNjU9N6kpbp
ZzCp/LZ2jRvnC3srS6foUfZ7p7PwX/fCKcodb+r1SmgeyvZUtQsfnJel2b6Ddir4x7LVaQvX4CRX
3oqW+CrHkMCKo7+MRhg5MWQpi8kXgiHBDKzQpE1ALAfT4nhQFkENa/FaVdD61YZobsOSE04VvwGu
EAIRHFBIRFd94AXnI2l5zmoA5X6OqcwPJCWJsg4jIOBHMZnA2Z7i0DcigJTogPvSSivtTsrBAraA
m/CZcGzkfrjFFhw2gMGU/bkGyOlj5p5/H0Gj1I2B0OwFBcYH69ySAO0CjNtxJ+Ky1t3PBNMPCc4u
09dtUOIWGp9CWoQLpnSnudpCbSKEWngYFQpRv1GPsFEcQTX3PABClOileLxJIBle2jfJLWmbKG9v
khJ01lcIdB4wAVj+FHtatDmKFL3hytO97n43DEPbzpTtb9VQFEQNoZbpC1uURS3ob062KlST5dd3
KfM8xPPrl+hm/RqnlHW4vY2jBs7jIWgAVy31T9VfwcVMKFdCh6tLOOO1l6/+pXydXbRoQ5Epung6
/6JyKAWOyro0vmeiU0AGX8+TdbLaTmZhyXg5LK+pID6cJ9JIToaodJnyOZYHksQmsRGbXBxj7IDb
B7DDX0kCEryAPLJcW72mbAtbaeiNuhTUNjgjpQ2BWbioTrmJRpD7QvSFo3R5YpOA0R3iz54x7adv
8LWaW9JFY/clSNtashTbJo5wPDXqmLCz5mhc4f7X8RpsZ5AIHjDDXH+fMThnq6Qtblq0Es4rm8hU
z8W5PS9Lsqk9ROAHJ5B8IinfcIP98BCHwZPJMDt9PCN3AyPJaOH/AITtqGemritSK/DNt+YiWPFF
2uwYLHWVVklFcW1RIHmZRJkgerJ2sJ+lQFfvTKZtrNVRYoc+VHi7OIwFCedNR2ethMsbPQcauJAN
oqGZ1NM1EOhT0vh/iDmdjuINOPwEe2ZbIyaVsR/ulmJK9bvn3MxihKrY/KvoYncC1pWvHmx6rJ3H
a2lt2/nUmdSx1vTeMWq/+CXrTqbuhs1NdC4bR30JoEBXJVuEyTn2BQhM9pjppK9gVnYpA2cct62T
EA3C7me2hYyYoU6AAJ04JY/r52uZq/J347LUs7vKFW2OpmEP930rgyntV2h2qfeuyBH9iJFeQ9u6
fQRyV/k3Hz9GoGh5TCkH5sglg91O/vir1T+wW5PR9/i1pPMmmM4DrxXikw03tz1Y0ntK7GBN5fGr
6IgylVgrso81HA0d4BwVjpu0ToVhwS3MmVu+rj/Jvus+4qR84MvLVy3JxX27vUW2Exk5AybklWsN
5eGqRLFew/YtbdjcVsF0oYXmTJAkUkoaFEfnqSvveh9+wEUoHfRX6bOE8qiCXRBykfhp9v7taUGU
6g776Tb1twlB+DXg3K7gjs4C/UcImozseShuoFHYMxKi0eFoZ5jlsEwY4pOf//6EwsnKoDKNP9a0
dPKThy/KNGAww7Jb5r6FTFxQmdB/IwhNBgcrymFb4BuufHcU39mN1QzfR5aDZLNsty2PyQ9zAHK9
5Srw4gSzEGldqIG01V1MNR9PK2hvV1mYQgwwSCiTUqrflQCZhH7q+u7Q0HiwKw0PLtqJpqnYahDS
xWswBF1lhkmEpf4mjPLzuB3pXOG4XXL3M6ZhxkYeJ6eeNvWj5NoTkBRd78sFGxrS4TrqTOsBeg34
0SEdXHbv7sz+h5AdwK610MwJNflpuvwucNFuu6IOO58ZC2k4sROUxcNSnmA9tHwmOUzNhbePe/Iq
wtaEtOpey48/SwmVvjIK64CL6LhNPWazbcY2OKZp97PFByVZVLhBvg5ju1ITZSL3ebItcCp1nca6
3oIsqYhgCRBfhlQlQELP9SKlbPeGCNGiXVFmCllkQZtw4lbzX8PeLkznif9cMGSqxiNy4g5LOODN
Ut/6XSbcoZvgPUotewcUm1ls1wrCouqn+I0NkhA4wXxvQmjF596urTCqNRCangYs6a21UY+Qi8vg
eQAE/0QitnYpxzm6KRMo0PrVFteYUHveXKUerNfhtV3uzocaf5aMeY6me7f3WII64imr5Njky+uK
kWhxrj9m0GR14T97L+RCyNRrzw3KAeex5IZJS+UZWjwvadcHIA1nXWflqodXVvwGFZsXuHOBfIMc
8JqB6lvp6v4gQq+P5LIBefBi5FfP/zN4UXdq1B0PdyfRpVj7ho6TDlARgeaH07o2kLGM3TjeUg0E
8S+5SNyl6Bud0hpP0Kq4/9UIkMZS0zcYfX6qOYq1YYh5V1ON0GsWYo0eakAc1lfq3ZBfVXs+iCLt
80/rOngkRMnmNB3dBaoihSIChVOtbj4sjJKfeRiTT/moJBY5FE1BnvoMcZ4bwnNbOWuBq9eEGVu7
yRC1rBYoJWlbBcHBqcn2TafEHSNNhMIzP7vM3W+HBjdSsZF+H1kirdeQB0cRw4YWuD/f7uzgfABA
l7guJgTHZ7WAn1lTkXsK4zRAnQdmGv3llH5RuGzjQ5gW3nRccgieV6k8bgFKrc29HUa/dGju1ouQ
xP/YPkaoGkIzZ0Q7LDMUNKOBT0hFuOQmeP29alwvtSoAquk/CuF06/wYnF0+cUaTEzciK68XGcwv
yIJ8wvm+iNlNxDXq/JF2toylnqFlPnUdVtPsyAlEXtROyk/G7XJ6cpCG+c/X9yarmzQ6OAxzt1Qf
8Xi7JSPpfo5lmPryg9+ZaZxEYqYCa4ENQIYmxCSkiKTphm7TMiw0Z1+sdrEJlYbLbjrkwh7z8Q7F
kBtI5WaJc0fiheVqDW9ll+2lrP2Fz/Su91SwsuYTBT+lrj9Fh5Ahb7u/UZn5PhHOtQRHRo1PKOlc
lDzX46ejBtoJg7CQWhqSV7YYBApYXgiW/cNoEmARDFRdqbIm2jcaWa+XDB+SfB8uEH/JNuaCNLxf
C+PeYCv2B0qAnVKWITUsgn6lo2kxICrH5kVVkwaXDBofjGwuHXTS3QmpBc58s3JoQr+H429bZxDV
fCtZkNIHh1HX4/JrizhFmQ/e1I6wl4WF3Wljrwob6A/gklt3S4frNFRKLgET4Z3DaogM/gepNFPh
LDYwTih8E8VjPY/D3ScqBZGQhMHIBAybpIx+uhsaHDx8px4gMo9tV+9GFMnahvbLK3FSc5Uhpsw1
0SY1M6/4UV7H9ToQvA9IYqbEwv2KVT2WND1HLX97e/Pd7kyfKKIXvQ48riyyzZJCE0q36fxnen2q
ibX7Yexeb7wCJlC78aCtKMLFdXDDVcPx2fbPcx9gfJRTFnPVCV55nvEMtmSktPfu5eqy3zn4TXuH
WjuEX7ekisCvxr//X0VucI3p/3Mdk4G4DFhFJb5VM+1PhJwsNVOsjyPQTEel1EBiobsukyOKwpBO
Yse1CC2rFvASWvA94tS6TQpU8SexMjWFPsbOuLAxWw4V5ttX5wlGOfRgMQwnhAzU8XRcbSuGd+Gl
Tnz8cEooLbcIY/Gcz+AVGuMbjo8FlFGGat/OOSQJtrJLfEm+f9TGUWK7C+dwAwKV7Kg71xK99hrW
kdv42d5ng+Oz+bJ8NaDLJp6jjlEyoz78J1GqrHr/bWQozUiaJOD01bTP9cL7tL4NWJRX9/r2vEmZ
K2B9s/elsZ5wTrO6/+Ev0CERPiEWz53mJzlwSGVePT9h00hN31ZErHm+t8jAEbkWBn1xWc5Q9irk
Gx6Fe6+6oFN59vXfj3OHgQSZh+YsX/LtTXHNfotmERJie3dk2abaAUHy36I/ZymXpwoTtgEV8d5o
fddkfG+VCYaEr8/tLEVOaXrXVuBMnsObX607OVCP2Vk0ixT8qseAdNInx9t0XomK/WP+GWuMbIaI
K2haZUEjxyrnpOvAE1clExc+svl0Ey4UI3gx+kS0in1ZOMiAPrxaxZdKB7ChljyW87yGhV6W9gKL
EWvHaTvoYMdmMMNAn4g0eymIN4o/DIC9L42jhnSottLs+q8wB9C9m4ICgGZkA8tsOhT6xAeFV89K
V5WbcGMtmOS+xK3O4jrZlId4vNwIb1Ul60Vy8T7Ll4AKpAoTqH+ODHwVPZxVBFZ1Fr5onxTzDMyw
jvwrH5YH93rjTvXE5s/Q0U4hiaH1cuosaUOp62uaMBs8fJVNqZislcYYccSZXUNPALtm8EkoQ0m7
fI5vmh0pkGrUc+8Dvwtdr/FhPbp76tAkw8gsXpjtGzNtaPEp1iuo2fZQ8pyKorjRGw6PAwG+jPdR
gsRPRek9QlZZXvWkVl2YOZr1bIozu9JdIUpvWA1JWfkyWO1KmGvq4qCE1S9Bilho1/gFcomH01vy
hqDVtzMiK2ydvH/mzgaPMJCI847S9WhJj5sDKPlT+1ydVZoXYnQxl1bJhWJ9OVPt1IrUZlbr+t97
4Q83DM8FGoVtdQ7ll9QRhv8aQo9YMFWdMOJcJW7nEBOWbyLYK4AjVCEBYoiAle9fsoc0q/ndz+Bp
0pTz628Gfzpwpj158xfy7tnP1DvtpxROBcrcDTl7mPoEJq8l+hR6i/79sa23LdTT5zHDoObkAwqW
dzK/3MllAryzOhxobn0K2ztOcXTEGIGzyeSF/ZX0Ftr0po+qvtNI9Y5iC6i/fmNLTuY4EjBU9FbU
/vNTHhjgKxFzOox9KfbJZilwpWnOo3ghgZkVmBaItOhC+1ZDQkbtU+c2FeEv0QseJDkbupOjhXKr
1L15jnSwqskqhZB3D/XTRO4Z3jT9mWtpjy/sm5XhV78iTfBHUL+hMuP/Sr1Lbi+/7lc8eTu6odIy
z2+htbKSXZwJa2WmxIA00vWMnwxhDHuwTBNwseWKEHGkgegGGYgOa9T2ueIW3Yurxn9wK9217bpe
XvC/M8ZptQJIz1Ftn4MwdUBJmEHG7TMth3Dr25e+AwLcWNBtF/+BB8QSH84BwcOdyRfPu5wJ9HlK
CsDVatHaZWM6BbR+6ir1ni4YGW8OgV0II2fUdwFdbULv+pZ9a7y0G/4I+pbDKN5gBSEAEDYhFvJf
wziiMKDbZcyXaWpZQVfDHkr7atP4EiVjTO7zKaeb/pB5xMcEqW6KsQCcQfR/qY/llN7oCoSGJ2Hk
GmQXRwF0Ov8KG7KZV2XyrEvUT5Q0enZGy52d9haVQdcExo+lcYGQwoClg0Zv7xO5YiHKzVM0qIz3
FFkOVjWYbq2L57YucpVucK6qbNZRIqlVlGB+lqoGeZT//kRhnQovT+OdOTrOGgkLAUgbARwc18iw
1MamMZd6rMkNpWpLqtARA0lgxby1wv0ftWo/CvlwD7cKwTftBasiKTdJoSmtxIbtZDGyW2OlDpoM
dACmynVn8YI5r5jfQMtXNw7rIkhlbfipn87zuFISBbyD71QWVwef4mth56oMe+lYYkoNicQCdWfY
zXR/Qw2ZGJlHlqi0PGluvp/3YdZYd+HtaiSCCfikLtteqjpMiTRrBAK5FYZo2j6/BZh0yioIvwXJ
eisWt6zw2i7rOZrJoR0B3CKGclmiy7MFDtNb3u1NEqSlSeNLY6VHdqLZhdwodOtZxY/Stl0cVLJt
ndwRG6Cl5YPvZJnLJZ01jDlsI81LHDzSAt1EIYN4jWHrSoJ4xCVZwHmij57Ovhj+iYKUA6uIbWY7
L8RyFNl4NC0N84YVGdtuUG8Z5rWb5ST+RwBCZ37SrCXEe5Rz1LfOIKqb7mBDJjPvJQPXc7XwNDOc
3LiuZo2v6wwizzqhiCA7Fjz/Fij7abMR2QLm9x6pkraC4V/LyRwjqUjj48VgS44M9uNEM95b1Wt0
btFV9gNKfWnhvLm4jg3V1xHkNrg3PnXSbugsj91Ped6DACojxbasWiY3nyKgspc8LP4vpprLQ/gS
IqDM3pKKzA1Icmvk7Njb51h7cD+mElbzLRmKE2wB5YyYzkOMD5TrC+7034OvhYkx4SexDk43fh9Z
CbFNmf+HaUbmJfih5iAY8BHpFj4wun5XaZgdFwl/0JKglVOnROCFZIy6qRzdB1271dQTbPIu8xIX
KHtLbPDiYYOXfR9nKTj085NBzlt1pfHeKxWNzutMesJgWX7ssKyAbXM9XF8OMQb9sXs0faLmgNnf
MzMWZFfRdk2iR5LMEU8lb90wpX2Tql64ShoCqTJePnpODKB9LTC9EH58WR3L2V/JthWveUALAXQQ
VNsjAgHk/xWfy4FJGIArqto49TOZI3fCAOB6xnvqfVJbmLgcIR3qGPW1PDe/Uj4qdHEyQGTJTWm0
zHK9SZjQZu3crf6UxTnp2uanLt/Uu7CB/za6c3cEM1sHCGnzVdNyKD5T41NuOtm9NtSLqQw39Aeu
ceTrP5g/YmfR+pDtpe7qgaMc0zso69u1l8vBqqEDFZX0DB95Ho/l/I+Mb1s9/ZAktsJIC3HYpONr
9oGyjWSv7GvDyqsLxH8mDmxeUX16kGo4o7CbSOp1GazNYtzcmCdAHz77a4Octekxj9NcoC671+mD
nsZ0gyAdaoOKEmey28YhItt30ZBNQhZ5O0nPAvnwUDaQZt3nbeM5rHA/Os6PeWoLrpePtlEWMeih
jVgWMzlq6XycM2ONCat0goCNgiTWNZwgGSZfIpg5otWBtMBpxkypZCcPBuGyajZhe26vM+cnR1rE
JJsXOb2RKuYEDT6ZydPoaQxpdf99mp63KPiHJEgUSXKAMILk1rrKysCUb4hFJNSSMwSo0i5Dugws
tjppOZJRH3bbn+ixienPBMiArU7UJtp5zWgIjdk7Kh6qwDdp+FlC+fc5jYwmgqj7VmLxr+QW9SX5
Ml4DeAR9/JrpooVLA+UAvwQOCH/owRCZXeAoI9Df/rQ0VgHvcUnxX0KLlKDXKR6HNPrHn7uc8GgH
Upb/89luEC9Kok9gXK14NpG8PsOmlZl04E14M0gHG6pekZvxc1sH0izjZ3PuB7u1MB+arovS5tuy
OPyrN2v23//U+hTxBE4HOso0FPc0FrhHk3G211oOtpJOTJGUjzv14U4bBuqZGa/9FnNIIFKjjuuv
wd7pYwSQS+LEHMncejm/oj1ZfHehTo7e4jOzyPSByVO8+iby7VZspJR3wSV9SZVgF1tBzBnAOWhh
B42kfGmQM/4RaNgoMBm4rB/HPgGBSMBEwbK7xQF+a14rzI7TFT4Ai6vT5jEvMDohHFBmdXelroRA
ibPHRkm62BRsxqe8smtiUazuIAkvrU33CaUdsvOwSLcD35Lgx8SmJpmBKhPhIBrVwxcoNHsFbMYN
jEiura/xct9ZN4tsjO3bHAS9Ii5OlCBRXca1iObgEvG+G33AhUyqtt2j+UK+/VpMCjXnH6KOnAk5
TEK8jvWKMERnft1f1pc655B+u8cUKyk30yl8II6eiQo3WHAXxC+oeHCmo2nmDlGVYHkQPgvhoAEe
s3ebn087GAqi6uJ56pH6sNw+/buMwI1LCKLbKoM5bBudKLDQhZx/DjkRtd1ZQNLoW2lstHAe2QYN
67pgRJWTl4mD0YWvzeA7cwEUjZ1o/Dy3x9J+FZlp841FpK50fj9c1Lx65O6BrX3qabIpVKoCMwPz
wez6cdgbwxNzLQoLkQSIver8cVxRHKWf7zjuIXRnzZxz7HwpwnEYaeVIMB7ckW9XwuD92+eP1GxX
6InY6TJNrQJJrX0N6242TEcdggKWGMuxC41qIcJgwl6EztrhEV7SkmrxsdT/evHd+cINhUrSilBS
pgZylS4K8DXBpUqNbBmF2d+U8yJxiDDjVsiU7f07KOb2wWS/teRXNVswnVo9yT9jxbJb2OEWBWH5
8fdquio20gYOU9m+uHjjBxGgn5z793phb0/ERK1KxO983lVQ5mCC0gR5oI6xAaiDKQxLgKycpYwJ
ZecJ5dEEScsNVEX2Ut/nF24e0daK6EhvEHytgalnzbqVidgIBDMXd/Sh/Pqf7XOVUDoPImKwubiW
hdjjqNQBvj3wcIh3X7RtnR+d6tEI/LuTulZNEE8/g93ArygNi8+mFbaC/oH9TytSKMCo2rXsIA2s
qD1KpANPswLxXd9f/iSbgkZ4ZSLbFhcjx0Bq7N1dhumTO4tgzZNOgHARBFexgYz3e7kKFmPdqz1R
oawWMqXEPm8GTiG5UlL8WdUVyEo4RxYoj4UbGUXL0p8+3yOw6s88ritbRajtkdJAB9vv9TXM+lyZ
OfqK1XuR0pDKJeq4vmbKEBX8VRvBZQGtxHKD/cWIHLNNN9OfkmXwmSiZr3tilIMhw3RPcPhEauCe
iSEelemYT5n+YlAzBXGYwV90iIET3DafYcVubVRbZzYE/EtI8Pylwongh3cgMtl66Ljd1kwllVHz
oiW1EA39IjbDSTg7vuSFW8x1D8qo5Q0wQkYMklkif+FYVFUoNxcNNJKSqoveLl7mqijTz9SgoqwR
6c1HhsTYckVxiIeYhPnVtdG6ACFOfYvvKSR2DPnSCHfreUj7nWEoJQsXWmZno5aqCrF7OU7731Xa
3zBDomUqYaGi4UxZ3FVPCQSIauHDYHsbczr6bj2WKmyQYdor7bIFvSPXL28y6IS+70AgSO+UvUKv
qQJ5c3B3Ia2C4CodhT978892dTx6ty+PKK+rYKQu2/06qhTyOcdecvQ+lc9U2NnA8DRRW5ym64jv
CHdzlFHBM7aDntLgKIZl97uiDm6nugl8NUN0vXF0cchpCCaPdvFhvR2KED+W3xtxt2eZWyXq0D8J
8pwFTmTEo3wQ36b+hyxj7xsgJjvfxqeuzk9mwJYE4sT9IwxEPpDWLipkFFocqLw/LLcxHLRdaePN
Y0RsddYr1YwzVDqBaJmRdGpbqQe1/pYyUrvGwrbb1zqThvJctdu2IFlG/WlH14Dz9QmiMgRqvMhB
lNwfFngv0YjDTaN0JS47KXQ4YBEZl/U5LPV0HjRT1d4ya9syDJYAdO8yqLbXGoZ1P6ogr/KAX0Qc
HcIa6Sjuf8nOfJwz1XkoULBU+liG5qdJ+b24nLxjw+6T9+H68wHEBzg11+viHkdNqP9XCqfDzgAH
wJEhYzDiM/LiQtkpUZG9T7ABDhCQMtIsg/sxELw2FPQosT/Dphev0aORhw+xI2D8FF8lCvcZuWUd
DnwurPPd3l6qfzTsd+xsWof/gVUUKCY6SanwPJ94dBwPi2bDXIrz+14KywrvUSu8Kn7hum8b+/rZ
rRFl6lmPNPR72LKPgPeJ1xIzYPhMLjPnLvqQjNKpUvp6WLL/C6YugTfUpHYVNUJysw53V3YK0SxP
Oprxk57qCjSnoXYJQdv/ujtTDkg6dm1yI9xPeQ1or5pK5ayJrdKMOSeAiyN6v2vlRHV091PKNd3P
FXGvjuJQ6e7tm4cmi19kwvCg0aXct8zRJj18CnXuz7TprtKOQzC99CGBcy26fgG1q3j9YI//rX0O
quhp2Ok3IV13oZwuceY5H7MZPl2/zkK7E4UbdBlw5ll7LeQHSShik7V5u2M9ZNbYc1F1Sq+PCz7r
4mtII+29roPHPxgeyei+Cjbgs5KpcPnL2askRyfjcy11C35WSC9nY34qEoWJ4mZwHfBeKM8NSlyq
9bY91EYJfoirVXWkbe0MU5Sg11Z0wS85ABbCpwPBwyVBsU3UIoB0rpZzLOKOSmH5oD891eUK17ji
UREW4h77/md3aoyflBAgbUNXnC5+jiq7g9qz1Ua2gvi6kLlvzc/ZSwEsSmY+965UjPctWQ5nKv3o
/6eKoEXF0Nw/hGPyrE+9qv7eWuoebUZJXOStkXJZJJRQOV7N9El01NEuJVex2AvWT24+P+RlsvMx
UE9JwUsf3W589uSVuYUz/iVXj2nTa6twm3x8Ek+Fx0iKzBCkrYh8MaoyvqP2llLbEzoa1zzZmbSM
egO1aX8igDocXKK7Ovz3hDks5f+TP2JpUlE4I7EAuzFni1aH+5+EYGLzfBip/kpNLX/HFCaZv/AR
9g87WaBFRuvvyY0DOA9apPJTHJlyCB81f8zlr1/rOPcdyTeCgoKMyyTb4jX6rHlnpjiAzozn5sAf
NPCMijR1alHGsMXmJxxQwHSY7SImV2m/pRP0bHW1dsYdHyWoJD76gvILBhg3qUb/mcudaSBo0YnD
GJHZ1++abWkNmapODbdHndDtOCvUaXezZdQNwLcJexEmZkr9NgFa7PCTAWtS5M4ZclYevuIYvNc5
ihERG193SiVk4HMU8b2VvUBg9IKw+BWpReggsHMXbUJmykj2qD57fVJCzTsglaawqeY2dgkPAi7j
+EkazQgCiRiMGpQZkeFlgrSUWB2b3KPM8E5XvGCAXg/ePByflaiOX3pSwGNlo1m33I3w6oMh1o++
ZLtsbXfvSqfCSyDxGrSq5PW1IJrH5oly4d7ZjOVCr4gmaGvTPEoiu6kpgghhYNvGD789Ar1vXC21
6OhKGbNzcT6Z2155l+DOww/fNDbtqf3iei71OsQ+JoFp3wPKrnS67UwXHqYd1rYkTFX+KwJVCeQY
Go7It1zIN6+Xr/xE6uYA53cqEEK6auiMLWYYCZOZcj9GERS0OteT68ANrjspwOwuimKtIjg/JHPw
MTHb0mulkL9i7OgNjByKCEw1xEuGBvl2skpwNKjBCLGloatPSuhkRJD00fz8p/Y9cxm59xUrByXv
YBXi4qLqCIB++scDl9cWTijEClMEVHNL/a555WarFDEcwfOHzS+VSW/Pxc6iMaLeTFdAZlL+BVqu
RkXf0wZhORKLTtVxZPF4VA/x983nQLHtOxdCMCXku/flteHsAvSCtCevdIGjPRGudhANUIMc28Yx
r7Aq+JFwF89melvZZJamB19gqI2YcGzVvUgC6CHKujlTKYh3z9N24rXcphnZn5JV2tuY3cuJyW8h
id38T3fPksJCcULIKCYLepR57bKIjLLMyCIF2qzKDgqCFQl7Ek3zgFVzEuZ2MN26CkCpKIq3m2Ki
5l9yoddKQoWdCRz1YHgjmxC/vUPsj2gNqByEO+7OlXf9cHdSUZxBEE1M6jMLH3CDPMgKN0+wnguB
tc6WIgPc29RgjtFkFWhZWVGUFpQoeA8WRQOfALzYnSD//4mULCKZiQM72kUXX8KcNCwBFlb8RqYX
796Uv/rb8e8v+i6+fFqKF5SEseDb4y3YeM5VpZf7PXUYtBxnIREjudIbNN+R8SONwIXx5J8keG6l
JgfsGqyRrTWpm2t+lwrCAGFUKZ/eb6LVVjwgj82Af6ry4fCO6Pm0exW6p+LXPVX8VDn5mLOA6N7r
/MMXUFEZeHKQXSabOGSak5yhGLEt6xHm0gVTsc9MVvJl2mQyUr5f63glM/3oMavg4nJS//JPapdS
b/VfmoWuzyVE0P0xD+PEkvHaIT6FaJ1MTFZ3M2j16knFktHcySR8jKsLYBAfVLUVa5ipMcAvCs1v
v+P5UnFOmLYclgEEIOVQBvdc2diLe/bHO9FWYWH9yC/FRxcHNvq/EIy29Z06HahcjKkF2mJicOoi
OtwYwmG1nuV2oYaqGBo9Ws+RhYDJlrJ31Mp+FMRx5N8cFLCyJ0JyCezOe+v4ViVvu1NGLAnjfO3g
UV+zEUr7AulCOo9hjIHc86nRXdG5lqqHfc5jq8+8SY282rDDQRhS9GuwI2+Z9esKr6fBXfxRRN2h
7hirSh9VVnN7+VdjUQohn70Kf5ZB6Yu6oGUSfKqDgxrOyl9LNij5FoXuyKrr0br3mTTnfcYgxChf
A8yeVWYucPkgnyaGu8x0pL7TE9F6GJNMoU3Nee5RNK6ZnNrXRRAkfeE8KTZjWrFStXHrIzybquN5
B/m+L2bAhztIcjZqf0r3Zm33Q5BQ4zn3KvtZqT68bEGiKOAPDK1V6R/EDSouawvj5SNPeIn+MZuc
CnPcE73t5EmUpIZPF7n+c2sB+7AyK0XAOi6Baak211EipbQDbwkHmQkjkRcA8hyF/TALpAtCZY0N
rR66HN9EJRJIqnGqUKFg/AfSWupHp5LFc9UT5MPPLNLCPEncFEw4yN6fNotTcLHYNB3rlmZ5a9cA
LlJ0TIUzQrvHrtlbY4ULkTzUcPX8qgHd7jRQxGouLG+/plqi5r5zo3uov5GRf7xtzLEFLhjOReVa
2ONgUeWtwVfP5WsU/+vM1j2XG4LuqiaiNqUeC8dtLWycMm7NOShlCToC6MSzAOg83fOVhMHgVf21
pqYXUakUzVvkLfIelUi6Nl2DozExLTZq1NS3DhueT2qjm3erebk1M+9Nn66QPNdD9ChUu1Jg1xp/
Bu67c4b37i9IBkulGTQ7c6T4h1cmUdOPauXGRtx2MISxQEcxsa/hVlwO41cPdpiJXdCJ+2dNmRb6
eK1IsBzvbgERDS8laDHhr82VsT9D56b8SQE4jolKrJWrqpfMn//SfmgCux6jW3OQQtpF5Gp3rmAP
vS24TNdFZWrfAqpuaBUl/23B2dfLtQmW1GXC68K//N1oZRVe72VBfly1A/LcyytSJLJ273J6rCAJ
DrMOF/Ux5rm3Q2JBX+BeG+CJzhT2aTQB6vj8PfjjWdSBRKSGqOW0cdroPnwrrCc+fzyVl1MKvjpz
8IkCUltGcFYJDtKT3Pjy7xv4KPmBrObFiA62HvNaqr9gZj4bWkj2oAikeELQI7u+I847PdNsUzW4
FtTZ/E5pIGQXNNcGGT/poqadFQaECB32fbDQZXHbp2V5Hfphk8004qeupoZkH6m/ltPgG0wb46sM
BnlHbqEwxooAPG+4N+A3Hhj0kjtk5ZM8AJdN+tRgVxyMWDP5wM2o8MDEehgxXXq2aqXcsrwuRZr8
spUxODlshrqJDzbA9Wztca/lyd3UCsfm3/1ae5qpxL5VkasGNx/eXPFgpKxk/3Vr86AC8Q6VO1AW
C87xwQ9Xb6/7nxgtunp3lOkbky4ohL7rRZB5uNglTLejGQjGC8poFDTGLux1O42HXVytk+NolFBd
offgYfbB68PzIUK6rH9jbqV6+lXbC54e42UqymaoOZSjNe0+OcCzilM8UEzG5DpRGwMhsriv/uoM
dFrR0aExJ0ngPMrP2SuudJ0hY09vcaA5v8/sZNHOPQxPwFWk4ms8hAW+PEIl6W29UclGda9Iwgz5
mVWbj/nHw6VRTiSY9/MCv/2fxy81r9bP+V3jjWWUEgrsiVXTrLK6uh7DSLBydUYE2XubukWVNLDV
H3qHjtqMzeJD5Ll0suCWiZDhujJSKHYrb+6Ls38tdtqbqxM7js0vqrX3xgOSI2539OschVUauS9g
0e7hf03PHW2820xuWw3A3SJfoLY/oUGWyePgG5WqgqUD37pP9+LiI5WiwIUrMw1zE0VFRmT3WYFu
EY/cQbddmRF9mdXWNQQqb5Vv5kHIKDIB78RFTXD+FaugXKOSuSRWYSa9Hx1PkqIaT1+hZOAqZBbZ
l8qCtKmPf4OOMJI+ctigdAnogC8nHbBvcaPvHR30We/MPsSJhkPMCMn3Q7foN5VARxs/c5cawp1/
UnNyLsmFYbOatijXoG1aXi7GK+r58GEhQiRxqPYRqRndtCYuzoXmp05VMPOxD4sPUckplCFCcOfE
+dXhyV1EasIlt1GS7Ifd6Ejatjnx6Si3JEJtPTLvVcYoI/MVgvMNAdnj7ddwwyKbZd50cC5QIQyh
MtPObZfyrouG6UZ1NYMYT7RoZkygUVvNKp56kKDPS7EftYyuOjQkaJOSbSw3pwKBSuLPf+S4OACj
dV2uPF2EK1YMmDX06WCNncJEU9qbXGFYdmPQxsXT0UutZUogMMuFOPkJ0KqwWD4mI1mzAsGEpb0a
v1AP91mfQaTYdFhcd8QY8hLBQvNVk7yn4uD1oXQbG6+j3qYdllcY9gJeKYm7BexmzTHvvM6QXtN8
Foo3CenDsPYpM7ctAN9e6+5/Th7YL0EZd86e96TQvt7GXv+5aYY714OALQujVorT3OTwbl605q0D
5Y4RyOPmdiro2W6xuUIouHOzX/KZfyHvUMDtTkQiaYAwtL5Zonq0MIHQMH/fP7GPNXDJB9142oPQ
PnwRLZG/CMtJEjS9mMBPs1NV5hIaVhqOi68BmwlwmVS0U7P86O7IH0v2PUMTGFyuMBk3aaIh8Yh+
FmDYtLgScHlEZ5e13CjEsaxgri3UIxMo3vnRxye3sPu+J6r0TjOAKR29C1A1OJjiM9Gv6QC5Kv9N
+8+bGactVweJBEf3K0MdvgU1r3i2keNyU280hrfPiND5efHjanV3NusFkP36/N1RIchr4XfEcF05
frK8clM3jUtID992bSiCe7vHaYbfOSRd2x8uouGEb7gc3rCjb2PClOQjyJtVOQCOhBj81MnIpil2
V+w32zuq402NXn7zbrvAEDIStcWUMYVKBOXPqNPaGYW/sXUgePjazqiS4rdgH1Xwt6YiLUfTxfVr
Zwi47WZ+KDI7+qzM7dY+ETdl9k+6LzhUoI3QG6eT5kE1nH2nKp75raAjMqkkYF3D3vwoEJiqniXf
AInvA8tqlwqkFOszMtzP+cxIOkE1v1JPLX93GsU4KNQ5TmUGbSoj5vlfNODSrSwt70QrU5uc8M/a
25NfK2ajCbe30FuCgjwqklCojM+yMgzgASF2To+XIUCJ1sTPuPrC2sI/X87FnCvTNvPj6iDSm1W3
Z6C0RZq0pYQJxt+gAvgfqEvJ5j6j4wxPTnjnFWDA5Yqld3c19M0Tl4b68yxiAeDjjTMeSBnwPGt+
zOmGb9APOj5k0C7E3onJnQ5f4NFlj1tx/nk50Ge4ix+vmkrpj8HCUvBvi931GS85lQesSLxnk7za
pRW0yp7SR1U2lbI7Z97wcfN/7u+t9je8Bh7rca/CMO/Vm2guj1jcAhzCn9wXBkRx4Wk8atKYEEMR
z+oz92M5iI4xVvuPS5fHQHUGeBRs2bjmyUTX7jR/qQ5YJFoBzk0OA7sWHkzs5Ju6XD30iCRx+cKG
H1aPpXOSYu6Q92vW603fxJwWt8Q+ajIpFVLh2UzkF7xCWVLNZihXsi9RVsdXx8U9yTa0xllwMO0h
YhyDfxVPxxtBt4QzgxaUF8zrl8F+veeNhDacEHOtsxUw3CIevfhgs9LyQR1rC+ZOdwViotQv533D
DQ06O3HvvwZavyI9ogviS29EFlrCy486/jZj7AxUsS4qeHzf9VPHnWhXgYPRK5xU0P9IuN4NkdFU
90T8Qg3jzUmff7dG1PLwiTDuLPkcko/TCkgHEBgz8IXpwWFYCtG8kIIO/K7qzaNivZ0GRMrk0AFg
k2rhErySD0dv0kvcTu+XYPWyA2/ErPfVdBpkkL4KXDUP8rTIT9KN06969428boq0u96SSt4Pxipd
kuaHUhwOQpP0DFcFaovOetIxP1Qlri2wzyUetFv/PEQYGXT5o1rsjXyKn9qn2HEr3Wt5j1KShQnj
CMgRADN4RrfC1/63gAlYCXoaeKUAvjXpD2OvMfUmngEMpqEI9dKErTEHzSpx00aepZh7MbItKF0l
1WH6RuYWdfwOLs/1tvH/88Mgjvb+dkTS3+6HlsaenEJSFDGfnJWsAOkgCnCIHEhAl7Irzwg7+2tC
iLHhZedTRqzmGKizPKjcAz3kM1jkFBHFQxyUKna4dHiFBfskMJDGFyzNvoPWuGhaSFMsj5TkTIxE
Xd9MzX0GAAWyv06zjaTvW4HG8/hhUZ1LvRnK3cr/UFPZ8UUUHRiAVo1mWJm7akAKfNHGd+qb7CGK
1vtWtpjRu6ZbrQ2W5jEueoWfvc9RfIHesZRwobzDU7D7/SuAm4lGYYSgNyudAF2xob+mdnq7S7/4
bctWGpj/yoZrqUTmgKlv1yr71zUd54FPt1DRynLOU8A1d8sNuAZLG/1NF/QfqtmcuZmR+vpy+swG
pBoIrUoK/Pjl/XmOjRsZJCCNf9G2nJSVOR8gzyHX8pYvWD/K4owxjoBEbE1JuQP/H4rOOEYMeFrH
ZdfEJjRllqj/1Urv3C+/cgOmLfa6q2LQt+wzT9GcaDrnOoozKfO0bbeucLVvDGvZIplLWlOWP1zy
4yo2EvrE3EsdRKRjh3BwIhBklYUNmpUuG8ebvd5BUJNO6YcRLyoAzuHlf7xxZBQhLvRjxY3cd05u
rZwW7YPBRCdKKPXJHEqCfwKqxKtSMFb/kOQ94B+0wYOR8pL4PAN/bmqx4MunASyt4N2oUCsMVc6n
a/NZr0gIWgX9f4AaVWFaDc5i7S/rbWkxB5iiRohMdkXoChx2ZZtP7vQ3eTZMTyS6Ru04f6ap6/fd
JayU1rc75ydmGgA4mBNlmEoqNoECnt1OuNRgVrv8DNdnsND6jwRgluqT4+C1hDKdhXAN69eo6mBz
ZJeqe4sMHxcu4ILjj3AzhI/ZkwtwlkN+MfK5Zwf1Drk7g1xTC02xm9gaw+IgHQpA+GlpXTJqpl4J
feDkuFc0dJOgabXWL0psR8kXUDORtIy4YAoekNBbm5w+REM+EGaSORrHoP7A3cfkV/Qrzkzxmw/r
cUpJjfMUb3fYTaCJklAj0j9zBh7wM/UR/i0Ct3wa5Yh09WH7A79TAH2NB+K9E/kNTOGrZi6monNf
GW8vh8ISGd5IoplrNn86p2q5GALHeJH/X2TT3gdsw9vctU2Bl1cjtfksxJVaXxj5AlNBMroo262V
tKikyn/lKvbaO6OlqAcpefqatZbt2wIFIJIZW3EIN8WBpuBOhXPXq5TsaIXGEo2RQ51GNoCZ3Xx5
nASZ2e4hunxOLJb/NztOlH9TiGkom0x6XdSzwWNr3sswqCpeesojecPRpmtMix0WLNm0CUVrfLv+
FUedBf8/7wvoevNIz9A5MJ/495adwHRcVFOQlIpMxDO2pu0n8r954BNx6b8WKh4jRISFjy6JEGXb
hkLl3QXFS38Nl5o4QziaP2/QBtVsPrBRU2g9RNteay4uyzUW0JH3sTtP5TmaT/K7/KIzs5vERrrD
jbzc6zMLHeTApNBZ72svpmZcCefqQFPBwwpPTidbZzYdQjAgnQdFVcWrMJla0yUkOpWtieu2xccR
ds1HVDe+HsODCR2V0R+8QZKu9WWFzqNFMbjiK3G50o91wOAI3Me7x90awWcNDs9pO0JXikfhw3HL
TcLldRd3fsx/9B3k46gBCBg3wNKpHPpitFom/yXPptzYwQXONSikGrMjFHE2mLXS7alWHFml5Tst
dxm3AJUasIbu0cIB3ApXU0g//rS2Th0l/+VA8pw3m0NogOIEVZ+DnNPA/kAEAteafM6jznToRCqc
yKLzTJkYsTqPmh7uS4iucl1nC6f8wCW8YAVE0TrTfZNPowYf7AOatPtrNX8tBCau+Wcb/KQgHYf2
Gcf3m37XeWirM+VJ/3M2Xk3fKLBFZMr1WqeZvsdt5ycNe0KoHgzNsTwr+T8zVhbhAn2WoIyj3yKJ
ROhwWvMrKbqJDDTG8E1u4/3dXY1EC9b+8VYcvNixcC34H7hAFqlMUDdFooPwOJU3unJZay8zfDPZ
3IiaUex2BTAUPdHl+SyU7mkF4YnK1q1PqFYWqs9Q+naE9Q/olVv5u+NMMqXJSFGgPaBvEgR61BoV
Z9TwCmpDF+n5hi2O+0FCnBOLgx9M/wXO6ZTtgIFtDPI4Xb8h5tjYgcB3NIwUL7D27oHAuM4x2Oa+
hm8EdIYEaklfm/L7MHYyPDszNOj6I7YXRkx419KAMUxrRWNJH/aGsceuiJUPfgdKFwjVdwQWZFJs
ZzO1z2TQLx7Bt/i0JKkOn2cWcIirmoktnzko5hW2vepj8u+RsQjAQ0u+z7tyrV9NWgoUNpquYS1k
MvNj9kIwpesTm/2Mn0DJcYuuceduMamkPB5s9RVxmGQOyZfvay8KvISO2mHjQ+WQ+y0e28km2eNC
quTJmoWDNQt+Du1+qwNK+dLHcUfLJVvuHHfXdrwEn6rRZtC0UEuUG8x7RVZNYThiqAAPVsLvXVWi
FLSAuuCGnb++VSt+Utuz+MUy9m8bxH2uFKepawAzHMOn2UpYrp/FgNy9Tnn8CZvwzm+mi+pskkVh
PYIq2L8q6R/B3Pu/UC7ZiKVwYrfUAeDHigNDJuvhFULIUAhHJaAOTrHYCAPBbN9uKAw6+/wCclIf
lhzFTrejSNCzm8krrHh0ZDAyxdcCOpwmlR3+NxhUBfUPWoNT9xSw7IOkTNJBZLb9GAlFRfsdo6E4
7ChKgUmvluNdUoZ+XpXzjLTXsJAdWVDamy//7E7RCl0gARtoCq6x4mO2hLRIa2TKNU9c5QJVTv3t
gNktFtEu83AcHDzIwTfXpOEreEsuLhiJdOXPHu3U3PPQxnI5ptTN503AHZXhDHhn/fyoB9uUEiSx
7UPPFy3d7QHIeSo0m3uEnTw3SL4AP6VQF9GGkBX0pwo/MpCWAfI0W9c+P0TNjtX0kQkDTLQFy8S4
pkAqcpDxS9k9fAn58wjh6rP3gxLURFUAz2qTCerlz0m/BJ3t5RclYtsc4gNxK+kVukxFj+F/VEJF
RD3eG1fvKhMdTRqzYwSP7wM5PRpy5LpYaiqiEe+HPQvB7QxO9W/Ipktv0IRPeAZr8vXRLH5GZLU5
8VBDVLDKNcTKo/dqg2nGiAQf7OHB2Nz8vJFmmv5aNR3mRucmx0brpSqXuenqQ4cTUdVctsnl736F
DELz7+73x8+2mDWE5mQNYxziFC7GRo3OVyPMha/XeCtcMVZMq2A04c6VJora/VG6My6Q50A87Mho
/irog+wE4x2MDi/07VX9+SgzC6RqCNOHMP/LBi09MG1GoGmowUNgBHq2u9YqsDC80jL3Lp7mE/Ps
6eU3R87YWt/xHniqwNaLVaOveo5MO6S9F6/UKUp8TfhrSHiOkR1tNXbUX8TNvOg84q1qqKghbSC4
3Ht7JvawgitDIV/ImBEJAyAnjDUR5d8SrUI7XOsnHZuiEyXR0iJ7OP0/lRbyRp8UVQ4V9h1agPiL
iHRxAZWLT9LB91Bedz/CxND2t8nZfp8YMPsUlRdxAm3ftqEHz42A/024KtRATP5JFVq9S2oOgFH5
dKXdHchx0fbGWRHtPiAxB2oPNxe+bk6OK/6W+h5zzz3hKGTZtyi/gvo4XjLXK8f37mvOdz4nOQLt
pfbbf33yNgwh7ZShMBvB1Ox0GcXLSO8VAVxFvvXIka6dylzY8q7YlE4UNt/q5xFlq5ZGXcsr8Eo8
lxN6GdeevwtM5B3IY+39cUUBs1rIAvXc9UchD8TZTu8DLmVZb4F2iyjpeDpKCLio00Zl49z1DbhF
jFqsPN3XDoNnlwQpX12bpE6Co1adU87tpNm+xBI2GoelIhsbmCkkgNMcjecEUaLDVLfOmTOtJYq+
gtxKU0jm+yYQw3zEr3jQGzIcY1Y9aTOOzvriLAaC88SWCvgwTBizBVHLiLc/+j73h1gOjVY560WY
X9hU1iiZlOZLM0k7uy5ndNRp2wzAM8z9CRufoLzH2quIlX38BpnrXE7Dd37QkyG+ISNf2gGrNvol
VKrjCFY1Sug7Fge50KjOerdvtE1ZBDhXqt2CkqowhX6APmwdYgOYJlHs6OnZcDQ39ctH3Vy4MIwO
VrlIUJ7V3y88pmOOde0lzGUveK+Vv+fifdUFvKYsGSNhinqnTnhppX9VBk/O9F/ghHDWlWTIgJaZ
Oh4J+MoacNeFSpaTHFZ4nUu9XIAcD1WHBloNGEMXsQmNCWmy102i79YHOqhj5fOFP6hM2UEOkG+i
lqLe/t+TF5mDN0sdZk9JV6iyw8wf/UzPteF+L89ZQCynKXpnAW5J7onPS/PZpr0V3ldfhdcrjPN4
Yw1akhaqkDtbSMYEf5DG94PaPqrxAQuX/AN3Mp1M/WUTpg1JUAeBCiZ6RlweVIBiCsKnxCEI0eQT
4AtFgR5FnPYUXDg8albaVhHXse8aMj/fbbpwLZ0Q0cG3nFgOFtN5plwfYPAxRpBGnV4fr5XW0eiG
nB28Sa3cNpIaPLpfDEGxtgLbu/KGCv8kWhzaXRqecnFsjcw71aAQBTBzXT2vtc0lTzkUzcffD0es
2T58LNYkspRz7y/Jwk/pv+5TiAH3F/KD1Yrd7IRvG9DzHeQ7ODRN129iHHyESFmpXnD91Egt7BNF
2Rr/P27b/IYW5hY7eayYoUD19Vu3iUvjNuK6GWPCh7HbhcT6FibVMUhKLXGUASW08or23Af0wLxF
R2A93rylvHAXgapQiJruKAqzYAh3N4CBo5sS/bdbNAbFPJQq6je79yY/UlPl+a0fCPK4BQv8HxTF
fHyZRWaJn8r9ozYYx0KQGXJDHyBbDHs6YgbR5vGNOeWhjwNG+o8AovCf54+ZFnsb6K4esH4CArrh
dwMvTjkoHvvoGYDU8rnnTVA5x48hoX+RcmUA2b/Wxi1yGqE5uYGNxIwh1rWaTuGOo0oyBA2t6d+o
WGuS+KxMbtBSoMaIZQF8b6UrPssCnEJfaQSphKKmmSolBR0kqW5B1VzHmeLVM2ZVL7ANPqikma7O
XrTKMR1mP2GaopbfeqDSlTMAoBlfJo7KwLh7lyMI/GDkRrUdVs1OT3SZakske29243hjak/Sdi10
XnA9e+kE4GPau44PrGjGBcONMnnmm0GRqBkJOuuMXsAXOmhdQzz6EZ/PtcEkZs9rLGKmQhcA+hZA
HcqgFP7qjT8GH+QyQKWvQVB2vLAXEvAh3ZuOxQFVNmDIeWOfM+ziNED5YqGqQ50YuRyalgj0ut0k
QM6nL03SQlxhcqmvTkVi28viEayqNbObV6HDTTnujHXmLzyhs+3tMq41SvWsLd3GXhxnZfSAyKcm
GohhAUt+t3Km8+hSlRQTLbPGsZSCHUqlsFZrtjXAioO+ZMj7eenbBZU/mq0amQnTbPnUfmktqIwp
6sArgzcynsiQwTOCFutKPe6XbK+Z66tX0E0R8WeTZzFXdJRFyXwKsIF1Eduhs0OekT+DjVsyzpT/
tgNJte1xmYfdTaZ6+Tblv09tLc4T+1Yo9MYm6VHZpA/PG+n/aqzi5UAGiBkIHEDrKK7e8wJwx1WZ
cFcv87BxZF7a2alZevO81E7R9irgq/VglOyFH5cdIAvTgqXtGFxAAqyeRR0TiTZAI4VFUMF554zZ
4tzp3n0r0692ETbuaxU7G6mys2SGvfgnGoPJ1Ikg0VuRV3cz5deu8Gx/PXWWB7BZGmrO7e+EtLAT
K9ImgO/VtTC3XMfhJb0tUgo/z2NSdePKdf3t6LpNp7eV6ShuQ3NK94DncD2lNqdSpY9gyfVg1M59
NO8DKHaxm9t3QzBXg8IldjpQOGZgtGv/k1gnykTIIfxPXudYtoGZaWz/U4ZLtx3Yr6MSqawkf4q8
ggdRuK4rlP93RTQvVjDSH/mDPWD9B3G8wenvrmLvOLS63tWuhW0s337X58/cdALBnA9oxiYKqb/w
p0WBhFh+xVUDQ2F92Vq7NB3qPUWbV+oDXuic5mdH+hIpjIo72xp0c8vbj73sj1Hd1sQTiAAy2S/y
Sl0GK/IazA1qOkjvdlOyK4FoUhsC8BMwYXr4h1yQhx8Mfawf8JuVefkWKe2ua2Di/XPYdijpfkKY
QzYqGqQm+E6vjBr/buVlKErJq4nFwqSyu3QfMt5/XxBL2xlwnYBiPfMyG/jZplHk2pPW9P1beGWp
qln/vJPO8LsZTHXLUjZyHhYc6oK1VBIbtkrdMaYPJz+o4HFRPZWNlOQpq5wvRMQYvVamPqPuUnGp
8NFtv14wwmWhNn0ABRgRrUZdAPWy28Qoq7w+v/w1ZDWVBXqe61/Bde7NqA98JHmNo5lAkMZ9iBBv
GS/H01wIfZBDBzIWh6iTJzKyxQQr6GrW4+kChMTNlnJWwn/QsqtJSgP1NRKnssRPi/RO1hKXsSNT
sMMezBp9qcpZnzeFAZlVDwAbasbzPkhceDrUYEyk9xsrqDwUwFDlWR7/3QgHjE5VmzCUipkXUqEa
gN0frkrQUfiryM2CP90MO3hlpPQ3be56xZnGjwxBabfkxnLOPQQD20rUrGlhVMJURBxMZq3S8d1J
Y9/33YL2IbeNM1/j7MMvHmK4BwYcimUHklXNRgzKM9827JOIq3ZbTzQGnb1+cz/B0zRCP0KrmVJ3
SFYT0UVF3biz7DJPeJppRcgO3yeuyobyGaI8xfkPi1acdzHFe/ye2RTsqLSUujh5dNMJDPLCrjo5
fykJG+1JMazHOua6KZhMsqsXmpCLrfgp8c6RYzOzazgqWTPBm1lfASkcOTkXItWGNjaeg5QyTM3S
mnrKl+5xaC1pOUds2YX9+xCpll9TIKo3p5zv9aG2F7L3Pco0HSK7T/1ROHdTvNyQXbK5wpzYBayW
F4bX+2ZOe01EPwPgzf0R6SREsx6y0jqua3fDpSKQZgUpEaA5Rz3/4OH05m42tMNEy6IdLjthHbjt
pBzJ12TI3PIZo2DY/eR138284g8BpHkI5E45hxUmx/t+Frp7BKnHslnOxYH/Yt5TTfSQxH8kAPV3
M4JCxl+Wd26OBj1kE2sAPYzNc9/dTeI1CMDwY2pZmrN2UMJ63K2qXa4bP98mZOs8ZshtFstEtmN/
Zm2hfbDlroTZmwG5J4+THlqfQMeQqCbwqCXlpp+kRZ9k1bx2Qa8GfTH6Y1SBrm0t8f5IBNwkjxOU
QOjc4CXx6leJE5op9u7dw1ARWknaM+gyUN8VxF+dZ+Tw9fEeWA7KEtaFeeSss03n1Fj5loXnU2sX
V44jBmJ3nzCllV7EW4M3Wel06oIr502awm4mUW6p29pf7cf5CdLmzG1LykZFPPtmVkGKVsHbovWh
8QqqYLxD7ZsVPxpwpjclKAve2sywa59EsDl9+tLq57Ywr7DuQ6tm/aBfgRAOlyKf/REw9B4ajAoz
Ahdo2CCXLrsB/dIL29jfHc/xjscnVsHKJqAl5fYDmN0p7DWcxJ/SQpl0O0Q1aTxzxVXhUq1lp4RX
QcFGMvSSi6iT3DQuFtbrmB02JHzLG/78MKzADYa9U9O5nxUG3C+dca5/nwOpta/ffIhTxHevcRJW
xDasDwRcHnSRVEnjChfGDrkSAbVhxcmJBsUCQ2QFSojCpZBxr3fqLRQlT+xfYWXfhfkq/ZPYVmuB
xR1wK+5zWEW8X39836nZ9Cfn+NmcegNMvv4P81SZO2W+l++DEyIkQ4Jy61cFJjD8myi5Sr560X0X
XN/59mkrXDb+U2vKCUIUXOYDHwGtUi+WQBHqLnH6velmsA9VIf+rPVjYwyJxYILoxwTtCpKBKwrY
KrdSdposWuSJ7v1Yq8aZ1SMe0VKRFEnz4WSImjdeopNSznMQgqHRFKSoR+RJtpjCwBkSNsfJAGF6
DogIaXrtjx5zTQZPBlcKQl6XxiJM0q0C4ELXA4pHx0Y2lESDg9H/rlhhVrIqJI3yvIV3wNY0ZOlr
bk2QoS1IuIvCUUg637pkhzDFI0da3TsRVxS4g1FqP2FzdpAoUMfVLSnsjw5DdVuAMnVcRPrd12jx
PU8bwSH1fLFdkChUCpTydesdcjxj34APRRA6Sp+BcIp8RollNALcH4YboeQQxQgyURddCiTjN4pJ
UZLtKBkd1nla4JyoUcTmiOP3+WZBkt3Hqa6EITS7vkJum5KmRmhvSf0zX8IcVPQagxFJj9fXHcbi
MmdnaKgZNgf0SDRN+5tCB9oGEoBwT50kbWsMy5wC/Sssc2hM4fK5bz2AhZ89g90HRUkGjGteHIBM
n9Cq1tm2fIsGjbceZ1Sx2OY2ROuDy4tjI9Vp7YQQgcgEm9x5td567AZEAbfW49HU1kZqMDYD1S6/
KI/qOqnZY3hoUtJ0h9893tV/Ze4ohZqWLyMXYntvaPlIvZ79zomvi4Xt6/VG7r2mkp341dlH8Lie
7JB0lcWPxW0qd3x1LbWu+LRHyn0mFyUrXNfWCeNHzhhOg3TrZpZgMc7Ib8bm5qinjgdxMPCD6uWM
jyqeGek9SLHE4jv8sZDkrSK9CdvGPfhbLlXmzQ1O2helpCTGMqEuWuUiwAheKeMfmegTBlV9KPe0
d7/4twhopzExjmdEHwGSY6rYhv3pPRQwwcE+PzlJZdxwseB69clgIu/dRS8Rb8fONAjU9HcyvL6Q
Hs3m8SWhc1jrmICS+kgbkOhIrtgwKAKj6NxoI6WD0xUY0TdiFPgHwTpossu/4T1NeJBe9M69+k/w
aOBCJNqiPjRwDQpMSc1YApXV+9MO1xKdjFq4m5l9wJdq4MY8MFxi6JfAjOAxK0gOpCAAaULlRCZU
Vodg5jzeswzGHszScgjbN7tUdZjtVp4LJsvA/cS061DzOUnKOHsVadEJXPTJqaAYhgQQIKAVyUdq
ORocx5ivdsxPimB6h1HaO5ntfKZABOXT3kp81gebu9KIgsmp9G+V8Yg6/Jy0Kh9ZIY1Ic54k1WK/
m3cF3PII4FM2G0uknVK6mU370k+XZ7bXr3t+TxvaAAdn6dbrJ2ulN9s9UNvdzzHIIY81BsgTqeLq
845DeKSQ+nNIbAaTKG4qiYBuUEqRu9gTH3iAVV7Hl5xHVsMLaLC+IXQF6J0NToDS1O+3qYPHBhLj
4ik2zzE9GKS6kZ5fW9CJ75wvy80gF7YknpHQRmWpT7xf1nX5Z+E4+dsdFtbaq9aIc+3IddlLETul
e67TCSyiKa5Dol3PhqNQczMpqM31Q2siEXh5iVmHUunamzP5XGU4ke9HYZP2zP6sfensE/cmckxA
3AggejptJ0+Dsg3rtB0AlHya1rtzN0irih/xsFyasBsZtTzRF573OvQCRzTt7cpRIAMrTssVJogJ
wyVDuWnLaG0W8IrY5FWkfsCvwuuQEdQCc5JSaHEK+DegYwvBFUQkv1Xx4psNtX7DI3V7o39M+WGM
C9GQr5ECZYDnHCKbwNWzCAH0gMqJ+8LP8WaPi2lkYnrmAmYdZ/fHib7ZEymtpG2f0W9W1J6CMUsz
E+KntdBRhY+fkjz1K/wDA1WSOHilknIP4/PjMvAykqRZXrS0dgVCiTkXJ5VkAoALAOG3d3G8yazZ
Xvoznz44oUHp0jQXghGGtxCxoFKojW2U8KLXwEPa9w0ndwlK7F9f6jQef2o56SUZmruRmYvPTGOr
jXB4zi+aMpa6jWlDLXpMIWciBMpU0ZiGeSP97fq1yoqT2yeBDEz325YTOTnZ2xF34KApqyj3qY1X
SFh9Mrn7d/vZfFZscpGetC3dN5jRlRcw9qofRhr7xL/cqoXafxCHJI3uUxkjy7gv5ZUYmfvDI0lQ
K618/cIAMHa566dqE1nK6KNtF7A2b7fG8iDkKcsOmOk3YbA80vzemki+nZhGAbu8Gq1kjJWuKmz5
2LUiVQs3k6BshjkEGQNcOLtZWZWBADGSk+rm8g0ZKlJy9l2cDyUUGt08Kp1d0j+EtrFuF+2rztxf
4Z8jtMWLblCf64ljEBrB+wvislJ1piTFyrrtIRrJjWwrPxHqbPuaT5wBVT7Mz5wZcm3wbKwRBspD
wM35JS+CJXGcXj0pocpQAjFJZcfWrWC/EOQD4Hx26uA61LWujERph2egpTvTVbjq/v2mSvetZzYe
h6lvuqgH/Gj2FDeUZJyasBfQI8PPRGu8w7rO2imIpLJts5/oFMVFR8WMMHG1LqnusxNIa9/kj8MT
JEvqh/4hMFMThbT5+2nobnWXiDjFPYlWrn61UpyiRQV2BJanIKST5YJ33erM5S9tAKX1l25Um2Ll
Cy1Gy0PnHkTd5UzO33Ahdbb7TQoHUD45lcHCJku26aeVfBVKqAbRpPrgeNwm9E3tAFAM1jK+uQrO
aLlAWbMsOlohnIHKpwTXY7z87F0Vkasaz+tR+9TyOy9ct2MSSEG77Yq1glEM1KeBvvi2pQMncoPz
UB3Jo1MY+JukDufLBvIqDIfluMtTtET4iYc8N3tU+msu1onn83yYuriGLDrHKePxKeE2Uc1Y7sVg
YJsAk5oHeBGKCYI04+GlMlz4JRbiThZ5CurBeIwjVaTFen2z41KKsEyR/siqbvmASH4CUz21vtAc
V91lkiZnrns5j2qkFuVl8Ot1SKUAWJw7KirI2zgZ5PP2dA5m2fllPH1DlVb6PasUUNuozADA8SN+
NT2Fm9nUO27jmQybHHBXFUMjGfkTYEDHX53rHxCzY++63m4mPW4PGTcNU2DfufXmyqWVHFO5wp8B
cdXdBqQt1WaDFf7DwWaCGHH2KOladVNlMQUIwmdmHOJajd9xYXX+ubsA/wRLA8eZb1VUOEtowM4r
527vCCa2GLfikANqiPENGoyjD0/ZHJlh7s8+XwIQARrfI9B8Z4AUF0ZLCOpH2g8bL6oObPrwv0vl
VRdUo3fbJYa8kWTyrxmUiMXWWqxuGX4eQ+3PaWjNpVQlRr+/9yqmKUpYOFjlFTU1UTtnISNqm0jG
GxOsgTNC2mqij+EOuErApZPfhU7YDquIaYFnATfR3lQ/25SMlD7VXBKSAQdUIGlqmG+3Tdej7dZI
2GFpjfHz8U7FLYFyEjrlNXvwKmejP9BtgurOh/nHbpHXJG6R4P5A392iR9Eqg75NdNK4yMc5YmjU
JcdWCuorBezhqN+PTSY4ZNC2lf0MJpP+xkBaDK4YHpwD/GobfLw/9s7YGM9FzUMjxoazkh0FG9lw
ZUAQq1Wu4Dd/oomdOGvnztOUWVGD7lInO+NuTF65GPEIYlbnoL0QyAmr/kARgK5CdM3VX9qNztPr
J/lzaySIZ/A4dSZ2ppmsQwZ98AL1gwxn6PjnUrLPD1gvYJ0CjEOkzBmWjHiltwZJ3uSZJUnhlbwj
tU+KCKnwkQiQUIdAkX1hjAyVIsTb+GbDnUbNr4i2ClQcSq8B3lf41Qy7wZuJ2eEzO8ukZM1ZYqgI
cZs5VvnuWdCgyyjcHOMMCSVDbE2ifQTGGDeHQpZoQLMMwNCtHtMkRnx5bUgVz9g/dXgUu1s7UrUW
Ds4dn5qZzAGjZz9We0Z7KrLqDFJmrBi6aAMsI3oFriBPHJAlCBrFP0E8MzQuvJIfwL2RkAL92C0I
s0JzZvwWFrbrCWQh7lPnQmd76ZBl0oQbYhh5gzk6hCOdu6IcDEJuMuvjRhkUGjyxha9mSgZbK+TM
zDinTXYqwNKbQsC9pxtyYOuSuW90dwFlWhECjd9MUEVD+w6CAvI8UjXJaeMNqM6khg2oFdU4BgqH
UuQpir6Xys3G5NE1FW8xBUhheQjqjqTMUM/MMaKqOP14VaZx3ZEVXC9MbVGPT675npps4r99Ot8u
yHO+pfKtHUvwno+QkOEvybcWquZrErh05tLNOINrI7+TuKhL/BaKwjmkTIDP08UMADhfZgMkqpoj
F/huxztrR7OGRZ5BMTjpvwJ0mXRDlK2/3IinT2gY7toUPGd7SV75UCAPymhLI1ECkQElxn/SAL3L
ypn9562eR8JwXx2EyU1qJmNDc/f+aRoBfzCY0ccLpbLMu45EsHmFhBWiYgXY2Gv9s5XL8HsPA1wZ
0Z4S814fARgT69fqcw56DYENxLgepS2faeNoF+lqW2S/R0qgg8J6KHGZZoFb0fLquwc3CC//bqBJ
g0EM0rWIjwwPKOGGk3CY33fvbG4EtEoXgMS8NRh7wbbX1gyu1AiskJe0u3V1yZX15rxbIcp6+hnb
9DLqeOaquz0zaEn+rzUy+KVfNxS4o/r6ger3/Lo6mlQG6kTNf3apqYJirKpXX8zA3v4cy54tD8Qc
BBw4C6QVzomW0QmzXLNaVO9kilTttHyTzhwCsPid0rlOuGWxi8+b39dpNRPo6OSZ862OLT1PxqlK
fyKk7OTQVxcGlVvLzgXCPo5v8OK3TzgnaMV41y+FJWvkhN6LqjgzQbY7jyXaJgzczbJyBwzhK2g3
0I/qRa3LL79AdTdK3wuw01vgEDLPg5F0W9Jl4dPvbKQVlMwbo8TdO3cGIP9ej8P43TcslOGEPNgC
cFBtPogHAJoRD9DxVunO0blF3gIEZZ/oo3JedTWrjZKABpHS9JkNoCEGkqvnbtvFuAzJMtFhG+m/
che4xvLFh72du7tsKoHa5Znu3DNCxk2U6LWecpYrTQ/b9df3uCgwI1C+vgt01POat/TSHIKS9uLF
RhJVxPNgDr63mZ60pj2hl0NY5OoDd4Py1aCgdYmMEWZFNpemKerJXNQOB6FOtiWZSFGH4VEWC337
2UswFJbIkIrzx/1RkwgllJkcDmRPPhFwYM/m8UhHu1vz1zfDVYnnpQicdQlF18aYSdY0VIc6R1BE
4our0GCZBAeGji/kckGiovbcDuEBwd/VHMrANT6iMYcv+UtGeHruXVISlMEnY8kzevV51T3JWJnV
rABsVlUjP8pVFZCHqIdfc5XTDu0NYz5NaFrCE8dkk4yuEjKflz6jz5hyfaka1rYu/ij2XKEU+64G
shDxPqJtl6FgNnGSd5qgHx71le6/Qs+iXDg2KBwOW3n3LDXS7jPC8BHB3qu35dKt4Smn7ks8Pymn
mzzyeZB88znrQim0/lrCgkDM1IavWpbn02DxvwSpysFjlxgusc/8bl0tMSiuPGuigyFRDqnbxVQS
uAhFroiVcc7vhgpfnFzO/WTktS8L+UCJZrGLO3AaCVoE1sK7zsR72Ztlr8J7tam4NLAtN+Kj/WJ1
mwL3IBLpAIvRnkktVvqMa22P2yzCIEKU3m1xSfyf06QdY3t29vse9lyyPi/T7Qsdb/gSi9PRdhJR
x3BQEEomGkzRAGITwW9AqBVnhaoUF4uKwHKbUQcTk8uICHMiA58B/6HSD9J8wiAM2VrYnyxZrauV
vX4qF8vqu/VN5XEoJuNIkDHOZyym8izOxfwmsBS2K7hHveCe5Yjko5W7yIW59PcXrpa0akcBp03n
WzF+euKgTel6jKyLJYkuMYiELLJ0w438knO0xuzOUByVoBnlGQs3srIo1CdXSzqB+8/yEtAHaWMC
tBA5a+2l93Cl76urhm/NM9BVjdfMoZ8xOUyOa4Wy4c69mQIfJK6a0PsgwkBbgJmS3dqTFHnIgbsi
3gfGhOfG/lTexslaw9ae9/0WpN+qIOyFcdxcieME3giU/IdE7N/KpX93PpJY1h0Kcj+2VAnA1FwU
bwoQ3xQMkBYGOAT8wx2mfX6U0gqFejtNYHpnnymjFY2AZPDDdKnCjUaH5XyFsHpDtuPno/sV83Y/
EbnAjRjBtxHjEuEoRGo9XzVomCfa0YK/taTxhJHzmQh9LPTXkvwZf7/r6zeLtH+U1adLhvzbjI+0
zfcNe76mK0dn9fJwk1NBp9tXlDSE0w7G4aH7WP0cLPMVIqE4PVDJgwOZARFZMxibmxFjp5/Y5jrC
HpwCNBhn1/4Wvqh3/0MC33Ix08RMm75Z9yhk8eVZN4b9BC4+J0yl3lhb1rsbBclaNc30XbUsGIRT
z3louwhcqaFFB2au108kx6EmYuaGPDvSE6sdyFfEHpcyiCtfKvBbfe2daFGBtwDoeSg7l633HMZ3
1yH4BSQR3EGpyCDECQ1Tc/N6NbL24vXm4VeaZ0NTSoKJmEEXmi/yQ/XkWRYTJLLf5kcxaiQ5nNM2
1Me5vDgNSYwP3pujaOUQUTpgq8Y+ecpsAZobKAQar+pqSUhxfqtJZXOGX5MDS1cxVsjbaNEOadH4
1t6fwDjCs5usvLG6nSakmKU1DUh51/MsFoBCdl+T4JE9uFfNZ/5szwBQFDIxRKjIm4O0JY95LUxm
ehso9aUT/7IE6xQnA9/R1DGmAuMNSTSZSW+lsUHklk9Y/IbnrnSh5Jh05fSOocAUnLmmerTAOJlG
P3q+MPvr3zY6kAdXdwa0cE5AauDcMUcWtMFpNmpwJxfPszwxCpTe47zHPweV3j/KB0URJWzVoI/b
ySM21QW2jzuvGe1s+AUyJIOE5oCbuT+i6+S73QxPAvgEiZJ8xWbQBS7FwdDATjtVIMj9qjuKPWKK
OTYcxvwqWxbwBta5sd3IIGdNJRE6V6VRb13cJeF9eb+yoxq5xDqr4KHHXZRUkJ45IH4FNdDyjhJp
75fd5tpb4HuQXmL9Dg4ovr3gd0/ZLUJD5x8DOVN4vCQhFhWzfQ9vfE6UH6abKe9TfRLmzW4Pc7Zl
H46ApcbD+bdhUQ5PvLWA1wUzy6Bq7jfXJV1KK7hLISMoLCQLaEJ6wR+Ccz8dnNb5praoNfN6NOjc
XElnL+YAZEOuHf6JHlWJ+szZjNh63EVAaJfwRnVAOiPGUrwS4lpAdRPV8666pteEWWEfBZUGQSED
3Tc5stemL/6S+ssYfYH46qtbk2y3D20jWRtBLYVChu6Z6ZrNehcJGh+aBtMxS9TOiYgOx7AIOvzk
lmiYN78nRDAlECRkbpXIif9BrqwGaq7xwfsYggzggUVYxId0ZMOt1l587TviImSVo8vX6Od7s71M
ZsZ9dVoKGVAXWPH2VaM/7ChI8WKoht/uZlGaN745qI+XesshGdaQJP9marFVMy7PNN9GtMTgNGbO
RIp1Z73P88xzhh4xGVZxULLYh6+x9pQWJP65fRk/8WCJ5FfHp/IV6o4I3Z4XpfNP1kMOifFg21xD
XGYwtD8tVSkLNolV3Jp6ZNgaridjwmLdjjqad4/B3EmIAIPtql+Am/WNztK7rgvSoWGsQyu7N4f5
ASD5TjZ584XW+b4aUO9cRgj83a+2AMxMvltWFi0h8jDU1o09O33IfxDk6MA51WHDm6vR/2jqlTGX
Sal2sMKFdTfNtvkKDGDZrCrR/v3GJ+hJT+VFXujkjoyoNNNiua1JasCwZsc/un6HQbGeVTYq7PEV
Lpwv+fbauC6DiZClYNxHlAdKM0bV4wbnYK7EUx6b/Xby+8jL+Q+Ylxx4S/GwVnH6vJDi8WFyCNAc
8kl4Iksi2lkCSMD+O7Dyti0lZBKdDekuiVY9F/oa//sN+RkG0d5PFYNagT0ZUzP2dAC8WeFyJxs/
SXczTQ7G2G0isC7RhGhqUIDzO03A9I8A3oUAmhVaoL64AvW2+AsNxyVP0MGJvN6ksRsdtRusZ0Jx
D1Oo8mNZ0H1OVHyKyJBh2FeCyUFn2U6yL/+jN/mGPw4yUhKP7aecmOwPWSiGoQOdeUz/OdVkW5ri
ua5c8Ys1E0t61zjqdlnBzOR9kRvUW4pcuyjfm6ihhtU+6oHvU+i7rWOPLxlAZTOCrDtykNhu2g9z
l20AB9IyKg8ZAu2OeQgs136Y8vMHj4wxcWZuUcuZLQH4Y+j8LraJmEf3GsUVxHCGW7a6v4UjbtsL
8gHdqDtm9jFYZZPbpfkI+81XDm8DFHPHPz0OmdnEZ5Kldpz1HtHMBVjUHk4sCYvgnOL57dcSio4T
E+drLFc7EkTmRZt7RxFXhdWibqAK0LAf2SBPwnOmPj8XjL2U+/rHwWbyfe2Bme7KFBLoADMh2z9f
s4MIcX/p16lR+w/gl7BMgivsSZpbhw+z6osz4T+gnJwxXl9ox6go7DJySuAuYqNm4uRT9fy/v79s
eMRVOuiu3UILutsJIBEMKxV8LmsAcGngBlxlZXSBnizkJr4xKTQVM9t8ZV2aSuo9Q/i/E0gSudTv
XLpwEosSF2Ufjuedmyjd19s4RTRy300zzaLjgIxCnm7uU6WBFDeAmgCIYPwggJhg9EltNGb1Bwlq
ZpbsQjGuPUC99d46Lt8M0f3IxRbetCaeRCCMSou4GuNytiv7CBXl3kUxXFf3/BbOsQ0xgcH6uVOq
ehKy3ETxZtTEJLFy2YPnDvWt6+Iqsj5U3DnQpGQ6bSOXDhSa7WEfFBUvLniqm+RFzxLcyGtRvpkO
eeomLPkIHR2OTNGtPLRErPO0nNJ5bnzH9RsHiT8xII0Db7R3dlnDaJF/LerBpeMAqV8jQ1wth5oy
S9tB6YV/XIQ8y2blJhKg7n8O0Mya6bLB8lXj5OW/hSZx+EPlVqkELiO8xL0AeWNjiSSt7A+F4pxQ
5VkuBwFDBmt0xhyLXbbwLKAbJMcqGr+3bg2rIkrmmE8oTHxcEr+gFJsz7QjBaa/a+H/tfxVWbPUt
31WUfZnK9LhQ3F1/wzWbQT2x9ee30qa1KoowIpaQFaimgV9xJV+qHidBQCf+lhHD9/dFgHp2gw6P
qU2F58CpAe0CvoEgyfIwXOa38SqtRKfAyEi98y/eS+mXEeW87BWJJCltl9Lk8CXH9FD/1fwQEJIB
TxHVdG1C8HsvWLb1zknCZ+OHZcHxEeIPKEDLiNTOSvk7/o1mBF6QkyAsFcX/nuV6AmQx2s3nbdhk
JgjGeLVym88aKa/KofGl9i9/pbFgbI4nAODUitny1slFMnPrpxd2TZq1m2FNtV0RXw4d8spQDyBB
bV6HR0EHaZLzuQLbm+xtpLRAG1ehVSgnIN3U/iwOD10auB5NccWQTCnRK3JT20irENBGi59FpQfs
HaQgeKuWvKt0mCvg2N3bwXBVii6VYpU0vnoHJLsb56+BmITTC366ZdZFiUfvGTo2LwfUDrVFvhvr
7jhZ8itpoiPcRdTr/jm/RVzbL1pJr2vSrxaojZWoNRBDh8Mp9YiIVpsNoLVS+O6tnFMUzS9vE//J
4Y6HDS9dsYSgy2b4E8Rw3OD5qaV3xCvIqcaDEASuxazFfknlUkUV41Qqm9KDdsJUKtzI6T3rFCH9
h51DCVhF3OWqv2PqOw1uBQdLtJcWWrJdZVsk3MtJ631bLzBUVpxXo6/6Fs+mCSIeEQR84f9hSe3j
1fQwXcRW+Kq9kEVMZ2FqTcxI3+PshSU7j0LdIkWXCLDT2cK0xruumc+YBWPeVLmZnsNzKJCF2rXt
lIZo8oaoEh+gVVKQXMLxCYMVKwMS6j5dVhH906rp7oiGJL4k8q7pW/B/sXKTclcspQRpkTKlVmFu
aPWHJLKfvKkaottyI58vE3M738SHb+evQ+/59soLkBBRHtetdY4KZn0MM/zuFCdJSERBIscOeLtf
WcabIFnayMADx0mlWds3j7n3k+E+9Ae4i42LX+RkEF2a4ymJxLiCAKWega8w9lkv2ry/yH1kQihl
F79DqtT44AkhJkNDo654bFmw+nXYIAVl+QkThESPb2Pnqc6t5MT7Q57az6ei/GkgRqklde2dY9ub
9nihSdH+Rmu8ZMj+txdvGv5FoE8r5iPMkRyrYlE/EPOjnuiccFrp5xuVS0j4IDph+tRO7YPg3GPk
xrhLXWh1GnmUbcpRJ3wLk6iXBipDz9Gw6n5P1KmDQl+b93xMeNtfBGuSKhssQhCO9r4mJQVfzEjg
J+t0rpq6aD5cK3kOf4CjvUHbiukOUtsQERodLDkPwKhstt4c2fBD1t3IEi1ZnuwICWKRGNcNooLv
hFaQDjLZEwl0G/4h1CWHCshd9VzkR4DAkbph7jXgN1PinceYpStKDho2HBlkdZYOUOHlJVjH3/fj
tt9Klc4QZI2Jw67f6orLnbLeypEb8YBJBaqZCx2bi0Ss7QR06ogeq0mfOt6HL3lEmB7knZV6DJvd
0jEveEJwfrnAxMLGtAj7THQDAEJZGV3CfASYaNQtLWaCDObYmh28PBEVTU/L1h39YSXma+e4IYSl
zClDRQagx92LpWc6S/5QPzvAeZ16XBlAPfO+xB2w7uI0cn7GhTah+5S1WaVva4Sxqyi5dIikSK1x
54gvlFkzMYpq7woVwWioSNx0CJcL9sRh3SZXoMNFtaD7ubQqtIwXWpj7FRqZq29nm8Qbk49aMSZk
nndyLfnMJFqATV5g39ZaFN0hm7RIbZRu9Lz/Y6Td7p97Q4WV4c6cQVdZlh3HcfUidqF/6uBfxKe7
rit6awP1MflaG9Pk/PZVRviNCDTIhjk8WdeCNcX6HVXnKJ8kzPPgcr1mizT9Du3RvWrQr3MTZjid
w7f1tTxnzUFh6jE5hG7l79CZHJnGk92DNaSzuiEDl8wGF4LeZfIU77RCR/kMGts5IRHRFiM6pS2J
DA5GrqT76ilBsXFm5SvzQytw3EvAgGHOQszJoANOIANeDvEE9VNOKpLhOsZoeLqZVD2aRGJp5Hy3
UwQVXBKTpOfjqyDQrVcMnVvofX+V/x403pbRapw+np28hD+5LtnFPw9YHnQdoOlNRqe/ohn/rGAP
u7U/1fAHMyAi91kkfuJUqyUJ0eFZtGLQU+mQ2vIEcKhy/RfVzi5kU2DXDVXC1N76flabUFAkmFrY
bktYwdjiksttI8nrvTa9dpSpxFmyrrEmVHcoylZdMtu8lsyfvyvkadO8OfGrbXAxY6VXLVFj1Vnt
G06iZ7gi4y8Ypb6zlOrRy7CitwETIC9osASoZUjJiD23edQklb45gP35tLl7GcfWfSJLafTd3184
4J4rYc2quOTrnKI0CIwRXoySQMiYYAos94LXJjI0hQM99LPMf5Yb0W76rI9YBmXmOgCyNLMVg4ab
Qcx8rvPW4JRgmGM6ZyuEPYOMNuVVhdzZ2G04t2pdt+weUwoL2YY8jp8eSykfL/hw1r3rW8KYGi9J
PkWB8JNVVOr8k4KMIAzHLUGTBKEGA08wtKM1A6wNsrPKs14asaq+EMUCrXeCbMMdWMFVCHOSaLW3
6/XDFPIFAKr7qQMqab4hHzry6Chbga1BPSDx+kOMmV1D8zfGEQa5BwsXTZs8l56tmS0mycSHbex5
5+bORGlnhQzAiJv5wSWV1wrPVK/xZrazgY18urvDbVtnaWPpz57nKv8Udxdzp3yvCVL7XJLKlWdD
zsctMpMT3g3YqtoGYgN6pxj4ymhWhwA0oIaN867Ts98NI9GaK/+KXzZNKSIEp04zL3TJ8RM6rMMH
wWzXA7eMY2AHpRKheFrcdh8rx585HmonC1Vbq7BO/aEyfImkAGtRs1agzwAtsPZdAv40B761DmQa
Pz4Nml20BrQv+swp5pYHLI9+fQ/miGczsWxKDeiTMK/nMXIL2ikgs/+9n1lHEa13JwKtuueTyu61
V5jGdQbao/5neYSsUOHajsgFVRyOb2o7FzGPvKzwf30W2G8Jab+2+pKvDfOAzjTC4/9Bly/X+UKd
imks24UPf/yKV9SeiTuyuewzhtG3hIzcgbkRmY332Yyf7ISFUtni9S0BwGwceeup8AzAZ6qIKLLc
z10waEbM0TdHOR3BThFukrJVMYXcKOUIV7RQb9dtYPjqiu5c8GDzJJEHvlQ07nTghM77gl6xYMPP
xdeRE7o+WLKp/Po8PpMypiaLf0cAxsSiWt1QbmO/ZUgsHF86h1rbPT4wef1jaXgoS/cEJYYic4X7
ofvmfs+ZAk2LZc4Q5nYw1X8YgMEghoUya3fm6yGCHnzDiG+UAO3HoxT4jwyWp9MBs81CgYlhwA6k
pEFbhVwjz04fnj2mYDNZfoKBn5qPVbF6PVWcIRqdna6RJHvYvCkDW5iAI38QqNJQdyFL2bN2yTK7
L8/Peawy020J/UlMURvvjH7O/3SZuHK9EDWJpROuQmrwkCj+2z/AvxbXbc9Xqr2pmnuonMfsJI6p
Y+4iVo6bb8lspEk9t8sL03qs9KfuAp2jPakYcg5l+0dsZeDGGIddT9b/FVdAqNYbIXFdCUSYrq7+
kh3saZ2SxxFpkQ8Ti8DDpx1Cfy8TM3kPOGLjw74SSqpLZpFPYxDmiiKS2KaQC4LxTmUOHbbrqp31
lqLMV1KPCZSNa18bN4mCDuthi5YZqKQrWLMKJ8gBzEf4I1thncC8jeYEUeYpio3xZupZDQbXqoaJ
39PwhNTGmovsX+WZl0gSLt2ig266pnujA1yEJYq7Y4guWb2GYpH/rWmCSHdwFgNDfcspesJU3aOt
stxMXY/UvX3XnNOAVBA/vZyoXbQVcjfDer0EYvPn1YsS2gq9MeYtrV5mmCZQeNWuzgDLz/vMsa1f
J6W5I1jz+VFYIF9fbp3AGuSzX6YNfScMblWAh9pTI6h0oZtAzIEDuxqXMU3wh2TFRLprWT1Hi60t
C6SKs20rJUeXnTO9GWfAkCiPdteUkPZO6cflCf6dLQ+sE4TZKOg/XGJRG/xwp0XaeQDkI8gPRVaC
yAzfzLgbs6xUraqlgHSOUNUqNb3EAs7+9MsXWpWnmFAlhSjT+VLEUkc4KUvTeQkZ8OyHhOMf86dw
ybA9l8DsY2BfNPcG1zFMNX0lLjqauLf448yqcR8ppcIs3KdVurlnOpsO94Wlu5rOXXeQO/141sS3
BiMT+KtB+hqTilz2xjqsZzPf1wkEyRhR8SuYAaqsWZ4H1i7GG8rP/XrAdGJ31t3orx8+GpUQ7t44
qFdUkK1r+m0QM2GTVs8COg0eb4Kjz8IFyb/zTn9dpoMs7bm1Kt6Hp1wXmcV8C61a9/RdOx1vG3rW
W3zeBfUHu9IGS/O0yUjjKAz0O0N57Hnw8wE14KjnHjf+Kr4KoRKeTCdO9NzC8CNziMAZLTGFEZIK
iJA4nT7VcKdMlgmp7Wh2a+6xd/HqBYpX2F+aEgZlRpoIGlhs9F2pktnKhrEsKVE6SJC0bknI5lwJ
DAwQhqs3g9N45VSXG9EfhOlOaGRo05REQnRjlQ1rZ50zCo7aY6mREBJno2xSneIWzWZtpV9tfbqS
q9pakLmDlP7NHUCdQwkxyW7KdKBTwA/y0h4puhlPFu+Qprej6bKDVt9zgXEzkt6/4m0HvzbVzZev
faPcnMqlC/jOP/MT9AUi1kJl8rf++eqQWjxxRi6slR6xEqM+yyYA/ibP3z05yIUoOWOKcqr+utVF
3tktF8LtyIjmKEyItQqeBu4Me9Yl2FdDV80ndFaoyHA7Vp9C2FdsdV/CL9C9u1BpkwB7idHQ1lwp
ExyrTkkLZqM+idp+gAj9YahtqN/SlCrCRTOL+ri3eDIJyzqUwmm0irDkxiLq+WZZAF87keGhLxJf
6K6CLyjPyr4gwSq25z3NqBmBun/FOA0cjBodDsbC91qAEin/0c7ArzjcVMsn5pYLQD5y38dZfkO7
etDkldXQU/hi1hFDyXFdwMfM6cgmAaiBNwtvxjCMGidKEHweUVfAtAVZvbtIB8z0sfULLT1taf9u
zUtditT9VuFkdqEuzKg7eLXnvhg6LiiL3s5joBNa0gef/FRHhXV0R1j6MkX6QpwSXMf9fCBStOwI
BqZP7ttSi61SNtQ2MD4Fn3Q8vjlh3j3TEW4xQJnjosRAxdRIG3bznfiF28wCrLHBtjyFJD9CBIG5
nJNjmgBb7IMXsrwz1B5b2htpnemEF9yOT1in8MR50Dz1FC4ORSwCAKkkF09rV7zrlYbXetup1wIv
TnbMFmj82l4Pgw56T5Pwo+u5oPfLZEK4Gmwkk17/5oVCAgVO73dvDEWMAttYyMy88kCp0tR1oNB/
iCZ1th4wX5U0uyWde8yYEJeYlTLQsEHP+9XhUwGAVb89wSfouRWeh3JSLZlhHRg1e4BoWKrZEsQc
K4yuVM4MHIHwOJ7tXeRrhtqaw2ocDwqfI5aVvPYaLUhBYhtTeFzMvsl5b/DHrWnGoOzAH1MopQhH
r5rfHYXrvSz4jJ/f7S5CI8SyZ3H9jFvfDE5i+Oh9+4sM8JmS1vWtRVWfBjVnRsxA7f5/Jbuv+A3e
AOtQXEODYY2V1S4spxagnvo1zk8HPms6JEZwbCjEbBm8/YzrXyRyM5QT2K+5qmbMXJmD3oMkqK/u
/3HzeWkWsi08tX+NjtuquLZH0p1qmVeCkkOPP/0lYWT9DynuK99PKK8jXTWmYx6mYcT2KU3pyFEk
lyPNWiGjMk2h+xeNcFMNnXAPCTwevfc9XZDmHpzt6dGt/ELW8mSOMctD2szsEQUq7sBfYXplcdxd
vfAFyogrFpuboctN8D2VprgUvLo+wGS1g8ZhVdzojuXd3e2P06fHTrL+a1cLoy8TvMsWOg9GlKPh
J94EqbCv29i+DJS+84AaDZ0d56xfNmt3z9iM9o4GZe522kHUcYxoRkGGXRxuRu1xTlggu0fm84yO
QlCSzzFkwcciIK6Yd/tdIW2cNuYTrCexP6OXDcYrV9fLy+0Y8m5nxWzlgoxrdf1bswGrKJib9z0Q
ovIZqFLQah6ET4oCGgLk2UCcJ614KyhUwuD8q4EHXTqrcgYKkf0WvHjcjtAO3twGPMLqqDHpgcTV
MJMqL8VXuplGz1aMPnHnosHEbAWw5Ajg/xGsEjUOChHHqsq8s83mIprfWqQfTLkycOsAAwhWNafH
3k0sf8s11ucAZu+Tr4UWc0xU/4idqGhklfNvGogxAgWsSXHr6MxGTLQO9uGATqHuznluh8GTmkTD
O/mMWeZc7b0OTRtZpY2kMsQTS28V68Kd+JwFMafkWQQfkCur+HLCaLbUdMydW5KEJXlnTxS+vLpa
h+w1Zxrr1Zu4C4UN2cARlF0yy57dcS6k7PqTU1NlS3QE04JbfrUVkC1E2M2Es5HUypuER8xG6N9h
Yc7UXQ9Wvl3MURF7yzxHJ9Kzc8tP4yU7GbRMziNgHzdKnOtOv9NcFYDKdgD5TCcLnNx7S8gctgKJ
UbvmV7/AND6U4cXmBzGP9BHF/PFPhpz+xWlv4eVuLJlXQkBQG8nQwCPGswcsSzXFQmuo89mH5wyg
1jPL/JccSEYpWH1kOYi0aK3IwtOAI8q13PzdTvg9IT10+EyCLWRyedQsbf29ua4ZG7ek5BoybS3z
4rLugIrnrO0+8pJxXRHmOsRAZkKGlL3jocKK0Q3CjCYOSsjexLoO6ajMVgc3zrIZzj7h8+dE5ir0
EKCJfYY6yzyqa+rBRMVr0H4+P2vGSCwcl73Q1E0872PHyCAlHPJ0xWRyDA3lCqbua/iAU98nUY6b
mkpq/BxUYPxga5XTZGue1NEMZjnayZcmHnf13JK0XlfEIYwD7d1rEaa/MfmroDTwZ5Ib0PwS4oXP
4axAdBFCalabBaUE4jjsbGVwXKYDNdyVAKV0lxtE9FW3GMH4yoG0pgN2NHZE/nR2JLgiG7IBsNBf
JSq68spwMrGndm/pXJnhIbA8/VOZYNvMPnzJazWhhYW3oBA81Vjg5RIdTT7Bem/GpA8Xp26KDcv9
Tl1jb0P+BFBHGlfClQelYfDjcbvtcvpg2YY2+BacL9SNmXNWH3niLe+6aVOOSAPM144DEPdWXnTL
JJ2L2YA7/BSD4ERFpu1DTV6VGYxr7RCgqJag9U1n90slIA1GWGk8euKUiSdAyM2Ugxb6R3qn8Loo
X2EC1D9AfMXkwgUoNGY6yo7Rv4la20SPht0JzgmMrxD8ZptfyM1R6donsU9sphZ5C/9bHSk3N5Q5
k5Ukv9JoyJdYcx4Q+5tn5TQC/EVuRCKt1exSBhJSn4Af9rz9tlJMKuJreWAScCxt9/VxFx9uuqfd
hR1nkDWevM9YuE9NWGYZ9V729R4IMzX+g1o3r5uyxNYtrugohe5tz22vvO9+lk6ams7DxwrmSs7F
bI7lyxgVq+qpwFPWG/3sD/aia7ipQpsu/jcn2MZCiCzHKpn5jN83RL/ijzWIgVlxo60tQGUri3hn
kM4d3FlQmM1d6hR6BRoh4s3R8VaLVYciRjOBGU9oazqALgfMOoJlKomqfmmWV+13ZKcatuIonX0E
4ztVeAFBrGlozDY4poR16uRVi/liy7GeZFBT8A6c0ATsGrGMgbpNsBIKVVTltpHwDRI+Ow37yXvd
6SLcISPdJkAPWBArzWhxvqC41azBXSXNkxhfRbj90v5Wpzb8/dHShove/skXsh+o7x5n9GXa6nr4
hPWiIuW5lJasiwxxCkqOrZEaMMrnAjXqdg7iPFqZQtlnRB5Mqk1xrMerbfAWrU7NZrziuVE8Lmpq
T14vjiYlXubRM2njXKlIjFXYvDENyfeOGu8SYvxtdG41htJbbKulYJ9c6vqzbmR/MQaWPIFngkxM
0p87b8WMjkbq1sXJ5Xg/PeAK4yqIL4VOfdeTKub2G1dkOMldb/yvkEBaWhe5qjN8b+LsU5N3tneT
b8CKmdNgD10hQD92ZdxYWGNNsHA1qBOCjaGGGKMTL8uIscUvlFO5zsGZWWT/vtBwOpzmc7evJMvV
gfELj5tgrEU5/8+l693yHZQv/Zu+pKhVCKukbegZcbkFkXByTN/MxUdzzlDFlQeNbpvDrh2b2Ph5
jjm6zVC6zwyV9Gg/EKhvV6i5SHaPC6zXz8LFPeDDvxK2ZOrU4VAUABqZCuMN5NefiF7SvRskfgXx
lu2ejEju6/surEpLB8/2YF3FZznaK/cFceuj7Wzf4E/38eO+YxIZHxkfnsvalrhnckx3DBmolXtH
itFYo6KDs0WIsvGCaCPeIlUTupKkmRaES9Qxb8Ep1xI7vnAjg1dnLF7whxiedZfmo8UBD2G3+lHA
scb7cYsn0GCFRFC+TGkUGmG0OCmcE2l7N+GeW8uD2+jq5MpDaV5AWZY23boxMssBuumYkVDAj31A
0HqHffn8Z8a89KsI//aMKT3aH7U4kj8BdoxXqlBIq6Ic6DuWLkLapaTYVhPMz12BrPjN7pN06K6k
4FR98RhckJeBb14vqPZ5IhUaFBJrZp/OZPaQaeO6GFAHRCtHcvOWCLCMdhrshNVmrLvRWkFZ0gja
yLwlIDexFP4+8WLCriFMB/sbN2l1s0aYZ9e4kuUcosty5XFj0e/Z4bdUhsFgRI7LBkfK79LLsoPd
NfNeUwtd8P/d4YOV+IP3H0Zm6K9mhSJapRoY3AAl/fqU7bg0sJi4EGOkrvX5FVlc9I+IUIbJ865M
I8J9TBZVQhIgKHZlxBRla832CmhuxLb+n03b7NvzQBgHXvsxAo0gw2BLBhkLQWa3nRBw9pqw1IWf
o0abK67xaAT/PsExzE3Nw6+zQGIObfg5688a/upuI+sMl/stM8542DB7Nxr8HhTX0YuZRH2xCRQL
IqLODJVVU8xtpW+Irah3aQxXjyAxswEgrw1Q5ZORFNANd96SLBZb9+QIUZrFAi4VxeAdJYah0o7/
xVuFUHUFZ2HftFryvm7LJ/Z9ao6DyOHQ5X62d8PWKPBrkD3W0Vn3O1Srjl4hAcRsumrJWlQftwBN
WvBzrdl77SKNbdasg+Q+gaLkFfv5y2OefhFDQwsUQPslO2rsxcQ8LINYh4n2W0z2NTDCbUzBPITm
X0dloo5jP9W1fNk5qq63UCp2Bzu+7/kPtlSfBOO0Te5yWLQY6mA839CAS/limK8KY31W8bCCjpew
1iTwd6OipkKzcWKINGBwCDEOEKrz1hR2r0Qbhm1HZcUA3tuLLn8d0hST9G2Ro1UwUZJC8ZXk0OxZ
Osudrt85j1Ig9vWZJtmhd7xIohgYFklAkw/mdblGXwuI0t3paHzizIesytIMAKaKpPSuzL+dJWsv
XBEDHwHAqBu7f/x7ZEvjyCPgy1ypW1ND52nnczlQUJfFaJ8SsShc3TD+B2IocgcQYBkW12feGAWj
RXQPWl295ktDe2Lz42IBl0wjUZFplypFpjfprgQrtf0o4r+Ake6ZpBn+r9G5fOqY9DfXmY5/s7fp
zzlfaegaKGv/Kkmp6rZCudHYR8NTeT1aYhe0FVUx/QMebPfo/FSCp057e9BM6oQDSSy2VqOntP/t
rY9/tYTF+uubfrO8C0gQ8lgMM6Fik9zJoy99HynIwIIFF5afBkK5NqUMYpqj4ctFmIbt8Upjd//s
BjuKdYNCmL64b9K1RMeDOIrVi5zybEPxwWMPgLEXuhSaQ6NHEVP0XMR1jos00SQpYv0kJ7tViv55
zOVQDRX4X1H3dPrbq+Kf5nJZImgfoRBT0sdkQn0CSjgCsnwt4U4PMFfpXeTKJ/aZII/t91xyPODF
ZGVd5IXCdP+ZqikKOELBMNWWjOviKD76+ejuLa/ongOFnwJSPcvjmbeohY6zM6JFA7/vueAiIH7Z
G4xVy4KINq/z7m95hkvWhd4xtZc0zmOsoM4BInl1x6ipZOrrYJ8bOEfJqFUZQSQ7KV1keVX7jv6K
x6HWQ3b/Vrfb3wQnukwhgeNCsGeGW63GswjUyfYwJsgrP+sv0rA7dYX/p3D6CHQ/cImDTX7ObuKo
8QRF8rwyF+Y7Xk0/HuTIl30/0XCJWG2WsXpgpxDlZYcMg+UAjMQZyQ2Jzhg+R9WD5IC+eq0X1M6j
eCuKdAbf49TwWsfaDUIKt6TB6miL00zIfm72Rx5+ZY3Pl9YfFtFH4Oy5EykchDeC3qD5EOOKs0ca
Cc+XEAr/NhyxjG1v6n1pQINPFo2YxHrRM2ZcsD/PVHjSiB52Wgn6g5lEKOeGL7wL3mEIdBuaQNxs
Dub5EoOkOAh22UNLfzjESAiuUHOq5LfHKI/x78nZCaMuytXWfdj1vQZxcVcya6erzrx4tVIPxZTp
r8lMFOyuAfcvoZ/rcajNFbnDfS7uAdmlzdHSxBsGtuiWuoH9W4a/1n+SIpT0y4+5eLvuOQBF4DoE
c1PZzKZJkIM6waaJyKOYYq0psl8ZINmdaAuiyj2dnUHvJujBtgiIi7NgAeVbgU6r+MdTO0trht9v
bElsV7UZHJR2/yZL0lJP7NQlJnkY/ZjkBZEKENG/yWbfYGva66CXhlFKGs8GM7ySUd2Lvj2vdy+u
6H2Aw7pmSYLX6gfkgEkQzA4lNnwv2EvRxZcwYLwI0sBN6w9Npqtc7Q+u0KjbXlZwUQy14cFIkolc
KkPMpFxgfDsjXT4aacTnJH7wZtMEJH5YbiSZxeilf3QE3i1zlUYBARK+l095Ua07KwO77h/VZTk0
wjWMkvfw0GtRi2aciqctRYE2Ri7WHZbvKLEmeF7FbkBcY2MSg90bTWHpNuk1uObQVodbIXpVI+ES
kEBAamYyoQNpYrAZJnccaH/vMOIi/40UfJo2z2T2zvV2TfiOb1jzh6HhVx4LmUQIwqohQ1DRvnB7
vnfqWsyZpeifQXiW3iRSbd2xCX1Xwid50CxKfCJKXtW2h1p58Zpdc0SF+HEMAFUXRthnJhIEhiF2
tPBzEl1yg+KbjBbWhpN19jcnF8HcXJpbAynPnfcp7KhnZtZ9BqpKhjAGFQkanj83SfpngczT08Za
6RmgFU0ubPTB59LGqx+BaJPDvLQBbLGIRP8ID25YRD0fsdSxIWdf2lXk1YOJDE7QLqaNSICIDyVZ
kUCAHsdRcTIQzKMd0iClVxCXKScXvXgw+EqL04RqIfamk7dUvibluPKXmBVvI/tuNLPpFUEwMFfk
vN7709IzgTza4jjhRJtGvmGXYpPJu+G+kGLPxzZzCl/XjqclAH8rVKllisK5O464M3yYZR+OCLMx
aTsoH0WR+Q3pj8e+FtjPUTX1GIri+1+qK2AXBBFOVZjMZocLX1j9HT1LF2tr2uzn1zQ80eqeROE2
TgbiQ0lxWylCZEHukJyTA9AVRv5fDmymp1K8tJlqclrRDF5dFdso7kbI4FkHz74nLtA03KzZL3Fm
3JvjX3IZctKwGJWj8agDHKUC+CzaKcpwJdoeh82M4uZxNnb5MtL+0VTmMZuxFAOwdL/EheneDlKK
UZdCF754madTxKhYsqw6HojcZDIb0wSR19IO+46aCpJO56Bt/V0+biEZ8F6uXX9h9OnBY6LILIZV
Vw3zxf8ZXH2wH6NMBCvwkkovmlXMLB4nT+1Jnlc3qovMR3z9G2RcdEARQsQIG5W5nUQky29tjBgj
/GO0fgHP8F9c89yLgegjt+mMwxIL8X4mpFTX9QbidzOvp8Do0Cp5DwbJi9rSEEbE9SQ3S01nTfhE
0spTdaTa7ULrZsKS/bLn/7SQdfFmmak/tGGAcNa2Y4phF0SjSQm/mV6FxAm5o2y8D1jev+5xG32r
R82/PV445+hDAnYHFvhVIP1Jam6FdkmNNNSQazMTYWaFzoo60GgMfZLH7kphIZcT+QEqHoDXoaj3
h+IpBa+ZwSXfmdQzWCpQEjTuZZmzIUq77MM4DjxVTzsvT+Mif2q8iNyZXYeESRCP0xEe1M7hwY80
AIsugnIJdCx86DisYY2cDbfzGfNTsHOS0iXoi8n1mdNkNbAz+9IlcSkoeY6zuO8iPXG6UsuzrdfR
xPTYorB2nPazoEkXtT5WxRi8P7g5fk5lZxNyxSc7Ra5GGW9CZ9P3lr6PXy8WezV5yJsMmvAUH1zJ
qeTvMKwbszlXV1dDuJ0YxM1WcYP3Fs388gPi6iC7rBosfwzmi80/LcQWdHd9fIbWK0dj6q+mgzo2
tKaLfHh7VuoHmx3KzpVvqQwGXy4EWy5YzScP6aAgbknOBAqNiEojqf6YHDBUFIAxPupDyYiOn6b4
uqlII2Dr/HULDRCiDePJQ/GdWlR44ifMFh0dKdNYDt+DqdqhlXgqgHbTMJtT9blnCx40fsO6ImgR
n+VKkVAU1ZCj/s4meumYV+0OQKeJ4oOn4FmGDBDv4IIYOQMwl17veZt75u4D5VCp2FLT7DMWL9D6
NnecYDzUGvlH13gZNWP07XxH5ovyoEa81h5ASg7R3V9XNlvo7h2JwmwS/y8EzgJEJStl60qtR44D
LpGUcvDs7bkX4jWue145wlJaHDhSa/qc72csRbpN4gMDhk4eHJTYX2nJOd3sod7TslTPVJFwEoKF
G5Bl6/ElTF5Pc0Y0enKAmX1wsIgTA3rXfsJX1/zgJGPXJJCfqovKy8tydYUECnzKpCSMpBLGgNnB
PKXq5O53azhpiGh/n9Gb73WfRgGoLyYfuINWXGEmseeCehQhlwPIqc2tyc0RrwMChXENQWant5oL
kLKRwDIBrAABPYYvtsE/e+1rKdR9ku0thNrPFiAeRVe2uBdlqhk5ltUMCPIQBIQadJdzsT330m6E
tu8dt9a/XLtNz5QfzBoU0VDZM0RRElG+fPO67k0KUHggghDwdToyqToB+xdy6SrJnFz+8y51Hdxd
itl8/i3Bnq1g4HKqc3En6j/7x9rFLYXLvL43v4yH5qRXzT7Q3E9YZnbYPhETNsHBx0Tergi1tlh8
SRPZyn9OpnMyU62o+0ONBXz+RWZr7C8YDZpZKxc7kO9FEx41O34WM2XHlyYIfvrAOPknGFAiSgzH
KRwjP2HTsyW2XPoEoIMtOHB2E8vMx9+kGVX1HI33vFaxSgmFdn2GJqWZEPk7VfDxod5qUnZcH6hP
Xy344JXtfmctdS81NYWU6D0OcFvN1xGb3jQ4ModrfX0EYuZeFSP5MYxTpZChq/gLlGkEY5PJC757
4e98XV4oWlNoPhSLa2efgVz62A17elvrzs0OUAgPGFbD38Ary4/CcAzz4HJy9+9kuwifUiyOU4DE
59BUEgi33BFnPt+7syR22MHwppYaqqKtPeD/E30D1i3al7Y4rgot84KowZqQBfvKgMExmknjgkqw
4+fN3EwGagDiK06onyIG8yEyvyDBb7RyUZjEQbdtNiAVGVrkoar8JfYzKpSmCWcbiZvWS3j5k9E0
5cDhgFO6YimV9/4aQ2jP64g9bQgAHN67ojSwXk3tjd8VErJuiJFltq25gGRsJoBtGO+Dlt+hUgzj
1/QDY+1xR4cnC4VVM5RiGa3ajFyZ7l0yXGVyf2t8kMjwOOfdggL76SoDCjzs61vLaU+SuhjI27dx
gw+CH3UWGU4H7t23RKyLppZ0uk/csLZD9vddrlDEJksu7rW1vaHmHMVBe9NgTl0TkRD3hoWkxJ36
7TYEepURyg9v8IpSjkt9u/EbDrVvqwFTUCj1JHJdAgqQAoOTOibaprW4RfaWOrXqbk7a61xSkgaz
IVZT7JuKgQLGob3k3WCyaqQfQVRTNITt9olZZSOIsqHDSJ6Zu9Yyt8RBMDK78R+4QJhWSVRyh2iy
6Nh9RodI0wwoNM9GEwhnyQ/D1c5oq9vSzjQMKwCPEaBGRqP26KCpxksxzamXmuQuoh0mOe5gYx95
RK3XCnBzuWT0eTF1csYF+3+l2AsWmYFk5H5pIarstCj8ZuQ11ltNg8Yjp+ic4nlSalQmgQelF0KA
7lK1zFB8I0FdsjYpUdPxcY9jp4kYdpsYQIA3mNZAq4z716odgIUmev/CYMsKi9JqEWnVAgiXc2cp
Oogg6sZvJI8TZplBDQ2CugwGxh8A1bMaBwiqN/th/GDsVkufEGapBVKUYlSojBJ5E1aeuEoTAXZV
VvdrXFUAeEuyH+YECS9KvpVb1P3zQI3YCMIcdrgXsEdxPpbV8RVCuGPTuu2JA/cfmyFCr3DjKBMS
xEToQsj4DL4ARPkYgYW52aAslzT6DKKMvHvnKYxINgLeJHGfT6/wYYu1DxbilcsobIi21tJEmCow
AHdMMkusXU6YAZ6Ij4b9HJ6TgngDEa7YSrEJaaZoIUCeu6VxG2dRnTantCAGEZhC4CZpOOBTDczW
sMqYxRmmlqPK4Rtk0QES0rCTxBI1kwbP5htDLLlYDY1tK8w3vZV/GBs4Vjdbis1jHBZv0IuqfjLq
D87T/0ha+m1Cek5GTA/qgbbRii1d71piHhQ4lv+/5z/VbMBsVIFg8UyMWFGcpKWkrIvUtZELP86R
UikOL7lXaUaV90JRNEo8OffhqFHrV899arKGW4CeZuWL9lB5Z6ZjI1IiN5+FMSZ7NqrL/t/eBZ7z
TaFIXqMD7xbNWUCQqhk9phIsuauB89TfS9tcHirOlLYW+wnOd15qdtThkvWNFPPkBZHl4tzE4bD0
oxxF5IYkvVl0Wrkcv/6wtV1+goRWBBOUADGGIDqx56TUp3mnN5V/zqz9F7e/FIzTMYVI+xn5xIPJ
xdIVwOtGiUKARb1Gdx800ggSLUkj14lbdruCrbTGGtv0cn4nkrCVTkpgmULMUAc4Zm2c1Nwv7ecP
tt6UBUuQsvvCbdjv7gk9H0CT1x1hyJcJwCdVlpTqXLjyZlGRpWCkLkhsl1Zpz2g8rAc7mzvDwMnG
q2pPPSGkDdBpWbVhhsPvtv0pAvaT0toq2MlSoIKx98cRBdw3Y89rIS4qnw6cUADFuYuLdXd63knD
igdDeaUbe5UCh2x+GHR0p8rmQQMLDDBQQMziytvfo654MwvjdXUcgi3a2wtayLz9+knq/7lY2BX+
MvjrTIIW6xKaPgR7l/SHEtjYpRgMXkFU8TgbuW0b3Q6FMFMJ0VIYpz2CHkMNgFUpTmSBXlHxv4cd
oetnaLASjZZ6XeYTCf86Ckyu2R1DY5xTLF115bBUAXhWQCJNED2yMiIWBkn/34g6/m79ocEpYIhX
orBi4aIKGfOhD40ft2Ilj/lFa5els2F0pSfX6GPeDqhWp8AqxITdz3FhjahYxXTnlvBeyfSH6h/v
gZXB7ShpOsqfGGhZQi6XUbqkb4Tg3wJ9YkpR6C+5+g1PK/OmxTteqTCROVLiGCIDOKQJRxLDDQK4
TZeR0M7t9jeeH3XFR9F8zh6zuWGm4szNuvn0OIzcG1MR3USTrFv/7o2iAS7Ud3ld/MPO35zbjWIn
k6YiM+vWkwWgV2uYOq1A0rBHmUbJyeNeXda49Vg10mdDGA5yZAqXpIh84TRtasMWSQV+oZ4CbOap
CivT4s2sL59DAL6xue1WlCafT6gyIaWY0Fj4E6erFut21ia7HpSD/I0onC9rwKl6cKphZ4DyFDQR
aCl0DUtO1iwpHm3UHQ09IUFZFXy44lVkoOFBthNp6IsOrOh+4i/AW0vtGZibtU9pEpbh4I6mLhHW
ccxmvnTGBg/43m6TjOCRpZabUHLU3G7Pa6XO3xxx+eTVyMxemn5ajAAxP1ryn4oQfkeM2+B/biTR
GlExYvEI6r8PyMhT7IF08+lZBriNxzQwi9KPjrSoPJMvErb9MObbXFSuFDrHsj8PnqVgHJdiJ2dQ
581oBrnP1zimFtQvqUbko5zh3mHKiqz5wQpq9alJF65fAlpfpdO9zG0E6TjHMY7/LnCVVAI5Gv5B
Z1n88ncFDcXeNL7lgyJxDbY0/yd+vizUCdK85ERgQBvxaturyjOj4oQ2937WSw4w3/X5d1fxXQmU
75tLLguWxb2xKPt6X7tlWV4PdTQg//UX4iCWyfqJE3hZ88Z8hNg9c3XVmeyHALWjWE3Le0LBeIj5
8Gqt2rEAZAKWfLAMsIivoINeYbFVrUZpYPUnOyDCweKJcZ/xJZom1smMRdF3o92/lOqZhT21tnuk
4v8zC3/GBLfTaE619TWg8fDdyUqQiIZXBi4toSPXU4svXeD2ZBXiX5f6FB/w/MjEN/sB+gNnlW/5
7O+A+lELSR2R5ItW0id2IYuLD7EwZC8rHntaLLbDXMgesko9sY42k9RuE9rDL25NvVw+S+Dtc221
ofsYLjEp3INHh2IlQhwNROfdAA0X6NtQSv8BRAVZtgpTzrjvmIhgm6mzIl0anRwAGRGTdwtSgnrm
B1Y2e5HuBLOXjJO0UVFoprZdW7ux8tmjNKSHpstPeaFp09t3bKVISEuSiIauKgqTgUjP0uU1qhUy
GbszX0qQFxoY7NpjYGC7qNuOUwwwakb/u6I6cDQgiYf4YCzActKXzEtMKprmpif2G4wyQcq+KGhW
nxZUPMXpqaAjFqvDwkH2BaOFwNwrA/uCBa6u8jgDbYxBT4ZVYgRkKvxqdqvyLKSSsEPaicHi9C/n
YX4gpoejc/4UY0dNb0M2/kWPHrSv2nTNxC/lRRwfThlemkmTCgB1qKk2VwZO1jShMpZPhLoi9Gqz
PIWNbct4y2eOb15KF/BMuodxKQQ8rwG9d0xvZiGBv9lATo/olaXXoyVIIXq9GxCUUYxJlsmE/2hD
Kao/dSaZ7F7xPUH7Z9MxfCGIQLm6Xy6X+1Nlwv/2+BOE9P9SNhcEPsnnkV5VlwX9uahfGtN/tLbm
dV6Jwz+/fB6Gd1UmXGivIIubqoWXHKroAkMP89ddkz3AJmBNMsq0x+qoqE1BXvDwDkhNlLcfgrxn
3Rf2nrnQx+j6uiuIvBxO5bWwmjmX8oNJG7s+dIxbyTl5p2nSULYblR563B/3H1Okp/kBrDjO44aA
zcf9m7mXOp+Na+JT/gPaFQGstJ5UTed7deyh5g4HJhpqY2Abyn6hfakTOxCMJNaayYadw8gCJbUz
a8hDp/R/Z2yE6adcQJXhFvLvH9EO/RbvTQSGi9dWQnUVGpsR7FPO746gBVXKdb0uNN33iBqQ8eP2
aLzCancWtc5z6MjJmzJT0FPCfwxULm0e5wAzZriH1uzCwFSSkrIXL8ELqObdqn7NCqMjyWVphZJW
8lM8hJXuAJqnyg4Fu8NNEhq/T6yjiPWkBEtxMnV2H0qAWRrMar1/tFY6X1SMpQeSvwwBll6JYa35
GzsDbB6DImmMgq/sf1i0C70AXlPcx+Y4fr8PwuBUDDIYMsIhyRiEFyg9D9nAE1aFz09Vmj+oXLKi
R16/7xxwWxlshILHO8/+Apcx4Xpo2kMfXPjDryw8PVaCvp1VI3b54bJAXO8KZPStiaF2djMe9pNC
rB043ditZGLg8CKws/tT8rGb2qEAjhrNLJ8N74V/SM1hKK5Tb4SJ9xJP9pPTP8k/Hv0W2jd6GJNG
Ed9994+eoyvIO0l5J6HKxrnK4mYXR/AZBDTy9rJsiIk0aUS+9K4v/zZ1Ne2dITL55rWPKGQs5b8y
l6O9g5Us1GQ2oDDdF+2jm8WDm09yvua4LoEmLqcGI6MxOAv5Gosz5QwvxhUaIRkvO07Nqhwe3pGZ
9BxtB6HlGOQWq1p3759pzkPjQ3UOceITSK6uteMHNPijIU9P9NTGxJ5GCRoIXjhNBKTQ8mr7IlEy
i1kFR+S+9waXyUKiVuoWsUY6RRIxRAqzxAw86qYT6swHbHZ8BCy7dligXXowvpkmczbHECN1d5Nb
OkS/F1Eu0j5Sy27yoYC0HmLjfdZ/6J4g5B7jthLpfDLiXWgFn4DBeLyvoSjhiG7AMncamgjaMDvy
52FwDV3sBtWxcpuKAMMv39EaZHPPmNz5Bj0Y1fvvat5wf5swbjz+te8XMr1tcUvxGwAQx3FlFO3E
yHfrJ9+u1FsGjvEHWylq+IwE3nU30mDYm2t/BS65UGfWgAFSfb3prMIiuC4ujHDDJskBanpzxBCe
2QtGq8obiWoFGC9+U1ToMkSd5oYvthWg0sI89jYtPG+qX/k4xCFQYlIRJS89/xPZhpfGpFxfWefo
LnrU8i5KaJ3t9rG76F+1PoaVMBSA0Sot1sNdgxsL3G1ZrM7AbMpMmyUfkqfNzMwr62VKi2DftduC
0MB8QTWwjQGY7j3nj3FZvppYIJCGern1Au8jTHZ0qG0OKIEJ4ZqYPw+JpKbgnD+QoAJ6JAlA4gO2
0MFhFK+6yQb2rf9tct0TzXCbH1WQjGXf9InM7o1BeaR/bOyNRF9OQx+7qUXk9nuQE5bYAfSa9ROo
eS2JmDq10wy9LXy/U3+88GxmzVASQGMoCuqbhRf0Goy3ZEq2PnfXP54x7yFHbm5wrf6DXbbL/wHc
XEf5CB8Ww3N4iuwQsQcXCj/SAZh+r2RleQmvbhUyeB1tYPKqipiKodVfQ47cpKG4QJjznMjWQN2s
VY8XEMwZUYL4hXUeFeSskV0kF7M75rpB0ifttfQCxTg5Kg0dsTKeF0iBHhnBP8ZHA/hqvMqhMDEG
d64DXw2JH9ru1F5ks9dHdKbqBONsYizPn2Yr/tgMKZcvpvw4GgsYjky4cqoSORw48Ix+vEMY9sQm
OqQSk3gQo4v3e+J7EzNCFhFz6+K6bM/uxGPF6HjcVXtTFtyDFd1KnWbFU3ty5+T0GHpYVFzkeJha
1XCk3RVK/pTig88R28YFAdek7qxttfdF2jyl9vpmsIUW0rNsAqhDG0JvG+1S5NMwVj2KYzYFyHNo
3T+bG9Q5qd2R+bmfdL25TJXl2FtaTt5/7LRHyqunPuY+gIrEXZLCJRoRswBoz2pHZgVL0UMtSVd+
Gt4DSwoKBUhhJk8wTflRe+ALKDshNVrEbNyOlz8Tf3enVv+ZWpzF/WqzzkcnVuwqMHXn9OYqfWqH
+Ai5OLsAEMxsL8unmlvfF/va1uyYV8YPiIKn7yFuyONA95iG5H/5usVv0wIjRV0z8dA+tgu6xTNB
6SDxNyMiqqzI/8Nnku2N9wyJmbFxzZhJhcP0O9qw3IIqIevoqqeKezWeEx6k83XBVeIyeQbYBgMF
Mk8+oXOg84GQLjAGCg2+FTa8QTGZcNn/RooUBeOJEVOQlj+1GFbK5m2ZcAuyyFew1REeo1UZLdAy
hvsi6KkwqEmsgZYAdHNXlqY2seXU02vVho5I29c6o5+eCxpPEmojg+GWXyTFbIa7eEQbb8po4VTz
mgpWEDsPXRfcZjyXh1sRGT4iKgrxC1zbXMR5oWtTROa3BCcAIswcRd5WiJ7le+U4kiC+tMt4D96r
WSsnG6pdvgzWthrp/LzZjGYX7yoFx1l2DRVXM2X6VBPuU0fIG10shWCse5o1xNN9r2VCPHNmVtI+
/ZLeHCuISwLVA7tc6Ykq68DRVqwMgSlQDyJJWB4pMicpSip9HT5psLSWKm/4m8xY2G3qSccFxTuu
AlvGh4KmZUTfIaFwaPxqAzTY1F3UhowHtDwSmgjHgJ89mBr/cBQCYWID9gfcQN/gR0ubRmlJnN3P
k0S7EmrRcwj76tDf8uZlfuhu/7vta83p9CPHGAkmnW5QCRydrxHtXsTPMlSp4TkLuuIyiEucLwqW
MJAr/inmzPoagCFhs4tD8p0ZChXjQvKR4UPjGZj2n1Fc0qaqNhIPWq3qy80Gn0QaKex+o6RL9anS
U9y6Qmnq7f0YA2Fzhi5PD6TJkk80CmNNBlCBAqZDAkUqaUF3xGaDy+RCBxBDg4atPEj60hcEXJSG
SxSWCaQEpVWIrjcq3VWsLaJsL7kp98oezXb6vbIDB6Ip2Fup3Wcoj0Tm0XKEX091ixoUSRkXW1E8
ZCTL4UKsE8gIogQt2r7T1CB5opwttZfz4rTI8nfQ84qFTatXsTImXas2m1KajsV0Ov6M8WZRlI5P
rAkbc1i8GwTzOq+qf4lnS92nzPT0TBHDL0dsiosOuYb1SAN+eH15QZrRLdwR25v/Y1PRqdSKGWOA
3LleqOaV8w4Uzyl50XNInMxKFZeWDZ7th6VNrY4/8CU++EVQgTo65q8xKzK/Xuuns9e5q8XF4gfW
68jMsxd+VHeEeGadgdvU+3O4td1BUoQZppK+TfTQTaG8RG4GNa//Vc4UFkWQZhDYc+AxCCCKWzz+
D/eX5hG+2TwaFQFwnYnYJbt4EYqIlq05QR3c8K8wOIsA6oULFAsGp2jpf13m7tN6TTIZ8Osb3C24
y39Xa26arkgzw2HRzvw3saVbqJddDDhANOaB+22cDELoXd+jXGn/saynz1vGpzHckAYm8vrC2Po1
ePJ7l+obQ3G/g1QuwQWa46a0DJfrrpi/ABdnkpsf7Kxu6DBe6iW4nYJ/TAwTlb5+Mq/xdF5DqZeR
ji5yLAzlR+Xf6c1fP2QXMeVmtWAWwBy8Q/XlLNAQKq8J5ZPzpqTSIVcdWe140Y65z6eVu+cUGPSX
3ZeEpa90Bu9JnHmP+YOD801xoVmXMpjRl4sw0Ue8kmUGvQ8HiOJbmVCaMFJjtgdsxTsWRkaFXolq
76h5Hw2euEBCxjZRBtgndhZNxZVmnob84y42IWytDHc1+niwgYUeJ7SImuhFzLpCrgdj3P/wlFh4
FtuU3dowkHLsZFffReQJaNRW2Vh8l8FwI9tKi5I0zeD7F+HNQp5S1sxPpqzA3iIAgMECgaB2ddLx
I8QzP3RUl2ssQcbMkaUT1+e0a1krREobKh+wICQUhFfWi0gE9nB4yb0mEqxWl0DhnQvxcHQDydru
hjA0ElGjlkGnBqEhmKt3N7cNu1t9M+8NM+J7W48vf5/nQU/NeVwLDep31F0CdXbxKGRo9Kj/6oFc
AX+yQLOwj7NMUpzR0vwUdZU5BM3x4j/ZZW0OBlGrGi5Sp9PpnBLZMzLkz/nJa+5bdj3ItfgihVWv
pF9utEcsgIhUE1/XsN/rOOVf/i3JQD4EjRy30k6gzThJdXWEDwlp7KRnv332kZij+/gl24yW0ZZa
YarAzsPvqe9DpqpSqCwg0CuD1MjOkeyZ/znSnRpRPS73ZwZmeHTDZXDqLiqFln6EccOpXUVml31a
rdUgyXs9qCsm26ldH9AuO3DIbRB/DYekaC1rrGZ96XoyrXQVxWQun1b8YAa6wfx3VGg4ARwquPmU
xX73rHxMqgEBccyxD7gE2ZxT1ddzG1/IdrOzR+tlQxoOE+TDivl1aeKxaDb3KckV1Afk5mq9ZTY4
4+hLnnN6xS9lQ3NL7xOxyOlXk9Lykn6fNgD9I1SxhTx8nNNnXflbFa8SsVf/FtpPuMvSFy2Nk/zy
wpyV3ib8JRfs9E8K1H4RRk1cFY/DzZcOjE1jF3KKC9Z7LKHOxSu768hSXhjNgJESDPK/YgC9CCbm
2Cmkl6VFaH8VVB7XLGKNZWzKlwg3Giu7Fm2IP9E51PDYwfPY7931a86oBxTFqAiUlpPSrj45V1O1
xfe2IVqStJUQPgyaMvg+67WiVXWgsLoxYvgD4J46cqFqnwbbZDXs9LIlJtblheCJXwN534/rpHZ1
oDgTlRexrt5ZCIKgqzK6WdkXUFGlPeVUdqMy81ZIrB/5OJM2YTdrZUCeB86OlTVoWGFeN+fWg06T
7DJIuut13luENuPz/5oQ2VKDm7utIXgD8FZ8NknRKJtk7N8vKPy3icMEw/AOdqJ257inXm6g6bir
yxY8tegSiy1PyN2jQoW+4N/HiqkfU+1dD+1Ky85qbdOQM75WNABcN59cOcGdK7W3jS0tNGMm7WTG
YZZEl7y0R0XFLnUd5p7jaJnbe6qJH0d0Nna3GhiEzjSO9cks73i8w98mDttDRZgq21I4YHNuP8d/
tmIFfCwOuhqmsiszw8iE2MRUuq5W5ouyOsCN45XA0A6673s0cP2eowdScv33zsSnlQ1V24H1ZAhG
OhGFgmKLontIhp9yDVbhAOVhFnlncddpYRJEYvfO4U4JfjZDtXcd3w2OPEhw0IIm5ze7aMdgC1hK
MtZ9NxacDs6tcCM0wRXSwJyhkXieWLrEGjnTkc20BFIQ1oBiQ0O8xatATx511Rg65s9JFyfbuLIl
23db769go/eBayYbS8QnaLedOuURR1gjiI1Bj0N+4iFt6H9rYmdMx5/CUCWyJbFpqjai0ZJHOyCU
W/rn3919zR94T+Zny4EjvkWjPwS6fnjnx98m0pdNgQg2jBVprI00xCgJMC8jjKb6kGbvLhWSt1mK
5DFx8pAIroPJWexLLjpGBNcxLXnt8XgtQBvGi5dmdLBO7I13KgHq2Mrh0HKRSfVylg6HaiyiORuY
UUMe4h6wq10n/NaZU7j2W0/RHjJNLx1sFOpYwf7jWoraJV9smPUWkdDaaQpXYz76d9uydanhn7wK
ydB3gFMa2JGuEgtgaykVJ29/j/QBsRquUa/d3QBjWEyLKjBD7WQbDTWiygAkdb3NueqyXxETVwEw
tNH6AfDYAnM139oIX7ujL6tE3a4SzDTMKB/Lww1CBhgTyFjVbo9dZPNtBL/+8+YP+C6AC6aAXsai
0EgyxKOQ+5R4XVXuQiDMAt2IfgLRlkPbFBLuDuXgb5yQFCXB/POYfrwCYq7aDiWxa3bdUJsKMTos
SGJaGWhlTEO2/4Sux6cx3pP9jM+4hkLZapoqOyitW0F+DvLa66BVc9KfHpHTcKCd2gOF5nU5y1l9
BWxoELipHh8tEa4sUZHV9a/SwA0zbUVsr7PrHBRMK8RViobXmZ89ub0guFUO2RNCexwpwUUADB7q
p+skFyKvPGxScsQ+CysimLBHm9wEbRLX6afneb23F8kTFEXRfmHYZzVEEq7vQ+Evy7GsuaNXvZZJ
Vlp8RZb+m0LXxpQ5FW3O01ndklF2xOtsfQ9CFxAXLx9NM/rX1p0oLDAYaEpS9Q4tzCVXRkFcrfQG
PY0WtczlJvEqBdS+esNM+/uejIVj7MFOkCnGA23SPzhUIAh7CDvh0UR8p9o95YE/xsQ5UoeahKvv
Fr2kRwrZidTt8GfUyIrslp4Z8QiImbwp5Zb60OstMPxiVQZAKJQjv3qDo6/h7vCsRYScZU8dImwU
gug7KAoweHV5+yw0nCzBLAngFJSaMTb2RnIK9jA24FqvjCHf/4K/a6ZKtxoFRhEiUl1bwL/Cz5ZA
5Wp2jFGkchqND9IS8xQHAALO+IQlwLxs3PQMrGLnV4utjLOhjumuS+itQIpoaF1Xvrxo75Z3K+TW
J0US0npknzc7enlPioS3S7xtlJWU2FdS3+ovvA0qO6+WIKhXVKUfYq0TJrFpn3xAxbaEcmk5XhY6
iitQa2epPPFeE8YohgmJnyYcQ0qiyWQKe5C9tMwM00q7xxfYT51J6krjrtK9bRtrbnmX6Rgw6lhm
WzagIwBKVFpBB9VMQyE59k0hpmRHTvGCdBDT5I+1n4NaPGVPCPZiHTlu4vjFwOWgE5FrcADnNw4E
eIHIAJys8BP5Hh74vZY0K+Qe6pHFJG/VbxV9k0/xDTueeXiXP4sTynRVTuvou7P1uFZDWKvGxBRj
yqkPKIvl98lWO76ooJsec2Etd/MiSFWZajc7q0LYWreN/MoyIi4GNcttrSC5ZnII8Y6UDX5anAOc
IFO/vF1XMs6etA7DlDj1im6iwFoqa41qtkt6IKIDtO+l20cTqI4u+YDZu6HoAUBzIwzxLZimhqAM
zQi3wmrahFU/o1dSxycs1//+7fvY5qw6BU1oOYX9uJK6ni8VgWI9SAneo38vaJTgsWmYskR5u/Rv
T/4VxnsfzaeZS4BO2vqQff9VG34inQktDur0CrO8ZI8vCJfcmSE7OFGLMGQ+ctW/cWiNaXuG0pfp
4xjAiLa9qJzAKO4FT4xUcBGdozDGOo2dqAegryHv1fTR/9Yzra++9JC7083goI1aQWyV6qtw8YvT
43Qq2xGggH/0XzT30CHEYGhkiiE1clro7Mrr4Q1v4KPBVphi4MXiQkrfXn68s9917H/iZ4hFthQi
sbJlj+GxkRpD9NGwKsS4qd4ETOURtmQlhixAs9Y/f6Rd4yxzK/s4CP4H93tTo8Q7GHZ08CScdfts
NozAaeYevXsy/Adx0mYOIe98rRSHVxaZokLqo0Fsv4+dvAbRH5lD38LhDI3iCvAMD6s/apHVhuho
zI2VGuJ+ODZnRbwANa/9ObyoI/Hc4JgzDFI2qVPu19yNGl4aSsZZP82TGE99Nn+98i/xEF+8+/S5
9ceP6lreS984BTlKMq7kHsZnE3ACzi/zypMeeM94eH2z529MAz869NFSwBfe7Og5YIazHI+jNbCy
31SBr3KPO7ozVR50RpL4dlsM8BVL/n99hPipPaYujPkFvaCnKrw4VYtKZi0Lt8rwX4Ot4fmMj+Zv
nIYMiNb7C0Cqz16a4idbVEKeUWWG5SYDnQu8CMK88BUd9SLFnDdyc30AlO7Qh43FQV3W53I+9gH4
dE02bGgaY3qFQbQ4xac1tPcVQhBeyonCBZgCZjq/we560BF5OEai+27PomEj28MEOg45MSEAeXd/
8T0Uuhlt2+zm2Go0DUFMPTugDo6/fIAeb/1N14sXMscFIb078RvlA6hG0UEuzOpPi/HV78IFdvjl
6v3TUzrRkYWvownhLzTPeteNy9zyTjaYvXofb3sXfZ0Lz1Ys5gTwuV1d2G+x+uxVrczM7VMCjnzZ
l1RlxOQt64fyVyC82ApoR9Ta9+42dq3lGWGE15a+rgQDIB1u2fexgZYRw/YtktVwpWP/nV8YwrNu
kfGT5QVxKtfNCdUaNntHqZdqiGJG2cH00zGycK+ZNeg5RKmbQZHrsQst+pNAW97oCAJwKcPO24cN
tuHDopsUbnd7hANtd2tAXFu5BI0Rye5lxJW8Mm4oFtoot+SpVsTov2zJBFb6kPt/GkrRcMgCe7CV
Q1AdDv4vB+K3fsS2NsdgCadadDvUaYSV6poLXuCh7ZsdHCWpSIotelhiDDqaU8P1VkINuywrAi/S
F5ulKQerDjcNbPLrw9lKx/eD/RwyD2D7SmAbbu2CiYBDW5vYUDtDy+lfkfu7rwnhIjRQ+fAfYVks
A6uqlmEQeFoq//rnBGNLnItZFU4E67Xfu4i+bXfbpU5LIcFIqa+D+ON/wnUPDzIiL/aUa7ngPM/C
jYUonxoWGvsa9sjCYmK00e7tnTlDWsMJRQ81OTat3yIo+wOpziZ7Kg4R65vrCW1KcQndFyM2UzVD
QcddPtPZZIOtot2CKSo+ezXpqcMUe6UdBghWxEtHx/t80i4N+LJmpqnPozY+HNH4HxDtwF4U43tn
muNfUYIqxgHWcnAu6L8DBb+M0BV/Vvxi4ZSdF+OOBHFm+AV915SLLOv5SxJnCmxyvjsXywD4eYTD
hfAOV1CrECsplAXlo4lFdzcoRBcaKVRl6yFN1dYfetbNRJ5/g3suX26Ge1H51hMsMLKKzHRRRUIm
vzgxjtP8bpTXgXJqDh1yJ3arQ6KsyWbtqs65tJ71JnjzpnBtzyQomjHBUaSD+eaOMTAZXSOb5wtO
K4feMo5JbQReM6132uR0mwS1TkgRYyOp2xCjBxWO0uDuWFvR3eoadZIcZkzb6+lt8w6+DF3Vn/A5
FjJiGYZWP9Ma8HsUca41e/7UYxH6wzJ93KV5D7DiREUGMVxXEn/N4qfiQcSESiAUc/7bpnTkibmg
aXgxbqs5WtEBjPLQv6Hg2uKhG5uxzUFr4rqr1NzzAD/DM4NiS7bHvQhSBeX7AXKudl8owMIkwAIr
a+AEGalSyzz01Uz410PBaJiST5yphQCNItH0dfyNfbiinhzrRj59dknI4i7hPOmGOUhJ6e+7ov7A
Quabe2TbkzQpPg0nfg6byDYuPVt6MafOk06Rg0aoQdVkltbFEQUKik8nj5/0CVqBA6KXVXlx66I6
9VZhCmpbEkxXDs1n0Gc/wUlC56N0DHsRpCToMhDSJ5tmfmNaMFtdlMY7Uz4YTMuFEUouTauI//nX
+j9rrclvgYqvugDe+M9HAeNyH4+wG5DGPL0ZB4IMgSId7wnx1NuMrDtLpwMNWE6K0FIQt/YkhdPY
IcH4zQkAkr6FjAqX9jjycUqQUg2Z/hkeEBr8LYqupxbA09qplQCAW1/uGr3P4A+ZzRwLHmMChXPc
Ip2pUp56/hF0BAOeNdQDzpnAGs90Csn+Gfrq3FZo8/qfjALrlhrFgQfoKcaOzeUd6+ymwqmE1lPe
0h0Yx83jwxP8Ey71Wj50Pf2fAmyymGP8XJBHoUKxvAQbA6WITSKFD2xSPDXkwQvx2IMijIP7SOo6
TASZdO2AYW1Jnd64wCxy1el3MWVefLPe8Qxe0YYSnyuHYhgW0cOJ80uF6mGmTaILPyaTy5sJu0Nb
IF8lMH6HLZ3CqIwOAF5oddj1H1LTSrFUDSL0k5D2swBptcZItY/UuZVaFOZ9SSDfeZWj10nWezJ9
E7WshJnd4I+MjnVoIU2vF8Jqux5oo4dBPypC+xLHeHisW8KJRbZSGjovPAq3ugBvrFTdOLrarmBf
NkEyrtvcuWG6JypMta4/qQ6z0leg0lPmu9KszABFHPyopu0aoRKg6HM4Z8O4QGXLHiTtpM3Mwvq8
kJmaz0aW0MRqVt8aGAEmtPnGXvl7RVoquAOtKX0+fajiEELMxsVKdeRe6GheSc3lNtW8SGQN/Ao/
BqlcG8rJdKZhN+kjcVtV+L/7pNRkq5lubMwu+nIbbmCQPYOmx4NpaW7Ee/B+zoA96rYIN4r2nnST
FFBWl/uGYygrgJxibPiSvysoywGKhHipVmwojVleo0oZRurZk5ZBUcRNFdK/W5D9P+CKtz+Jxczc
kBnLy4RQB75szVD3M/AklnEhokiNza38zca29MoZuRHeK72mfzpdJ/Yd3MOKDoOti4UjB/CzIC81
gn6GMDxCPRsaQkpIghWbZShxNEbQBtQjAi39+Gyozc3LXywoeynxURb53FCgLGp1ZbBtBnR3fzw4
fuUZONfY2a/PjSK/Ci44Jx3EjV00VXltH3v3V3CDcnKg/XHvK91r7XvuVSWz/8MZIisqlJsnQkZv
jqJVnsukPT+djKkDPXrM2xrqf9Swl2RbYnYDcin5gyXJH85y0bBJezqgCqFLmxG5aYq11PAD44oB
itfFhGm2XXJPf6DxTZO2quUxZBTnA9UvVOdQ7R0XKKEy9IuXf6FwDhGyc0eJbcMCEYIOiw0LGwhT
cd1+bxTViHDDskL0SjGsoGUjjrpsceN/fOXHEGqacDHx8WsEuS+Ua9u5LX8zMwPqpM4PkdjAf4N7
j6JA74R5WFIIGJxJXSuk1rExNblU5yTCTdcmvCcGVtQ6xG5mS763xh9nZEtMPOe63VUs34XzAWxb
TYnvN03pn22GmGTZETzpYjEKP0FeGyjfJeeVP/ibMSqlCA0NyiJ2SlamJE2CYb4PhgF3oS1nIGlA
zqX7okArum5YvX4dhEqL7DdsWu27sbgR0UfEzgBODVaJLjcXSIRrxu0J7fhndyiM19vmsZ4NCKFp
x7vwypDYzMVE4TyqMdAy4LwUqSamwN2oMT33qQ6T/G+2cDuYTFE0+k6f6+7Fv1vmo/Z2aeBcLJBY
/QvuDt/7fnXlfC6lrUqRBadZ6q/3DsHN1XSzzAEdsYpAHKpSWr/NSeCV8RGxL5vAyO2TT46Ca78a
j8zg1Z8n1l0r4Sebbz8fqXAurcFwsKc/j9lH/6RjQH7YZonbNZvVobZ5VYFZd68zWOIkMgmRbZgu
nXHr9nMBgsWzfrNm20xdPuWuOzP7CN20wFCSu59rPd0HT8ezyAm0imKFj5K+VH5Jv7rNnn0tK5WE
zIe9A4LK2ttMBfQWyL6sxkotVLUbnei4hNvWDxSoRsnddaHNgk0vcB9a1ou4vmsCB9TJ+1kuxaY8
xScQanGL2SoGO1yTVv0P76YsHZbjdAC4rnbdIxfB/1wQY27LlfEyg7bYiMg9KYmXIjJrmxR04fEA
GDdcDjWshrE7bAgvGnyxT/MpGxXT2o+6oGF4F5aUwKSPuIhyG0ctvJJcTBn9rkb+n0m6vOjGQNHq
gkbCymlZFgxNRq6atLy/QtbU5CPo1/wfG7WBq44kKSdE7h7dNC5rezO/fYQSTWpoF1C6xTsh/L39
XHg//ebS2zCtjxOs6SxlH2x+EeqgEjEZeFsayTer2pZSlECTjeK3smjzUbqhJvqKtIVO1RgUT9/I
LSK02umVBcCCmmXTXM46j1cmpk970MlMe3FvwgePJzjzf5rSTXoxNGXIvaCNb4mOcOZKC8Yn085P
Dx7kyPSIMmTKb0Rn/wIXnydbTqvT0ElX5pCTnsF2o9W8S+PKtrb3KhFBd+0trc++RpGBz/JnklRv
uo9f4IYs5cwSdNn95dN8UMppYYfK6tZnCVny0Y4LurTBKjpypyeIUOqTSvx0/Se4/aGlPLnzDIZO
feWla0WJT600nXZ09EbogdL4QYk9x4fc5md/Ci3/n8ekEP/ZrKMBUgNzy4IuWi2Mn0p6I8efRPn3
5/ItjhNrezgb/vzHsmarb+uLUfEUdsIj5spXxJVBUX5HioluQZO/3nUQdYRslj3uRLKrj7Xh3Lj3
U7jMKAezLURDyQnoHuYwUcuz8FW5KzJJ3JoeqHMNMTfGwM7UHGZ800Vkau2nV16nlcGVXU7tluGD
C8nI81HB8IhOLCypSbN6vyU9qRYXRzxhe7DpZvIyVLrSZfBERiT4V4h62822ZQ74BT6zpqwU/pbx
wMfKiZUzI+nutKoqPakiyZVghmpWs8yj7rp8vsjyYlReU4lll53HyTre5C6Ik4WdugRu2oV5KJbT
1tw7ED8px82fpSfLIYQHAdvgdElTl0x8N+diywWi3Ln2HyXmWgcevScJiYWEafi40CgKmIjbv20h
MTwej8rVvjYSN1SyKijfTF8isdAnaLqDJFyG/XfCIDtLUtrVIVC9Rwsy9eIAz9uU5Yi8RcaozePZ
6LLHiHuyhImMPi0YSW+sovgOPIEVgN32RsKDR3Si7BEYKuLj40sIEV4MBxmrKFfPLB6JgcFnykNr
Qk+o09U7zU6riEqdpxbeBY+Q9JSFnjrGamfkhQd4rQqq/F1uXZxUY7s0NJElvsQYH+qkbLdRmQl6
rd/rowy2QBmjHF9YAWvBdhdNPTarKVj+T2ztPr/VgBWteY/maVsrgyV7HMtXIZ2FLbyTYTUjcD+T
0MzHlcLAf2wnqemfiXUnEiDKmtvsRK8JNl5KEIfopLtgr54tSzRO/GALEcTRj58bVdVXi2qhgg4R
FjxqUBOElP/A67S1IvudrKqUTDn/eUa/pPKvYYO8lsyuob//goF3iQpct9HLquDwIBKxxMknRY/T
elAvXo5OKp1YyjFm7u0WTJZOoDCbWxq1H67tkJ4bGnXKbOXXoRXK0ggKCsgl9Lz/bSNKtqwzXtso
YJpBMNrKrEEZUvLwQPwlyP/ZDaHuGtLW7vW0ddnQgvI+DFodqT7vJhA8p65KMpAsaJhAA7rUtjnk
fp470H9MQFWFUColYEpHN/rt9llasb7o6aEiYdjN5VZHWcsiQnQJ1s6PZgQlQHIW6wA70mJAzd3W
1QxFj745dRgFOhNDUzNhVf83Wlvjnx90Ri2k5KNwCgW1rwiLfhfisCiKIMwh7c4rYrn9SuORevul
8rlEyINhhndhn0GwQq1GkDYlF1MI6ZXB6MFgQtJ/VUJPvYPCLv22+KNgSfl5FtaYvMgjTsSB49mM
A9cHLEldDyvktauZws+36DmTYAE7VcyXEIcdistsMuk4+3U2hY/MZdGawUk715Mb+MZyqI7uD+M1
yNXRz+IE7RNkMWNtO/teil5S/j2lZRI6xwyGk1WUvHyQ7wRTq996HNsqayDS97y/sml5pdu0Uw34
bajZkeVd7lkrmezyzgVgQ4nANe3/AvgDEo/7BMEZeE5YBiJ3+4Kra+FRdG7BZMHAJur1N7ZhA7fJ
w4m/zavZouWgguuGjiPdwxIe2cvhZftNVBKXBrK/DBRb/3TWD18m8JP0UDDvvqFD3VOsCZr9Av6l
jHYNtLu60VvBDH1xKBjuC6HxtVHWf0Habni8Km/5+8nz6IGlBTbZGPmJ3qzSfewz3Uql6VPPNlXY
WQa6NB6tzi/Xii8b2PWCnk8AZAfSO4sGCTJeWYo4EbENnpa/UHq8XbeADVIuHZdAcj31znxhTHOh
mA7NAL3bESC5oXQ/s78QHh6Qsj3MOcqdWeJ4wFoFbPlS9uj9dOgpoBZ/NmmC/EhGkvQSWLDkmhZS
5qAS8eFg6tzAP4EY0RfpLUFmSKk4qWo/Y8hjbJyjldD7WYAJ6iV1jB/Z+oLrr6sAD9uVw0kTQ4kO
ULrr07HJ+bjfe/y6lYtDGSW/bgqZeVp4T9KQADIkjrwLF7umEx/qxwOsoJ4injXYu418nUDXBaMY
nywkWnLR28jhVC1NwVGGPE1OEq5x/XBMODkZQjPk/Gi1sfYQPaDk18V4lVGlzYamKoZMqZSgrDd0
9IMXkNQtl3Rhofl0SsoA1/61jDgzqZ5uRZMYFP2yhunT9x+H+TJs0OLCZRZFGBT4SK258zEogdI1
EvFq0jMhCNQtf42hSO+6ewpWu5953OKgf1jvlDlXKAbILmlEfk1MMse3KWog2Hy/PqqtRC2YQ1s7
nxalQmOxC7YrQemi8ULFADX2jxVJdO1E5eE6VEzbe6bpQ8fuQTYwJGvoIjHsFxy5yMZlqxhPp4kK
kBOIAI9NHB6E3700R19NKA4juRsOc3PSGH0wVv7LmDUoGCvu+0vge5GkD/Sp+/fSXNknaV8rxFNT
vv6WgMSLvGrOeeDARJPp61v6ffg5dYNcMfld3mmYkg/E/C1RfDRGtCYX+1pzBCLSfcrvYmMHncN9
PjTGe9F+MuXQAujYHba+A0sv0DH/FqvW9f81uiLZfAstYi1MWVMfzwIQUB0RBCHy3NDYz/MqjDPK
dg8KC6pxJlDKbC5KnTnuvgexVQvOwS2nDpagPZc7Qp5KQ4Op7k8QtIPuuf8X4pyyQYgfznj46cFa
mp2X98RvQED7plz1pvmte1890vE27SzKK8prR+ZLw9G/LYv/N123VFQDnc3SrrMt3zYOXL4eok5r
qjiPxyvXVDTTx4rkABvElS9fgq81r8si065HyfVYGwYL1UcwnXhe7RLQi5rrasLKhEPSvPDSQjjg
7OhP1Qj9STPEVIN+2issqY4QAflpWXyrbi7k0KBSNVQXJ2sGKhxtnl495jU85PDdytO/xvn6RTso
IrSbKpCPImryZ7XUgJxD9TOgGDdkbWDe+TEdVwN+KuJeIryYLtJxEa4tODmzNDbQndBAV4gIqHGN
gJ19wVf67qGk1xoarc+vlIQo8YHD34YVltLmEzwROseiE9+A+Xof9poQ8LmF+7qvO4qOFurPhIsi
LXKphnPEEF72fgphtQGCXMPPsXp3UXxIBa6uPVWMhg1/8WC3kjbGy93KpYGMLaIF1ry9JdOQnmHt
/pNQmezOpLIoghFvdiCPZjIYb/dkYnGJc3WDZSGnJORRrqHPgxEdgYc8WOeZtrERxcV5s+FBQ/7C
m6zxNnIx99Kq1tp1ybjHiXXvqsWblOWfE6Jc43dfd18524DJHjlTJK2wiMQBZLF1jCJKmXsysqIC
AuL0rl8jX6wgG8WByiDACeBNZEBI78pMhT8+MWF0aPoCmnaHFX/vCy+IDUlCc70hEoosVn/9RrVo
vFAwGNIpv5geLlHCXka/wtsvJetaU2YnXwlynKVUM8Hqekkno5tAt4FNyrB6SAm2C7s4UXeNyuJ0
guFs/zZN2ddv1XoyPKZ+bAn4PvfnNx/1D46+xKAjn3M+kqWwRYMsI9KGjER2ImroGovOLXasdd8m
1xNpgesmuDbIMh6TKr2x0SyUWWUZsVoUjxwr8VZ0fpBwBhL2r9C8HULlOs2WDU7ZQ5J/bOTFSnDa
gar1TRLyhadaroV90BpfuxnFG4r8oOtl2f/5pyXmfJSNvtZ790HroGeKqsS2ruW+q4pvCspkttaZ
ConiD7H3AQ1H3k1MhG4iJ+1LCYJ12tcMSdh9asgb3g3IiMh1rKjYCEsjrLz64M+nYX01tWbq005a
per1lfGO8Iyz/yvQg1WojqMBZcjM7RsqP2OjrBsvjkUdbpclhZksbfb8v5/DT1JemAj4vhndiCj9
YXd1WoivlayNKj7qn2auVa7+K3vsUgBT6iJhkKKX6XEQQqgYjBURtJgKm6mODN230iQGoYbuuH74
mNkCNxwJTrJ1U2l5RsdEv54FT3ALpdbgFSpRZVPOBpHNhTLdJQQniwZTIRupaUivEZmMTJ7eqCfI
nhL4/64KbK0fW7d0ITMzrd37PE2e+BFlHMDnPs58+ROuO7ilH/z5YAR/Dy0FSFZtDQgwzK34UoeN
K15N75GjDE99jP/OEDv7gwUrXsQYeexkLoYXBZpEUvEe+ZH5OzccW8YdvemW+v/TwS8AR1e2HHlL
K8HV8uxg3QvtlRWIiswg4h+Swvy4EWgk05qO8Mo+sXWJNd4LmE+hc+0X1JavyNcnkBE64tZOvnaI
L0fWRHnMM2dRr6pXURRa60a6tyPAUOHo1qZD/VU/WBEjsNDYbVCYU3WcBHVQLb81Tr8HKn2HTb0f
OQzctrwkCKb9/qFpJ5vFlgpa8gnqnmjXs5nVWIXoAOKxONMVYtU6xeIopd/wn1QzFXsl18eHIBSO
c6G0bek9BeAwbKqtf5kLTjc8AKHPffNnMS6jhz93DdI9drmtxLKiuUBXps3Q4Tp3H6haqIUDqYG0
ke0cSKWPA+Aq08IkHZZVVLsYl0HoIw4vzSeiAlfJ56KCumuaLQJ7Pvj8v80JsvKq9KKzHbvnGBq0
r7ILTgG7nJYVoT2TcQ6Q33p3+P9C5ajFwjXkq2nlK8I/DWW6oByiddbDzQakhXZ1eDkNiJl25u3q
0YKE5A+voHWT8ZLOwy6qEW18/7J/iiuQbJAw8NFgOs2cqpbHgGtK/Dg9/JmhIfI7MnxXFFkxJHT6
V3wpMbEElXGox6fUAsiH9eC6lMC1hv/cxv0i0a2kvpxwBEUej4uzPO5DtwGvHvTTuLvkeTPo9s7t
v1TdjVm6x/Whx6cvwbRV4bQfCIrytvGfpoZPEj9oNzcX5BNqjCKxyP+XcXXdBQpEU7M0cLLyv6LR
i7OOOV0eqIhJgTxB81w5PjSTdGz07SNoNHKbXDZEUewaus+WEG3sxS/0IzWpdjvumcM1dk4QWhgF
+u62nK/7NhckjTIQoHBS7grykZR6sTGTpngczilx/7QkBxhO9wWBzodR2JtMbbXXVLnPVGetsyJY
5ZbwlSsiUB1m5h+gHcQ22G1D7Gb48qNSOUiyBBvdAd7+zf6RXPGnyWfV/Nid1sAYFEbWs4YtIDBH
4qn4MqBeNA1ygar//fANxuxh2/UCsmgtTsFDXI9/2VEHm79LgeFsa5VBCgToD0ZFPIixrs1BOoTU
zsu+rtIHYf8S6J/Lc5IEDmPRwyWEO9aFz2p+zNpPI6sDlR73rW5rOBOp63TY3LFDloRKrWsJwJ3t
fbsuOkBIrLY1tZrRgzveGWI3BtYSBkWxFlPDadcvNK2yNx2pZjELpkh/cjhqhQgFgUioIngmS6ZQ
/dL9jPcClAU/KI8t0X9kW7OwevgBU4JE6XjGyrTFhNNUdlMDc8HeZsUFtw9+PrT6Glvp6aPKG0wb
LjrpJkUUg87Udg/+dO01O3XNwhoQQUJCWsSu49FPYIH6bQUH+AB3MZ6NsMQ5OIaw/hatzH53sE7M
EhWEAKfisHL/v9VK0sXO7y2JWcdC26o6uwRzGP8BMTMg9I/c0/wnXMugFCy538gkQA4xmRWzUqWL
vTphpRANE/PaYlg/RqTarkblkY95/zlWvgGNOvqcndhpBMt3aX5BptldKX/NoCmEG/tGd6t1QW2w
fa5C/xC7xWCcHGFo7VlFmiqI2TCcMqAMDtwhjdCF0dvwllAolSgzBZYEPMpoVsaTWBRCHiAwZgKG
7vX3Ydb6my/+sNKJOLtwH9yUo8xCje3H2h2Rk9AkBl6I+pH5Lm8DcfduE+/itKOSnd1xOh1kHrx2
O9KcIFZOKFKlZ8pvlmHD8V9DsdfQXqfe6dtQf7pKMYciAD12OTQMrTlvwc9oIT3OjPtK2DLE5M9I
rbz4LZCUi3OcTl/OBFUVjspGHpQQKUVjHiUd9RBE+h5VTHKKOCKHjYRe4ynJrtxxxowNMvJiC1Gu
MA8pJFKrI7IiOOv6y84n+FEDsFY1fp9PYIUgycD+Qlk97kBr/POviMIjshkQpTvauqLh28SQWp6N
LfJnGureRJcIbvOvMSLNcODjz2aMjCyU8pXm1TfDPe2KSwPA94YERXLgZWWcnngSn88JZkhf+KtV
6OezR3WZWBC4mqvVLLRYiYEqMFKJyHZQtNFdNoeUyV+J9uxJ725Rnki2Fyh9y7SgEURg17Yki36d
i03xaDmXJSiX+0nqA7JtcUL0uzcSHinoBPDM0kX3dHAX1xDgooNGaNGNN2CaahjK7eBeIAHnIavs
g9iAEr2gfSPjnlLM4ahHYIa7Axj8Cc7kA1UFEKFuRNIj0oTdRHJxGMv3IoGdN8MSVdQOi8HaUXct
0NyYa8J5SlU1v2wsKDBvQ9iNqdZhVmWdmXPMTYuTQhF4rYLvQMXUo1DBIq0fxqbT9ZZt74KE55Ci
yHik6E1+6Y8v4I/W974frNE8yWAr4XwfbQB0H8+wS2EK0vRwLOT30pPHDbDMhVo2h5s8pUy8pbhG
fkLJTjp+BgP1tWy3PzXAnppkAuCWUyWDSVcGFHR7s1yL1sxutLhH/jDpKVF3f+3enLXtEjY6N4i/
VgFFaDPDPAnsOQ06KC1mOTzA8wqXpJur2GHeTDDPVf1vNxC2eBnPIaU0eivlMoCrnAjONNPqxJuv
9dYSZrdcmWAv/HRMT5De+3tSckwHuFVTu9ohqhZm3O0vYkYzLZbfp21Me5rVxg6oIC+fzhoyP2xu
PQxn/GPOum/lnfmm7o5U4O/KhS8WN4iPlg+kT5c6J9Z8UuBHwPMnPTur7nwYFW9RLcqxl32BQnVE
hOD9jweqP5wiW+f+VoCiakOkUJ6tpBCjf6Q5bzZVjhGKrjg7Z9pbC97YM/XVuD7/lFZ3yVuTL2/6
PnpnhkLkAO5u2RcbuAnzxAkOjXAp/1o5MKCmpzIrAuMHOdJnOn36H0WHpHaXi9+vkPvSZiPzLbF/
2V6GojtFB2D5ALss1hJ/qheWx6NAVqRDFw7USKdAjnthefUpp1TjzQud1l+j60UDWKBV/3XIMhvH
PB3tuWXXRPpxITfCVdZFlTt5QsN0sX1DfVea36rUvKvmUCWlqKJ2Nt2wzLDAJXoMhjzxvXqTIt/J
2djqt9AD2G3lOvaeNUslzvUfUSfkuWWkkFFRKNIR6gbDwhKME61MzQJnMR0Y+AGTo/FFaGkfZcbQ
1ESOF9aA06sRLyKjdqTDgXh3Enfdq/3QX7Vc324mzlpP1LWOUosdGZ/0Z8pU3vwfF/w6W7Pyf3O4
pBZmCbgHySQQlWj0Jr2xp39mFNBPq2IyhC7g2Fn+s0z/KKCa5TUOUIz5GQNGaydt0J6MPnhEoqt0
Swsmhq//3eiYX8w2w8Jc/pRNt5bNX8u1bDw79uusFuGfPRa95o0V55OH57G/untgbyXMLgDy/aRx
pWT3iKDUFk5JQQgKVPzc1aTkPyaUzV5FEho5tNBHuwgZk1SgAiItcr5vXUkvWJqnoVffQHdttKCK
3QqpumXKG3SZqRLnxU0fufRMxUaNHmdd0r/rB9aS/d53or+BV79N7XlSLJUpL0H3PWsU6yTd0coI
yizhkNWEtsd9yi26QjrkQ+kpcHbhc0X0rJ+V3BopOY/ryqpsALC5SdN7QCxu3wHQ4c/Ga+uyUsBq
lO08oOEDISDP/WmIYXu9HIkgErp8Bz08m7ZIZS8kM3SdQ2Sj+w5aj8tDOtVUw9J0t8+M76WpH23H
iaBKoy/nIXCR/J3KXX4WEYHCXFM0RAcbOH8/Y5bMpQsJkMqRThaouDOv3C6qtHfyaLmdvR3yBvKR
ZFCSIZAyHZw9p7XzqKQHxTmaO18PShGK30AMf2cJz0zNRJvu0BR86Yx3z3ZBHjorALxBD/SYoQsy
21QFJ4k8sh1tLZQQDCmTzX4OkxHrUFOs0wtEOT5G4CXveMV0l3ak2rgS+JUx1Vgme7Aq0xVRBCwS
Aa38CNaALQ+N2Lx5L7uwnd6PNNquWybiirK5pO/P77iLM/4BBq1tEyfAjoJ/EFvJ+1uV1rDZAN4F
ZTdGwMNJz5bMOa+wxRBUs0r7iDtESGCSEinPZSlE6axqWjbMzHVayoETm0UEtcFClqTBpldi+ItU
O1iUHiOf7isqyZMria+h//kYCe2Kt3Ks3Ttm9Oe6ZIbWW8t17WeJ129v4oSLxBDQgHjnDVErZW05
bTQxw8CgvBzgS0Y/Zsg8AAmWQDlgET7aqZn2cKGC5KhPWvvSZxChmO7OGbzzl/Q9s2FblXdsjIEM
7ko/ZlqWgPNq3FUVvhqIugJxa8A0+ZxYE/zjWkE2LTiyyUFxJ7f/uD6FhT0AZbQ1/5GN2aADHHE+
zeJE4s8EdjrPv0NfVPj5vpxnDhaaDNaNk/dzS5cPvVqclgwgsQ1cwV3QOn+0VPSjO70AInLECIyk
1V2LavEWVLuJxamGxIQhMQS9C2y2z2nWRIua4sksddanXdvq54hziyKqLKkZF95TkpYKjl/Hz3hN
YcGZVpvNOWvg33myIouHh8pVQ86FcNJdBh6+Dm1T+wQznFPolpP/sZYp4F9yEpXrzT7LaF05Nj0+
4TwNd96OhHsBkChJYQ7jVr3OD6ScSzv93ud+qLbHwVGvnsFhYh3m4S99m0bjhFilFHqR8X33IlHq
SSxm3bgKew12zVI3VRiIkfH+cbtXpgUaf2VTx9JX8/b5Jo7RvLhMyhYI3yvYywu+JcVGnEveXOgF
EMhkS5KkH6DVZRqWi2UrGgTgOMoTNXP95/9QgLxDIquDxKu7KLfUocX/YjKeOS39aJ8OPwug2jcr
0j9abvJGQQa8oafp9GtHyzCZ9xxLugqyA7n+x/pKnXIaFKQvronrQnJOkd1uTLnOk2wgl2J9QSge
fVzvH5DUEAXqBXI1X5ZpvUS6TL9Fq/kiAc6+WGrIJur7z3Xez5QDbSRnMxo0KWL+sFb8UBHs6Tfa
nMIJbECGWgoFVdH3w3pjhVvPasjgkksCrx2MzSW7JLFNLeD1O6w0hYWxN6x8qAt2myWC/V7zkl3z
BF3+b4pAQ4pE6I2uOci23tOwn81QzLkkH8YXgfuurvEOS/fZ2HEP4C7JFvMjRMT18+dwjb/PcwY2
f+M5a7FTSsOJlX62wG40KXVB8MGbqnreUIXwzt/M02WIobAd6X6O3K0x9hDmMBevuu/kmuue9iwN
vsjL49LOKXqi2fBXLYEuAsZhP6J4aVVEbHLN3Yr2bG3lxqQGrNZQmTIXgahk+x2wUu6ED74tj7VT
FaP3Z1swh1Lfqc8Qy/frD5qzU/mlyQbNsfB+QPBntc3M5EqPuP5mSq4F8c6GAFhZ0S1QTxRj18Ao
esz4TJEN2LRmYN0aOZK16hrLDlgAlLsi35bszXXu+2/hIMiOw9HfYrNqMHNno3RLvuUV1JP9ZGdp
EFS/vzRiNOhNifYQUMmt8zW7eaNTQNWix1Kw7uNtM0IPe7H0crGeY4XRMkZ22WDPJ5eZleo90Suy
lDtWrqBP348GHfT8LeF9kFF8l3LwGR2EZysNGATSo6qPjQJhs0ct4sb2IM7g6hmmftaF5YpnmMjQ
gO8eDfJ2zZYqtmq7aEZ+FHNnB/aveLQ0u4cz+iEAMfAlSFrsXEGLQkbYhgkmgd9xdb1eJ3xSXDdt
eUYnk73Th7pYO+0yIyNvM/7p5Kkbg/GBZwhhZzCaXbGYL4JkHvIizqGjenRSmqoNXKjwq0EiQhuw
tB8cypJwHKQb2MGxvBFwQ6s4gCsIux7yXe2Ic6oPJhI0gMXgahpFq0rAf0pvCx4j8ZDpRnhTeJE3
5L9eikh4EFw0fc7YgKJZCGSf+Qn7UAuBBHoMYQdpk+zM11ygcOZ/4GaqpEQW0McVrCvrPlyPbhnN
YJH8CJzdnxzMx5J/LD6+ExTlrjTfUTvwspCPFhVK2MQsFtNQjxY+AMLUDBNIAriQ4qkODbWMETFi
xAwZZ//H7q3rcFIgN2PfZdZ90buZNiVwMggYO/qOfKTvpjIgaYVXsTfXBqv6XK6oEpsL/TSvNdOh
S3laVVvXY2AsghCQ/8sUXeG5MHIOSv7J0WEG2CV3VBNB/PO+FBFh2qnKtWmF9Y93QvUfg/VzcrWu
Du7sEsZ5g2BTWKi1ScxngUzH188QpmKEEa+xCk3qU/AU+3uDO+799jWQNz05ZK5vl9Mhz08+Z1ye
UeATK34hs1YIGEvxIF/GHeiE/CwwAxldhtODfmHNpsJ3zZlL1y++dku0aA35rEcxG1mAg2soTxxz
YHuLc9WGhs1Wb8ZpoohSwAnV8bu7PHmTGKONR2y4o4I1yz81043FdCEB0oEx4ZRQfSBjX7IOwnvl
ch4gA6TI7dVXlrAN29TnOzcpfe6jFPsbTUnB1qrlOpeQpRtnIfAAh4SBAZ7NHj/JgLZ9nmhZuLNI
x7IQQjGpIsqDTzWNwZ7HbnRuKEIcEeEbfGz7eP3CVUTXk60bNCG3PeK9BwAOximSb3KG1f7Z0fl4
K4JB8DOK7dONAP5iGqkNORlUeWJ3IJf3CvBAXIhOknDYtOADBt1aSSuJky6suGphZKzSnl06TUu/
xLlLEZSmbaP2aCmYwb+zfmVgIhfXDSx6yBtJOZgbVbpurcOPvk3CjCgNblB+yDor6FUEIGN6Btv3
IrwakCu3JdfyWM7VT1a3kVRBqkgA/lxfhHyroZv9mJerNXRaB9Lint0v0AgFtoe+TbBirTmByj2y
M6uP5hmneqDfJBEKmxbB16JtpDU8JOBJdtEH9BFrRmtPW6na/jEDVWYbbwhKGkReNhcscbsb0v19
hNPll4TVsOOxoj0f0gVBHrKyq/gst/BXCL+2qQ06yRsDNYsEw3zJ6xazrzg1dzclgcSz9aLAqZ+E
dEIRZ0PxBGXNcPEHH6I/YHsfNaG/sJHjV4elAVA2lDyTVGwVKDcg3aQlI+NTkxR7AfOQJlcwZ27n
3bz4vJc/6PnGQi36H6510isRGOgx41UgkH1/al/cB4y0GFFw0iiYC5ujUdcicutYC3Wdwm2LSuyM
1RrijCmMlSEsOCLXHA1jnL2Nzasa7YZXEQS+E2npZ8eGFIL7j/Irciy2Dv3KQ3GgarAGQ76LYz1o
AucFZRsi3+8DJXoexQwfIRJ6kglfJYOjbkrJaYcgT/sIPrgwxBMDuiwxQRF9Zqx/C48n5kthgPMm
k08HYuSwofu6XWEKvsCkl3dy4MTh2xHYfsmN63KFQUcko8egT0yqfpZAMTIJAKN+ax/e57AH26PS
lZrPvgaZeJBPcgPwjBL6uCOUdvbDr5jrPj6YxUarZBGSHcXnCDp3onaWmJSi4GCrA+c234uGzWlk
+leD6jvnrIgXQ5JMNLmhPt7opubkVUxJ0V9OnmkGrBr9GH7KYxSWpIwN8YiQ4KRapoCRKSFwRqUK
ftWYFSvpBt0ue6ePXeiIDQ46nGN8gADtEleIAn/dZIrOO2fT3JzdYED87/Rpw2BUGRv5hebZjp8Y
/ZDZqAg/ajLa5XJOp5uKK7RHkICTRlHY+YTqpB2VlMBa55E5vQxtj+hG7zVDQQbqM12CcRLE2oPt
8TJOrj5perZ6ZvzNbgkfsOXI+7qL6eTiIPyJ2UgmCgOgTq2fn+ZAX6vwzHhzI40M1WllOBrj9AuD
n4b/vAp4UWZWi+vxXGpF/QyUcu645FzxbJhGRWWYA0SQJMB9eRhRkg2CS7kp0wfI6iwfCLqeodfg
e4rxwJumbmZin1e1znalfR6H69l1OZ9i6dxHWNayEQCxAzzCtatCdb5ZpLl5SfiTUQQ3s0ZYdZVe
2r49Yvb1kJPM+2eVfKnCImok72wGCw0UP4nBty+znqbS+SCnSrElkK/SoNeFvvvNi1wscL1oWdxb
82yOSlrj/ezxHFebYZVFdS56ZsOfZkFCWVQHrWZYjhCA1F5PmdBxqytgJk96JJPfJ9VHLA4sJv8z
BmUl3joD/UL0P+LFK1srYzYJ1AQBmzXNjF7/pnEvYBHxpuL02y+asCD/zXGoMdAkTdeGMs3HevUc
CTdbYXMNUnsd3Ymwmrnnh8CVdxpdOQwt6JiCbYWra6/lA9sb7guFLX+DhMhQPIAfiVDh6p0eHR8T
2fhbAd9aaAIs40TSkkSepzf59M6fl3xF7l+BJCRhh5xv5BHI2gxnoK4x1lxKZVfDm2PYx44fo7KX
jMWcN/4DjauR3Aa7KSB4mIpvSbykodwZPBailZb+2THjYeLoMHSqc46Iaz6XF38Np5RSHM1ws/iQ
l6V5zOvpiOiZaOOi9ZUzhN3/lrXez0LLBlxE4nC/7qzqm9HjpzYOaVwThvrdRXBsMfi4y+kpHq63
2G0G41Wv+yZNBaPcVnoBzSocUFLbVMZI2R7M3QZdH6W1n4mdi7k29cUR5y2LuMKJz8a2x/ZkW+FC
Tu6waPSI00fnrkvXAY4eCfsl9qSRRrvQumjYi/BLEBiKnP1+5TTAsDfjltBQ7tsx9PL7VBmJJJ82
gJ1DP4a8doN0yMMtC8hzDWT3yGK6buZUC3o2xGM+/rM+qLhcxQBVfKbMzzRxmSibD2o+84ocngRc
coanwaPI4EowCb9d1iX0V7HtkjBXYZka/E5fq/WrBtYtT6sSEDP9TyD2MVze6e7cT5eWSi9dWLA9
gTZxYqF+phFs7DR5aMYydyzPt1R+BBP91mjxo2tetEWjuorlziNE05fyNsL3Ic11tf08uk0l/VUc
MPFsovg9Ywk6obopC/0Mcg52bePi1afPAx0kL+xbXvX9epn8l1ekC/hlHxELYNR6+zgDnZtG433Y
gKm/7EQR7nGnBhIXo7Dm+s0R07uu8I2dvG1ZpG+25u/NK78kt3cO8KoBWVQREyH4WIfUOZejT4VF
wb3iX1XwUNl0VbfnTFY9hTNgXObXQ7TkHhXLTxX8U4MLeX3WuLsv50b78USI9NADWbscevY4pEh5
RGLYp6/JHjchS4Yo/1zujrpTYB8j5QUYq8J4lrfEgou29g4qoyG8+QHip8xOz0vfUBcQ6L3W8+eW
75tP40A4fKHThEyA0Hlwtd1ddqZZPGkisVO1u2L5m68BT67SBEoDW6Tq1JlDmmW6wdoLCVtEnl/T
e+OyVKvTZpuIgBYqhs7AQEE8S0/UdM9BzzLy3XWZsQcdIC5G+B8QS+ySW+eBJgFgA95H11WipMU5
jNlSACYzfJFimXct4lZNQG0O3GoU9vFsAg6PtAP0zoSgf363g9n6aof5CUW0hbpFRpjxAyujvsLN
xPVG95n6uan9E/adxx5gp5Qwn4ZVePIxA/StZCA7IOlN1VoL8VGKl4KbJ7JCtrzWAIxB9CkAAG7k
N2XpeSFHaQpoNQTz1fuX91lgT+zWaNP36A2oGSOMyh22It50UjAK4IE47Zv00Kdg/6ub+F2tn8UD
H1+YxIsDQB8jstxwG9CgEg48xFwqjndX+mlH5MqU3AUqMPDf6mXb7bPjQJtK4RaeL/sztpP8v9au
51512d+ULGsKJTP+weKu6XLYMqGB5JxnEAIxtlhPvFz9kgfsGQgAI2HOMBUPm2ZzaxAzScxVzFgy
bWUZBiJs9cgR401M14DyLwaaWjMwC6k+QCCJ4arez+Rhzesp3maSaog2LjOg5/x70TWEhiCvtgaa
Wx/9D6VZR0b/7nJxSHY53//Cfv9lmLSsXdjx6Nv/h3gw5xwEvSjoTTDOD3R7BYP5CgH5HEAqn/Ck
FJfcnjN/WezUk1NiimZ24GflNXOmpmCacKbfrRYResaghG+O314bZajwr6kRUpATJL7z2VDAFqx/
nTA/F3pvMYMRCbxIqdcasuMlZVszkx9LRpVnbDlamnSIAkDT16RUXD8XU2UJaSNMNP+KZKRqsERO
cUQCiTWhKuE8iClnf6QUy/FLKUtEFoeHqPWTX7cKkrtbMXmKnVjr4nyEKMxZjVcshWEnS7y8oMGS
IO5SX0uPg8Aq9ziasx74yJyoHga1/Zopf+7OJ4yhDsH017kYTLWohPdzNpTn52lD0tQ0nCQXC1wB
bo7W2tC8Jzftx3r9VA+noo697z5XTYkG85C0E/hUHHwWXJUhhJxBUB51Bma6YaYCqaOUao8zWY5p
pABhugE8/WPzqmSphyDaOQz/37dLA5eqDVEFs3LRTKocvdCD5ux81rTvLl18XKZkB2b4mlFzF5jf
KUTbwaqH70Qulfbw5yfBueKpWN3dJ77aneGwfk8TMvFrhx6D4fUpQGN1fmhQYewk8xB8XwD9c0Vo
qImTivSzoZ0dxpDCHgrvLhdUzm2GYJ85Ov9YGPyB8VWc60RSQWk5QjIcrpJER6txwRXjmYLQcVCd
cwxkbbULgKtDk6ef066Yut952sU1HbKUqH4chN1kTdO1OHmQyBLXXi5WH5e77FNsGJaRrrsSvw76
06cwWdhnJd8BRHXMN7kjAf07hkmChnxNLeAnzNpW9CNAO5K3LENDzHuYrWwHMR5InnAriN2ZM0ck
nE96S+DBMOua5/vjk82hvdIbqcPY9OWNo8mZOFPqzNYRdT6mSxIjxRSgxjIQCKySnv8kVAlt8EMy
hipkjWesC8ykiQB1vzH5qJqJV8wOIXG0IUGu4MPkT4otok/ipfpC/GUsaKJ3hBxES7TKzSfwjoBJ
mf65LRVF7SAJOwVnbLcoMLFcWRAVn54GdiNGUpXdjJT/9VP2LXLGmWBKdDsdqRRmL9LF1KfUV6Nb
xu2L7sUhxeokIf2cZRminXIoZ0t7Q272WlHNVjGwqtKu6OmpCAbAb5GvToaaZ/k4Pxv/d/UTZjE3
yXD9Re3zVFNlHfo7jdgCjSNusIGN/JeWF8ya+h4YaknlF3hGA+U1zHfayNQvrk5JwOwO6tWoVSmL
cZxuOtyD1+2+CfS/0+mOIkNTQcFl+fAm6ptGEwgVn9J5IWo/qVYUW/Uag5fEsv4SnX262pLHduRr
SQm6gTV194WRJ/nJCf0Fz0ue3hLVsZPuGrDEt5bsZ0VemVtIcXWX9kpGQ6B3OklheeJMolXv1L1f
bNq8lvrtvQHkr2hG+spudcTg/EV3oJymAkXlwAtLnHXRjKY3JZ1C00bniowP9LCdHK5Lh0S099zN
9x5QWCrzhKks9X/1JIrdmxR1MbdGzwry9EEi9ENGVl7pizYCC0kWmicIoOx3x2J2XoiXfk2cVBJ9
n3Wr2cYmSDXkRwfLi+TGSK4tqJFun5ZSrpc+cZCM0rA1KRjucXRPvjyBiMBDt8oLXEnG06AhCBJV
B57xyDKRFDzbGn+qTvwta2ITHdpR+H4Dx86iEeF+Y+lg1s6YlHGPisJIoL90BOPedn2SJH+rr+Jn
KQ3nGVMbajIAOozOBk5X0JFBCVgdjGDc2irLLY/vuEjMwO2WOoXXRZ95UZ2P14I2yz8H1GB3sJNR
HnjTbC1xdRMuiFqYM28a1Zq+38nCgEqNFnQAJQtEbJ9vSCBO7XXfOXcuTB7yZy4q9IpdmUCLepzL
sE/IDe4YHSfRBWsPVv5Nv5p4m8HkmVhNH/lBSCQOOjJJyYIN22JKUzXg1/JfZsUk9/CqqVgEZEkA
aTmp2nkxug/Xq2L5eTIU+3atM0X0Yhx84mkAdJZ/btA4sttFC3yZMFntb5q+PSybs8fyCmaAT42r
P2Ptxrt6LIbu0tW1+M5IC7gzRqsgBSQGbWicONJZ/fNYnNkMmKwQAaTarFooXr/yksHRXcsSpRQm
t6BJkVnr7S/yrDKkST5zNL1DgvLhMBqlIo28aFh7PqP2YTG+AIr4zSn1aLeqF6rzYpJuKakkDizw
deyJL4QOOtntvqGuoukkHfo4CW70nLeRuZpq1r5bgqV1/tloulYMoJ+IZPGSCae5yAMpaNoOYJ08
r19KdosZPl5FrIKBeO+GCUt8a0zUGRCvM/hN+1rx4iF8jJy6HhrXYvpXdYGbNwmUE2WXJffJ10wQ
8vbodfz/sN+jGy98V15o7bo2Qxj3JZOkYqChcJdGsWmwO5b3lbkNL+sWeUufweGHgP9cpnsozG1T
Pk+UAwhdQoBBpN5pqOkOKvRqurNPKh4KmE2F3enATB1QZozxX5p9KgeFfpsEEed+q8IUlUtfis0k
GimtR18AIGVt+xKz0XMB+NG/T5Pvw3sXbt+bWWljbQNCP8vfmWHmNiUIU2GY6UFJAbHTRIsE4iGr
EehO79dGFx1gzHoVv0Dp4Bi4TUA8dlZlxlApzqK3DKVJ1opAhRVJTPr55YMdb0NJi3Yp5+c10D8L
qaYwTmnBUJLH8hsUaSJJaWwoh/LBQec6VIBgQoac+VnApChMXyqEvS+L5iH+tWd/PEo/vIG6IsFI
GolXP6Y1rocFOIIEYVrcZBZpDaTBqgT2k0PLytpwUqzkrmFgWwk+uViFqPdAt6IXPvhRNRG4wyhT
RDkJv9G76l4jPzeBifz0sj/UCoeFBC/lObW5A2BzmfwttpbSuLFNx0sJpqDsdqRUKK4lZTUvOrHo
k30SX6CZz8NGgcMg7+KoUsmcl7GOnahM0p4KgH746h/6HDltSbuCqsf9+bfYrNWJAc/5KNVvlFC8
RiqRJ3Vf9wA7VxuZI+WIzVrLc5X2GkVtfbTrHzvwA7KrTNqX4CmJa/bJOkGlYhV5sBHR7Fq+9ETN
op540C8Zfc+adrhRsjiRZQ6kSmTwacp5YORCOeECIgw4s2cC7FJTDJuYCBMzu5ok4tuwRHGxJER3
r6W/FRYJ0YMToVHLFG9B8fCCBNmFLInrsrFJ1eSj4HBvZW3Vj6pXN+4pfDFq1FSJmNbRpwF/z8uD
CT6UA6rCJOfzwzo60Ntl1wXem2+nvSYoKvFc3QwlaXygY58bSH1IeWUBH5UMvOKqarUZs+6UXID3
VuhjyXJtLV+j452G3Ej73MCn+lGxfKud9iv/ir4ieSQx3bpqnVz2VeZR4qOcY7EX3wnsMO7qiGKn
wIwmwp61qARaxhfz/lnSi83NcIfwff66u2q3VqinEUHrmonueVikOp11t2VEyjjpzgDrlAxGDIcG
vB8OgyaZ1dctoBFMVieVaAi8ubd5ZnokPgg/Wk4e6X4B5lHqtVAzfJdm+zrpEWYrwaqexQj5jmZM
81NIc5i1vKcMm4ZYvITO5b+w1toHvCuN9XzRf96cfjo1CgbnbWysQ/8hLSVQ6QhgkYpYYwrSCHEm
gsxqkfv/ElAev8Gu1JEpVPATEBjvNN4/6aOVu37LzeR86sduSf+nmpVJUO5KMUUlQAopCYkqjU0H
im99czmtosMqrer8h4x1qley6aHDh1CRjNIYkJBxclCoSTvnraKuK4a//tyMRqynioTnnveYJ/xw
PW5xrJdaJeUF8TZcKQL5OI0oJWgfpf/mbADW4GsZadbmdyLY08iS8vdyeNDykVc9WT3g0whGH0OF
eiG+9yuyBcMcOJky6e+a++489pOh7oYw8VrlB9MHYi8BIM47rlhqqgqkSm0HhSN5aXP/dv6Dug5a
IaMlViE/pstRhPw+Y1f8QiWFSNMI1RtF6Vcqv6A8O9kmcv4OFMF4U3Dkqp/rIcBglYi0SdwEqlgQ
hPgfSe4QugthBrlXXuRSPP5ySchKd3570b7ReCRw5A4tG2BA9ByhtdgOPD/HVeKJAwB83UIDqw1n
2b2wLPc4bk9h9JErN4XRec+f+CSgW3/oMZ+gj5bo8ErS4JaNa6PkadnBvzyJ0kJkxknsy1GURzmO
Nzs8UI5/R0IvJbGFcPwW6UE/Qx1uQ/1CuhpUTWFEql4OMjTa0TtfjyQB/mzpbzLuHwcGYkHWtQvL
pgd9TjEOBMHQLyvIrQaM50w+5w2fF7Gvk536SU2PqLkb6QcPynRQxzkHWGz6zSbTQ8DRJ59Ve3Zc
9u8hqe1hD7eazc7P/ypFiaLXLXRuuPm8q5hTIVAuUPklGfMiIiPeidRV1XJq3Lq7wSjBkTClkOWU
NqQDJoIZWMgyJUUFOVN1XXoesh2O/1a9eQywsi2dBhnVFiJeN1qTR+DeQPwNlgUgB/lqgCiWl0o1
AmYko5SVW6nTtqsPoZ+dubYKsXkDP5uBfgXAQqWTPJhkRRc5BtgIl44Idocu+rGq5IDk3blt6bt7
XBpHX5F/LsfRFPd8RP8LiCMkNByuyvqtZDn/Vcc+CD+ur/GNudoaXCKyysv6Zzx3i4KUDDJtkRe+
+olQoHcfQxUiJFCdaw9rO1wkzxEEY/nzujO4tNcSU541xtKzXXTFEKALdJGPVeFMynNeT+BkVssN
CmV7JVTCFmebcWSG6nAqQOhxOG5fiEXC9YUAHGMeG15V8gYcebjTpVkGCmpJ10USfjz5VzdXlJK8
YqB5pVf1vOBwjx5+eN4MU3i4/6LlmmI1ZFvqe55BHtREQDyxw5VDPxQLbQg8+3nYUAYTihBE+Iba
ASQE31XRgS52DyT84K9ibqkRh+DsYD7/VLrqvCPaMAiduiC2mIYB+oGMDuIl05jUnExYLedx/jP3
gUQNmPAZn+wCNz2JNBK4wjY9FQOOzVYCrEHFsug8NySWGbbV9DhKSihWt2cWNXT0hV8+vdyXgGmv
JA1mqh3n3FsqeQVhaBwvoQMonOkxSCn/Fet4EvhGfP/0kgAY75al18jn/UpT0uBafjstxWhrcGlm
gMgB7h5IN2ybkdJEF56YgMYYWT1UWWYBVfzXWj+3CV6LWDLyrBxdXSZ16G2qb/NDjqItIvvmfXlJ
lT79eDR7pSeR4IXq/OHEbEo+TenwwUZo5tq8cx32gB9HtTVYfKHz2dektTAvx3mokg4pde3JR38m
uwMDS1k0q4m3N03RSbWOi3sRPn3FuAFFd5QN5q2wOu+Ixmz5TwEmWn57jEi6axaHQIToetM57PAi
JKaXFohYHDAOH6yDx0AQY1OPmwuVcp8rgfDMEkPNVw52mHAEXGLrsWDJuaGQYQMapvjLbAmaX4TG
NEqSrAiqW7x4XdSiWnvxYBpb9mDaGs6ipYtmaBCauPbkVVfa+jL9yKclJLxuqXuKCJNKf5jlLuZc
qaqclTh9pRgC5WE9rMOA5hGJOObanUYRGjk2I26qzz8X1+IimdhQvZU7PtIwSQLnJJCI9jq47awu
V7Rwv6+jmPG0D39EzotbcfR3HEpk3bFzzITkKoUzJ21WxApqZ/BzwAGGi3ZNJz1bZ4qtdNPH1nvl
kQ5/9iUP/gmnUY3bnAEfGlwlp/wZgyWk//nMfsbliMSWLavyam0KIUpqp7XP0uDPNy4lWzFWH9uP
rAJGrsJmPiwkQ6CzY3Y60P507PCB1vo9nVHfKLN7zfSMTCuRJhlw52vDH24UzFeASArnSMRTS0H5
MtFpffdKS/FtmRV+zSxCgo2u+gvboZ/S2pisQO96rU/hjKjRLglNZfvcvgdNcfm76+TPSyodh8+k
OIXh7AMmMR9Hd8y/sUCKWSeQb8qtT3xA5zCRTFYNV9M6bboZf5yPWapa2kz4Y38WmcNWxoRcjV5j
9u4WnL+QpauFZPFFB8gznp5//rvGQs0x2lMQZTLhG2Nzw8UKBO2MXvM7F15TMrlGZy17cjwjMwIE
VU2afqtqNZDgflVRZofzDUJ2ZVFo4mJGJKbtjle0Hj9B2GUrcLPqu0Bi6TitnLr9CendsdzVXM4d
AMZq2fQeEf15hrkp+oaD6ReGrcedOzvlAvMCb7w4NXKsUEievvkk5RV/A3vEQbldZuUhk+9Q0xMf
jR1VGK1B2OSVBlKO+2VNcjrRM/hmAVK6nutri45MxWcwc5J9FCyp+TOHkwp7KdGjbldLfMVGLBRQ
7DlHgohQGs5gAitlsO1f4xwdNGLGXAA0rRS2jYr8QVAilWN23pxq23XIWoW+akfLulPO/vKMDn4b
cA3ypllz9BZYsRxL1ZeMH5tG1gJoYs1Tvp+TH3OBDa0EQvrGxQ0DxqttBbuANM9id1zwFprFA0xe
Lq1yZiT0HGpqR/iqR+bCSG0qwqebF/SygzR72VS5PAlAXI5xQ/RkNIAPhpIHiIBMjuATPhoClncu
FdRSyPF5QbKbMUU9ndMiozxu3l26BKNS/OVDWiSDlzWj6UUUXqhtS4STtsClDFhURfRgn82hW6Zw
k3xh69SXo7yQSJM0gEliidkbiMDGjSysrbpuoYHNwv1qQ2UpNxzAL9ToR1MqNfV4dVHRWdBFAiJh
qQ2Z7jnsoL2++3KoxGuMXdYyqrKMpItWJzrdlPMAObe9YGUFvODY+TDHv4QlyYvlofxA6NeBVV+E
wGrCPCCCSdJVkEVxQyn9e1mMnlCEnhEPIca5OCwuyOXJmz6i/RJazmiNsFDSWduFOc5lcOpJzSJj
LeHvAoKigBK3I7mHqYF45k3bRxBv26JnJ9ZcbvlWDo1ofZ5wgtsehj2XSz6mnxmYmiweMLiyL8WO
5w/F5wt7jq4BUHV307//YLJ9zT7m/uFkT8PLhkRcL4zWIPXtO0yO2rQRNlROPyUXOq4OXdsOySBF
cJHaSo+afFdIP+8gkx1aIFCh+4U8h8lbGFu2fI42Ini8IomZmxeDNfZ60kvEnwMOsG7tIlTACmuR
iA6LtagYDRT+fzIngbyXWu0n5W4b+F98xXE0sm/qgQjG0n80FyTeR+AMansI2ol5tjq8Z3ch4fsV
R/JzKw8DeaXpxgdsVi4eb+Y1hMK5VpSHIWQuNGwDTZU7pgPkVNlSK380XS0tfMQ2KoX0Z3D/9zIk
e5ur8Bbpr/1tbHWxtbZrhyDEeBazcvxOOpSLI3SVbs3VwAnGKdI52OKCp+sbu9y2KEHG9k7YH+ma
zhx2aG++zEA8cLiwnk0JQTCK72OBccw+bOk/f7tcUHPa3yiDrNLUHuw8joNh7s96Vz1fhJ+l7m5Y
eKn7qyvRC9fOZg/zgr+FG4C1XuSMruXxKp/rzaleRlAi/P4fIJxlHScd61SX241H4LSUAu2EzwBD
mar1OsDUhlXN6t5JPO1I9aApa6KjIe/JRd6hh1twmGzoQ5gntLgVyI2Jai8JM30eq+1x4f0GLIwt
DEisSMx6GLptO9nWjeMROevdv2tm/WF6hwFGGh4IIqblQwPyEhbCB6quYtqHEGESSAgwxlm1sRm0
zZFiUo7QzGVAQq4cbrBGaWYBFBlODcY6pDVpalMzoPLuYb4g/sHSf611fmzNAof7pvjA4EnbuWlI
s93+ToLz7Z2RWglCj1P7FKXQDcXQHO3C8qiReuqSBJnUqK5fwCgDkFmPxMlIfR+gs53H2BM59btW
v5FXhxC9LvDyEcYBFBHhOkDROLqPKgpv2L+iaGemaAvdWs08h0DQfBL0gmdKW1Y91NirD/gqUyLZ
gU9w6PgGOQbLYsSDXNu9/PwL324YGBfbVflGeCO6AOZfKSRs3peHLzF/U8o31QNNHVBSq0yKXPRh
sEIxaujcrbzJ+4Kyp5dIWJLie3UwJUf5RN9vy7JUZQyER7Id0nsECa+JHDDw16nq2d5F7a586XKv
hPM0IOsVFV0gcJVHiHxVPn/BtVYcFXcvvHYbNrU2tdo1gxmAg9g2HrS2kL6E1kfTli+xFl+tPzv9
pqwDDkfS5apNASd4IucDU8RL2ESBqK3ALsR8ohK+RrDwtgl2MPsV7lW1+HudczrrfsdQuZdYdoKD
jSEI5xvg0C96cAgwNO9ULqDkHrN7lOs7FUW2dHIf1UHWDJYoxvSTCSsv+3O56V5zsxJ59mrSVaH8
GUJbX5SHkTtFaYZyTfhvPsrD0LOMxPGlui9qKpBSEUTFL7qweLbvG5a/ll4asZCnEXHifqI0Xw7r
6FM+QNTBDBhMYgY8pHgrT9eMqZgra1LLWVmsjdwMSgVfxVFGTMnIFrxQHWRzMBR9LcpumFT9WmRT
txsYDhblq/BAe0+HobhjIrGcXSqb0C0AWSqZW/OQAzBQ+gNX4V+zLqPg5lBgbDrvCJASzFV0OeQV
z+kImDN/mpI91cEL8SZYz3gqF64iMjCXAGrvtyf4wQessC1zN6VgwYcEWwx0r1Jzt7Hq7v9rfgNc
Cyzw22Aj3rFT/2boqihUPO3FcogmAuWP3YuJkNdz3BfNoVEu+ZKnPDQ3+QfLT2Vau/NQaeJ78jml
sIH5T3mRC+qKOd8rm6wDDTaHgZz+ACU199KY8HTeHzYwNlE/q1l1FSVvULSSuiMiV1rggk42yYz4
I1i2yIZB2QdLqr8SRZdNNauY0j+DSHMnGRmmZDd1Tpxz5yA6F+kQqJmGRrQ1RAKRKCO/ketOAQa+
yAQnRijUgtANp4DyV5PqqFfzGRC9AcUqhmTmtEEBg+AZIk8pyAMD/XOdK7jQ4armIIg75atFyh5e
0rkHwVQJMJn68KAZ45FH04OnN27GM5ilczbA4aTxQGGNBf72XG1H05ikFRYXMkPBEpvE7oLhdw7C
M6ijGDdTmvIJzESE5QbbmfrEnwkGSxaL+LyeX1097IKZEjlmaQo7SGjmZkP94yUDpqP8ndnYEdEB
wlOXRmTrexhS1YAT5QRtRaq4GnQsAsL9vp75fuPok/4ILuKwdqxMOMShdYQtr0wp3jyUoNGSGI33
vYQ+Y2ZsNa0Bq6nuPfXFDYATOOaiKNHwf5CT7QHsWn9dtt2zJTQZYz8+OyoYIQp70mPRp9TqyloQ
3cMXlCxJ1wUh6e4wzCKV3ccA7VOY5zgjj6XX/j/kzGH7SOXkM/GRZBVlYG6XRw4UXYp5SGBo7O7g
rjxnEBECT4nzpVGVdloJJXckytheQh/IeEJLUTCc2FdRtkE2wQA8BJpWZ4BMpt8v6MQQNN84+9ds
YhxzjmD/XiMMsQkMezEuwG5CrDfcRVxxSWwoAbqenfH92NMQ9WCGr+6H05UOXwK9M+T+ObTZU5hh
tmcP54PBwVf0pcJx+fxWSnhBbRs4sy60dU5pAsmZQ4aafppEPPxQaQ6K25J2/at+ZCjkfETJ4DYo
uqxEu7Za3BkirPUWbxyOftLPdBnqksHxuMRJzgFwZLQfxbDGVlaGqqUhtNCPNEOgzdm81wz+CBj+
k/1oNaDiVmpk5QDY0vTFiva1vnO6bWSewSm18gGUBFgkTfNSPj5b51BfSQAKsyHy0WNBgmIT2uF+
CYG+GmWJoyIQPTxgd79WLB+31e5st9MO8ftpHLtMrjJ4X7cg3I+yKkMww/P02UO3SP3a9q/E1qyM
w90al2u1b1PE5hgl5B+NOc8iqoD2C+Y2PF0TEj7wYnH7VGTmYtTcxorJfWdBdr6A31MKEjSKeCOv
lc3lqdzMSH5aZMMly6aRwtL3ML2lL5exORPOTXTfQXhGIE1MXfjvlMojj6p94i6+Y28VdXEeXTDJ
yjj5DMSn1Bey8UxMTQvDEgG2rPuZYlo5a5xdZEXdJTkgu6QnnHcqon/evkXFIoW4L9lBt+0d6HYl
cyR6W8c8ighGoM1hH//AySj+LeDbnt89mujJnnh9apH6b0yT5T2zDzwfU5RFOQdWzsQr3XARnUZ1
IsBKKmZpsqKxLLVQlIoDxt19joPbYnYD9n+j6VF9d9vJ7pHii5oclH6IixDS0d50qwTVdTlKLklP
lFxAEZwQ4XS5ndeM61SNJspwxNV5nXlbIMWTf/7H3aYZmOrtsZVO9MDy2HruJCk95ILqkFInsIok
x8givVi/FoRH4hkDIj76N2kFUF5TfUsT2/OTE+Qnmunb9RnO/n9p5Uevsi5QlTCSmp9z/h4oZJ0R
2Vpk8HWpUITUIGeVIOIFvCkW69ONUAJeYrREsy+V7exAFT5sq9xubcf5J0cQwedGF4sADKy50cGH
cbGtR8B2UDA+6GK5X2i7J20SQgfW7ZfO6+2M/pRHj9QIXs1F94OtZyt7XWkVH6/VRrszwJ6b91ck
gkmxO+S3DTUIRV/AxsaDFrsxq3rx17+sZgzsq5eM0EvQmS5J7P6cQIxFbq7T4oJQNAiOCHY0B8wd
wNOZfUCtCqKXuKBWqH2jAYP5OVSECtPRTZ0o00YQfmf52gdf45dBalQ68M72cGBc2Hizc2xJxnFi
fkhUAd0rmx0UMVA29GQaB5w5Ojo3/JFmmOivHJHa3I+8tBdBGbu4qZPOKoLUEKcZkM/JcXkMbiYj
jwZer0HIMZgBpdaCyPcnKkDL5/5BGB04qZcUJKt98CSyMyQzfVBgP9xbiaPmtmlwSDCQuwN86saw
1dWPk6Mxmo5JDILzZ8ySaYJn8K5RpDWxwj+VqbYMYLN8YOkvayESO/jUReLB0zzy6c20DdN2z9Wy
pvvEg4gH63ePEjdNWhkut5FW4+hoO8TjN2XXhWMcnrWYuyvSGjMq+v9dfJn5EuEXaG0BNGM3tO/h
zXlQzZXWwKpE3DjBHSRRUGXKFsrdoNfvbQTldCNCAXKMYUvI/JorSzOLSNJSvxNXcqep4nVqu+xP
hlh3GZMuPMINOoRV7gQJo9ipeLy2i41pc39yr0bf7E0aMgAlt1l6Aa9SyWdWZ3JZ29dwks289aiq
j+UJE+BorGLWc7SQ8BsvYeUtZy6w0Y665/Oy21yX4+opWI7+EnoWfdcc179WoFGJ3x9PmPEfbY8V
TzGGk6SH65HHIu+YsBt7Iq2g39pSjLrYfDJOWqSwpE4BtPaz4jxYHAUtudYs8BFAfipnfdpjXmop
L4/oOpTcSVoPtujAsRsr5dI+nDMtBQgkRmBRhvMtcdVgynLASw33cY0dF6VZ77yL1dwFjN47xIW8
VrmWSAfvJERHIKN6gokBNrMJvM8EaqT4l6bS0P0mhTEhmcb02imkEgHKlhPR9NtTZrFPt4nmVEqB
vSFBjGVQt8Kf7UVS/qDRo1PuPOdCL5yIYQtswCuhaKN/KkKn1DUgD4k92sEApiUmamSxdgI5gWcx
ff4Ft6plEGxxnIOAj+biKd5yKYPV/+/ubK/DMNPqK8XbhOm2zUN7z4hL3BJB9ZMHcXQ40cWLx6mH
7Sq/Gz8yUC89gYhOviDOzA0/qcYhDKVlG7D1E9UKwJ8mJdPwr4MGw3sEPT3sqnmfZUtKQYDbFarq
Pt/45oW6hqrlFwdAtwHjNJQ454CXlKpGZGFv0pCugi55lVjGmCmYGhjChjmbVPMr7MCpP7Aj6WLg
0+DRSf+9Dx3eTe+QSjfHQE9RZyWMnHjcDCI6unnf+fGo1Riny599B0My/TriTRd0cEwv/PmcJln7
crwGA8u38H9dyMNbyliJlOSVa2XaiDsOU7k+rwYnUpBki54huarORl/xGo8UqcKozQ5zBAM2Os2s
M/5PNyaOPtv9Qwx3InsGULasqJKzjz991vlZZk8VSzSPw3aoNFWegKYIUfxwbv+gtkXuHOQbyIpW
iAZMKhUVD6NK5zjpqRRnzXf3d5yeruxGCqHPdUmHXEBkpYFS4Pe3BU+sKuRJWyUDfyln6Z+fX3ef
3TmJy+4GFu6j55qMs58m6sjCCagogmMEXd7HJjkggg5+ANGuW0GmpIUHRDJcLaQSzk8rEa8xKC48
VztR/UNw/HUYUqT9d8BQqmwYDjYWxOFpfRADSvINciNVaUEsP1cehCTfQZTdvGyWvESFbo4+oc/q
VJyZdik4sZUwjUn7Bu1///RvXRgxO6gWmiPYZUB88bp5LI8e+YvDrLsWpa56D6nBIrmCs6eNe7FF
QbzKaHa3pxsne9VnxFNBP5tE+WCa5jEdZbaFmPftj0wJoPUUKvFF2mtiYWXH3z8VrNI0Zdhd5hDL
CErsKeAAggztwVCIPjlsppk7cBIjAeqCtM1cwHyBtZ8cNXqM4jtPgJqgRXWisMfAtuEYnZ9fO7NI
9zEomo0jI5KCVVGn8AniM0/mNMB0U0/brYE+W/CzvO41qT1jxHX1GQFkUj4ZhjobzdPGuU8DIDIW
lK3E9FCcmBXfXL51dZzn+Pqm8TqAtDDpozX52JmspLmkqdSvgmii9PPQ9Uu2Jtns+3uRAXbplG5L
2fZ3igfHrm0eR7tWWGGbno/TVvAmrnHpP2cFksSsF8CyW8GkJkhi6I7DcYEB12o+snUWQMVKHhCt
z4JgwVAwI3ieUy46PFAi07RU2A5yZr8yFrZaZMaFOa7Mhjn2Lv1A5BLuF7kyWf/iaFtpQFefVqbz
bQfI1BtLN9EUjQNGr6b8TxMCEXygV6mMA6EQa8ORVvrD0WpeWd1gf1bGldDIo3rY+mZ8S2OOR3gb
mltIJgmnLjt278WyusPtFMq7tDeIXtAA+ZviXOW1Ev8Cu6KJ6ufm98gQNI2R0cRTh5AzfkERtGNG
9nnhKKS4qVKCMA7ZBoew2eDYVk2FzOjybgVVY4SLV2DuIwaIt6bX6nXhXRYz6PrNYnxX+KLs870N
LvWrI8lkTCqEv+5Qe992O6BC8xdS+QCj62ByFI6kA5iWl1cx66XKYPoYRb6vAe2jeNZajmYZ0UWH
4lOTu8C1Ie2vjCPOk8OjcViGD3WFVt423Z8iVP8Df+TpXm6eyIFVpDjvZ7e7TxghIRcGPL3hDdX8
Bhtp08yH43tjypCJwdr4dGBs/HqZs1HRHdEZ16jIL8pv+K4jJWQI/Ktcjqi6J+XEdYy8lp2Cor0S
a2NvIZGbv0jF//m8SzxzJHiYijaYelF0mhvj8hDQh3v88ss9qiZajBcnKuFYsU7BHk1EGDLs68FK
Vn+7tQqgNyRqwsJ7Z+Ia+/tCz375/YFogaiwKdHXWSKnzdqbpoWxU8o7Gl2M4xIPpc3wG6fletOf
mgNay1r2kiIEMq3AmUnfposKE0l7IITZvJS3K9JA7cZrvw3u+KUf7UXABzfuf9Fh8S2v9zSt20r9
PO5D3G0/1z0TipS3xuMVq6ztfsKF+3PRm4TXxLgjpem7IRMUIUBThNDq/BkjNLFDBlMvMIlJoNwI
0kbdD+yPVZIe4R3JOFzgToLDmSOZjZ1Y8vBZS3fF2U7fJtzc+cfUdf6qdGWl+3rXudYIVA3EARyU
OPY7G7S6xtVpxCXFWLlRfwPGrS/6ZcYuYmwC7vgZRSPtrWbx/v1V3KiYtsdSOjY2Z0v3bSg3F/3v
U5QP6NJAmg/FgzcnUB5QwoNZjb3KBNIx0SAcjLhrwzRsJiyCM5NpD2rpkZUNnrd+qODGAB272w4U
rnKBH0Wldgo9e5fSFPZIPu7ZJl8ZyrJWQ9rERpFW0vInUa1ipDCGlXp1JPxnEzpJnKmPO6QVbIZK
VcFoYIfW42ReunOVAbWbj/sgVmtBzuOjkkh+0z617UoIWd87kvsahnIHTNfqR3N3J1bZw6FbkVum
WSH0Y+eOILgcT98OCGP6Bm9W4gOCIsxJ7UUdjohDZ1ST4ozY7ArbJV814V+dGGjAm8Gc8iZeowIb
8+VmhgrS5OcfEOFr4oGBHTCX7la+7tvOY8CYPTYdLttwQwwO5HWQI8wKZPEO6PW2xoozwsKi3wvE
BFFUfsW0d9pips/HoF5cjpNHS8nP5s/z8I8ENPZsI3uNnKbrh6CuYS4h1Pt2BVTyY++1zmAYII2K
XWwUT5m8ACsgxe9OhcVfrDeQhNcjOgOZPByPj7MxrDyxuTr6IwSM/sRsNhX5I072+Uqp2v2ZsCU/
U+w8GTARmEslMO7/MaBJV9yYAkvrQufbHZ3227NTzCj8s4+PQOYVTM3xhCSoM/mhfXni5l1nyjO0
Mq8oltdEE5J3OTAlC2O3fxsZdwitA4ceG2kffFSceIqoxcVSowTr63YCVVnQBTjM7jD7C5ujfH8K
N8xd8606+jDAkITBFXaY2TKLh07AXJYAxjPEnlII4F/38+3Hc7XDDZ8M5kYdc1Hldso6ghYOSrfe
2AOkU9FpDIWWnIw/XL7QFUMzomhnZsTrV1EIxK/J0gkZ5WAtguT+L2/yYOALMQTieOS/No6wlwir
rfQ/EU1mKZOwnBuhihzsgbpnUKuScQpbzYwnjuFZzBOExRZT+1FCUS4h2vnjWbF1DW9W3JM1TOf+
D9QLvNX2q2zlOA0BOsFaho0yzXwPk1rKXXda9b5mdAwtn7hTTl6f874SD2ThMDUKQlhFTf6iyhhy
RtFyhr4Qk6S7IttvPsz2WuRGvwURO2lxSkfBlSjwmhIXUEin/dAeu2p9lqzWJj5z4xxHUkgaYn/6
FDFsM0Am0IjuSqhg5hlxt7IOh4yFztrx/ROAskNKAepThApK8kyZUz/zqcBzYkNJUcl3IsY1PnQI
AjBDwy6RmzxVXn7cmqXy/77a7noxHzMso2TidHXsb8P56PbLJeNHUiOPk+NU3pmRNMRdUNGJKML9
yt/cg53PpQTXAm3DyIlht7EtPSDQXNoKgyM7p3U7vVVSw6CaNb3lj/q90dKuE9kPjMT2gn6TinDQ
ZDDKjdTFMsv0Br6uNA1Yu18zlcPe1gUki/9454I6TS2CglagnA0Th590VpPef1hV8aeG/BR1sEOY
ZUCyA0sx7pxhvux6bKX5gne5JgnllHeLLSfjW+4IDpmhTjMhPJQGdT4PC1bWVDP3fAYv4bI6G5cs
Uteb0OWemjDCERJUdpUJqMoBVEV33O8CAPZsOTM4oLKXXyvOkh1nXzYkMHplBzkgOiAgp1+KIBhV
a7wUrd0p5jWKrF8jfqNavDfYMbBLEw5q3rWAGLLuP/acMHalCQ/Q7Qhv9rYBLdWY1XXZg8Ivg6kV
cNGjUh7SNcX3auAGdEhcq7FFb90s4k1grP20Zgbrr8z/QD7qd0aQHYQu2ae+EqVqsliRKJgk9vci
YYzpnN9IXj4kQPbiJFLTRF+LLnqV2zgxrGAEa8+sOdpxmt0FbwA8bLfoV5bXLFZzOG9vtJRsb+Jq
vLdi9rcskJoS8pHTkaFNpc2/NTPaWcYJmNWS9xMrk9TXB6+XS0qbHSe6ATwNCpHse3HnwkbFLoks
iQRGfjSSOjPDGECf/deXuWA60e+F5/TWOsEjRZkh56Aa9Z/FDD/fDkAc+azgUnl9x709rxvNib4t
ot4x+oRVyOPMKMqOHmnFmXxi6a8YDcjFrDfn31fVfvffuhepUvjScQJ4dPYZvzEDaTT+RAIt4GVv
dkqlcwvr12u47Xa9sQkuFI/aq/l6sb1ASrTM0nLK0vHKMG9xPGbqSNNm/hh/t/SYNB2865piIBGQ
HdfkSiMu+oikoZWZXFo10jtJCE5UgosL6U09BtgHIqmmhKyjYKyWnq2ssgs7E6RiIQjxOkvyrI7V
ZGnAgWg+hyn+dpU3Pm77TsXJfC1F0E2N3adSb2xRMnsjMwchJm8Hh7mplRaSRmTenEQTeihH0lRH
Qj3t3beO4RF7sMeK0beUCQjI7MUqIDRAAmITLPxXsnuZIqXqbbAdcLeZepRh/cGVEix1K4wbrc1f
TjUnIz0uhXmw0VPA31p4CRb0FbKGxNQxkfa4kv2/ToOYoP+ipHkm9wGjlYYvvlXKpvU9ZaRDR/Z8
iEYw2+3Jtpcm3RrWShA0Hsj17hrwWrQHyKaNoMiPQPs9j+6mrwRey6VOXmDNmbhyachnQcXCRbMY
CJgN2u41VAhwx59pMxCTpp6Fmn3WGnWzhKs4n1q3LfvCxhiURzhQ2M6g5rlZk8touowPINYtdPoi
RBIRIDEep7oVfuHFyLFlsTd8deHdndnYjjvmZ/3VE8bf8XPGwCYxOxCDcVhEujdDTMg6/Veuf5YE
qYPvFhBQcVHXmjyboe5FToRVcPA0nGxaLEQoDZtQWWHnC8dmXQvM/BJFMR1K3bFhIfZRUf6WTRPG
KR4lEzDUxPjtUQl7yGmEwEWWil4GNJOmtDs+UNspB7cwiWSTlneeZmZPIxmqmO8V88b0s8+4sg7k
jIMkGWGWHnsVvx0X+BRh9ztoZJayaOWpBshpwxbj4gtvL5P5E33HokMj7qqTkgrKAbuhbrbA5PL2
5Xu/iILlZ51GhCO3eAPL0xsycSa5cymhF+ym8yEjdtXemzcbN6HGqjzJS55JO1u9WjnvpyCmY6dV
UC8STjAPCPL96Q6FfZMNjZ3QaGpb/XKs77MIFlz+95ROT1sJQXRnFGulW+lTqNq/RNnr8RZ1Mtl1
rhlj1lFaDuyyTuFY5z7jRu5zGWfor2DrHl+U/vPNSdrIj/15GumE41BTYs9ssK0D6zJdqPxum4hq
cfCp/PeU9SggH6/4A5sIf8T6eS5LBXqgmWiRCB2HUAZ7rBSU31oCvLgGJrXh2FJEHjpb+gBo4ivV
R1gAbEqFh7S7wVIORl6ENw6hkPKdz6ULS3qIKvoz9tr9TdOnPzVclaXuFQ8KNUR7C+NGOAJM6rcK
Lote1dLCsVzvr1APHz7TauvIQFCW+iPrQIY1Jors1sPJKe+GqWEuMc3HbTcn/DHIu2Gq/pkGFsC5
76GI48b2bOMP83MkKEz9RjX4pXxE5C72fthbw81HXUHkg7qxHFLnr4wOnwFvjej2zEvZGDqJEa85
JGyqtZ17Q/1UM7jhvibRyOcqm15CktD/XaRhpG2/zJGIb9GtroU4v0xmLeAGLFN62zHU/qvsMFX0
T28v1pXn9dQMQlC0Z+W+wv8VCcV6oPAt/NflX5k7McQ7Rs6AjHdlWH9LFhbrqGfJg6b5iEBDds4S
+Nnaeh3YTKdvoQe4teDBDIrHEGjKylmLYs+7Z9/NYtORcqw3yyJDZAYFYR8NfKcvfZjxm6iJE5lH
Q+kCItsLpE80HKBY+YMG1EWnbUAURN6MG6EUDlzf54XOdf002tYBvDMqLG762oiKBg+SoKppYwUJ
D1eWOkeMxBPBfXuVSBi75corZLuxaRZyCb+EDZTBx8RPl5GaNhJvk6+yRskJZOgCCSFOEl1ek/YV
KSqLEqT8Z3luf59eybdm42wsUXgFCQxCav+irP4DieXNfWXtuz+b2qCDDywr0AdOWXw8dS9cnurF
Od95vSlPNFCUHEud/KSlde1zScspRi41XJ8Z5lKtsJQpIBMGCYNnPBxioJoAwFDquscH6nMCFrXi
q8tJIefrWB+Re2tZh11kaefB4nI08Zv5GM89BcNaIngPsxX0+gEV12qS2ndlwu3zOHq5TDCvuJyc
l6zXc03b5GZ695zzqbmS0gUwDBOoCb2+dtfbUPZSK0noIHQ6tZ53BM8fbI4ebDUV1MFrluSGMOWE
7rJ57WYH3EIzzEUHNMhidnWE1ugMiSayr8vH5cydyT16FzluVvvllHmwDl+uVMn3tN9/2+7o/iW2
Vz+9MUHmLI2fpkhHrwl36nSiFd8MtkMeDCk0o26VflWzJqyMEAHTunAf0lGJFDkFStmQ+KWCFu9U
KUym3ioe3svBF9MitUjj2enIH7ZsAivZ7ob//D6v+0pwiNSO0mE4It25whZf3O5U9R05UrEyobc7
kvYRku6Cs+9tAZZTSqDqq1PXznkvmU4CbgjH89epF1brafqmh93Qf+tMmm7DM45lSpgu5LaP1AxW
teLN0HlQyuEaTUei9CHYo9f1ZXWY3KWwzoZE/hs4I7/9YALBge5+vfszidWgGC4c4VjhXxE5Dl28
+9B9TyhkWmQNkuzjjyF5rpWfV3LC+LQxEcHKOBShZ+LpOIV1Ao+VJtpyopWFOUJKqkjyFfL7zG6+
nD61Xr90UStqHvDOMSdpBGWBvq9pNfGtb3cHsKFIFPVNO6Uud5a9UjbzzuP+pbJbWl0QaiWqD7Wr
pOusYpgQnNkE1PAwWc9ucLwftU4G3JPPyWWQ3OfHBmgn9JCNRsXq5EtbHrk6HB7XhN53xonC3p1d
joVVLhwxsb5kzm/xnVV5YyRNBqfy8ts8ht8DBzMdkUGo/O1BRHBKtQNvfy0MTTYmli/13ys/hNGz
En1JREog8zU1kNRC0GZ3Uz8XWidyYvMUNrUH83cgSFemPkVgI2L4ZzUQZaSauKKlxPb5BDHGG8zP
D029Jii8zp+WxPT/PLjBadmYMZJyApCrzcTk73ErcB/cJJkx0qNQ1eIWnpWq5Pa+lm+EzzxMO6BF
M5U7/kdOdBIV6TKwmystx5kJqOdoBpjzXujNb50nhylB76jHjdZghMrqCq9QMjBhMKA5vlLgYaYS
SbqxDYxkMayIw4QSE8ehJUDPT6XBFDANzzOneASnIWYJCW//l+HXY70VOF/0CalrymLf7L36yYOl
oUC5Ipy+gpkyQmKsw88mJLcT6TdvYLHXV4kWeJ2LlQCymRhPw0LXFp8dfxcBloCoxCiq1G9ffl8Z
P0Ojfl/6mNwg7/4DwHFzWuOqM9lRf8CAwNkiwSYLNRdWa7lQ12JJITJJZewE366s2MFRPAgEBk4f
m/SfCRCApRpe7iSM0GigWRQez27q8ynpRu9MGqvopJ3FP81/a9+FRzIWZ1T30P+2tpdHP4TB4mbT
9kJo4e3acFwam4k0MY+XZHp1dnX83LG2ElM8iMiybBmupJoFpIhajXw1X+rTSLMWA7Pvaxyqgugw
D+W05SsaO5gtxW7kJfhiU+f2Dh3jX5uNtroD40Z4C8GoC0DuPyFz9NyYkM27f/aely9LB0LWkMpH
2Ik+D5IEllsvBKHhybCehmW79hWXpfJ3bfZNIXVVZY+Byk5rR/B+iA1BV/QRe9IqQTyzfQMNgU4L
aJ+vYpkzVSM6q9h7l66l2x07p39Ip37dKQ7+lgjImqgQt7RLrTxdRWKD4eY1d7z1M22dZve9Cwno
4d5OZgOUjGUVKO2LnaSwaQOUxAgcpiQz2rWS2s3lVOH4zDwlw9QNurc8lP7Gh7QnLiI9YToeWPCg
00j9VVhqV+H/8z7+nGlBT6n+9DOBnxUN/P7TBBwYvdKzceq418SU6h/qiVf8ZwJRoQZqoqWalWEC
DP58pp6HdzsIc6cCHz4dT++TFipG0GAP3hccNaqhVgEVab8UaJrzWAhc0auTubFER8RdZ6HXxMKU
G2yeTThMvT8Qf/P/6mijEPEcOFRZyvHsqifIgE+CRxpt9imDGbGPPy9vpNCZop+HrV0Dk1A1rltA
QXfiUBvrfWDBUXT+g7jI5YEg0QIVHsfLFVqkwmIagmUASGmvjbEfA1Tnlr2wsVUH6WYjdp014amm
bPP3Wkf2qA1J7zkuh1HTns9JttpUJXfedGTTUZdB24onwBhVcSNkC1RIYvau5FQMriVlfnrTUgGo
2IzXeZCeu4x1+ts5zyZKch8jntoQ9IcVi2siLffvTVgnZKjUEzZbGltwzfDx5AajTqiwM7Foctua
YdcNJd4A6lnc3Khqf25O0ppV01ggchzrvTCxRXj6NQdqzjOMSGTV2yNKSgvC4QmoM0YiQE2NollQ
FytekxN0DBu5BR1VXridgSls+AKFQud9iz0WeoAX20ajH18YR5DCqAcT+MsygaJXthlLz8R6Mrb9
kignilvJNAiSfzfYA3sj1gGkQIrSL4AtSwGHi0k/6G49v8s3vv1xJLtRTTujkgszfrXW970FxpTT
6gEEoMVr/rgR6aTtuoB2IFwnWV6W2LlwU9KgYngyYA4tTj8jblyCFl9qin9lxjIqmGoNWhX2cVbT
q190Ws21gMT4KmAY6ZLL8KybuhMIVoMrSuAv/oruImQ/2wLQ5+fXEkItCw9jJPfgX3NVZcvEj68D
0AL2E+CZtvwiUDabrKCPDMVgLoyxGpRZLu4z/dyoz3V0nOzexNePtljdqTGUyLFo/FeZz3QrTFh4
S9Y/ekUT0XHEx3/qJzt/JMOpqydj9JJlY3q79drtlHtsaKtroTg9x1ZsMr9N+OvdtWWA0e256a7i
nsIXjUQaej3+zY0yySf2Hqm+K4V5MNIVKONwwCS0AWhyW8xkLZwKG1IPxRm7mbLkP6W7q8iOE+OQ
P/ScMVu8BLi6R3nrkiuUpkPKNhJXjbxcMKabFJNpE9zCPsr1cqfHbWOtpzE4MnoiTHcNuyGZl0cU
FSpXk3lBGHIcX7ekHPAKrCzQowC+9LrWIFCpOy2nXqanichwAWpchCW4Q8Wmk3t2LmWrlD0SeIzm
HJ0S42YOnADVy+yA7QIkt/SG9XGyzly7R4C0GBmXmP7638VitfoC7pZbKHxEbTO2XwGrcg7uHOxL
HLB/MqSAQ/yAli4BfyffpZukNF010ryxcSxJC7T50awvgBo9mU0EpN3dj2JThZo5KLB+rovcbw0M
BR4fFTzrjEjWfV2b/w8rkV4PJo9563gU4cRU08vG+wkPzK2yP2GO4irMRtkTLCW3Xz06eKR2NvKy
zBJTPpEoD2jToTJZDC/8bCjBnqPir1Z1Kq2F2AZBr6NqVFyoujVxUwsfZWIwt98KY1FF9OiYslL1
cwMaDa7DtbMnYgIxXiphKJs8hdR2/o1mr5NNb4sLq/sLPx/WO78Azx67EpwIdlPEtXold6E+jbs5
2HrN1OyPNaoJcBXEhz/rfPsuErTikoYQm8gZ3UvPawy2IjYCxjdNzr+wcWYGXT601y2JQlAxlRyp
oAMQ6AQOq99RQ65SKHm3IASaAtx8L4s8+GhrTcWZvEQtq68UdR2KHczXM7NYH/nGhe+WZZ6FOVZ9
3BezG5VNG1uHR5V2Kqf62OdNWE1MkH10I8yI5OTABphoUWkLNAPc+zGcvF2u9OpJkvauKsIK1fy7
P2mDJ7XbpkD9z45IUIOZ+67qyFdH48IUJXUNEiRcQlqy/69LAZmXnKl607AjitNZAnaTaZt5wxhr
futa8KAsfp/vdD74BWHqYEMWtFlcEtSY5v0QfrmQEvCAahd+97W40XgUiQkJ1ZHxy2ShyEJPESgc
4gqJU8byUZZwTjnyoQxLjcBkUYrPJ9sEv+gWvvd2JhZsKgqVKtMBAg1/JR6HPUJ5A6VqRUQ47Esj
uALKJcWEdJZfuaHX5gZNcY9uoxxxriDD1/khyTtILzIzB+ofhpkRQ1sUyC0IwMBLeO7DfivR0Oq+
lBcbZSKo5k/16bFj/nYlIfaBIgIZA7t4aXcHKFQc0xhJARpsDmjSRagJmiaeNlUHafp7FWfhx86C
W5aTOPPjLCM86Mp6JrbjX975nZqw/m3AlNAIhAVtZcB3j93FhYOQ6TWOpXYBPasfSW8Zcduw/UiO
cjQPDKoeqMggQx4JAO6XNBZGAAi7e5jcS5ajO6axm2iuC33NL62JyAcMps4X06NobEfkEMEAf7bg
lkTvZBlf9Cri8M8bZr+iv1hFNAydTceqnGgov294vttwj+bJlAVH9X7EaL/XJOg03QD+kOXRxMM8
YKNDLBDo+MtwU3+SX8SshroQSET3D16iNXQY9N6cXUp30SruSxg9HqpBXOj0er8FsVXiyqw/i1/7
0foZfgApStJ+W/sAvfQDIV3HC6DZ3l0sJGyM1QkFx//FvV3Sdp5RPRaa3TSzWlCJHdvoJv9bR943
tR+qEDrRQR8GHHhNFZpiMqOMuGCYBm2/39S0l70eh/nNrU8ucDVWxX+fn2vq7jbDSss0oSvdAJZV
TP4EAEyT/ljtxWbb6Wye1PraXwOGhPxhNjC1xxDXPVDLxeFPdphfsFe7QhkhfzwCVodhDnzQN3/q
qiIero+thuA2s7rqCDPnTKcAh+e2j9s/e03V7Ecx6+OYSHRQY+X+d7sAOS0fy8XU2KAKwciPfG6N
2X5rgsvGDDF0UtN8po9BhCN1Tch+uYlYwPviSk0OLw8b0rlPYqg3ZgfEwE9FmmqSRe+bSC7zodjU
lqdI6QzvwiO8JhfbZZ8Te1PTzvv8IJkQuyeJXEfFAYCs8h7sgmxy83T+FE8SeL7EqqUsPExfES/l
aoW5BTaYBc+CBxCOSXa/CE1XW6LQd3sjd18BjbLjnT/o8EL8/I4FxPw1V0ZhpqjKdZtK4fYl4AFK
BHuFp89M5YOjlI6qXZ1D2+xmDKjw46vAmZmOcvpZ6xql7KtOfc6MpZv6HBU9pdKxvgl3sNjkHYRS
piXHkOjmSNE/j2cBCOBOEZ99xQ23zwuYqIWTrxm+dnM7eQIMXj2k4NgwetwfFdWfpL2i3RxzuRBq
Fs+sKsTvuxlohmez9hk8fyIh/gJ2bHh/uPjWcffex8ten3m3FzMxWCSAnZI6RhjBG0BI113up4Wr
hIcjmCiCKfu6tCBL8kS0rSpum4k536NleWoWea1/Nunp5pibBPwPT4W3RGLLbyInKVf8jVooahBf
4ir/WzIpze4niCI2OqhhG4+jwzGISTucraIRRiJ2l6uisXsLFY4Z0ywbpxXpuZS5wk5JpIAFXv0R
4paYv48aRWd0j9iP/tcWhxonay5Rac70a3si0Oi8pEnKmywfzP5WvK9nsOWKDLwYLpVEGJpI5gxQ
F1PUcsFFNLrHivVshpRQMHeWaNulyn9/3k4pG+ySdntDBfLqcvRmWtnG5s4tyWbJun58vheAxyru
QMet5vjZO/DXLIqIAJLMzUTH44kawKrtgrbyJM4WNwFd7VEFffS/KEDQ+qPBFRgHkTLSqurfEM1M
SXmy66W2aHmtR0IijzRKT3EcfijrGrU7yTJIDkjo3F81zg8EepuDMeBPEl/Y0fzaX3+4xoZvm0Yo
no2l0EUkPoCWsnSww/70jdj6blVwT7hPgWF2njB6n211cpf4cTYOm5oSabj03RsrqoBUmBi3kd6L
m0ayciDNh8KjvhgD9EePCE7C2Gpk6/qDl6fYJ2YXNoiUTeWKx6XqVJg7ufhNrkDdtq02ev16eY+6
fW2ucapK/KahbehIB5/AOjwH6Ug3g4Z+tubQiPu9V24w31QTHcGnGd/UUt6AsxBWTr63WACQszAT
xJWEkwe0kOb6FfnisraHJfHT4SkPT+OwdPqAIYHenusliGSNCX0xOBVD+zTQb8kL6T9Z+Jo330YI
UU8TSbnkXu9NJ6G9uMGIJStukXjy7pIzUKgkYKfruuJldmQrRtCnUwYyIME+klkIPuKMtUvLyS57
8t1pJpBL6EhLRyPg/er2wtehoBcpF+naM5RiO1OPHXacwEv1E4tCGnDo2360o0k4KyhZcfzNRLRw
q4USzbZSwBxoe4nFEqNOHWIm6SWHVEYfMQpxAIdqwwj4y6y0KIAIRIAgEiWc619k2plZ8UtksRGu
pSEYU+vr6E2HntjrTa3HmvSpvy3oc4G6g0mkYdtjboIgE8OUTCq0H+VJPYLrUKqXq36fqV5kUZ5W
7F05k51IvDWpkpnSguFHBoXTEq08nMW17i7R92YXgNxtOp5ZtSln4crif6Ewrq8OH8zsTSBxhc3r
7Y56fSubrOt7RluUlQpDb8aTTxhg+y2iiwwN0qVWQL1mB5Hia8YfiYUA8XXEctWM957OOte4g+GK
Ati62eslR3MWQ1vGSdIC18MNr3ux3QNXH54rZ5pnc1CjwHhESNMAH0nv3qVyWNNZAGdND8j4di9l
FjmUOZQUaJ9T+9LNlMMGZL+Yb1uPOuFheWbjLwGBCboNSZcH8r1vshh6FzOcc6LngjO+AcPAB/g7
1SLfL/4MgfVOIXAGmSjhIVhTK0mtxjoNEBkh9QNBN4Iy1HAT93gAxaMRN3ecxQ8YskIGfxkuFmkz
HRwOdLHR7RPtl58HBUFGWFms3JY1205bR95CZVxQ2Vbs/gty0s7UkNBm0+wX641oyTqNOob49Zga
vCvHKPneflDfkbzZlg6iac9ft1uSQxPYfyzldh62Q07WqIiY/MpV3WbhXJsvQdMXiF26pwqDZcxV
3Up+knd2FIUzHAfzaucOizUqCj68lzsVYSIKwvBfqD+DPS2qSJ6UrkgS3s93u9+Wl1qIsPasLh3Y
fpGW4g2KdSTQXqt9raMAA6KqlL8b2o/e/VPbzu9xrpC8p7A9iebzSa7gg+je8b1mfeFcOOwsIXTC
2vjEYR548B846HqY6STAZ3s+oGdvRwYlV+7UY++h8hTNCyB9Wl8O+GbzjaVwUsXWucx4DDuw4jX8
vpXkg6omnwCg7fXNzZFKHMxOPndRng1GJlmR9oPCl7va5AqFvKAN5hgf5kZXOfhcaM7O7GH8NVDf
MIvQxxWsCM5td5f6oYSA+sBQX+eZJjXtXa9plcrbFxD+dekONJlW7pE1Zsed27x/Dkd4svvIeES3
99vljnQ7JqNffE4Cw1KR80EqyYZZWFOmPOB997IYXOKd4OijepRl/7QagPaTn75GmkrantZdXhxs
iHAjbWnKutub9yEHWHN5OzGpbhNN63WJ8pfRBj49OdRVN2MveHKOgMjowhazx/0WqCco8SkJWVgs
ekj70TnGrvVNu4GO65QCVpa7fZrsWoLOTDCO7hZIjbu4u9KoudiZbb0OIM/vOIE/C8bm9X/HfanW
BS4xlmYfDHfbZcsy48s2Hdw5Hvfe+MEL+nXY9TnMUDEXPhvwBWEHkIHE5IvQSKN0pC9q8GDGxbAt
WB0lja+r/i5kdJzIy99A2PAO6bdcWoA/mNEovoH6+P55QltNMXaNtPWX0FTtP7Csu74z+e0rin+J
qaZTki9UvK8MEJnh+W4aP4tQeh61vr6H5KWKgMrYYla2KrEtZgH0HL+Zf8ej5y3x0QBupUBCatD9
5xkx7c3WZl1/sptaGO0FOYcEljxdIHdkUVab1tou6OmcI5Z+LOeE61aXnqZRUFNWw+H9NCwPpOSg
uZ7GRrpIrnAMuAXI45J8hvdNefpTIEqHjLU3sDbQQHssTMqB3T42Wm4bDFYCE9YaRLxraKBsHlqx
Obl/Mr6uqTJzUTniJFMLliQEdEu7MbQf66E3HF7qV9FYrZeeIJv35tstTab07eWFKwTl/qDHx9U6
iWAJv9jPwdJ/Zz76ANWD11WPBQiRwV5WLCWPL0rEhQNP9Rv9tKvUGeJRhr+Heog0IqPO6z6r/qGi
99fR2xE2zmReZeD8UyRbBs8CnDCEFrWF0er95J/LPeuhNLzbDfT+WjIoeBZiNU3puU/yuzdEcGXL
pHop1KLrvMmbfyuu1KPKRu1fqCGdOgeo7v1JGEg/Wv7B1Wk6rcBx9kO1xsJgnYoIaysdnD+DMTBS
UIDi6jkIlD5qMMYqcPmw350elWDobB0UXcEig6oxvm48kSaDLuUlekAa79sqj2xwRMNGXTuQhTPO
0Ho3k9q1OG9AgxUp8m2kg9jnL+Q1WFB5qOKaI565ARAE/bTe7sTyd168Y17dckEww/i42m60sMEE
/BAQEryDw5XDJhHcDMptZJcYXJbRHKrnfkAPgT/pNInnX9Z94hEeuxOogtWDLSXwnYWfyKgSxZPk
Zi+qeHxxsowLdrKNr9nCBp6zGUNnlqhzOlZeycW/UaehWuSWJEkJJoQJ1fcxTeLoGklPnEHt5PXC
i9x+beF01xm8DuFMZ2JpynrZkjQ+mh85EkhBIAPcuhEUzLWwfbhp9Wc0k31Y1EACGKYcztJY4kqQ
A817bPGJLLxzsgpCMpat3YNyz7h4vdMeI18U/KvHmL9IPPGvAs9NTChArKIzlg3Ep+cMlgBkJPgR
NvJZQaFAjltcBSHBvmUp/yJuGbLdkmU7eout9RGrenX97lJMahY0cQ5GiI49h132Zs2j+1m+G0Ht
NITisFlKh79/YB48/pvYirxpnw3z78gwD9d8i+rbfuJwv47v8t/hdst9OxiV2iOirMsAgmQK1dZR
AE8dRNIGBpwPjjZkOlJyg79ZhammyfSd5G4AVjr5RcbjrRu4VkBUKKFRqrm5Tzgo7bCCHYJ+WNdx
c/I/w7J7tJQXDt36lQRj8Xen77d42ot+cEKpa06o4Mr3jUlRj+dK6cq6Za6/0MKXvETzZhFYk7rv
gyq47sOUbJbjo5ripyFZ1FAuqlW2Rt3BTgr1fX4oJWsJ2+VEFQDb8HMfJRE6LR4ao0jRjBMnsa1G
Jt+IwRfTGaNchctqsrO2lhTMJ4MOPBReLgEyytoVTDX1f7QeCFbV/qtk5iW7fM4MtaRekL/fei1K
CYWyiWQXkFOIvXpYcPCgu60LrewdraKIlygxEtNUkvp3v3ZPdpme4vcy5r55/alm5nT93gbV8PNK
UU9IlwqHKjXyhy3L03XGiGorGrmT1+kN3fzJrT1HG+5mKFPDbe5gn/n9Fzb5enPUOJOfto/yTzWz
IIRJFxRtjLmiLIwsXG02CFxO3GkoxmYw8fW7xDaPX8OAbjmn9xdlCpbOvqfe/xS4FU8UbFa6BKyV
3xudvF8eGJLiB/LlpCp+sSwlbTzIS+oG+D5NRI5AATd7FQSdvAI6ehiyxXYejTH9FMGLOWXISf1I
NmVgMMwFa14zA4xdr03adhcLSdh8ChqPnYG1Za6ceID/0hj2BCW1+hhy9MsVv/dnH8kJUUkBySjw
GK970zv+Rf+2gejO8dgiSFq+QX787PgJQmrY1EcLW1ZaqAyIiBfflbBxr0wcjPSVyiahA3bUuM0q
AiFicLMRlhWDmA/nU+NKbiwRo57rw+5t7oR5+uzd9skiyrR8rtzkCZTUQMuswSxKTXG/iY9On2GY
iwlHyd69s/N0OGg+hFls0HxvjVVOSEbnBkcZL4Qn9Gz01NAO9J+nnflNdGyPXkGt90Zr7kFzfQQ8
8h+0fMOWDVF3IxEtnvrQ8GA/jnl/1hD0y8CnlC3Ts/X5kauxfGndBoucv1nuiFIuQqK9+1Bvu/ZT
xVR6GOiV7uCvVsz4AV+/j1tiVqBPGGgUGncod6zZchWrbvFix1V9vutqypBEfFYYGGE9kydXi4hL
dpzscDXQhY9UEshi7J4bk3Cr+VxqhfKuv2oRpz6GiFqmi2cbQ5dKGnP7/M4P+qkNAnIE9vC/7OCs
X6vHYK7gichpIlAivIeQecf/dL/vIqjvk2wVW0H5IgrKojMqgLlFhcOD8uWDsNWlS4aPUd7RJgZa
rvKHDdZLMvifigLm5o98MmNxrGywECLWMBGiNGiY3YXE7O+EJ8DZ5m6zv3BCXYzpfdxyaMTx72lL
YQIfnnpgs6K7ZGeUa+y7wnrYPpoV9mzsZ3XbaFpPcS10IR7LitZVrTDCY+QZaz0PokNl43MKyCx5
guAPBrO2m1CXq5zLiGsnE32rtNmf+42L0k2ZWzBknw2qADw5OLoL10TqEuyTDr/zEOag5XBrBJSO
R+00wl1kexVXdMkQfupqe3ROWte6jblFn5Rs3Nbc76eFigRdo7D7K2dkRCg9XntAfKSZqAL1f5nK
7VWd+NAtosWy3cDSKU8vAhTAZKJjt/CW4WqcfRRqTubOxa/c7eXtk0qQEhUuYyuo22JVvacWpZ+p
D7+gvgQMzGj0jUJ/t0cd6mC7/dumx28axg0svopCcLLplT5o9rQgpU5IqDhkR0cNdoRxydMRjq7T
Dqr+CxdbTyF+pJJhFHbFLIVmyz3NZQOG+Ds8vN152fIZesz54CG+CTPLXPg1QT2OFNICUxH3WOzx
N9xH9RvRKvFT8Q81j98uZajM/+Qr6uKcC2dhnGVMtFCGsAFB8n8EoKdgEK3sCRmLx8rkuRskw6BJ
tPwbUH18SfZXw02BzpbX1Y1yewq2yN9f2RANKYOInzuVpWU/00dxgW29Rbrf9dHM1VnazsQueZD3
bORX4B4Eqbynnd8VFO4Kt85wK7LhAXG2L68IBOA2p0cORSUhpeS/bL2fV1Ulr8Dk3EoKJ9N4uBwe
KNibjhbN38Yws+BpLRsf8K5VDuXOynGm12BwX6rfZZJ7Q96IWH15nr1Y08lRSZobv100LO0E5q1t
k/77aStdZands3quSoRLz1eJBnbgWNfb1DmLxuJgXWZ0ab30E3I8UsGP4i7biS5WmQ4wBJr3r4iC
MgHramWxP58t95VWWyqEn8zJ68rAeF31NPAC2PGmx0suyf7bIF/wSTJCrVdBWddjcw2p5szrLevA
cpsckXfSNmJ+dcH8sBS35M5kzP7aMXFl3XuYEae5J0wzDO99TrWoGU9FJO4hkttvplCDPOkLTppK
AnGV+Tn9zmBhUcNSbUeDbioyHP4UceL8JmI/2jNLZhBFHLkgM6HfNQDuL4oP5cL1vi3dk+wmFh5x
hvOupnpOFakb9Udqf8RZBR0MAVauoVdKe6+ZG8Tt+Pt23/p1CNJiH9Uvy3cU7YNPwcLOhTP5pJ1m
gGIZIwN69hP928FlWBG8iraxiDOEtxYY2Y5rzF/8bY5QwdzcUHnqRIo9+zKjgcPPivHd3ZYoPX02
U/fNjMOgN3yYn5ZMI6Uj+ZrLh+N4Pat9kPoaJMqcnB5VA4dt+vb8/CuHLFyvAfu41knx6aNvGdl3
Awc/m4aERGAq9VzfjBY24gSCUposus2ofCCZciuuKU/O5RtaNNUoy2ng6glFJvH0v5npRTJPizEx
8SRrBPwd8BYusKhT9nsLSwFs/BfN/FmGb50o2yrVoFcCkhtbYpRcpPON64d5T/3lGcQIFQYlxGMD
KGAxbVspOKmJhdcKp8lVal8eSW5LMbWlrIS3u6xfEvwbjdJ4cOok4MRoxSsE8bft86wWfJ3JdbwI
UCsOwrdwXz0krAlJn7ywSPDNCI/uFy3El/iKuWPHI+ero9QOwySe6ErDB2V/r3240Cc2BoyKBtN9
uhKYfNdVVAjKiUTpAHOYJjxF+U5TSRvO8lksc+Qzd2ua3rSrgQH5YrSM2n2WGlzkERhFRdLRx9pQ
EUirYIPoxp89lKmYzNmGGmj0l2hR39YME8IuQTxOylIqZWOEtGYTuU//MxsB15sFtHB3bL5gjYMv
oK1NQ7Z4dwTibUikJ9QeUz3H5tMFN1bn2gzMivOhteNBs7X5s6O7s5xhYqqHJCKsgo9Shk3N1GUj
NJP/RMTqxfbpy0L9rC+uGB4b+ruwPX/u1pItbGgVw6ZsAzLPfkmmrx0dLqS1NfZ49pN+OMAJfHGe
QHwowSseLc5U5D9tNsdWsKLutVpDWZFe0S59PJgPY9X8rfp56eqD45v5nX8x4jADHU2G/VgaU5JG
n2q2Rs7Up9AsYVNPJAYDWJcfsWTlMuafiYzMvJSZ6nn1qt3yO3dldhpnB1JMg5g0h8LCfk8qYNLU
zUqwDKVtKxMjPGrJa6Bvs8L3LKZqfmn7dtTZPcfdjmXnCfiz7jjzCZ4E7Fpnt8yxWNVx9tExTfsN
JuQCmc9HCulG5W87vUGbFOGOmH8wpPZza5PZ2s7+zSn2bxwNoMYnNVJf2JmxqiQQyPNTIyG2aSTc
6DkTmIHlDOwdPJur7NSVQwttYK5p/uhuVglDuFMy+usjqvD4VIuQUpgm8YkHG0nY5qcmRAsM2R4h
8XZUFL/bG/MY1mz79WORw8GvhdR0m0YJJl1JPduD/p/Re1YhkmOOqFco/8z2F/tt7T0tOE3ctfK1
DqdsZ2oBey0ZJuNoSorPs8LOxsd50ru13jgx62NrBK4cc81g8VJfkp4so6+lfK38QFy+ohPXkfX3
ccOAJn+JEJRnWJRZKZKvp+puZpx7H8aq1iWL3mVjBcSMztGeWoVg1AvrQ9/eSVx3ejAtl3sCN3d+
+BBZjLrWY/GPhniB01xgUxaT/LL4BpDPKF0Itv1JdpPrY/3lq+aA+aGo9pMNrlfRmgy/0iBDfFQK
2lqOB324dk1y1EfgL82yVfIxoG9gXsrdHra3KTI5cH23P0QUULZ9WCAAZh6RbLPzZRtB1AzpUkXx
M+6bAMHg1VSg33cFaxss0jnSnY/f19zSkewNKMMer8YnXWl4mONo060ROY08n9EBAf3ecINq1KX0
aIjDyS+bjXtspIJuL424LUuCzzIghHTlSr+0n9p0obOt8mplN4ZT0xJfM9mDJcCR72TL0YSGtrEi
oCz0va7mk2KPMv0ZD827bZ+G92p/K/x7Dil29NOhMZOE7IubQ8jtv+yy4t17LupjFrdKuozpInxI
5544eYgvApcZJ7E/3kJVW6enWZt+B8cJ9cS/qT04G480rcsOKx8jZdQJymDgcrB2qLEWhbEs7s+m
ToZbqzuqMMc9g3a+H07ZC81gGi7xknLVKv1XRSpIrP5DGaLEUFjVV5+S5MO+6cfByKiqIrnNnycd
peZZx6VjvY7sq3cZMTXFdJZxpWmekoCFFgfNmbRTZ3dlZLn6CKUHnq3OIfpVVmG1VezPwiqHAK13
XThRzkCyt/VzzSQNhEzCf6ttHl/Ox6ZPeuI/w8FbWJAUDY+hLj1lhoypPPvkUZ7vUuGC43+0FLcD
/JYdx2reinPCNVp7PiCoUQV+og7I484IYREEe0+lrKL0lkEizbw7rhfBd1LeEMD+a2FfYl96OsRa
lj4aCmalhebx9q/1pVvdgcwSbwPj2j/PYEskgWIQvTDT+r1vBtH+kbjaaV2v1QD4idF1wjVvmc3e
7BQx1ORELV7D9zLaXke45pL3VVgxp9tOKeWtPlOaxEekPWLHJszJHPpz1ToZrWDBC+z6v4ewDrjT
TnEVpeKZuQQccUDaWEUH3cvK6lxr6dL250II7Hk7gaiEfarAc+1c0Zie9cTh3t/PxUUlbIfay125
OBvzHydp0Wx9A3xSA4ABgjx//8Mw2ZNX2xHrkhxvtz9AK6Jn/+011EPT6h/85BRPGH7K2JD3cu4v
TIHvsMeAjPdxr3Kjcfr0PBY03cORM+EEkn/IKaGEVSaYhEsO6kHan7gaszSnDo86vKudKat0NCCX
aNTy+NZ9JOVDRRB1XWshWyuk5CfX/RZCDzxA/obt3mif1oPGG7y50T+5KM/dpkGZUMKRNxIPXs33
8D+i6S+3XtBbkWpqZGI812Edp16ODagz/7Rp7CNzDAqrCi8MEdJYO9JvEuv9Eu7k0r7aJ2WdfAeJ
cZQsZtXOB3POe4m+tIozg1cDmqkNCAj5cRfbuGuddAKyZZ7ix7l5jg0utVs4cLjrdawDBq6QMEPn
aNloOuPkXR1DaHfVN07g9LHLbNHcg24iQGhx4Z8aGIwWwn5/eOH27pQjqHL+SwhOWb8E73Nt/1BM
EgGySJhwBqBGxCk9p+wDJqPOllYgJvOjhS6sFZP5CsJEUrEQ3KoBaxb3k99rqQY9XogZRBmL2fOk
Lxq4tgW3+1wRaaeltGhhx7GNOY0LChrzYhmPC8f+zvN6z1LUofVbMBhVHPnB4/M0pK4E6y/sMDAD
/EdYNJi/z6RV+SA+hIAF2lykums8sdad7I7696k4CWCS2tE7A7yKyansbJ4gXUKs/5D0ryPfRsxB
VPuAZK4cmlV1//djHonwP8fvO2O21nFnfLfjHgsjnBCUL1Yl5Fmij3U+ejMBFt+tNDZOufvvF8tF
cyfEikkU7bktDrtUTn2T7C6tYpGHsiwA+7UDHAoDQ9HJ7t2jtHWV+wWNooQphTZUNL5tsWcuNMeT
lcgU69XYEEMS8qTofEGlrqGaZH75nAnRsw1xZ2xUwjSNkaaIs+YB8LIcxv9Ml1KN/tpIrGqNQgxp
gxAuJS/5uqdeQoUeJDhkiEtDC4EQZJWhj8b2xSOsXBtQC/7TkPjuPqBpkOnRz6pnIWA1dWqklO64
N67Q8fmqb5/v1HA8wqWeBi/p8uIfrpC1WUCxd+K7Wh8jjSHyRonRgDs/Bx4iDxcE4c4e1EF1uxAi
7Ais9jaGDCEXm1i/cBJchJRDTSWL1olE0nnZNNOXyc3Wl9dXFiNdyepvkhKc6AfMIVe/GXJkMkhX
GSD9GHbJGyrQ8XjBNEMHNt5pIFzLvBHj6zIGq9WOF1dRYiRIcVk73V3uaI8HpXcZSAmHTic5b5gV
SRUPXFONHMm9gTPOVX1bnoKa9nRss4nL9y4GT60cDD96DweoAmfNX5PGYxqPjjE0IL2UJYulvouL
8H4OpS5OoRR5fj+e13gzcMHyqgxbcR8ubugM8NCmpZcga2CHpcnvHnxRxlQhIxKBZVDC4voEJFNI
/wx2ccJ/yta19ZXd34Tqj0PS5iSktnjQNPKjIGKLr3011/E2ubdsyUblssykCO4js6yyZdfRXkMq
XaID+o31Gt/rtMkmAR3EhKEpPcX7pgnyi1zAR5T0hpNgdFqHoBg23tsel8O5K0WPmE7IkA3eqUzT
GyTy8NJCje9x1y56Nx0GMQ7fOrw8/R8QN5COEkOzlObTZyhwqroHBla5v1FAH50vNLZuKmiJ6Fi/
rp6DSSLOrCmSqM8dqa5cnNQOl18qy+IGQmhdyUjsqNf5ZfyLvDwij7/nnYFDRNkksuVjTM3o0OtN
l2y/V9pW9TxEGahS7Nt85fAn1XIcF4FgeXjCNvESOWBM08/osq2uJOYN/XXPoWFmlHosyge1lC3D
vHyEcjO55cIFnDjSG4YVMmrdH3yRVqEwai5oEZItlQZAEhsYA+BYdnockX8C1mKaItF3FOxNTc5w
7bLNGtUwWnX7lgWFUKSjnP9vyfwlTi+aMC+P+Nb+vMoRoid2tHuN2bTB+3cXHbNtWyYl1IYii8Ef
K2YoRjtbTHJXFUfgkleU2iWQNEshGEdKk+rzaFuR+rMjDPbTe2hl4WSYnItYDcbvAk9yrV+sMbMs
tl37wOOSYZfgMCiuQwkzVVak1BiM2M29BG37huUxfw8AEW/b+2FaYhsfKhTcOKjw1OBovSA1hQe2
KDMJhMRSd8I9bHujCkJp/feTqJT1C3t1WM/NsaBy7MBTjqcT2OlHhScDin6rv1eCljceGNHRb9cc
tMIyZhdD+0r863J95LGCAGzZ0HeMrAQpntIVocmwcHSJVpRBJvBvx61fVQCqwjVl2n6urud5Zbnq
8G2H6VbfTuzZNGdoiVOj4Yf7BWVGZF9ray5PriYMnG4wg3o+jDCIdErkkIZ2Gwi946CAj5lRxXnQ
xndIkwX3fmd3ulIGZDXm9Iyro/taBNdNiNOEtbNBNx5etbGRJXAlxBuBq6yjMSNwbOVYI+Srrq7E
YoxTq3EZCaPq2Fc67niuT3If64jIUKjw5PcHe+9DNwjZLq11H5O/Z91ico+yQ9gmdoh2Bl53paUn
aagzqLHZ4Em6TG6n009D7grVFwKdPa0fCHtITaWevEDd+rMoSR6JoFLkJomDsA9vWUcY6F9SqBAl
b8ZtK6nHl9ebu5w6O8qhUIBYnmcSt9KASFIT4+snx0VEohwlF9LxYFCuXrWwqJsfYJMSoIxg4lCF
/hUj8kfTBYVLYvCYMcCLcG+tb/vBGQOC6hn4ttnIz0qAMo2F3M2WULJUDgUDm7rBuXQfpFH4PG1i
Q5rylOULdAgl1xLj6KRAEvZ4PneXoicBOEcCiw44Ng60XrhlKuT5AM/gjj6PxtM1Ta2gYGKbeGYk
ZYPKP607mHVdS2GVSEIlTBzo2oziGEcF1Ig+SqMYxx6+TbjQiYctd7kr+n5JjtWu/2bAHwZ8hdOl
O5laYewrwu+i1zQZimrrG0CTGhIE7bN3Eewb6xG/XcJkHSAqDeCgPD3Z6CHy3E02UK5oFYvZcqaA
lNx0aOh1yx82qNyrgKYIBVewOqVFbUAp+8boOdvGqdLDlzQbSI4k+pUgwMhfQdmjdjsBCmdRhNCe
exJ46EuwCYUvNB7RFl6hm7hLlvQwr8AFya3iiyuJDTTSrGdCE2M1SalKGsa6PMjS+T0s2HzH+VPe
55wPSvy6YWaNadxFpdCPMaPNGUpt0f0OUKCKH5NU++Osr4uDquZ6ldqHFEWKYZgGttHPgbKmv04a
srpuoqqggNpvqqOIegJ/7mfxdp7yPc9sjUMaSGjd1c7ho9jwYH1rL5iwt6FPxmulxwX3G5lhrFSn
iEMxJc9qYbH4LZKtglC0m9BM2OW0wHkSPrRUQYTsF21WZbk/A9kRBYu28U6X5fzGFL27qqA06q1g
kUBypZ/MBmQKwLENW7OtImjWSrPKJ1lvL2uZ7C2hcJBvjbtEnv+idFMRLS6cgxGGdj8NeVfDapGR
dyRA9I3EE5DLtNHS5fZ5hbNaDNw6p/Sifvx1TCGE45Qjzk6MdYKkjxZXhWXUiGi6RSe3SwwxPNkO
OzVrCpdT1M0W7w557VRFExM/kgP/CAvDNMvxP988nIcpAd04JNpiEw81wAORY9+l2dLuriM0wY8A
Jd8NrEBWu/432nE2nuNXbxHYgcVNhl2+BI3XHwqZFNUxWkdtB8inFWUZ7U4iplLmy3JNpJHNkkJ9
ckVv2vBwy+pvSmo3oKn2Z8/CFQikrQY6g+CyIs7JSjwauDriEfQmNAKA0ztzWjYvf+crQMYtsxsL
5+YUnY0HvVZ9OvVSGcPaw8iWGLyhrRInh7sS+XD/cuMzUtX1NGiAlM/RXAQ1CGR9cdq/JScctnXI
JZkEOofok4vwHzZvAvAPAxAcqvdE5ZdV4JwnOOpITRA6Ekh5BXWgV4xEDdFTUAKm5HGHCPR7ClPs
MaiLlDgqm8BfZd8aqEs02IHcb1pX4OxKdpFXdyNrQ/1aLf4e/I1LXGi60dL3dqsNCLBdUheLY+w/
Z1FTFMW12Tzhd/5YWtpQmBl41bcJLX/Pyc5wdyrv+eEzgGRBZR6fJyCmy4TMO/NjtpMQwabGP1PI
AaKSl7YJeVrDwQNQWCfgkMzPAgISuTKCp1vkFE7yIy6etuBqogyp1uMn283mX8hFQiBfEKGp9XWu
3BFGQXseFsQFMDcSlh/FZAAHscETkSkqSmMTasBeROuuGDAaBtFXXdKUTTUR7OoTQQfyB1TweTyi
/uyhDkqNDnk1F0jxiI3WtaCxwGtrZmE+rGlnCxrtFjE1cvNEyqrCcWd7Kz2/P3chkpIt+UonNDbP
HBXPJze8eLAFfQlrhbAhXwrAinYwOCYFX8w4M5Jo3Be/Q2P7KnaCKo9/ENNDdYc2AjtEEroUrREm
r5TpU0L3afbMBI+AfhfOd4DUfs8KHnhFdDoAC/4z7Su3g+UWZI6zDJAccdObiC0s7ltke6thtmIP
RDTpm74YMfzTwuGcOyfjxDeH6KxHgfGEA4WxNWbwnwMKR9w9j9s4m/saPI5M6ac5Wlgg0ncSGBaT
vPZAps16ArlDl2oNTKq+a170ulZxxYGomXRsCjeCTcuEFzgOlWa7HW8o2T56Cq947uVxzIaY95oh
Xha5U71tUG1SbMc6fB6vbGRjaRynb9FUhTNmayrIP0bTjIVrE2Ive9fK/ep5VMgf7yQiY8uQNKHu
uwCCNT/RhWP2gss9FKlobifWmFECEr61U02KdxpZegis78b4Sl05WuTCxcyHoJV6e28KV/nWWRzo
6kh0873/W9RFIkKf15WXH6IADy1es7P44TR6omMuRYsTOzdKCphVzV5pnE5JGejuYCzBCjwdex5a
jQsSfO5qo+plA4CMMGrKpboNGWzlgkopX5teEzAOMFmv5YWQsoLWcM1qHXrPJyO3cDVAxQ2WnACL
5vmZJ6uz35dCEu7iEmWe7b29PE/ZP9icD8+0w0BDUoa8/T9Zwb1L3GGguwH5uZjxgO0RUDbNcQ6T
LEtaQ69ID/tHNTgDptASTwXZWy73JbvzWu3seT6ELGYpYpFVkfb+rwa8MPNX9y8U2Vg7IpDqUaVT
G7flcg6R9u1CITaJxD1XQVtjDMA2MFQ7rSzD3y7PxiMyxwaM5z2seUP9YaoXtjsfjMDeIXfZtGjx
q70XCB7M0n4DWeNK2AXrctfR18PQZSzx9hooYrEOfFMefw1b3WOKOxPVUcWO0+pUdrXEYoZrqVZD
y5mw5XDrjYmrxx9aaOp+We7e/K1aOmmwB5JfcLUMCFJ0pNYyVU44cj0dXfsCKH/mgWSpLou/qewT
XPG+LTFOxXf6PyLTebRBBLa70L/WKGE209SmqFtMUR8BKaBWmZiVkD4Cqe9+RkDLeW688MWkcQKA
0K8MXvynBf427AoxHeJCkK7U2Hnd22iXSQOYzL+t2GoHpcHsKDfavV0OqUeU0ExJkqoxn29334HO
wz1BaibCvNLRvFSwcYAO1ZJQC4wO9KLR8hjse+XDRWZxuYAhe2/0qneWBFQXkaA4XXrRpaKBqgwN
x6rJJeRMBpmSXXFZgDYLjtWnzv/1hBa17zXAJJnN8BCa/CKSX31vQKv3AP5ZU2eBZN3oL3jdiDSy
WTvnT3AL09Y0x22uNOsIfLQvrFNma69jDkbhpXp07e7WQQJfCfSnGmUmjL81erDlUR7jjcZZ8I7b
/l6NIbdAp1dHaMGs1yxPnu0cgTwc81ziN1jbKAJRvje1+VIXV4EVGRyDX8y4z27SiPFSnKhWJ+6f
DaJOciVahT7uTMzIIjS/gpZS5pY1wfkto3znhj6ISHGAbIgdJqHCkeSc9ufupe8gTNzSJZc+o8Iv
FqWIizdaJ7bqLFjGrYFPqhMkwGwq6VBA0p/a/sKAodOwgmu3koPavvA5D2G0JtW+N4zbW/RisaZ8
Y1/g7yeu8mK64Q+gnwN2X1aDh62yiJU0MdK9CUB0hs2s8qVQFUYlYRnqc6rREtOYOGppcBu0U1e6
gFLlFRgsQJrEbn5ggdq85Ien281ms/yCVyLtHU6/y+5DyfsgsNdyVKuCZAzMKUC3KB7S1jop4UO0
Fwalb8tX3OedhDuUPHSw9keF8V9GxvEKCb6NBFrMJvMCi6IdtwGvRRtagPYnAHGFanbNGOTUIl0j
cSns+TVhpCYtDE4dFBp3Ew/P8CME5QPtt4GZJxL1zZm2tiHPtTRbfpK6VpQEugJWAt0Ab7Hz86Wa
kG7/slStgGWrgsp7Ny19xgwtMEpKCB9fmncI5MeihIo6OYDlqlzjMyGh9lwG3TNclS+1wuozAl4j
ZzZSnYCy2P+/gB33LnJw7hINA4/3ZwbXHsNgnJI+pID4MS1GqDlyQoLn4c9cLr516Y24E9HI2eA9
jxpQCzmxbCy897iY5XIGuFuKY9GKrb5l6ZrKNSWERPhJMqCbI2oox6TE1ylmQ5ZDt8aJ8g0OYrJy
VpPXtpCcrjXPlnr7PPSdGsuOhFXIDdUZu1cr0slGawydxZr20h1XFLmF6Qzk7n/T84oMDrPFbIMj
aSauPML3Do79gcOXdfIn0Gl3NT0V9qJP2yC1H2l3jaZ5SVQ8bkDHyZb7xuulTHEok/sljtMmj9WW
vLJaF5nZwXhipXrCgXbCyVhU87IB0n4991UHexRtjCO3aUIRBJvXtHyKuJmXdP9VXtwJ5wW8Z/Kh
9SLcE2BVGZp3eGPXcMvvMSw6/hv2uVTv8yVh3DjVuhZWnuFm+a4ogibqXzRy8fbT/NO6QIekQ39w
AxVIeIFpy/IFcXtia8dBLxFE3l5e/niljrbCLryuRzQIzeEROXXyY2AVxaR/LQcXeQv+yBnwRkMJ
rXfCFHrfqUXftXjKpUHREbniMeomh7wSGL8Cr6tt9vvOEk983n7jprI+oPLoDv4K+XhT/FKkgkjW
h0WmEK26mkJXPQyyxxxg/qL+GxTjn/7FskNdYN4ODJs9hpO3xz76oKw9GK5ELH6DZ4koIzYjl7Pb
fe0QpvWBj4nlPkVUiThh+6cD+WddR1DdC/e+8jOi6x6aqRNb49WpsTMRAK7WPjaEtnbqfHayt10W
KfRAQ3o0xwbXbrFk9/3dwUhi430FdzaZkMQgZBGDHkxgWoEFcoZRWLCyUHjTsxsZ0FXOdd3VPWGD
xstqZt8AIo/6LIWDLjghnzJGIgvYECVbhFulOBbsh6B7qvBAzpsmCdmeM4rwnEBNnUAATrlkSqjK
Bi071WU5t56zSvF00YkQHcLCmAmijJXxzi4WjBrhqKu9BZoMylWXEbHbOfLQVCLS38dRGZ7c9QhC
7QbejOMH4nryX4lstb1pO4CI4ID12L76pABxRYeWJxDcXvWBmNhy6oma1MIYOgGn15aASArMRkx6
GQQKSaGmdNchEMehjsZx6QvZPIv+eqhhXLq3BzCHt7nxMDbXzGNu/BL2T1nrEbTbR0fkEe6ppdIz
08Lw39ydYBZIMfYJLP8eUg0mq44d3p6aber6wymm9+EpX/O2GGJizGFi2tQnBe8W33uOokpMnrJY
4N1tBqm1ALtD3NbC77A8tKGMzIDDXSR0HifnkldJok/zm5d/piyTjLuZX25cwxn9JLT1TII5aEvL
ebzUDj2Zc8IEOAYZe6iuNUtH0V3tNWc0gwn1TJCAf9ZowXGHraI4CzKqZRVVVWLGbbsa1imwDlCv
q7LN0P7ZMttclX8CjZY/IW+TtPzh1jqPCt28+yAa3tluMwgpQlbZzFxpw9UGcitV8Xalfg3aXAjW
l/sZTfsabH3nZWGnviajVxBcuSH36cgRxdOY71dYjyE9KSKTnUvX+p/S1Kwe/2Tx7whZTdwPxbsp
q1uvi0osNYp3KTn3+af1k5Yiwu8IHZPqcatSXvG4wQusSvOShP+UdA3jMVJpUjK0S0gl4q6ELTw6
KvmYpzMWTSBEN8n534qgTS4MI9w11I8niA+Ftu0eSnlC2trJfs04+40GU4bR63gHkhqfWEyM/2uA
c4p0iUoePU2Xk1xwd6IvJhVmQH8sLYDy//zJXze04B9ezmYQ9Az+9nrLjatC2hALp16uaM+U49IC
/YB5O1N0YG1ng/VOi7lrsagAhsdjokJ6IvVb0qNa/bjEjmA5JpiW3PGs0q7mGFXi3HrMZib9peb0
PC+fX88n6ijZurV45YIFOc/nzuXSE5RpvY1iijQsQbsbkzQX+BROnv8dMg0Tfm61FYOKqk0vf2I1
xR5EmoeNY+woqidoXo9FLiOX2eUCLwwB62aFeqCv7/+a7GmPIpOklq4+zcNqWpzfxmZhGItAhe+f
y0QCMPWYNNTw6DvHavm6/2gJhyfHEnnKAYnaVzMO9cBUHnpvPQW9O3etQsGFBW6Ykz76BoBSd9LG
ZSbFI1s0PBi1+nZ/eWn04QeWT2xZCWhvXB0B8IP2zF1mfL18AcIor4Sp9ACcuLt3J/Lbx+bsazWd
b3pYoWUqPNvw+xDBtc6lIpJu9x0ul1B8MjOycZdx/2csFyEf22K7QGOOAqKFrW9w3hzsHP1d97h1
DxZnl9zSi1cRmlw1vN11Q8VzyBJp5Lr7GJZXmznc5L2x675XL7OnBFNND+ao0AlyL+gXRVi8Ntgm
OPC6pnweWcnQFZdcbpVYoIDVa+29So0rpYHQ1DYEkzQp1PQChymD5hKX9WEzszbioyG9lcCMfcQe
rLYT8ay5ikc7XoYwgPsRnkvQqWqZOZ8FX6n3bpg6uSV1Ca/F3jHbHZfdAKofmSivMLxh74qVBbT2
e0C1oxCiooVIv5RFRkXE88d857BMhWkJRQbJ0qAzY86X4IRwVubJlxNUgb5rnlKxt+QHCQB9oIK3
kuGwrZBdQGrWaJYdd9kVSo95vozcD375939FyAHcF9rXInDAKXK7qZuT8yYYEVy97zhT80uIh1o+
SiF9+gOUpOBizCNOX5B89xT94Tp5vfnFZ9yxFnI/N980FLjC+cpw+t4x9ZuClNl7OTKSDIFbRq6B
MRcR8h9aihE8cnbyWpeau0sPqo7SADvauk4Nkq/auElC+xP3R5n9a9/vnMbzFTy9Df5Iyrauo9kk
qlra755PAdduoBnaoWho/4ejCGfv2vIDvTe0PA2gK2YSucFw+Du9N28IJQyhYj6X3mF5oaFU6u9e
xXgznylLnldFaF0gprJFZlHyhaJJGRnflOhUYrsfL7WeIGrmF3SaIFDRuojFYEUGW2pS5ylo2spF
v/vF3sZVvNjbWYOVMDciFNmJWeJnyFJYQJvCETxsw2+8HDLIc9TKUUrtlf04L14tkbfyGt3v4eSU
ZfGI1Fc45zAyuFvd4hv6rBb5wEInJxzu3WL131haoHITMtru+u8QfuPmkkEKO66Tn1mQZ02Nd8Td
pGl1/9zXO/6Aw/wNf160jIDfodh84XmCivDHvt9/FKU3O/q7ea2VCRXJvT29kcc03KBsNd4V8KnL
/s68fgpCigXlKii5aipMpwDDUi8C7op0nzANCQ/7C1wXag3mBJMDZwNj18Ekl6+EEhGPusTTCnG/
n1N9r/jFsi6Lq1zNYvBYcZIx6Y/qAteuGS5J8bvrCLCO0KXpyw6ThqGnvU57JRsIBxQ2l6lKkUnw
VWxkuErAStctUjjpSFvW5JA/XY+mCYIxoWNiYUl8mw+wK89iuacX9WREoidOCpZcaZDGs1eXCe0d
5dKFTDCavf5EvMI8xuzvAAA/xjjbO8tauSBX9EILFBoo9500TzD59VHvU/M1zmZP9dCG9iX0sYm5
aeiOLyCRECGxFep4sP8VDRwl6gAeNaZKsCdJRG/mbiwHe7j32Bu77cD2rJ/7hXWmxmToQZjJnDnS
800stZWqDgA+dT4ZRht2403EG8bCfU6cFSgnRwumWsiB49MvtZUHeN9/iVcwvnb+gIUybZubFpD+
/pfIAmFvqkf1lwd/7+eG5f6i2V+x1L3UKvFxFrrP7gg9FRCV1s4XSFTXRsaXrnPxO6wq7Q2+u2gz
fwtFNBM+vvKn8NM5+FLOZG2dBaC2DVr6niwrO7GL7j4Xvebe9aLnHAUBk3Ufv8b5IqG/znqHC4tN
WhEyWgeYWEDMPVdYRt2PIlEBnDXlxIZt+bk5hR2V13xuWDgOT2mo0ZzOsL8Cbh/5Am84G3LDMual
10fuQjlvlwHL1fu3duvs+Gi7a/InlKE3QcN3sgxwWtsvRJtjhgoboaM2VoM6g9B5Yr/XfvGvMAfF
dBdXlpx0tgjlW0qt4fFwOsXd6lH946OfPJvuOuh1UYItzuVAwX2XeVRBRj6Nl/ksyDXL9cAcSN0Q
MUkOjTCF4hCv0qsby/43nfbm3W/004N1aGSEXpHdf5bjfHpnA+Xr2LnVIpXx94ZMaScVZPA5Yryo
VXFlMwrNnJJHw9AjvAzozbO7rWQZq6Ek7rE6HNZxsjT8wcxdwb8cE9p+Ogb/DB2nwbg5VIzcXvTK
Mk5DJO9y5VFvFisr9BMtF11VjyVdYj0yer7685A7vdeUFx9ejhXqXMlQOOSt5IiWNuJWwZ4WvBhB
sbJMsTiSRNFVVX1cQhdzHXSa7cJoYjYckdcB2OiMsWqVQYVeAYV/d1KFcHHO0dkJICpHR+sm7ZY6
/x55jEBEmHXfdwUoVEdkf27Kkcqdfu+9QmpPGPukUoeHuK3h5vYwSBWYtFQ0+qd6b4YF8Hn2UJyR
FfGpUg42ejuUmFLnwVvnkqQe4ROMoewo3muj5F7jPmSWrz+V891Wi1ZEYKSPRWaqOJetjgywmZq/
GIkBhSSui1Y0qLZq9yluIPVXKTEqomqh4J0fcLXWQrLaowL2oeBbkn1SDuciupSaVB4858ijCBDz
UQ6KPD4NCKQDJ3vNWxFoP/Jn8s0ooFjJthgTfjVnI483Hs0t7DcLU1FJgr2XJT43oXIGZwxLw6nj
GFD6nzqcUqD1Gi18208aB30WvvDRhrpyrpJvHFwylswm/0GmaDsuosU2twcveWlAFvhCvPd1Fm7d
8WrJkF2Mrul+E7v7CFbUsZ/NTVIQnOOlKZp3OgbHclivklI7R9LrG/miMNxCLUIfwvlTTikgZ/Vw
NdLnXepbLQlzwspAw79VuOhE58P1vGqCDyJUAvhKHeHz66M84nW+vnYCks3dVULqh4S2JTc7mM6j
UwK4wDgigv6Lj0o1E4PxfNPM8SXHrpmsavJeQ0oNFydIRCGeL/EOQ4b/Vf1SHOk+BrfEBDKCa8l1
lIYVDFJI+aR5ibRHN273Hx03lrtgtwAFXl2SIC3spDj1ldMsgbM71a9hNdGu8sMtpzruhsdkWpxs
wobXMKD03/Ez49JGyNk3VtHR01rhrk1ow83AD2fc0KxfC0qA4HfZ0+y/9gWzNC0FUSqqqeB8AbtN
vUuNQB79HwmiMSa9/iczbpeYo4TcsvtPDpyGCgz5CqKPrxdw1+EdVmXJ2SZ4lZvZbBA8AgiaF9e2
L3vD5j9GzY0P0jbnCwj5ETmVyUPjx0LH/lwe5S/1WfNZ5uFZGj14FCeWkhAgvi3Kn/X6FkbB7UPq
A0diPjaPY9/pqjFSzUyLCJreoKsVoMZCp/CarNPuU6IRUfqFCSFBlL65QkgyjLrwkmDmt33YCmdh
OfoPk5T6FCXFee4MlPBwtWCIHwMKxdWIoDTG9LU4r5NZAp1q6tpLSn0ZsCv4hb7xR7INMvD/f0O+
JVA3TXKwYu3v4pCT+FmN9Dc6a4gPn+1luQ+UE/f9uVD0QR1tp795zzOEyqj/5/Tq0cBxuJCYTbde
hr9luJjPpoQjKRQFB+YAN4gt4+9SIWfrn30kbjGsS/zUIH9P18983WcJGzFfXa6Q2gd/hnL+tewq
YpeLw9tiqupbKvCeL/6bZWxNCoSzmD47FIcdXYUXzmdGK+yUdglVnxF5uqndPWSdzk6ujrqjrKrC
HlB/Zs35fkTO1NHRQVg3IwLIVpz5EdAHE53u3NRxJGCjh8BBNOB3f+gClgX6AUimBFy40mjhRv7G
kjyC8H5NfIgRxxBCBKDu1WeP3guBjipW5Og/Dvq+XyEB/+HrN/DvkdZAa6eFZL1yrCFY9LG5PZ85
vg6DtLJSHkfKsl5Aj/x4fqPBlhCPzpTXSX2xGpnVUhIOm2T3BdMtgZ9vVOovCIyuWohpIrIqBjzC
b2tvNOm9tzrzdYI4nRm3Di1CesKKLqmUQpHy/5XRcPzV5av5NXQoWBLeMiHF06G9CQRcaOM/tDhb
qN1X6iPTxUjUj/LMOE2kgwzTR+X6zZKkp2xrj5KGr6R5myxXhokbXKp6lEXLg8PevpWBWg/uOw5+
WM9JSsNPY7lVLw1LPnJzbaligW7MWzP0YfNvGStrCZM9hlHq+rmOeiQNWAveN+wp97xr4dG2rkKd
0zijHU2JEMQPRLGvHonY++WtXjd53Wz8YuKnSPmZ6zLQTKq2TfGqqnsP04ewmHInTdqdqgseo1/c
+5xpy6A+mqX2E/Bs9spcWMPgs+jGJjaq/Q18xAl5XIGEA6YAstEcQVBdjPItMC4VeTxXjCfzHLcu
DGfhcbvhUxi+vS6Rrx6QPRcJkusgV3k1h7N779dJBEIvzHlNkkbmMRfMnxa1EU8bKhlMw5CjSEIj
n0RU5K5IeHVLvB5FgKuzun1OyhKkOqMqWARKbG5wHsaKnluzNDcLHcB+8adNSQ5oajALlOmaAaZ1
ENDSmNKR5IuExyvtJVv+EW+Yy1qT0D67ajc4Qs6eZXWHzLHv2ON8s7gmTWoJyPi3ZcWDFTHcCdKJ
nUMwA//GV7CuDzmi3b0L39XvP+DZEET4CRClJ4Wqb8Oxfl3JUgKtCqQvvGwp8ptk9IWUrQn1CNrJ
47+BVet8abT0CaGxqbbt6ZH8J5xzSNUcU2AVKSPgqgoWQzA2s/kx23mqmqgtERinl3Kg2lT3yY+r
06NXd+KEYFUWgbpMlueWEa8pTLe8l8Erse4e5BK9rAqS7wf7iGcOVQBF7s4f2RfA8MJP5X0auTjj
eMPe4aYrmlldUB6/Ij58rFVrHIoSnvhMW836SQKmUn5fd0KVOgZZJ1iI4THaSUdFjurSRzrgZpPT
8UMEjdyKBrXw1vG9vT54Ye3ZtlsnLhAMTSqAG8nDitc/g8z+NsGyNUV2LcOeJ2cTBwW84YgmcdQs
UCpYPwFMio0DnrJwxgAtEta3IGtMvDZD0XWuJmTLyYk0H0NfQdax/AoEkthqm61T+7VVKJJSbUMb
0wwjgsMQP5fn1MiSMF+WrydlI0n4SXLW0Qg3Sw7VWSxuHZ3W6zLCRk9mUCJrmMfOaAz0Ldss7chQ
zC4gMLdc/aI6PT89bRtijke/OvKwBMqOjfKm7trSaG9UDX2pvgeyJavhZc7TpPD4IUh3ZglVMx3q
q9z/kYSlOIRuA1C+9Nk3SPKV4ZDgB2rnNYMUeJVhuh1lKjfZLJELhX2ms31b+qZEwh2zKa8ylnnG
PTdEoHWtIBF3mYyCzR/j5yYL7CWYvLhQ1rYLzqJ9BNbr93RowvhgmX7E54VRH/y/0xaIEhbdu+k+
QIhfH6FtN93Sthicj61cyR515OopB4dnFcnvZpwLM4YANmB+F0iA88RbBHrm8U/ocx8uVMcJijev
7ZnVge3Jci744kmzR1VmQLcbb4Y7Qy9pk9R8yMf+Xf9jr60yJKgfkPY0ZIOFD6cnSp74syjMTHwY
eau31Zli6ZeJUdFmVfFcDPBqfgq0M5rXOIMj3fiySK3cuoBZCV1vaggewU2QSGC5Oljwg+5KIFMB
JhK7YHwjf3fRv1dDxNlHLMrOs1kfcP3yvn+sbWRI1tovJJJUZ23K7TYyGGtY0a91eKGppB25aeDn
m/imKCE+SdaWgzOmFfwH1b3axnzMxqE+klJqWigbvQQwIsHHxz1f/oNx2ranGHUtUjFDpUhRDEDa
W3tGWu1r2UIeiEY4gR2zIkwpIeDw30Vt/s1iyiOOImcFBUHV5JZrDwsHIzQmM6RIvtlZEtr5oRtB
FIUoNXP4j591sT4lwqe9exnSAmdnURXaDT4CcyA+Fnr9bbLoVwf14ixxqrLCt75maEVjQnz4QD3R
x5JxIRB+X865Ne8AZzELSSz2mTO1J4b7XfJM4+6/Zjkw8nFRc/fztuLhqRtAVrVYJcD9S9iU1gZs
bERX7n9gApfE8/L5qPTJN+PsBA+S8N15HNRjSPbu9JMx+cH0IGzKOj9CmViv2e1guEckNA/D/8ZA
vvXkW7ggHcEo9FnyGd+0y1WmHiMkS4vKdvPcad13CMsmKzydFfYtjIgBLtmabfNe+1gMsM/4UBmV
IJthMONtk8+rTgdS2JfCbyb8uYHQOfibau6yNl2DJdxkNEIT/YaTK/oVZOENqhBzM6Z5jQ/3a43w
8pluwZnEKvBln8FhLv23C//AWzXu3w0q6xKwW+6wEnkCLIJNN5cyAG33QNumBKUI71x6wDVBNeAO
tBr+SX6Ns0kBFfT6ZIZ5m/nB+9NAx5VVFirGD88S46PkLQaEjIbV/WAXS6jOlq8ni50q0IXDGj0W
+0Fes54EKTAQ0hOCBJKmwSQ0DVUn8n3clz17rj3A+VpTMG33V3oDXFXxaK/8dwPOW1XCAYur8WPv
ZOwC3q446AqmDwAeusA6RryWARxYueNQLJqPqsvN9Gor9s4hqJ7iOR7agc1cEDHdUUeeTGPRIxSO
N5h+DJIe6iD1Rj2u0bbOppYhMLfiDxF6knE3hC224qam7yjg4NHCoqtt9wuxtErcgHmPCSNcVpXm
HswojZJam1YCLwzIjuKVT/WH0FK9Ym2wbCEjB5VT94vuUa3WxU6OKXf6OMvUpETj6tU+d3sJIJa4
FPNZ96OdiFoGigB3Dum3YI+v8d2E1Cd8YAp7MyE5ykSlwTNbUk3mhRLtV88AEJ4sPtSp/4iUeYhe
gRAVA2zNibEIpf4TC7s2r382SMQ9UVk/qE/3v/41e6w/xyFBshzPpafsF2x1fw+r2RHkVmQrEZza
Igjthd0dvlCuCZMHoRELtE57HK4nRexQ7El0mcb7uxxsbgvVx1CyT0HXRYR2aIr4CAdaC8FqZVW5
i/uDNT6OkS6KlCWCiNm/D/Y+aTd79Z1TuWd6VcFjvfEq0eafii02afCULGiyugNtmkvwhNuFRDeX
umNl0jMhcrhgxtYVNRYQaN4kAXc//8FJCxJNWRGwZb4nq3K5iymsxODZY6tHOoWwjbEO8uUNG7dx
g2lH7YGCNLdbaQvy4CU9Jl1Ia+jbr+6PcaOINYxCyIdA78vnUdPPRp7Za3rajpXfNwgzez6bzCzd
kPfKTaZGkv1YTal415yAm4HHkOlo8l1Iye+EsKbiOHhlJ4486S7vCm9wJCToEvr+ZtWHM9zJ/Cy9
w+bO1Zq7Mv16y+3qOSzoARpMb+rzFPflmTXvs8waWx2k8jSF9aK3OPNkb/VsMw8dKjsV/7QtvxyW
b7MRGMAI2NqnboUdoEsxrJyIXlxQvvyHc2ur+c/44YHIvgaOy3f/w75EiGdwpyOnosCuOP6jpkAQ
w68+rcC15mDPkJ2kNQKJz0s3M3AOn9RZAyhzXU/RIpGy0HYVb0WVAMQSyX9G1QgEnfIF8f1mKMEh
8hXVMXx0NJqSYOn7J2gEyzw//7h7FazC1KDx9W51QLJVF1fEfibnXtGAwLb2OH5FTGx9Iut84/fv
vja+hsHPIPUeqf09I4mO+xvd7wbu9VFJeED1mb7XPHJhXr0vbDJOCK0Tvg9jqJTnNmSiVbnbeSSb
z74ASYRuEtF1vm8gFchI+qRnwJlpLbYHfRNcI+yWyXcuEDZO5zqUQfv/l7ZBa5wkJfHnHjM8OEzf
B3CTFqmwqYSSLLueQftVadVP2k4qGUOEC50cOc34w6JTzrXFC7zxr5A48vs9hrQbuyDK8VUTqDMd
WD3CaYtTvQ3s7mMvUzvFODeeFidd/li6His2WE8ZU7bG6pJyqMPXF0p0Vw20bb9YUQ/laz20f662
taDSoEyx73SdOS/mxgLXJoPjEZ4nGoHZYn7WhFElc5aaAg3HUGAI9xMa+ttnHvx/f/EZMWylGbFc
AoWyXaAl2HM4MZzln5sPRfSFusFqUvUb1oCkA/pUhGAD1pYdi6m6qJPaP6033sFD0TjgLNOaDnad
eCApGsD7bELI+pxPOnsCMhTAM7Myh3PlUFmkfjEaHwW8SsTHERfCyb2QbMWNj5QCmUq39QtkPrAW
OsM3otfVT84ecpO9M/Ob8ZwUG+MGwc2G9SWQI3KjqpdDnOfT3NB+69BYoC8YC5lk/L9U8v74YSbK
O9gUyczUh6xwVpwERIBUMXcIlE/KtMfGcCcQEI5uBfoNq+BMzoMoQRntDIV8ptzkHMNOScuPTcev
Rs+aCzqCoaMKYOZqIUwG19agMu/uWCgI7Y0K1IY2KHQ+KaYXM7BVVlzRN198eAHGSRMyPU0QKOqS
J9Famn/pvZVnqyB4x277SO8yR6IJrys+lCt7x8ua8zsYSe+kjCH3r0LCp0wNx1WXoqzg4RjSMuhO
FPoHDRPzjaHnQKywupMaeLe2oTCnbZyScZ5NUxK3LzS/74GdellDb8cnAnhc9Gv4Yk3sbija41ER
WNN+zjXHxgkdyHW7fRurwjA6gQIUgBqlmK3M+jJXE5PqUCX1x73qeTl2aXu43WQMkjUydRAOfI7y
IoX6eQFoQ0WeIkh/pI/vYktXgVFsu40rmLwxdbyts97m7BVPRcrLlSu5fYrNDRnlZD7jFLfsJd71
6szvpyl+yBDK2YGUP2ZQQfszCDNVLFCvvrizka9QtOtcT3p1sVpMi1CrYiYrhXAOSSXnV33c1txq
P7ntKXqjGlHhG/51bAACoCu0yWJ4cZojI9OLJ1oBGwjOtBEFVmJnnGP4h/SL+QX0qjxIKZ701odt
mttvtNzri/MjeXeSOyqeF1sypPz7+b82+TC9KfNVp/pHLy39WSN/BTyZYCeCFDPFtbwkQEqnLxzs
v50gls5PIDlejwRhTLpku/0bjRhpsTLob6pxBJYBXtjcF9JAovA0B4ySB/YPmEQFV/tzkm4HW1s6
FeTIgfTmo66tYYmHFZJ5sOUI5RrDXFQCwzRTTIGG09w2jBSxtNo9U1qhb+6lW8yeF60rK8Fq1Um2
uNwpE7D7Lbi/fWx+Q/9m8CcKqUGVVty20OgjFl4g8NTUZ2WNoGDyoRc4coZJqzxhuMW9iEEmH6jj
qx6+iEoMrnNvA5w8hBdbZmRSEb/wZHwW6k//gjKrthqAMY13wyqrh1UbUTIba96rFvJTuAGuye+u
nZNaVJkvRQuK6QLBbKfAr2Q5t2tD06YgEDCX0pjsxOK0eJWMDNmhyIrfcAlwl887z/U2dyPHuErz
TnGvzNfFhjqcIG8mvX+jH9wqD3m/7yAaj0SJQfFf6sndkKB9QbXE7lmOwKu68HFXELsUTg6Nau6g
Xc3P+yvJKAkqFcPz7Rf2n1khAyDha60jmz3VJi66d2Bf5+Br+tzlNe8f+ophbCJV1iz4fBZyJHGj
WLWTHfgWtX7lzTPUxDqcCz7BGdIUBdjtpayHrF/yElEdRtkhRR/h47ODkdu0DrNC2gyygaMJve+Q
CW6OjkJGq2aj/QgD8N5lIFdJ/+BmuSNN0RfPKlM8vlZVjT5v9Nh1w0IqJghTCS7/OLFPkq6fGSrG
F+6k0h24QiafiZIATGmaMFQtwmHFNKAUkvkTpcoAMb7UHFNo4l9/gPWJbjCjOJgHD/h372rAR6KX
YT3emDk48t39A+ibNYyI5QWOpcE7dL6iAlDBFqhGaCKfMYj5tGt6PkCGVOoqwXySTlsha6QTi7CU
G7BNEqovsHP6H9DISz3iJbUWylnm05eSRDpyGAq6CEPQvjO0OmRRaKikTXw8SX6X6O3t9xN1sO7o
4z4xrti8M67t6Dl1vBGYSlJNK5859BXDXLbnjAAAPs3naPtIAMIH232OvoYYwh8HZtZUj0ExxlA1
py1DAYKXG7eMQ3qtcU4dHHPc+gDHF8X2RdQohjWqknd43mdUmhpJSEHBrhRKcreg28ezFhecZG13
COPe6Rl2zstNLigFJr9AsRZKQjliq8jhAnPUruyW18B7ecBRXADIYMAe0Af1v14Zv5Cq6G3ftNs9
edNMQZRekWfkHthdEwj3NpI6jLNZJoE10E+BBjAJtFLDtJbdH7xSoBEZ4sihPV7TLVF7VC4AKqEw
i3kizkf0kY8m96YRP9Bp+bUCJh4O+Ws9KqQTQsGfZvz95Gx72TPmmM4Ck/vcZKh3JURgIxupDHQU
Nhx128kob+MTYcnMleON4ACuUG55vGNnSVD5NfsSUkWue0rA6hPS7sueB4YC01B/8gRaR0uPqKMR
cOQG8J1bKJ2USjuzQIXvxofJuEzN7A0wTp1Ve7ONk0xs8bg3BrJYt+TiNjRSwOaQLfyjLf2cJsLN
7dgDvee/CbtWXkDAdqE/Y5ic0gdMyn6B1tbgNdOqlFoXjwpsXSVZrWDow5fHr3TaE2sYKuaHuvjy
nL5r277ihGUUxCzgRpLB0nDnLujbiXmwnHMmDeuzV6Ej3zFuWRW6VPsO6NA1c6ox3W+x9yHIxKX1
1EOM+dXdkPhezFybNMEiL/lnfaxfWU0IhcPq0jDHu7WGtZxRhXw6hzwOCgxhm709Jh3bc5kr9VUE
8IqF68uv5aIn2WiqA4/BNaAF72WrDv+dPKxG7kvbEZun9QPbUzDp4G5a6SqU/Ji9pzrWR8l+yr2v
fGARhieRxrVd2cVCbk8fAfP4iks7yqSHD7IgfTHcTCyv/PJrlG7l3gSBJ9dlQZYlDafO0Kqg+li1
UHrOmEKHrX3WQ5Q0w+oTKUt3t5ri5f29pUKMrSo913mxgzs0PiwEgzvxvU9I5+JZ5kaBH0RooKa4
0VTEm2ZOJv/yZ099HI4YSo22CjyDMrQ/m63wKVBbyhyc/SCR/Eql6LT6W32uuGlx9GBkY4H7ZcN6
qouzdolRIc5Jle7a95To8zZ0NnpGAy1vpXzg7X4IIxqPnyyERwbYs4tc3Ub2w6DJYSRkXCqv3wAz
+CSKmhPBR7gW3nqkjA7yg+nQ7t01Jd6blx/j8W6gj2N1djsCxEl8ZrA28DMzMqKUfsdBCXA+EtWQ
y/gh3Y/9vybpX/t7Ia/NmJaE2v1OpI2dfnqOfulQ8rh/XduDQDaz+cFkptl2jiQqnntbVgLLkdIj
ZC3ZWNwTRZ9vU1eqyCu7b+3zvRI0saueg9QgPrUokB28lhY9n/tk3kwgyJRuJmXyMOosIZsTM/BA
NE1HEmQ3w3M+0tDMiRaEadlVMVVeMDZCFLFitqaMre2j33MqWNsRwILphFV3vrxcNSmkBRXV4V0s
HJ+/AGEDx2obpWgeB4aQRnPO3yIzU0/waLl6l/aTw0FzxL9Yhyv7FJRGy6al8fhV6sOPgSFwfEk7
BpcHLJrdjWkGt157FJ+dJEF2undDVxI7V6mzBVwKvZ4aGakNA126g4mIQ9OfkJBS2ECjtTNRBNV3
b3elcInr6HzfwPTONI4kDqtlW7Ov3pvNX3pJ50UjD2myXgItTHgdOjEqHuNJnu80kW5/p8cKFDyi
QAE3/pwmQWNpzarnFCm43KZHIZSQy3k8zRcPNjTEIx8c9cnNfULjFQ1hNlFm3/9q4ag0xDjWqfVp
68SWplCPQS7g7z5zI/BSvTxgc2ZqmGxyCAQeXnXrhuNVkNcer7/1wx06eWfUc/tEJE+CmvD5GHOG
Ap3ZjeP93RT/RsSGp6F8ctYiZWK9DxyXIwJ0X/bTLhXMH7r5zZgfoBNSIZpxqPoi9Z/cpcx8Eyqx
A6+JHbymqbSxjV4Sf0mWrI9y2zWH3C+FklqLbwdIzdW+f7qzPchX/MhCc9fOdTk9Z2q3dg1fUSPM
6HXuXNADxHDrXqB4Ba+hyN/p7/xjtSxCj8/9KFBVSPSe7XGZQMH8zi6oPo1UPC3VE62k3jhFsj+g
jTG3GBRuh9pagCDMxm+utAjhDWDeTax1gnb8M9XkenH8ofYoIyW81IEtTgniFXmrwIOEslPn8yx6
u1WTlITzJxrK6dxLsnHOmoSfJutBYeowdKrm3inaQlya05vS4yYGgVTHwjcYrHR0VIG++AdxJOLW
uK1VZBAqjcn+x7kYtG4phynKZ44oQd0BdOPLKDWTKes/Lv3Vs368ND1eXwbfrGfqmkSsB08tips0
2vGGHQZoZkPn3pUwL8f+Zs6zkqEqruCmUdpXDchskmSd6fc0jrofFRWfZncsMMGRqyrFNprjC4PA
XFQZT+KA+fJH9RhFIzprOXmMZ6nybpom43lw4HI1OgW++B4TkM81DeJTZK4u0CT2cjQdNNgmJUm0
CgdS7AfV+Q5xjWHmgY02FO3i1mLP1Q84eyH/L695MKCTipwnqY5Zl057BAaw32U2vPzqUbprmfSw
Nt4q7deOlaYeXWYV7l7rwfdHf5M1BVW8P3hTip3s4JBXXFOkG+NEFgvdcI0MoKCCKXfGrEFanEkA
mDnAbbh4g5ANid/LAEO9gaE28PO0ynlqj4Q3ybtCB56SR2aTDb/vzAoh8cuLdq2u7ESGOUYBo3KW
7RpsP2WAPiaUl/5XCwOwxOFajG1yQZ4wbmgZJlY8gbY+CyE+ORQVBCGAjpGgkCre8PakD/CzagqW
8t/G2C52Or1bkkF+ImXVg0O1hd6SSOGbF8Pr6N4KvX4tjWwmjQLLiLAoIPCh+xmeOqmBO7lkBYZg
iLB76wt4olBW1my7FKY4SIPOthGwNpuZxF0e+38Pivd2Mj5Jp2AJ3UzNd7pKaSa65tVgG5KEaW7c
aID4jsOhyG64F40X6sQg0cEJF//RjExnccqP6XWPxlPfCy+nUiF5v79jquo/DaavpD+JDh8Hh3Qt
8+FMtkkJgHK+q2ZNEFgB4jWqUJYyf8GFxn1LVJuqSXMX1diht82LSZjcFbVabT+eTtg/RfL8Bpzx
E2RkyuHTWwyfKFjmoreOiQ0nRLFAHL6Q0fuE6qCR4trfbYaRGrg+oTKpruIRthatGky1C59wCzXy
nL16mPpUp4/qGIw3rc+0FwB7D5e/Z7vxLR9dvUeCEe7Y0d2K4NzW9aFkfmwmUnVLVqyID8DiFEQi
/jBn2SDaRyiU4XY+afky+KIKxSVtPcuS2F5f563qmdutULAKNVjSfTtVJ1jyXJaMGjye7xnA6GTS
8YCUiPhHQWLq2FTH5rcPgRHG96VNF2W0nhC/t5/hv5NzRwsvNXkw8ruWU9/ihxJVekDN2AZpwFeB
+rU8bHvl1UtuMXhrAcyhezPvQQAZRL3fLW6X4aKtM7hagA1GiH5cn0MH26hbp2qJ/jr6Q60HzsjA
yRipQeFU35P2hcA5N0A1Wlg1HKjg9pmzSqAxmWk1F1XLAjy1mlFFsOaSC56UthponwWRSbGQVbDQ
wvSlBi9J/lxpyna6U/c5rEBdFIXD66bfpSUxBddtZIF4xR4R0TBggkwDcjw4ECWUkC7ZpH1Wxol+
28PO15wgIfUC/GcQv2G4NQVvnLuI5gXJOyNKoQtXl3cxxhuaueD4CuhIMUlEYPIBLLJyyMgcO02X
iPxxgkRHOPjKCTDWuqTXmMOpdy7Qhvf2MNlxFOGCgnO+zaF2OrzZvocr0uY9h5eFnUJijAiVPlfF
Lb6N4fXpZVUoZs2wPfnd89M9KFTXbmlcuPTUESDQkFdMzpxKSyry5S5Klkl3JisdHRPjDCAizmpI
/TV9yiq3FCgEU17K3Hex+qTuGG+4DWFkpVpqrxBTQsc6Sa7qLWHTTvsPgbyBKeLB+oDIGWr+1guY
U6tRqv/wI8wJcDnrQq4RSyEf+kLpOetPMv91pCHykwqgZblvkMSFawl/xFle87P1YmRTTrNGgUsZ
XcSFbZWqJNIJNmR8hIXYkrQ1Rwmsf14jLdiAFJzOCMzgF2alshhtmkgXFWLOkVXSPVfrGaP6n8g5
735WwgLlHZXg4QGbn/X0vO3KgTJR7ahjo4IsoCErpPY/PySkjAQxx19gAoSzhK2L+Gj48I9tjIwQ
vrGx/7ouc8BWOsG8aXcS1qsEKzUa6/pec9BQdNpoq2RVV4QAuW1qRQObmpfEpNtvylAQo+sWqSho
AfiH+zvZrybFJxj14GQkQtPn2YN9YnoPMos8Yw+pXjptHirltNjuiezkEVlF0D0t9O9P9IQvJGOg
Fz7QY9wbOfcczZAu0tKWwBdzQjVJmiLHHHE3Z6DtKwBqvdFjbOvqOw00+/rP1GsYaK3rv7U6v0+6
L7rz7JV29KbXMdfwsmfn+7gAYX92cK53SRHlVDSf164mc347eW63ex/dxMh7R15EZ5sam3ffBh0v
b2dUIqEYOSul/NeezuORKgmrVzMc9/MA6T1RJimlGVnQSOuz8IjNZukH0FlpmPWMkI22Mj/aZms3
jurvCn0gsDe8Hue6GSW4c3+kESqzI63h1kCR1A8A5W51GsbqeWOCTK9OqHBXGWfXW+D+Zf9OtEPR
rKkSc4qBPpO70DQzDEwOHJxipY8JpomliruiYXITuqSQaBoH7BOZbEBUQ0Yi/6x56p/Ef7Ffmcr/
z5nXydsPuLS47gAm6GOQgT3ckv8bGh/zciy2JeWDSpgpcghu322VtZxnAxGy3S/VHA2mCKoD+JtG
YnckQY6Hth1fxZ7qelKeFcLeS7WYedaqTqPEeRpUrrFmB2IjI7BHqVc+w9vFM3ZYUzOp+LRsahqq
kuwAvUvHtLFMdoNHbKAHDHzStk7OYCwDKxEkfILuGS4MfkPMZsoKvfMEC62fy2godVU5CrGdxN6H
oVSgOvHwLawBuVOeeNqNOz0NnO/i4wrbUeDaNYZdimfYtfwMRAGOvsPq2vp2qlVI5Eq/ltH4JnBY
yauHcrE8DAWY2hm7jVj1nCO+MoZHoXu3WH5sa7eb8XaAdRbCqUtO6EcC6AhY0Gc44HodWuFBv92J
jwQP2pbPxarDZqWJpYBiyWS2aBtNYCEjHm/k6Cu++n+lFDCtQ4tWmi9JZp69NDK3S+PmXiNICc8t
GRiX86jOk/Juo6AP1+ZaHeOpansgc6iYW9Tlr/IRWLkLovDJUS0bL1+7UatZPU6qzUAKnLaN4mhF
6itNhSTUrLn2pD+Cuxla706HT5u64gU2nPGyaQ+cDNP9SI+y8k3v5EdjeiSs+NpanInEf/bEMAsb
y7U20zZT2IyVBXRiIgH/NwKd4D4p61DQtMHqM5XLZbFa6UrnfklJ+jeQXll6r3kBe0rQNKIBsXKM
5h0dOTm8vLaJSoj0Qs+Ea156SQhyAKMuL0RmayvrcFE401dD5BKcWvq3qocoRb54xXbeNCqoHkxe
7h+pZqOsFOUkfrVVSyvyrmxGlahrPqpyl/l6B6P9b0s/s1tI3TInWyHUy/fU473NoQmOGHQ6ocNH
gv/Saj+CVai+mbRfczCeCL5DWFFu/B2DPDU6T4ZAxn5sEAWMbkQE1T/OzpXLhJBQ7pfk9JuZh8z1
EDF5xLy2ftJxsX5+a24TmmrThAhCq2uN8OL+XugZJiKRIIcCcOxIY4kpF3nOCda9SldXdHQtwmgz
JJDJWHePR3ISCz5IVfPdEN8qrckF/sDXrYu7wJ5HcOT3Uo3Trre7Nvnrlatha1nJgh6XNsidOFJ9
yVFELqpwI/7/Ghnf27+NYf8T9ZOSzJ0j4x/xY/3dQhF1qc+jj2QLhtd1HsaDbx+bPkWq5I5TDiO4
ZHQohY2fgjg4YFPzNG7CQ3bvsBZqf4OPoROFqFgu7hDemer8M2tY4JyP3vnv+MKQhfMrCZ4Qv0mp
yQcViatHO3A7Qurx9EgAjlb+jOwPUXnX5rlGTnIESMB7IBM+soK8i164qYecg6JylRPD/Vj2IAev
5M6zsufoFxwCWUT8WavhFf7U+Gmp1omGJu1JGukQ1ANV9dtnTOyXYAqZNkSMahwD1ezJR8V2d5Mz
TWAgC9Wd/mhK4eqSQ+PKw9C4ohHHvtxG8bpnLZkB1vvle196mFJb0Aonf3trJSKxg7H+Pohg3kiR
Dh/EQIpqOZW79MhewYuntpLPB2IJPJ38npWM6DaapZhJiY2BuepidovWMFdPCacGco+0NAW53qmF
jA/Xc+/Q1q4pzfGfGMQQrKPwG7ePiWMWS2/wp2FhojNULqPNPlkPG/vbJS1G8PgdZVQYZBqwh4Ik
mvd5rwTmKi2QCT1JdPoEjVHR85GiEA3bGo2i0I2nffgBcgZUUA6PEWwLd8oAEHckxuYhQCgOO2Ge
3ZrCGvUhOnoPDtnt19l5j37BkrfoBrERFl7q88M2iLWCnVhowE++kgfpKSSxRUpnGQpEmx3I37zP
tiU46MFdajBS7P343mxgTlb4wwI+TRvpG+Ax7zIMcPAz3YjuuO6pI9Cz2mRjkoafnIQroKm43owO
5CSk7lq2igSeTWZnCZNjGM+tDKmq6uJDeBwiHrCDD9Hj34RoBu6lojnHgLE5wbc/bTGEFxCwv/FN
q9wZBQQTTiLRi8g9TD+eIaZUutQGXrenUHFmR3m7rxeP51iuJtLYLBIs0uHuvDbJKH/4ENBsJ3FP
Hh5Sd09mtoh+xA97H3ZSJmeQ9bnnnHo2PUf7JxVF43V1gBH5A6HOkDb4t3yDhiq5jUwwc6RONFZ3
F8HV9XIEZb0bkE/MFOo8h55UNEelk6DpuaGv88FTMLPUisWZIdktL2j2OR3ZzI424ZSX+6+T5Iq/
yWKqKFNPScOAmxVSA9doDkh7k0pcOo3cvvAELFdcAm6f0mqXxlhTT0inGQ1yHmEJxWJnTjNm+aJR
CCuNrTR+2G9s7zfake72BsXe11I4y/WfFlpmJ2l2k1mWtfZXKUN7kwGVskAp6KY/Dnfx7nNtnRTt
YfP4ey9tEeO0XDyRS8X96vpGBK91W8L79fdWdE+3cp+/ZEboqlvkj2QHKfZq85pMwUvd5sFCeHry
PWzNZp5DqstUDWtNWFiVOrdthsjVEyC7d6BTMT0kKCV95ddcWq4h2M0m2J36NStE6ZS/h9I+Itfr
53LkC/JUtjwQS5Nmn7V3+7cjlXtPYCvsXpiVk/nmcNcftqBjjmILaM1gS1WN2zOmELsm4m1Bt4N2
9Fs6izDsDEv1PuAgjw2dlA09VEaP4mD4HRLGeOQby1HqHDp69A/w3fV6qZ2tAtCKb0F94UFdSyO+
8SwSfzMnp/0qMwktTzBLZBxGRs6wqeuQqh4FdgS9xJnXzAEPsV75gzO/0JAe6ufwoGONt8X2gqDU
ALw0kI2BsxzR2PJ4891ZxZHVQnZ0/g2cafyt0P5T9f7rvxB8sjSj4ZvYHaO2GINQPeL1+HQz6PWS
FMrUXeZDfKNdg3mdaIc8Z7KETKhA+9eaVV27CsqHwUm2iWSX+VCn5jHHTQ6un5nZfgB54u6iZ+fG
Sl6lnaMDCWe1uPZpplojluckVdedTz9XDLkLgwEiDBYbuyueqDsf2/zmI7xZMhhEZUHG6L9dAk/E
W6uZVy/ju3lBGHksOZuxiuDtRPqaF/hqFs3VnXZ2FJZ+lB6NPSu5slq5Ki82HcC/q2sTeC6ZicHD
rfvG5vcTjKgJPP4qpPdBU65QaTxIOMF9w2YR0FuZHtIBH3v1fEiiN7bM/iF+JHgcKHbdekmS1/Rc
leimZe/22XJ3c+uw/U0Uoav+9u7Y2dgL3V69Ox9cdyCgSTCl7FlhgXkMbDasO6df5Zuyibg2wVuw
E+Y01VQK57qoWlChvAvRnt09b93Ws7vT7uW2bMgLpGNF4M/GCuLf0+UoP69DWh47lgbVmF1PaI6l
z98XqBdSuxljp7bbjhNzOWG2SQK0iwwImDupi60fpNe59FDVqC0haMXB+uxzizWdq6ggqWB5PQlR
AWMWPSH/Lpua25SeCcfkr2/H+palimRu7eB+tnk2WrX+gKTXHcy5VwXzt0r4+ZCG1+tjzF7zmes8
fYpYZiSSyMmX/8G6reewkWEcOwM1skFL7dUYQ3J1R0SwRzT/4lO3a3veXMfOWJEAWW/YbSZ+JcRv
CMZJ4Rv6PMtz4Nffa9qSafiReurxnEoijSBy6cPWVDWEALHfjm4DlxWGpil21scHtg3niuDFszCo
oCCRcusH6ggvF1+6H1/xmblMTuTouCb2scYJhI4s4tMSdRK+wQrc+i5aIDcQIs1xMiQCKcomnm40
3iwf/LfG+PiZFrd1JVaEHSz/veXADTo8htxSYveSykfh6aAetASbWJnLKJwbATYBxJ7IszL5MXCK
QMVayJ7hAG4owj8Bz8x0slCpRcqxWTfG/dysTVv0dD6510nWshbSa1jWTtIJl4qi0rAWDLo+6uzS
1ClVul9dIxdeu4peX3RU/UFlbrd2bHgiFjpK/CSbJBtFJRHDlefNRmQp63yA2x5hxwjzKigpBgpX
cU42Es0n+MWMUw/Jk2tkP4AhwcY72yKzwkzSSfvCVAiLu08DAoRVS2taGlCoIabwfOMxFJYuT/LQ
nCoiQh7uy62I9gVG0TfSQro8EsyttEjgF7BSPk7Rv2Pws3XIgwW1VFpD9f1LUq8Fyjm5va1wq2hM
OT81XSs0xGojhoVKoAmQdo4ZIeYM3cWv6Q+swWHc+BzEUZM+r8dKb52rSmyp2OEs+feZGHpl3Uog
M1T7BY1w3rilOpe1EHi4UB6FAftbCdzx1hqhQkfkXotshCd5NWNeX169pVujhCmtL3jCgjQ0h3VW
NqwDX7ubXMOrWyr7v/MIFYBUUTXw1MZdaRsb7YDBVz3H2DlF1X/cqND4cf9gUtKaGHNTCvX+d3G5
eLauMkdQN8mGGY6eVfubQ4D9Sy60vJJWWwv7M4LE2eJAnea+Pkz/DtmMXwahxDtPIx9Ih30iBHR/
iHfoyWrVfiIfE5qOFijwiFw3cQHWD6W/jukW1Yf00Z4fUTwLwb/iQ5Ln7++STQq/D/NBcNwRKUQi
kAG0MICwxLHSGvslihxzptxI2/7kX/u6uWS67dRJlajpF6GP6k5myYoass0dIgolE6bIhkVT5+U/
Xi50gJY3DWy1K8PSiduOtKqgKhreEVYC2DlqLnRlX17M0jQkCBo0QVUzyCSSkoziHcLv5mybDGcS
4XtO7Lp4101mT1HKN1xrshM/jaqJWLGVEemq1CvtzIf8h8cnYNjFKJ0ovCZldUmjGoktDoxg4fJf
ndb5PopN48LcqTHDdeODr53Txc7UXzRMnEQXya6bAh6oSVWtapqeWBEgNNE+eBkCx45Q5v0jF1ks
P19KE+qaGdzsxZiYNJ07lyxFit81WReZocMetdvtTyoAItMPNuy3v8nIxCnREXmr1WImN+1FBoCW
X/oq+sp00ExT/+JXAFHkjdOUDdZU9RkuAeDb/3BdKueyKgGfdZXmY6G4TwLNGRih0bediIEyvl9b
WD4GuLucKB4ry1ATT59XBIOhqI+7tnExcwirmxUQxmHwk7kMB0hG3eRY/JUErdKbw6a5fq57B5/5
OsvlK27rinmSikVVqbvYDe+JDfkeh7qY0R1oBWiD6lZLXxyxhvfZCWOzDJmztGQHTbZ0d7H1LR/J
NRf3HOW/AAZORrhvWrCXfXFRyT3Rfak0X4sN832y0xrHoFSl+uOe7Dkn8Sevse3Tme/nZpNIBVC/
P93Ktt0h5dPOlvBKNf2molCouc2gO+bqWU9GdoJqV6flFzD/AdfsWvVn5SaJoxyT6iu961GuVP36
EGRTbPmW+p3oxz6NYSno1TPRdEwIdmJbNMjgfqi4qOnHwZNBq3W8yfQl150ONUqS/r8CG60b4zV5
3XjOgpuH4OAxxdXbBzV3Dhp56Ii69YLpaD3n19cNs8TlQlGZwHUZoE7L+jmk27ZyNZEeZmpED8yK
7eKY+Mjj/Blxl7wo/aE1IRFDeOxKIlvz+m5T/Iwzgw27XwyDFwWppK/PVpZZnhpf9xhBDGmr3wlS
+a680GE3PbLmsJgQjWSVcwZlxa5Cd412d1qWLXebQGinaciossWiZsXImEJVzjLTMXV2FHMVl676
lYPoU/uiS068pgQoUcuRo3UfjgwlBcWJRWgcVxd9hZw9ItmRM+1VmQInPHv68/iWZWsqx/I/CZoa
BzU5Vg9Qx4TpnfEkFhSb0MmbtQnwekzCv6DFQFXo7Yog9w+j+C8ceUJkTamqlMc/XYfJLLEZeWn4
PfNH1DXHupwFQVoW14ScuTnLhOL34NSrOttyqyJxlpiPpS89n8XvklhdQMJ+m9rDUBxEbFsDpIPI
0dEa+zcsaE65LRDWZrQu2/9y3QAoarfHFDotL52R54E+VuEjUgEcyEo9hJAu25QBWIe36daPMruT
Zfhz7rL1DBnbNeoEbwpwYnD1QPApTSjxmp+MQCMUb3cQ0KsDb9mQSAZ+09bz/vdoqcyIB/Se7beM
OOuZavBvQ7QIk2/NbaatzcoW/Cvz2oy3CG2aIULUQtsooAsGABEJWDmyYg8Qwb0iMHFUG7f/DKBP
vPlX466PXDX2K8XJ/mBFk9igYGzckTNQJRHjZC6NO0E0ZTgak3N8eA2xh6FeZ8F99HQJtLlH/PqV
BudbYWqf2bMDPJ/K4AA8H3EIoiUnZKa8w64eQ7or8oaTmLnHwqeuUUrctUV33SwOpsW9oPVHDoYH
4EGTqQps3KETNiqpoPEeX18v6OtBcxeOusBwHXggaJBapBP61j5ugmRumC45MZpsfSs1oSh/3oqs
8MLJulubFrPMMnnlL4YsxciiT2WjEMVeR4bhM4V3PB2NeKQqQWUiY4u2KkyLGYPOoQdSv2Yaj4ZE
NjSfQtilXq+BpUhDHPdeZqFUMktVWO0/up2/yiy5u4TBJQ+XAnvEawWGDrarVipkHFEvtnWOpF1c
QF0ATSe4iZDMpZ0gKoyFDzBnNNqfxUlH1emjd4tc/h5gOVhCeXRUtdR4qFRUTcrU509AV4xiiIZd
VISrRQRPEUY/eojHdy/DHWlwHN4h98gHwvv/ItbAP7uzJ+zDvj7N4krS77Umb73JXnvDizxUh6gu
DKVhrJbR5Ulg8DC4TRshaJUKudFKj+SrMpDakhwAn5vYhbfdu/QJFGlNFOQTefIXmnaI6/U0DcdC
0JoHBykUrQ/PFMXkDnhyF0ex/eTuDOGXxy57R7r9Cdu09Sra3mq955KgNFa158GhW+XeYWV69gQ/
fSLXN6J9qwk+7d4gnLZsNIJR/jMaSYBMEJKCk5ysE4K6TTMR9vLFKQr+Ybf+5KWKitYaQJ1T6F/2
FFg3YOH3wmifjrdS1CUDM0lkQuY6cIuPVL6fuZ5d6Y4EjXNIufDse+UhXs5u7I733gGkflL5vZoO
a75ZQm7kmujChwrpBLDX9W6IhOvzsoBkWRSCbdGdp6ObwIl7pTGx2TotiPwnPku3S0YmwR/c7bDW
Cr+N7cuqfVQJNWLy1L6zXotcG4pJP7+x12vJ0yOgbndq2Jn4Yt3q+ZgkWN1sdHl0B95ZfFe7ukEI
B5B9m5jggpNWVdbN3AjQwU4zNnxKJStm9DEJuLjHpxnUmTAzUgsnSZOqK2ztf/SBvvESblWW4KOx
XqFOBI00/X52nmtOZQh1i/KJLq1/3BzG3hSpO0xlY+ZwnwuSoQNrZQnlbBwgXqN3M2Y7GjWWS+AH
vJyfEZHIwqqSf7fbNN7lRr3NAfApXxq2OP/02pszU+955etDoeZC32Lb/+raCzfLqik7yadbDtMu
w4/sjiVjjFKl9i5XqIPUObib1ZkRQ0DjbYoddZb+i4SaPm6brdcicG1PiKSSLYP9B58ceawq2IZ/
qI70leez0peqL+PGLKhrfpMqdQQOZLtOE70NpkYCXcm63SQVoAf5h1kUt3ocU+RhOkEy+VfQ5g06
P48f0gbgefL++4CSvqe6ICWYMklJzqRy9SmJL2hEqsD9MwsXPGacKEIlQLgwJ1FRzZSdnAJCSkeD
EyZK6QFqKzJsOxZG7990UF84Y3t69zhg//roJpgkwVL9nnsjcpKuTERn17a2BPTtJwGD3kJLl9+F
i1lu4Bbl2y/6H6Q3m8Mmp0C4s4M7eNc8E78hJvKKyBIRYMOkqn8fCDtOMG5UARpyDH97SB93l1f6
+lOP1kETAHLGowWG2ShCKhxF7Xh6R/VIUaszLNZbixjNfz8iCrQLRkif1yKg/nDJljz+nfnBb2ph
vZdkMEFcX6j2ldFDwDDBmypoMTby0zIn3qQBFG1Mp8dB6nQmkM3A2DnErdzriimMizoh/1LOwxYY
H0/Ovg4FkbGZXJaCIXyKqkoLZczpx9MWWw7rVfqfAoJAvadzA4hpS/Jq9bdHp5jyVzTmzyUFvq7M
m6YCiuVbxXxWblmCq/b+/cAJ71GjTaqHDbaDMovCUT0suaSCZ3A3ZvOhJG+A3G+WlSoHudGpUZEr
Gri9wqxlEgIu8He3COt47dV7dyW1qzr+G4QB5+tX8ys18kNwHVCVSFJayHt7crrpbkXJOYnS340F
lQfvi609HbpECdtAxP0ENtuEfecyiH6WVvXTU0KzpsXWk6c9ihWhmK3c/LRFVweV/iiboRxmdrf/
lzQDK2oz2AT1N0xHq55wKbaKRWvKnfBoHCdMeQ6xGMWevREQ9yAidZmtuRhL/OTcERY4+PuPM5Cn
bmrw3XqLw5rfOdsDgq3fL2W1MkNoRDWD3P2mUgJeTtp9fkksh3yGXEjRuuHJVqmDxop7xMBIpYaG
+DqvX2No99G3BWaRt5odfPevTh8tZjvfolvReDjADKf4LTGftzO7TFBsC6VHFfkaoxv+XvVwn6eD
iFCN6qtPCf+CDus/D6u+5moLxwfyw94w3ISPxqAz5G7UQOBDgDpV6NrB8g9RdSicYU5lbJp4CMDM
xHUtWO30RrxtmRBjrt9ejkCg5iRNaoRwikCu4WCE+IBwU3nPYbGVKy1Gwf/ReJ25PeeLe3569mil
ZcbXiuTcwyXHgXbLaLnDmAjI5Xj583+c8TF1VXDqRT2MB/e8PbH2JaYe3ROqO64xO1h+lDbNJzJ4
7rGrXlur87+8GFQ/Lqukkhm6F/bhiwrhNa8jrcrVSb7zbzIJMIYsHSRjKpIHN7h6BrvoAUkgv22D
zdMQfD9yepfPpxIPGOOkr/KpIgrVyq4454vbHxIvFRxyL2G8vjPW9sLNdzctot+rBLBpj5daG2Iu
fUVHYpcF3zNCfjLVHpTb9PjxJp6W7UPkoN27wxibG/+p5DFDjGfAhAr79CGmNAbMqza9x38ibnbA
98/r8A29QUW/AIphKvXzynQ6FOCcwVusWjf9UREo+Wz8Icdj7MDFcvYObur50mcNBA71Bo1B9r4w
/Qd0TKVyapmkPAhP1RB88WcM8VfspaTC21cacyV4QbPlsN+ki4iyrrFtKDScX08LNvhDMVRjvKxJ
hprWPLSIkNCvzFCG89Dkg8p5TXbaIAd032X8h31DH7oEGPhbfPHf1sLdj+sBY4BcpPGlzx+EPSpL
Vr8Dxxd8rMbB7amuUrBncgBMKEnC4TkuPlnXCQOBzZI0edsicLm0RyiRrrdbDGL4woeTQ5ERgwtq
Az80vBkodXUgFITEbR9O91iuNEoePwat3ZtmFJHAW/sgAeWzcMa8MP6e76xHKobs6YqHLSb/YaMY
p+/iZipTpafc8HHXZ1voeqsJFeVMZaw1KLdrxaoVm9XPsAT4admBu8wTVWm2Q/SmRM3/zswvOHp8
SZ2k16l8nc83aR1lWmf+Vcv4eZQCeEdZ9D1uC2Nl8P5/77HjNw4bjSHHOk83rySzPkLRXfKAiZe+
++SxbGuco/oS4tML4Xv3j/4JzAOMEpx1P3N+4MVmdMwKBKOq3pEiNRuUJRd9MeEdmdxR9mkNwv2Q
QQAGuAojvi2t2X4AxEoHr3Ns/k1vI2WuF27MYKFQQdChabfmAA/MLqir7zHVMxEPeX16gPdPXxxm
/odPV0iH4r6leqL5/fDUSUS0M7iCTj08DnyvwXo1ubPg1Whzk78vTuY0S62q54HKnjyHcuoXMxSr
H23RJJpY5nCLEQmPmW8VR20PXDV0/zaRf7kJrBTUkZxaLPVH+uVUU16fPx9ZDP7lM9IqQF4i/8pk
z0u8hX/HtsfBQk4m22cieKW1SxOU2LrctodGmYul6f6LpVY7h42edfPfjLg8ne6ysHF1QVZJYVe+
UViPUQBzy3+9AT60Eje4jyjjWtzbHA8q+pyTb3f6L7Tqw4M6QgIaMyqv7GuU5OcBYGP+Ab5ZLLFz
NKYXZN4vU0ai9MTENdwTNmznb1vQCB+9vZbqu5nkKym0vjd7YNnpyipOqaNFPDOh2eYgJs8ksfSt
gzQ8l17bkyGKLDhIxl6MNXkLc0Vxl7uXDe+ZAvMqXbESgQkCuJ7Q7gUATRNzIF9Di3VcG3s8EtUe
GtDPo5AlZ4zvMx7sdx1PtDio/qCqADCmc/WD0Ejjqz6BaElVmHY7J/G8lCPz25wviWCxfjBasp5b
ygWUse1gUqdpP1jzzXvQVrbRAaCuPL3/Rws8QWmZc8RRsmQWIfVvOLmG9ES2ft+n1qTj4HSUFt8l
kGH6sMCB3fz8HhXyNfq6tbeRSoK/BSIcKAURdNzno38mG4cD4hMmSQZBV3rcvs2WufUNYoFspV8d
AyCSD2nursYIlBYYtOrlhBtgo1wfoi6HiLhBFEEL3wz61qPl8bsFJqgRyzYNWj82+fkRk9FzUJMp
pQLklSXCAU25reY4tSP0d0T9/Drx9/Sbq8o9vbLrufrcc9CmCM5VG3DcMQrXdBzQLzFyIZyNiQZ3
VNqz9hz/4k6FbmFBANulrR+IJuSfLTv8MMeNuJ4KURqt3JwZ1ExVZCTT2g9iHaCehF/JSfbDouNZ
kvq0BSPbu4rEbr6Eb8Aq9XPxmfUFFLiBezQtWfCokQb4XomkVJqLEY4L79ipl8jo8IrtDTnsDPYm
6uaXYIF1+3EzeXU+ZH6jEt7Cy/PjGu/Idowr4oDnj/3Y5olncUXh1DKT8RF3ltq2+5Ehjgsx9U+2
YlR7GYhSmouXzwN+iSUav0FsvpxUmYyzoIZl7epeQgfHABUlcdyAYi0fn7+OnC5Hw64OkU4qGY1D
bYsUD6cBUQSIZWXnb/sFK+/iUdI9oVDugqnekXYfA2Iz0ntZZsDQPpwMjSpGaQcrjRMuMIZbyi4Q
dd9AOIl3i/gGCtkaxyMmN9+TdRythXA46DINpyrX8EsECrsEd5B3IbumhOH1gNqjjWPHEVDdbhYZ
xEzamqmDDQ9wskx7ZXbMAJkPB7XSuYIaWUtQy6LTCrolLTv15DO9VOyYYtngB+uQSGo1H0JXDEcl
C6h4LVEuGEJqxRW8RZBSy27SQ1agXUMqUAC/S8+cBcbA0JY4IIltWH6njYKVDrk8V4S4Jr3YK36J
olEmtdgYg300gjd2d9zVc9P4yRLZxMZj7kwtkVyihFz+thAc439tuth2e7zdpQvilg/s1ApxGMHC
uysBMQcro2bnrr/2dExFZ/xsp4bvShx9VGmVxXnGIpwzJhpfDcr1aa/1y9iJT8Vt1Rt+/8isAuL6
LuoytjsC1WJr4SeO8wRlieuDuMa1LLoMMmXRvDI8tN+3vSXYxH2rP7eqKWStNU+NCsNsTi8zB8Et
diUNXBwOMO1mgIe3Br1oM7lm216nKMJvb4pu59GF6CH2ItsD54kynqiXwhOTLO4U4DgIYG8n7QkY
h82I5bkHbD9ED7RJoi8lu4g+l/5yezrrnN+nCjRVtZ9BP7OzogEj8VreK2krpkt+MAGBF8yYPdiL
g/r0EdkEnVhAkKQRGqM2xhWAuRyjIdQlxWtPrDFwD0taSSbBG+ZCwht9hVHOjPrLgkigWz1nXi09
olftvRaEnBonLjaLdoDRjfLrMrKfuftCjtDkfrTENBYex3IU7Rj8827IQ3BXDoTNPGWdQUnO4Rj3
WctoVRpkchl/vv9f3X7TLMvGnJWsR598NoQEcN25VEXySPAV2sMJqyORIptongapMCQ6ubegp0Jh
wpWons92ZYIvwANksgquwk7a4jUWOzDQ/ZORWY7mkvthw3l466k0tvMbvOFpoQTeStwSAJnp4hMZ
eE26OSgXYA+2UFe3KuK4oK6BqJ8ucvvFzLmYy+Y9hfN/o6KvV5cg76Ak8RssBw2xHBfcmKLZ+1y8
YHVxadH4UYO3mtP0bDvlJmeKsZ4vdPJERTmtPFiODLMQCNZ2bZzL5avq9BgzbqywXjLR2SbQ8+uN
wHUSUMRL4N+Sn2rqe9QnhJyg8HJfLsGlhciazEzL/D8zTKdY+SzJSvV9F9rgIIWGs3vE5sfAUlMc
MV31Ixhz6WR0ztgCKD5JWDH2IpdP8Q8jfaEy5u3SZFVXaD1EKvIjNVgQagbEh9LNJMtB2Zk9rEoC
whPsMVW5huOw6yHdnwQOheyQx1mXXqUwjQ1zvwtxO0nZxlIjAo0VERnQXdRCJHWcVPYqzqsCDOsh
R5aN3t1KDOlqrEQGtm3gGUmbKB0Wu+1VlpjWiWEh+HVVpyxWiHUfyyxMaB77rJux9nJvhLAmFqFI
xJDweBIsgsdPEsSZP4KzK8y+C/mQhlSpoHvbaZPMj8Ijdzykzix1tKvG5XIZMpKTk4Ywh0H/353i
uMGkU4xEkKZcAMIZJ7KXJFqhxwgK+x1osK/tkOhDOUCUckttbXgUDedoUZN5rEpJxAfWSmE9u4sV
qaeMDZXtvCQcWlGR/YpzOg3r0QEgKaoauLNAMTbDYs2hXR3UG8B3ScJw9WavGxu+oiTFtupjyXJy
h1OGF6brBlxgkKGcHCw5RVzICGuH2eLShOzrjmtRakTam7G0ZhEPn+YhZ8OeUaQIVMAYc6nkF2tN
ZeDqhQHkgeCFIn0hxj7FWu1iR7qWpuRpGoV5MaVog+N874Fh8vy++K8Nu8sYpQF4UoqPy138khWH
Ikl2V8uf+HwGqy3mUy+S6d8Vgzg2fzDpmvSLz/JuQd3KhCFKG4rvO6oJFEGBvYopHL32MU0lpeC+
8IySd0sKc4lae3/imvTFueXz1Sc8S6wqemSnQMPwkdXLKhxegnovcuzA4BHHYwlExqKZVF7kUh+g
Ce/6CK4Vx18P6qUmF6WzF+5gLuxqZb06UR98JhxDQhXxJFYfeCk49cO67g32hhdzqKws6vVrq6MA
mTAyKUJAtdVdQxQGxcCuY8Mzbhk9TXCnSYNpH/DyvM3y2Uzx4VS/ZUMg2D5b8Oq/A5egLN1UxUbB
uiyv7rsxByHcZp7vp82u9PDw0by89jBSXN93zQO+CwNatEKWXSAcEXgf+a+OqbB6dZEgsxy1sxTj
81A8jHbpOCVfXPVndo6pqb5JesDPl6ykjEZCxmwJ70fXB65HqHo8BFL4+Ub+ThO2unVoUhFE7CD9
l4BjUfFq6/GbsAcHTcRKZ/NmUx7PwRM2Q8p4ALK6i7q1zlxGaGZuFW8B5FiLvWEnonpMSLG0zfg0
LZsF/yswf2GL/U7Uyt1jGJ8bNaryDFr2BXf+brws+s12tchmHKAJn71BtS4H+pZVeexyLKug25YN
Uq8aO4xGA+YwyfGGqP2IkdiZ3GT18++QejSIFzXrnjtQI8z6EnKUbGuz6wbEPg8TRal0Tw+SQ60e
HpI3+LNQrn7/U1NhezviT75jerlhw+liIvUXJC4l48a79eNYBwz/LQG1HP3mitELFbAGO2FgXfTo
UktPFtjkdMEm8I4EFkeIqXOxAQNxy0azbxMHdCc2J6xgNMfS1042epKupkmeJu9BehIoNyBkhZXe
ES5iuzLvKBCsOwgGNbpS1o/yxhv9EzYo8onolQgYvWIxAZ79YjVtyKaMqofydkxkwm/u9nzA8gb1
fE3h+M0ZPKz5xe+misAXN1hQA1zHnqy0Bppp9x2I4Qpm7qKKbJ5m2rJqQClx8wkww9bIRbbwmXlB
nzKEwoDHnjMbLT39lFaerELHkn9He8QwLrArB/QR7YUTodSok/Zwn5WePYWw99IPBrrZbhhztgyN
4OAA8242aPOStEbukfTLv3IGF7g5A/9KcMKJ2GPXxkzpYOZBGQ3aHj8ykjEOB2IJPfKfzLRW6a7/
7NtuPyeUIFLVoM4xcmGUiOKceo9iiKACyaazOuoqe11ssUJIaGek6VLihg6MAZhDF/9m7ulLuR9K
YVKxPm4sR2DoXyzEiIXoscW7/Pn2yxaWch1u3v5kHHCI7gUU7a12RWV+ddvD4KjXOplNFL6N9GXS
r1Pv3zbZoqS96XqTT7BECWlcGpB8iaX99qhKeGsIqzNQjnahrlg7nz3/Na5m5yF08VfBxbcJn+wA
4tm3HoungGfJUxdMrl1BscQ0YBRhSfKEhoU8paSM87W6Jd7VCQimqX+CgBoo+wNDBb0vCR5aqjyQ
0DDvleSd1vS0N//561vyuOX0yIeeegyGYJ/3SgPpqAZbhHbYly7pc5xrUSRgaToyLm++g7xb4NAN
rEQILyY+oyPld5I37EP5eSJRnjXM8u/ZAAl45ukfjgq1PJOCoPqZCE6n/2cEjR+azHR1d9n4EXbu
lU2q1lusLg22krme0uxF9joXqZyqrn2WGYZgwu+snMJPfaMBDSf+JGyrvw1vpQOheZoNinAobc8n
1TDLgNah8rRk/N1chXMAFuJIpJlY0gFpCPwtEXcS0/BzXZRAimqN4hGK1m8P2Xm7nEQh2uPaPGSM
ytPUM8P92MHL6UehNq4gKQizweoZv6PPF2kQsiUe0wnqL74qC8odV4141thBO5FqY7ZZQGhkXM6a
mYvhzASnT0gjNzccIVisIWRE6ZAKJFlcxlFCCDir2FkTSbQUhghWuXjRHNG724vx/7/d52L1m9cE
FesxBtdcL6VvTsK4YP1np5Ut8uttG85VZuef83aNmv4N0E6moJ0ZqzFjgueZexaHnYOoSt5Ofjhj
iIMLohgQ9nqKkVYk44+ubrT0eSi3u8/uYP071qSmQoKMDLHyVzD4+SXcbI/fOpuE4SwkTmFWIgsa
uBHAbt/i12fbleNKwAf6z5/odlYElKtBGagjIDIGJcUZxt2EtRazKqXvkcOkysir9QFV9XDHyo7T
JhG5IDFYpxXC+GDkd3YYh/yl48swZZbANByXIFMbZKMvVj6h8YlqVSZ/mlN9FxwGAyFJ3mLgzX2v
LbSeVhS0+kSoc4HpEbR2M0et+5XQVsPNhrFHSEcg1upJfb29tgP8WOis56bTqzElZgXcNCcmth/E
42ke/XSPw0tFlJBzjE4o4axwxYoX7tAiMbPDOGx6sHo2HbsZECtGx4MkWoCujHcuyEcbExKlnFPg
MoeYIFuXE8SgCnAvyZUwyD4B7pEcmJ8xs8bsXPCq+qEWse2ncRnvJzAsAAF0on5zzm7vby91GZdg
/mOeMDt+oORfOIA9Cq5ocf4IziHNVn9l8vTUJ3142FYEqOYhbLpMh5ibxitjBbmTgeSgeq52CW6i
WMXtmqWrM8w6OtSBRr/q8x3fXeJ9TtPoYVlhN4umoE/sTGUH7CdreRC+JcI9Pbm406/b3Fb0UGck
rePgJ4bvv5lPf7Uvys8rbPDBgrjinGzijnDxoKbypUKLpoX0apgYa6wPIzJIsPIYUAmmTLwt9iN1
n9gRf3CJCg+M9Ew/LcFvy5e6IosN8cI4BnI4O13da93JpztMnr47aIp+7AuLusx8gPSqh74dwqC6
fpecuIlxIccZgXZZLga6Jwv+GqUckK5zo+eZn8Z4IiYIt+TLKjIQ0VQK7qd5/SpEJjJaKx4ERtVE
fKrdzxAXU+/je+/TTs19oOUZ4k39JW7Kdl3xx5DJLT071wSAIdZRUz/goPREjkf9TezaVuJazmFQ
r9UqeCxlc+b6H7NJxd5GeRmRLBYkEAX35c9LAgGmjEkv5/g/EDo1ITcze/7JWhRbQHbLMaIDh4r0
0yMVBCHDIELpCOdm+R2U94QELKTg6eZ205bLE5IcCUZCbdSFe663fWKWES3YONa750IjK+0iiImD
Xk/jOQLtjED1nPE0GE3ZLDExfZmrLrJ2MdnMumBzt9FHXDWP/3ZrpzYHLM8xcmg6Z7NZOSQ4bmQv
03jxvDvwO71lIkuDGKtHG05OYTL0SO23LenD8JbGD2Moq5/q+RHVVP4soPKKF14DNtoNdW4oF1Qp
ZTemMcTrr5xI0cllOglv3FE8mp1vzUhnLM0XOmFlgXBKICwFMjFCOqIbz0TS6R3ldo46ju1lmB2X
VUDw58k5GY14wJ9R/uJJYRbPumHH7xR+ORt1hUuLLK8rLcIP7dei9rkSAOMb81g38ofGzh0sp5Wq
9z8s3AGF5xeOv7YZsWM1TIRyK15OTnrRyF/5zQeuRzl1NsuU5XO3Hvwk49yMAulJ8IAje/Y64B5f
kzWyTcWBXHzzKqzQtfih3ht/P1rFLBbxeyHwvHOJ8mOGMoLCykresiXUX831w/dp5i/RpIH5wqR4
kbzS3dnKEzz79lmMFniSro8m0Zqbz/v2LKT++xnYCoQdBhNsWoycl2NGAEwgSMt0BkveLX91CX23
Z6e6AELEfY0ymKJ/7fKdY85kf4ypdbeAipeQd6yATiMLGrwtDQ/18753Sj7waSZHeNj8nVuKbuhF
DAKgbxOtK8l8njELLyQEFK/jDT/EKUtMfmWQKy4yCt0moWFE0mL3jzf6vMBbIWcr/xvte/OsLUKo
/ieGQL7xgCKpvpFM21HXtFK2W/q01vxqsyu0qUpTyTUrUYxaZ85Y8/Y7xBkMLuN40NNHVx2iqWCv
k6OhCx1oXpGVFidooc+K1lceZ+E8Y1UjYSCxGfWBLt5DWJX5/p00YiXLidYrbGxIyz7UOJ0FfEfW
OtU2IeMUGRnTeyrv9hZcrH0l6v/X+9RbKP/fr94fiM6BlzWp4V5ucZKc7H3f9NYWnCvFrq2tXkdb
63idf9P2QFhJIvg/zSUX09rDbXlT1VWBebyDy9GgHJ54UrwAlg7mG70M188dqSiMpEhVwh/20ifb
nU71U5WEgd+VK9usT3liGVQlL4igg9PPj0B589+yqkVFdNtkmuxJswoA/M8/RtnrO2GDGbvtOZJl
4ueebfeWINXgp5hRwSg/7qB0mpndRj6EoZ/saOb/K554WOkBzXVbYEYGt3Gp/4DNet7AYkJXQLDP
D6DIQ4MYWhrQiV13ZdwLp/0wkqx2P4/RQi+PKUlXrKHAHdgaSyJL6/yTMvEz+fTAjDKAGlAl5wnp
9Is19VCB/7bLL0jGoQRzk+7uuDm4JrYpV3XBEL0QIbmzZNKH1nxwPG/daXENr5jO1SkTgsQDqjA+
xLOK/TkNMs5N1Dc2zWQzjiuSVyxN79JoYwa3RkcPZasATL5OBl++gDN4RyvrVa08MFUw+yRyqb0J
2Go9JrcgsIjEu43qNluhKGcEo81pJJKtcJfE8MRiWL4PGgCZ8+j7p8/h9JKVgL1fUhQ3BDYIDcIG
dSdyLJvXfGsJ1i2YK8Y9ulTugop4hzcDYMmpeST4b3crl02As8G09xw8EYsZQlp1XEqOGhnhkUde
51u22EDdsujxe9+13hoAW2TYrC6VoBt2sq5YwseD8EW/vXLsvPKwCOpqEB7BLB36S7b36RghTBnY
gDsvPe2wHoA/iCIYo7MgNHtiwvoXdZ4r37UkkB/fixuXTzGw5p3xEQgY3IG9cYhNZ0Ax3BYYc2x6
uj2uvfKnLM4/L6LT5FbfMg7M9EGSbgcTeOBaCoGWeC+lBHn42TxyIvVJ0TE0NgOX9ZtjsHIfB2MX
knLr1i31RaoZ8lGVV/8G+qh/f+50Xedt+zTDZcFpXT66TVoOdybVI2ulBVISxlt90DxyEutaYduC
Q6zH2R9ZKLLfNsV37UqWtySN/esjzTesyaBeu5Wp/HOITFtzIGFaF0N04BhVzmuUyoEMS62knFlP
GgLEmM7oelB9grqZ+7Zr3rZdBPetpbF6SmX94/HhXP4VLNraomrMk2ULku+eBXEHO3rbePoUhp6S
crmvoIFneBd+xvq6KyYUBxG7GxoQX6+rLM+1aOOIkU8nbBM5C8IR5GlfncN8H/NfpW4PK72CKnYA
iK/uUkOz1iR39qDga2DU1ZekxqSjIvNgF9DU5tthI9z9qCayJQ1EroCHGF6HhF3JKaSJQljfW7LM
hKLQjbw2w4c6ZTgfXLGAeaF0c60+kEVM05OK5vUADcDIb1BWhidqntmggsXszVP7uc6/fSIvgnt1
qprU1pavIW3q4sXhfa3igovIFGrgRYLZltZ8gEiR849TrhmjeUYXeVlullhdspDI6LFv6l0Po9IB
9iuoA6EpDi2riz5+CmIh68+cEnnGe+7R2h78TDjHQaDCrKPC2cA5/nWXXroCO8yV8/VEFvNpTZ4m
GmM5YlAgKSBuLa/s62YO1OW72Vce9hPOPf5OxiN91PKSyp5Wg6IR/1BbYHFc855eTT7snFvY7w5f
aaq4F5Noc6bJ7M+tFqhMVIrRJspxVV5Z4Iytn/DEfpiRKKRpQYK0iSAZSDa8DvwMyW56kxdtDSCu
mcXtrKKcMgTQDp+/4W8zqe09SUIEpSJL3ufKiv4Gr8NRmFuuSvjLHEUOrnVSoqluRw4I4Pi0n8Ip
PMCxkXrBIZnxNQL5qzFw04IrHILfpoZELJDoemIXEy45OtF7Nt84ONufhP0ML1SheF7QGVE4B90N
c+xk1fhGIv9bA3wb8O83mBMuczA9IEYD24HuwR5rdYWcOirK3yc+RHPcn2NJ93CT2RKRqNMFJ2V2
M3N5mNBiQjFw9U+vxtJTVey/7aMPpr8EB30cK9NPTlklOsiAdmmeqERZfe47DipSqYZRCua08Zxd
CoYZfixEvf8JWmHzIgdavmvcyvVZ7G7BrnqfQuNgZ6EcK6g/aqErjOCHj3kfX74cm8ND2l8t/jWu
XWDDtaHbRglM26+XoKmPbwrFKz3z8uSK8A4HafGiers0E59yWAzzPuJPdtbybzMr5zk7Rvg8RaEo
RPRVDYET2ESX41KeepB1zw8teEKok/juiRB6/h4zs9YNil3qYacoaamqjzeHKkxSX6mGxf+6X0Uj
75+5sg+Kb1YlP2Cj+JvctlWAoEdiQ7HCo7CKCjA5uBJ4VHseLVqB2/qTaH4q+VG4w18CvjN9aVWU
Ey4gvaWgyYOk65wbDDwYYFPARWHBkmpi2uZ5EjbIWscfm3GwbdwN2Y5drVAphqPBIHoSPIQjjznY
sBatWIu/QE+r9oeBXk262XXs6o8qsLPKEatdzGR8UA1VcgwUJTFIyymrKZDV77LGBJD34AZ1mb9B
W0HVnvv5lulJgRcL5VJmgjWFTBj2JAq23IJpBYsqCb+ZfIk1xJ4jhLpJFATIrG6btgNSgWFipnMg
hwQ2gUlPb8zzEIVsBj4JmZErWEcy0eEpDEoDLTUqhECxuPi3hKIyeKE0OB7jCbNzVS+GzOwl8A6I
jF41cR5NZVPAcZiVzOSaT5mPodD4NjOeiucjN0e0eSYzSQrVpElGP4HsDei182mDUHgs7SixCFtz
FTDXhvZIx6pntiskzmAP8xPKoWbTCSigJ2WVlCXLauRYpdWFmwNWtZm0klVCciZbRLdyoJiNkw/L
5c+7VY20PaZqmkXG2hegLaBolXpzZQjeT5DFnhYKQhJswbZS6Fy7L1UO6SsRHM6Lf92neWNydDIo
LchtSh7JdEk1z50CAgt5ln6l7FM+JAc8pDQI6KOteg83rYIIlvXA6hDciuuiJDMK56IsMR1FijxP
XOmaou0UZVEwIJOp+on0Aq8wUs+QzMHmI35pMx4UDkbN8UHQji/9tSybnTG870VfzC+FUjcoOT7i
tFFl7MyAImjc4+K3dGCRXOFjeLS1Ql946INextd0+xpMdxh1f9NMOpZwx1mov2sXOOyMobrzu5HQ
dFkF/d8hGX50zK9Uk77AlKFabAE4f1gAVib45YyfXJYPiOWklxkMgXWLgSRU9hF12OF8MXE8WA80
iQXNjKKtgvJxgRY0KFiMuMAOdhf6PAnrBo9Ivm+PTNLsZPahwuJBp0JRPY41XZmcfr6pZ2d24em9
YFmyd5uwViGVPF18C2E+rBTk33IAtwWLAXywYzVqT0xMT2ZIDFodQ49SuwN8mE1Eu6zRiWVoyKEw
rDyfQWzxTMTvNYwHaz2O/psK+q/eNDrQn7BhUQzdZlKIIM4n3Go6Jn26+eOhOrLnvMqrMRQ1Byak
ev6H5AOQ0c8M1o5MnsfSoYe84Xq7GvZVJr67Q8zQlryjMKf5tK5rhQBFCvFfuBg6si9Z4z5a20DP
jNLDnbetp8c7uwdPGIo0ExLRRlhMCxkpU4gz+kaBa8yUWo5Lp2J6Dhe6Wt/2CM3NS3xpYw+vi1Hs
D5EwpMhz5oMOBmYRDPuTwpCi+Aw14w+8g8NIJVBV2598TdW2YZ515BlTgXktIXzL0qvuk87cnGYE
i3UWYWNI+/cMPqx3k8KQcHZ2zqKoTb8N3VueuxuQ4J6wSMUtO2hi7kO29hdydswJo/BgR/owdyzk
dOwZGopQIG5KYPEu7uGU07LPEh0CaM3SDqNGTQZ9QbMTky9TbkKIc/f5iV2AimwLY4wwVQdakh4j
1g/X5tjBJj3UuTdX00Q0Nbp7wn0DNTwLTkZQ+knSBye9RwfNoID1pIgj5WhSmsTHxYv5wrWSBoH9
fv56hpyLPF+viMliq5vZ75GGjDYHnPai5l9GyTDc/TIDwo1wejnqTdGVKywrtxBp8XofuqQNze6i
J4LD1zmHg5w1k7C2Kw4uod6iugLHz9xV1nMPN63JZh4edoxIsG7LAbcOfkR0N2tXRMhqhekwn+mP
5NWo67VpOa/HhNMV0BLbfFfVO1QlunguaGYI60YG4oovqWg6x9m3G9ovCbDHT1fNdMihdlSjEmIp
1ca/dOWftfc1V8srzzxTFcrMsnfthqSBLi70p1AnfBkYEzL2Tvf8YsqT2J1i7tzeGoqs23CE4dpa
ygBaDTqAVjS+FBmD1poaSD4AdU+j7UBriuHMXQe23XPWc9FmrNtzWSVtbP5zqy3/2Tk5k2DIDvih
FpjP6il3p1tTN94bJkotPg7P4UciLHXa3sFoPP4U4MXMM+uz6s/kcS9+T9bN843GtEKsgej+v54k
Bjonj+QI1cjQcZ6KbWJYqlUBlBn8SdJanZikbheURVlISJPh8IpG15uDIyQbpz6GzxCY2/+qMmXi
ia8Rr159eIvo7oDxuDtfMw5qiS+gYxh/v/0XJXenkHZhljuYq9yZB2GMKNjKxswVk57XWdF8Xkef
4OUiB5Mz07ZPTudJD35K+QwLA6f5sTfQWBR8L1FtRPOUEYcE10EyVYgVIIhTWQ+sReGpEQR1TIXj
g32DXBJmbwOoFRNEvlxa6A/F2LuDvH9OztF+HwB670aMlHXZ8ThJ7tnU/W6SJ9PdT7mmXBBY9/v0
b4MnKSRUCKjwpm6d2YjiY1aUWjqcpCoj1aMx3aC0ec6sYhtkCqUgD9UlSVObULynkef7swivtsTO
EZxUEOK0MfjkXfKy6Em5EfMSGbGGmeWaSLdNR59hiW8Udt3WUjlDlBUqzffd4T135Pw0HROLNnd1
KGHI9o8mc6v7/Hv+b1XxQkQnw/cMYuOHCKx7ZbyqtgoRAajcInB4OJS096x2tFZ0cT9tpDTGuaGt
A+DzZY/YJZSdulHPBZGK/MIQscCJePvhtFFMIVPFYucsiWnVI4pphTIRvBE2zIb8JVnzXfw5mqwj
bN0vwm2vnFzPErvRxDvMJx3PEL1iGrbD/JCJdXUHeFIei7yZ9r87U+0Z04BVQBk8R64dTj4hEqQx
OoEE/lkAzaPPFzhD9jAvX/5jDSRWkhvwRPkOrAw1dp0uIqt7lma53KE25WLHWyXAVDEhbYsv7Qhf
KV6SzHPt0cezE+D2nywp4vY7xrm27P+xiDgUhhDA1/kol2rtJGvt9inoAUS2d9u6eUgBmKvkEgBq
jEst8AFR4m0NC+/2TMorBSnj3mSLZTIzDokq9ob7GYRr0bTGIDs7NVAu7kcUsCKVGguzR4vNfx68
TWhWaDR6LHNGRm3sE7XuzI4mHnI4wD0zI99kPqqBnqVhLHRrQSrC4ufld8D99oQc3jNPBhpgdJE8
BhLOUL6uV4v+lsdgK8d0fDvMAfMfg4h4DaCV9We4TQ8db987Y23LWv3PJ4xLpyPfS2S3iaKPpuOa
XpRXEatkmwhWacGUzutJfJr4MtlzJcO7WPgMc1X0nqZILDUYw0IgmbcYgotZPPd6DF70qgkoD/Ux
5xpaqz7eixN8ECf6oAGj3ib+c8hqc9XlG/DbDBvQEy9LiYSRnlZYglX0NDA40z3xUWlPYDPfbsko
C9TnDTKBGc87m7dWnzTOhxpnnqoxQpCvdw2lzGVe5Ok1MVhWN6D9WQbW5UqSPtJ4I6FN/rk8WFwH
PrSdQTTkF4uYHRhj4SFy5dGc0zxi59oUegJbc7z88xYJKOLX3AdH3crAcY1VmwJKfZLDkEq0C5tc
uQQof/KCiMCdT0drnv87zd1r9q2vq7EKDj1Lk0qo8MazvVbSuqT0qJ0PQAqmPg3fKBEtCv7WV8lg
HXLriP8++5xeiZFK6JVcifOeQ8lBbIGsrWIipZSL3XZff1FKlsT4Snu/I+5t+AYay7Ns6c5vnPDq
Tz+DQyfgLsWXhQ0DD0OWx4AZdOmB7AXs5Nxy3rCfo0sXm33ri3OKuR3Up9IRum7Cy6CGNI+yTu05
vC+1mz/Mly/UE3ErluEnl5G5vVe9uYZYF0DmIqLP/f5PSTPRddi1vlJKoiaKjS84SS7EfjvKWJE2
AXPCzTte8l/t1THH4YSCU/fRibQxFVkIgDi0wVjgTqgsDIkJ2pGy6umIMsBRQWHI+rkZEuYcvIgD
ng4uubWQsLBmEFagiMUII72jpDzySgHcZmvVWzfGJv/yqzKaZDHEv1RV0xtprTX4fLhVGR1S5xzS
se6565JxAmheJfpVly8x3Z/UmCJNpymQAAQJMR6gXEIwjWoAuHVLgxhVQdY8xLZ2hEbdk0kfWppx
Q/1BJ+R71xNi+CKo77fIhMw84p3YdUhcILBccWC3NNop4Z3c6qPzS+OzBAom2M2/HS6hQTDbq3ii
jYa0hBCS/G1NlXhrGgEHMOEJOdUmnLghecqkcSSxs5VUtfYV3/csbfOGj7wTGv0ZGnjX8vAip5VZ
/AV8KKCN+AEickwx++1YRB3NA+bNC7PymwEGDwKkaatYWIkSFAKlIyvt9eVMEpk5fPf0Yz/EfhMr
9girSZb7NISS5JAlo6A6/dHRTpww4p0/rSshs2zRqlxYAXxYDZ6mIEMdpSJbcaKuteBBhwSDuvqL
hSFO6m7Byuwqn6cQVkE+Xs10RPUZugM1UXM1ARoQ3bDR7SgHu+t5MOFpbaRgYwBu37hagvSK6Ydq
VoTCNmoBzbfnNjnGe3bYF5a0s9gVNQlFbm1iCixnX+cwIrf+dxHcsqs9tTJoOIYBmBhiYJh8BeqH
4qtGrynhYaf7ZlYSpznxtbcfDsIL2TLclhX8rfqfA1cN8AUVeAXZA+whsJftS7Xi/SgSrtQK4+Vx
ByiF1E3YhIobO3FmkL8lEtlqn3oOUXZo8A41ZPFkdHzl5nLXAz7VJSSq0IPPWn/VuvUWS8mghP71
X7i+BMlL7k2Nt7uqKgY1otSoa+hdhBLXB5IiUxMYLFJXIUFPjQ5Ya4KprFyuRsxL3MgJuYbAvLgZ
YkQmdT5a98yXCuq78sSTLd9sBlNxSbGJ4/RGcWFiotNeYbo07AOTfgAORasn6LUJtKKy3pLWcKFh
Nmxrc6vJ/VASAjVCrgRDM2jcsPiy2egoXiNR1vA5Jn7juMtMTJjIbhUCrEm7iYtc1Kj9R2Jkidet
VQnNajlC+VH7DxTd5MOD9yxedSG09bor0eZOiQF0kfA+6dHoNlbhKk2M7xyBBoCKVj/kqIL5XyB0
Ekv3AVR77YdbTi1HJ0gmwpg7hNBGTwLiIEmjT8Jliy1XJFTRxG6xRMKqA7jzHBYiCaF4zVbTcwuC
6ZgWFN/EA7lS1HMZZrWVc9lLF4mt+Tl2lbpmI9/qQ6W8/9WgmQPQPt9OrPx5Bt/kO5uWUMjhAhK2
m0N5EUHFuVrKrOypvGUuT0W+pLLWTqcH5hNQBEWU5R9kVSFU1xmXDCGlZ3tvebgoVnNjLB676ZGG
qp41yyAQr9+r0Ly4hH8xkS8kjCxelQUmaEHsHmWcL9dgIF0ioSQK03JUcKQaB7TohIXI30rJ0PVq
3dBpeQKvwM2S5JJE0zut5xmYJDetFpSjsjKBby9loW7E/urIZiWeZvk80qF5+aX/3QkSufkQOt5q
7E3D6pGifF1fITmlJBQzONuNfwIb6Q6sT1G475594rtqKFHKNhUDbFkLt86510KlJMj+Nh1vXyz0
gmKygVsVvj6hXROBiFhS1CgZge/3RXO0exNHOVD8cfhfIsegVBoW4HepX2uh5jSF8+TCFtrtwYv9
0ksOxeXF1Qe3EUlhCmlMkqHBN+nRqaMy02GQ0OvKnFgSLH9MW69SjIdMaV3SIBD+xpaqmQ4e0e2m
p6z57bx3tTbRMDssZrHXCa1jUqrHDrXooljdlzCZSy9ll/pnNPvps33Z6AhenRzyV+VafE3FHo2j
ythF9mvHblVWszwBbPKobBX1tgK1Tp/hCdCuMbgpAN6ChPd4FifWJnct7X8YK3I+sOCscDR6uzmc
hjGE8BdP/wL2mh/XgQV9yPOiDUnyAzmwKaVrXHc4hq71pvkKUdFkkXydwtMZxPXXi3L31IaX8we+
sRVsQdt0oS8g2VodsG7SZMPP8ItCMhgKDNcAFkH2M4QOuW9Xwj4WAfMEC5S3Uuu3e0K2/lIxeRyo
0K600weR/QQQ3OlHZbF+L3B4++REFpfX8gMxOc/oRF126Rcq+0erO6IRJ+jtqZZwH2ff+Pxq84Lc
nY0p+FLyCIQaHeWoP9uSQVV3x3c1BBSaMN4+xgIOhuAMrV3K2wrvyCcUoByui1KbFE2VwH1LkzMz
VbAvGiRISM9hGSSV8QsDK9+XjienkjOtM6+S2HFSUqytzXMhEtuF6e8VI96OhK/x+eytQaPwdhLV
+vQMnBiZMBfEofTD6UC2G9But5u3IepihfxOYUKx9NPKDWHQjyhOEEhQ3/VhuRgM6xGyQpoXN5Ny
1oNZ6RzXA/mvr3R/gJD3A8yj7FgKMUvozIO0agu5graIE55eWggmh6P55qARq6lin4MJ4A40rxmO
GNtKNG4913zawIVmpNGlmOHDFFpZzLPcLQRSdspxglqJa0d8r6aWDP5TUdA2XsbYxoRxt8Lo3+kN
m8HbldhHip4xEiIDpIVAsqETdwXAIh6fLKiDlzKBDWVv1KSfyDZBQuRC/j95xRfu7WUftFs2UUc9
5CTzcTDFzayoOt+/k2GEbORrIa1FI7fj/31loXANmDAjJcAJN7K++hoQgc/t3uLjY5ltQFJbFIZs
1vt8FInxlMYJ2XSlPbuW5YQgmXfdIq20dPIRJ/eSKUaVMpW68WoepYuS3T/aEkEkiM2vCxmxQAjR
tsehphXA8S2Holj2vAiGPKSvRnrQ3nDOeczbWNdxpzoyxN5P0dn2YQN0+SMQ1JtnGb9QzuBL5/fh
DRQf0JW2EuqqG7j69OY2C9mLCGCdeoekiN9613R78qt4k2lUr8eooijOVs/iYMJhNdLBpF0oWfaL
17LAipb7IvzLbHudtjzkr3nXml3hvxg2TVujexKv67p1NWCHj3DMeUBYSmR1KCcn9XcwSbDIYs/0
DYl9i3P1v0Iff4e9L+CEF2nlrSzaWjVYDHXutPSdpo8J7CCQFTpZQFnuyoiJR9Bj9FPvWzudQAOf
OZFHqQHpzC0t+fwiNchZ27bMaHcVH3m+24G4dgqlvDy0loLs/dsGV6TQ4x4ZvOLpV51pxXwPQ/JV
1bOFFa+Ah6MI8cf3rF73De4XLcZniBv2NutxZjYCPfnPFNlxCTAPxuEDevaevcZs9FvGvWk8jfbs
7X+hGT9SlPasfHxKQ7Qg1rYm2yWVd5UXdYp6ad/n2o/MgejVArLv+StVLElmYXSnoHtPrVar3Olk
7WK3SEJaJ60VzMzdWQaWfmIvWig/AYIAJaDHdtsowQ5xF+34ShTuaC6AeTLxjfdjz0nFH0la6x53
muhQtXcGKike7aBCSMGyymgcYTI8guw+pbydKZKpttmQlGTQVjpAzk9mIkz0SwCTmBNnbOsbR65x
WfnvwBlQ+MhLPN4Wy+nL+wlb3Rnv+qlBi96sGqj2WoL7xym5W/YEpgyEJ0pxLKn4JZERd4RU04a2
snTiLJTDDrsKKjzkzRnyPUxXWRkxrhLYHNxqWcCdfCHvrBSJwnRn4fyue1xUzZUuCi3+rI3XbEoh
67mcmlapTz3/tUZK8b7ocuKlSyEsQRTyNhpP7nxnUuc+XFx/4dwMHl0tS+tD0lrXI7JNZ+65zpW/
6r2xte5ZKuhVJhZA2IJAnMv5J45m9PTSYgcb4Y2ZRHIRL1xvKsYZxuMSl31whVolRn2SWGfHN7QF
CaZXbXeiQI0QQedwPKd7U9lma6jtita9Fl2mosj9tcM+h+WcIH2CXeDAw65HczcuKC8EiFKOx7sB
ryauz2qboSZx6DSuWHquBzCFxvqHYY/gi5HNwgftx/pJfIc1CmBfaFD/xMestaGJSlNWKj/8m74o
bgnkA92gCG7FYUxNq+HUuC8pJowVARmbzm/lGM+6BXvm1ndWOjLT8mowbZWp8cfOLnltwR24vNU9
a7MRjwknyqg3vemViGRnczL3LYJ7n0MR/pk1zcai+Vcr3WBKx+1DFHQI/VJpxmCrxUtfMuLo48dm
Sr3he8FYIt+IIhaJUd5mavVuXy1BY+zYRBeUalQs/rm0S73OJMnn/WGoOBV/T2vHbugFBzqRTnLh
7KtYcX6zRkyt/mYZAQq9inh9gTUfdpVTyF6++389W2YMGnEEgsmH8NxWIFiL80XDM6dblc5W5gBK
PfRfK4f+oTF6RXZVx4Kj65pH/a9V5OIMeNnBgIXS2jVx+CViPOK8Z0TWctFCx2u0JFN6LTB48M+2
GUK1ZbzOkkj0GsYruDg37wLXq4uugofclgx5nTo3JevrdwcwMuBWevba7pExLgdoW/LmZ2ra+ziC
St4hiAya0o276CPgLdDeZmBEWmJoYVw3Y9vEdFbS+Dgn4+4kuPUAJ9pOl0bhrYXS6Vuiv8qiIvRD
+ZnwhLngoKfmCl15cVNJd1ciwNhd/zFfOhjbZ2v7Q+B2+h2n2He4PWvsOALro12TTlMHVslQt47r
zS3umwYDcQbEE784X8A6MSGJFSkO9xR2HpH0GZZW4slQdMjgj8Gs5Y3pYONZFV4TVoGZDIvQum1c
Bo79lz80MNJooZQEXMTLszkvx2m0ZUhpepXKns2EWcRl39vayEZvyE71tRf6U3YNhtg0r3l81NIL
5BU4xnFf0wLJA1TFTiT2QSRtzgXPSU5h6Zc8HHWVDSAo7lKN9wzB0bS+GmNeUUc4NHsIiK1gqVWT
irMT2d3cvXH2w/H/MDvYYBMDlU2/kiekRYD7c5XeWE27SUTEn+JYnpt6EhWeOCkJhtezLuuDWl7V
9Pl0ZwBiHZAtu231KH7sbCUQLZ3rwLGLoIwt6fWOjZc6RvXQQ0sOo+BiS/19H+7wmWjP7Xvivkex
ucG8dHGcvPqj9bsmIw1HBpgY4EnW5u7jeXXUb6DSX9hd05Gvddc3zxsYIPgC1E1I7wsGm53q5OUU
2uhASFboJcRdvTWCVRHTqfLHCI0+nGwiK4U42hiOhsqjOBHvfGLkv8GH/E/Ok7xPMjUcB/utHU1n
r3sLJmurKuKaOsDTn+UaAy3C7RS/qIt6BB+iR87YY8RA3qi2Li6Lho1goOkNW+ZILwAUEkx3QV8z
dUyH7kAkfSe6awDykVHWfAcoV8pndzMaVkkJHMHJ5aaxz5gbcwuLT7D7e0mK76P6OAy5yNCEACJp
4bw8n9T9DqlK+KAVhuGaQkyIXCJQuZqZ+LO2hjnb214lwZwDVS+zCE1ihIHm6yQkd2AG4+rSYQk7
Xfz5ec0bVxWUvMVRahhOTRt2Xv8fbxjG1OeEAXypC1FVzFznWdptL2jCQ9jcgkMCS8WE69i3Mb2Q
Nf10WhumjfJOS3ECnvxng4HMiMdggf0FIdx3cBmuXyNsHUPx5xjx6Y5DZSrA474xDZ24KuEkRN3t
KCe3NTsEbE2cME64vPJZfT5uWCe6kuMyd15uvKC84PAW52PzKH44qU6PLtfIywF49PAUMvuqX1Ss
k7UufRCEfpM4ut/crjcpk/2joVZLfl6mnRuLc0ih2rsYwVoHHREFz+iDC2Y9q/cJwdjFEkHw3DnL
OonOKG8cSQGBZbSp1whguV/umXxO7d6a1o8dKHUvPJhxRRloQBvTE6wcZ0q6Vx5sarbT5t9hvHIy
ejsR4tnmEaWgVq54n+XF05RKM/OIdPkI4wolfwVd5c2xeZD+XMDAVNN4JoIagMuayB1mKDpZWnAc
/FIjGeX17FAKs5nPW3InP/wmpgBt5+L1N6/dLiEnWgVCs3/pSwXnAOXmyb68Gpvoa/vcNIrIcM4j
qzoC53ko+Q56OesSbtN970SGdCfScxP4vAWzh3YecvluIs/VTK4iRTip3AmxGaw1MJsFxqES9K3v
LMVSaZcLNxX1p2eOLLBDqwOWb4bUWWZLV1a40xYpWeRxhH9KWxcZx+fqaq5t9UM05mDVHOyFh2zE
KNbb5qYB640gNH1QDkHZjJYCA/JIWd9g7M7eW3oyh6MJVhD1ako7zihI8LElsEMEr66O75hXpuZg
9l2GZWHw+M119HbDcpfjTJQczxfKjPdfWtxslD4XbNlpBzK+2wdxPgtSZjeUv6x1iq6UMRLkSkoV
Ipc1jY/N8oKOCVn0XCpc2/nuYsfQRKLwz4Q15XksJErXYfxmzZn2eD4gXD/uI/qbS20WhHcZwUbq
Fhx1qjSK3XdiIjTxtY6Ag6jKtOqYOxCcGbSbbsrqc8rXRn7J8MORWuUS63Q/Sru779pZ5BxD37pb
WXJnwD95m7vUwgmdGFgTkRWKMRRzEK5uT7uh5qHSyxSkyz7L4NSQvP2L8ZXb/3LGMMgn+4KgXDvQ
UaiFWwuLs34+uZTpwgsbXn6JlHJ+GCQmLg9cwe4jOFRsOtqeuAauk6IllG6T/gCrHo65U3EC40Y+
9LLe/ng6ldwiO9RLVE+CQLZgXbR1yTo7ptFb7kRrMIU3GfNnVcxxkUT8SzwkUYC2w5FDP8imcBko
QCML7h6eGxg8t7fu3rp0H16wDib0QcgEB9JDyZeBFLISdWMnhEWH2AeviTRV2Dn0GG3PfrFAm6mH
JMVu0gacddwTLlG4Gsd4KYcg9yiTY7kuuav2U/vhOimzoUZ2BHLbDJSX0piAuAOM2YFhCwgkfYiD
itAlMPsmTOHfapac9tT9cR+oPq8XF45QI/L8lJ10aViIpim03+++nX5RFuNK40nthhHzpeY7BDNk
2HMv+OuvkVwaofiRxEOMKoQM493/8bTgtPYdJOg8/nOuyC1KKQeeZShTcOo7/EOTB+3e81okFShR
wDwzKEDnws3bahB8ZuhaH073fIztWdZ6W+Js4y5dH5ig0IBjwdwrcvNijSGePnm2amxibROy/Nh8
3pKGqjrikO0LRPEeGw5obh66kIWfITmKGHTIPkzFpY7EJnnS8QWTkYAfP0FMlzWuAwEMt832Lj2W
gyMsaisk3q9mK0mW/5/3k0nAJo1mrX1VH36rVoiE5WbCJY6NBFXoFKJYJbVP5nmPqcBFilXf/xuu
ujz+YdoZ6gzXxdsBmOx2VAxHgBrAbDYEDj4QvS9kQGKvx17/wFQYtpQq8EIC2sBKHcOVjXlBYOJD
oPINw+blRxlr3hZZ6J4A734XMKNXK4X6/3WjT9Lto8bB6lqDtE/lTMiFyDzoDrD1+MNjtNfAv1Ta
Du+HKnUqou2NF9CvHAel1TBfHhaM4aX85fStyrKqSQTHneAk/2tQezHwkiy5fiZXFNSfWyx6Nu6M
z15XNpc4HsXWassbaS3D88s/HjkqagChJ/05uO0qYrulp5m/NLvn+dhx+bxh8tWYFxZ1f30EbRjl
x0nQipbQ6CX9ZG4UETJenpnNUvwGGmknO9m8CVeRLArdUGycgNiuEaGL1PPGai+GK4tULaUL3ubi
d6Ny1+zEvKsjpB/A+tM1APgrGL8ZBa84G0O+l5p9/3YCU158ehIzPnuyqFo3SR1dITDvjPy5oiss
bzwU/FY1DIITByAJaqAiVWrOr/HDsXGeshnjbON5vusDqUJtBHH5Tbcrkpe9UFKqiS+kNtSviuvB
UbJ7dKLgTvnG3JPARqZe71zPPBefPtH5+WM9benWCJm0kPBb8Iv5XzI0NlyA6MKfOMpCfoqvC4oF
+j7GFfqA4Vr78JlLTvo7w0u9wSVPmhcqRdZs6ZCOtZtJy7miGvOh8KSNQhTs+0FWlLWiVfNuwPui
bkqFsB3hWWgrZ1v/CVelSwTPxPTAAeLFDR2Q6STuzxeim/Js/E3KdklE2eOknLCMmy+LxOf+XjdA
KAi+Rmwmg0S8oItyEOQ/isgiSWc7oYybBcEyvjOYlzEcnckIdefc3d3tpWLz7BeJoyvYvk4+prEo
+NbRP+fKN6P2Se+TFGRDSiakY7RTrQv2BQh5iW4/vuj6h7xcMzTObDuloXuHmm0HqfaSKccc4eSW
iDippJAQDhWUDZPnT/dUQYb8qIHiaU3vCQboWcIg6tJbU+TfiusbJYphjdNmwPc05/j0b5Q0HFVK
pYAOofnL0lkjuzpyBNUDwTZfqJO4BdXK8fOERiYsIGviUFLyGUjjs3d0/DBtG6ev369QBccS1btW
HaDAEu7B5nOaY30Ppw6P9Gp2E2gse6+GP2jq4Kob03QpsSUPrIVfbj+MJ9k819iRcImUpNiqQLPe
+bvmC5KPFmnBc+u1gFJVrJMDqeqAcyfgm4mN5x2+UBcHFDPDeCWnCYjQqgKI9jbUyH2IGg6CPixR
GA8mvF9Akf0nL+GKDz3M8yZGRWA9iifZ2lAzdvKXPXgI6gzhMtktHGrcHCBuD4YDOiBTX9B+AHdL
LvV/mp9cK/7a80MOWnREbmFxBvBpIElCOKp1NFuYgQcd4Jv3wsD3Kzc6EiXUSePsGLZE7B3wZbLl
oiuF+W/B4iXxK3o3Fp9YgZYYKEBKnJ0RIDYQIb1nFRlXPpURTewAl20gSvNQRKCn6q6pbOuZIckz
W/Tvo6LQiIqjCiMwe8PX8kgnLRUuaMov+J6T64QRucInl6DYCESLOqHBJNfpeBHYIg/cB4es487Q
1wTphoge7jLBvndS18sBs7IvcDj3j95KBC5nMOaXB7Q8vv+LqrPl9K6qhJBhISS/zx1q67HtxUOl
pp6bWqzBE+Yxf4LyuZfNiSP5EwpuSXJmoqfXCUFR2rE+uENY/kqehMN3qILsmJs0N92gFrh/alwg
Qb16mpRVf375/oXI8qM6ZUtMur0nddykK4RUUOOx9RHbGLACeno6dlTnOIXvS4LSkAx0VAE6uQu8
X3dBTDmPCYffSa4uAYa5cC1JekIEjGJ0v7rO0qWFLQbgr64XXK7C4iQKhGNaBMpnRB+dqHozfD86
9o/mZUsipdE9jDWNfXzQi0YY7jlkZuIUrC6h0DJDvodH3VcYsdPcKkwufr2e2mCctEbZ/+oPp/5U
V/GyqwpvC6AY9OT/rSviCsggkrfJklUkycWffRtRMRF75x2BA3Xfe6RkA2BjqGuns1a42uKB08eq
zcZuuFO53Pa+wTwk1fFJZ2qGYyiiIsr6HvY7A7F2J6ci3F697uWv/wXzwkN39CmPrDOln5WjsyKL
k683mv5Z2dt9bwD4lRQZQJj+vTBjxa+J1H7onhQmQsWyaqrGks9j7S7sjfrl5v0ZF18ias/phw/M
OzbGzZmMn6YfiRQP6RyLFJc4+0pH4GhP4RxBN8n1aDb2esB1apvtlJFpd0dQI/0tIo5hjtORyeiO
hhIo4iCyRTOwpUeyYM69niT4x4GB39+tZi6+PpcSDNQHaRhOp2UXmTLJRX0IM4YYHsc+dhhZ/Kg5
A478lKS/7lcP08QxbuoqSGApm7XIP6LuVDkDDUDex9ojoUG7nTgsP6PRQ5KSW+Knceo+nSnpN33A
ojgMT3b84yh3eJSkTpZ1dTwZTLnwNl4E9+U5HXvtM1LGqc1SqW8yIE6K1OEKP/T2qKDbOXACjrhQ
6eYXkIwxCXlotMWLqlyowu1s5Ld3vfKBq9MgPdlBdd/0PxFHwWDRXwIu5uMdnGzaz+64olFLWUzh
izefUovptUufNkArT4Yxgo1lq6N6XB69wqWbrw8wS/ORPGHKgafLV+fD00twIATAgQPgFN2jUffa
cFxLYWOXeAP+IZ/c1D9yKuvpJtHfZx3WuMXUil0Dx6RaSZD6+jqUkzk7EOSI7EMV8YJ08O9yDePf
rc1RjKLzrvIlpZrLJoEhjd2gQfR5ZE77lNtUy0wSKVvOjBNnDpf6Cb22iex5aPPcKxFfWC02h9iM
2Vkn5kAwj0CZnoEp5nYl9sazbfnV70EZ0f8ZBW3FfY++11Tj9dZRoPnWIsm6P1q//jlq5d+Iar0A
sWr8EmkJyE9kY8C2a84YJVc5Q7aSYH572HPJsiSPbI84YLlMUig3gMnBYFyadCHhXuyBwZe1qCuK
fhbilHTSlB3C4MfWASzj+TRrnq+Xm9RHN29L0trzoEOCHigXPAHllt3BKfmv3WjlIUwburX1rm9Q
djqROkN4IUs1ru5cvzX+CzVsF59HGFUIXltZ7EZHaggqbeY4UEH4bsHjh6A7GlouFgd69a7t0/+5
TEQ2uPMKiNh19fWL+7JutD6oZErLmZCQVWUYaRMYK5XLRNvlRUumOcCQBok+MB8SUSqgD2/ZVfFN
TseDKRU2rodv+TCOiuO8cueiPDyQVShbaVnC4plWt7r5phu83x5aWX8AUdBdOGcD43WF1V8Z4cQW
uNM4i1yf676eD+LAGHgGc5DmJ+pVfe+9oojjOQsQrJk7LjhcG99ZJaXpInKMHA4gVtdtba7UARnx
fqr9FK5DIMAtHrgUJM4KFrXG+77ZLPNb0hAh6hdxvweDR7OyFEfCDjZ9VPtBIUF8uyd3CZBS0XFI
33Ye2Rl+AYSWT5hTr3xTZZBxNTwmC7oMWXwuWtGsQlEniqWj8EJl2Vfo8a2wkbhbjOoQ0dMCfY62
xusPyBuMy/2bWrM4BiXz4xU8cJWU8spac0Brsn910mU+X9ndI4zuNG6MDPHRX3JGGUMxRUCdlgzd
uzYnNKR2bvaPgprIUzLJp9X8AZUz1jm2RQBBQMvXXDPIAUn2amHXgKD/Zi3zxRmlW2cMw2yFiLw2
IpPEjGHKtqcEgQmLq43AywtlbCpgivZXP1P05XoSI14sTAbBgmytvMurghzuO+g2HzJyLy+PUt97
rKltsm/FNGb3Hp3sJTXyjTnkZknqnplNe9G6K2gg/9eUG4QCAzpjlGDJGT8BQOw6cj0nxvp82faV
2w/12+wOZtolwNvLBior4sNiA8LZi126CDAZQnSqN/Rzjip+PJwt/wc1buHng3/Ny9JCTFL1aZqN
y9gao82+WpQZ/byDfNn2QU+I/dXrGf4pBR2vHdm0VfPDKl4FtHKTA4+fsFx8ViB2zHPGzGcfPs4M
rtyZH2gZz5j6w2Vh6l823s5hnbb+NIg/J6NMkrs6bnTi8IK+V6DLbHpkbdrFekPEgUtwZ5tdu7IS
NS++SdO6oWXuQSMZQWPgrq7bJ7WW/fvrkU6/3UyTomt4CcRRcyy5w71YQNaDfP9xhpThczNTyR9B
38HuTH2iEvdlN7x9yh3ALXmGgqr9WQ6oMwxBzTq8DRH2FTa1TTN10slbtxv8a5VMdI1hDm8FNDT8
oniP10T4prd9+zExKkiMJgnlddXT3ditqI+45LEcl3Xt08qwusxYaWRC9IUftfJnmpECr04+c44O
s696fiks7OTzmtGSdE22qIA3YJc04epH7zjH1Gzcn2vy6G7vsXS5BjT2jposoK1xWqhXrqoy8Kfa
NICPmJFynXArtHMy2LJELg0E+XwgXMBQ76zV2yeMAJs/v55IEp3Hpq/etizfF8icJe8CrwAegY8z
AIHxqHNyNnZWXF+9f4WPb3ZHek3JFsOB85oXmOjb34+YXRTLfQH55W0RzC+n7dquDH2SqV4Y2OBm
9rcbwD3A6VIXXeT/5EctJuWROE3NGfHrQXtXYTjeGiRL6hguSyYKjnBjHC0nLSLTGrIEb2SxOQ5L
KwYoB1DJo/AD3/L4ixQ4tye3l3s/purqAKQ1st82ZkJZ+sT1tG4wPr7LuNZ8eCMZd1zW8Ku3KT2O
TNuyKUQTp/KTcsE+uzaiKeffB4LbZ/bgoqLJBtvjxLYaavpwm2tOIIFpXpvbHSMw/WItz5gNPHuy
fDibEv84gyjztzXlYZj+9n3qEQEzYBco9xsJ0sca9MrCo3tQ2KEmz9byw8sf8IcA0K3lQcF5+GdF
SVg0P/6u7gx4GhCakmF+KGo+XhHatQ8fIFD7/fdqz4QbSzn5y8HZtQ8v9kTLuR43tfwwQcmXQ+Fw
Nrevzw/xe+2ZfZj1bQOujolS20jpQ2OGlNA3HFW5Mg23i72Kf+subA1A/l+6zuDNYE/m1CSDJMQ0
lDzg3zjVp2M6c1SB3jwae/zUYIed5/C1ZClK0J2JgtjEBIAMNVj4v5WWlkWVDt96jy5JIY3YNfbr
t1SJ95sDdt04BuEhJ8uTQm9CqwccuS3BwQT5KJDJ68E195lKLH/bLZqii0U2UE16NWLI5pB+xwGM
DziV23feeY6HA0T951OXID6PbVrG2JOuyCHgz2IY8XbjnruGUmfTkRqa10wudtEinL9K/NYfP/SU
xzkW/wmE35XI024D3qOtIPQCo/8KU+f/j6QI35wWGKQUMlgPHt7Yh3RWw5blP2KB+DAjq0BMpihE
7ZD0tPb8GMWkzlV/MgvulP6gYouLpC62kXPX7YnBcZYc/SGPlYGEYo09aIhEPeaZqItsFdMqsuQf
JEMb1DEw1M9B9104k7YQWgUwZDkWjJsdb8M0hGC5ywqrstQMvyDMZ67Kt0CN3/Rlvlg/z++wf0Ya
49HaMVG7J1I79RCvJpfqQbLfH4LjKdcbuIVMf2RAvZil0Wv98hRofe3o3FmGSNqw5p6CasMielgN
7TTl5gQRxxflhq9+YlVl9DsF00XPy4/92GdjoEpOBvnUtMm4xC+i/jChXvwwolRuWqeokZlBTooI
bL5FyNJYvgpbOkuBNqhLNLaU1FZP1ybYW0jAmJ6QTHUSfRjpp/e+2GWAtjjcblndR7KkuOanK8bi
ssH8n1+nOqIUAwIF+/TY/rUb75kCfhURdSb8Ys2pM34evex9wRytscN/LiRGEGUuz0DYwXso/x7+
C5ZVEFSFgsL1sAAun7sAPzqMvHYHV0ldp0ORtVdvyzA62ovmMtTE4fbei27MN+/JzgIWSe+mpfW1
kkj/7CZt0eOzm6kq89e3gt8Pz/7dok6VwDOYukXJRszJWNRKW2/m0H83R6OhKRWxKEVsQLLbAtAa
XU0reij3k6/swDyQ4UOlMjD5EfQKwN3UXxAMvyOmYhQr0j+jKzC9GaAyZeTVrw09+teKwxom5gZS
BoMYHRQ/jLzRz4us8of6t3SO31pJMeIRfJVxkB3r3qz6JIbMfU5M5eyMlo2mZhd/mcwq4s1oDPo2
rpWkabKc6zwfaqwPuoLiLhsgXsCHIUfBoxWuYaq6zJKMvPLxMOPwpj7htNnNo3eDC7EMDhYWhjYd
dCdufe0LzzvKH/9yJPq2IYGcxFZe/crL8ALRBKomlUYf/sD32KXWYuByDt2urPjvYNLSR0TXi3Te
htUocCTdZe3ynyuPMl3Ky5xK5ISFBtbROwdooVz1JH/tcm6AgU3+676s0bCAJoUITjZ5Xi9uOzn8
v6jYPMDjGys4TX0KauId94pKBvDqtLGLoAThcPtJTs0mUbx3GOkr1/0N24RZb0BP34Z8xTOQ/IoX
YZFkNTxGlmJdGWHyJG0ALh5w+17V/h51lulT630eXnrVlI86Ud+5Bza69d0HYuVZqd6rIAROQ9ke
UCV0HcUwf1Nhx+pxvT4XOIROhu70147u/lq31+6aG3TawxaxX/dcfakZ1qQqpt4wxrp80ZWxj0/d
Vpgoc0Ld1/paWQYIbHGN0YP/jbq6TmGvxls/9OiZdmjf/7xHJizayuOD7PkdquVjVuLr5RH4aBZ6
jEDH7qrENyASvqCEgYvG+qdbXOGyNOfoFfcvGo6d33tG1MSMFyWpA5G63i8KBpELQc3ZxxSfTYa7
4vdCxv1WdQpix0UoycyX9uAEZYS2m67LXAx9lFanNJtE4WFTx/kBde17sXxoulncfV6NXZGP3Xjj
tAxY3/AEJA8+BFntEjFjtuuvPCa4irZvegyQsS0+GGp8DEafrHREEDY+BlwKoBzbMyb+b6CXT1Xj
SBIVMxZ9HlHzjHFSfw/th2tE0mzFhjDA+ThHVblXgT2IF1WU5iXJElLiTlu1hmvS4fc27SKSqhV4
Cu+Ro9C5KENDvQyGJtnMM1gtST2ufZmCGiKqCNGV1gn9V39w8mJQWD+4/97mSPm0CeRzHhndjOTT
cHx7HwUkndhNC1tegg8pSq0QJ5T3xmc6Pat3jvA4DCT/SQVBMCo89CW+uAywjbeDfLtS7akQjkzM
8BbXVmQJyxgDfV1B+vbFhrxCxo1StYIVTk4h6JukAIPwA+TyLddmdteuKyk/XdwHRRmPpAGMeqtf
Vh3Wzc4Sj52fJOnJe5wggDaqtoMDX9NHGCqnT1XanTzJms27ey9M8x2IL7dAQat2hjO+wgSeKG/B
FDCDN6DKrGqt5gLKbp9DuGvBcAmFrrmksPYzNtFcNYwutL47CuMd5F5U8JulRl9my21SLkHMNa8O
8Lq2ZMMvST4py1dhyedHSetMpjJwYYr/rkhqer39Ir3w5CIN/XX0WIl0QFE8hYl+2uwUd2KUL+o+
RA1Bw5d5MQa+xTm4/WHAGs72dbg7CUEQxVhRSHwE6TowrG9e7eKbcLjYLHPyQNxqriEm+iHyY8HI
XjbCsIIj4RW6T4bAkBQLZDjSsmQpgJTOwXwNUu2pLC+zPeETdHa5OEJRaeSXkR85PYzoduISwvnE
pd4eN2+GapZ9YMN022zMpyd6CmGv3/5XsASRo98GI58BYhY00fMqNofD3tKz+9ZlAwZfRfGfZ0QB
iD3DZ9rdocoraoeIQo4pCwo44FHcn8TDsPnyxZ8B+45fZkUtevWmZyvWoHbfT7kS6eutkdFU/Fmn
32FdulZUDrHKScYpjzkZVqL0RjaH7Vq93ufRh7CDkzs98NVscI9cSNlNBDiXfrrGurjBl0uafzuK
xkyYdRKiYtkGuV6AnL5lgh3oPhj9/XVxWQeGauREySixp4dZUSOjUqlghfvVkOJo0Q/Ao3f4K5JJ
wa3JSv9NqueNWfi/FVHoje/oOf8qq1A9RSx2k54MwoqWw5FO8I1j+tRVSYoKvnM3gTXEUNR3lrVw
l2AjpTsx33eJ+Qkl/Jf1zkbIDAHpObvpEQ9yQy7yZVpWUHcvkECsNek7KhzcwS/264HxAa4uP/lM
tELxOPdEvokpwGxLwSDayXa5eatTWL0faKSJ4SpcRpbRV3CRmbG0C/Mhc5rmoxRIINEdiDbT1mv+
LhWmSxjBgR7qOJvcoIKiG5oENP/q4ZbFEV8yZBk+y9/7f8ugZrSeFpT5vukXPNWNYl0W49UJkPjB
HEQ7rpYYGSBlnR4i1q0oNmRLaqy6vQ0vd3pJNgYOCZn/aAGPrx3Z/yoLA/E+1EzFnBe11fozY9bo
W8F3B7snsuhi5SCwun5Y9M50tCqjMAxWnsTAsgxQqkWnppxMxRcolfv5OEU93PubdjfsVTbrsutH
KUoZ37SM1DXibLWfPs5cT3+/835xMNT64pofQM6mTDflipM9PxyfqK3YYhZjt4NSVJ9yROeRaQRR
bUjSAj8SxiGmu4n+1zzKzg33vCA5iElXsCJ0odz18JUaAD7EAIizBXs67sNwN9eiPtSb7FQh9w6w
R4mC8Sz3Rxbmx3oQ/2q24Wuq4ldJZRSlsrKvW2QGXVbOF6feybaCKYtVv8e/I0nYV3UyVJk4uCXh
jcEI0ggn52ujyaUl4buH2BZc32msH359JJL3Jw5zMZOhOeoGoiJschC1aBS0r11oWQNeZtR2WCwm
AiDk0Sv1Z1GHVtEF6OJAGp9OZViS2BLfR0AXValUoqH1IhgPlNhXPyHTBIAgwfzpRuS2mklaubLz
CtpDk7jkpWQ9Ou6i93UmEkQ51jU/qWWJoTmW7AA+11trApE4jVKgL4QPhjVDSg8b8x9VD5D32Nu1
WtQRHcjflTvB//5BEKnoD0hoipeIwCj0oOIC3udMlsNiC2kB+I2INv0MbN1qZo6vsqbDXYasUhia
XSC5axlMWETGXuLi4NRgM5bW3A7pur59iCTdV+/vSjwPY53Siak3OJvzgRkIz6qMFwFQXqid8gfA
+qK7r1ZUY1uF2MZoCEThJGF3wh3QPYvysPrLa/JMxOro/sFJcp2Q0CK8rNAbQCpF6CXGDiqU+N8L
/d3kg3Udz5u2xLa34f1hoyOvdeK4QS8+hemJ1WzQzRWO9nN5oRF22uM20EQznhfNSqVY8yqiyTNK
ma3kw5/vht4qd7s0LCQLzgKmBzu5S4Mf1A0IhXotr4ofLG9B46/jzjt7vMhhE2rnc4svj6O5gjcX
l2xpH/vxodSrAbv4UaisLtOpB+L35Y8NHuKTEyhP+jB7+IOr///srBTEcG6inUHD8parFCNAKdr4
Hjn5YfPBdu6s1r38I1/P9PErUgcVfuXpWCzbisulsN3eqANQU6aFvhRnf4+QhtYIPgBZHkW1fQVy
TgRpt3J4h48oqbg8n01Z7B94+C6RPYDqaTJY0JmuWlQWSdKA5z+9dcTKL1b4l+0P/u0/HO0DyupA
0NyUZga19CAwKs2Wp+6sDiWNijc/8UMdFVPJWX64srf8K8HFmbKAnLUJbCCerKZpVMgn8dAo5gbm
QvmdW5ilnSdeEhlxkQnRNpTMChxUDVvbHjLfEfCq0cwZ3w7QabqaE2MPxjBWpn3lQgUi8UUylkOg
ph/IK8Tr01Wmi8higyt5qHkQf+lHoFPKN5tMRyfQCUQ8X52sa7Iw0rZq6/YQ2y34q5Wrky8tOIFe
IAeaiwLaTjXd2OMGyYh60hb99Kw0TM2SZIZ0ySIUK6atOtB51vs9QBB5sXX0uRSpzPrqLN8hmbZ1
mGEFcKL+4ILpbgaPswGLpPdNfqlAqoBuLtHQJtla5d9YzOyHO9TcdPTQBlw80vg26+AAw6z4lv5P
3Oz/omD+nuT+/vtt89ayWc2CgpvqL20KFnjhoyp88CmBzO7ITMi6CfdLQPFNOaB1xNjgXxiNl1YV
mpmjBV9WACHGAL9FNILbk8+GPE6cLPkQ74/aic+4I2MIA+96H9MhEVuHMA40A5oMUfr9WEiplO4M
Y5AeznDGRfSKc6vTqG6dut5uQpHfOa4sqf3/FruaE3nTRzI5KG6QnCna5Awr7hn9o1hSuvdGwVtY
KKQ/R/cPX4YP3b84Lw9pawP7/ebtAHbFih1nceQ6tm0juFmSkTvh+AFacqGzq3vL4WaT9YYKS2Fi
JOjyXgXbSlYJ4tf3dBimXElFeyUpTjjuP5ejqIHoL1vHkoxDUsvs7Y47shMqg5E8NQlKj65+fXdE
xmPmOGkKa0xBJW2Zas6lzEhccjkzJXY5PkTwu2ulpx4wXEAZGVy/zrh3itumQ6XWPnpgxKdMk8Ab
dU/TGhG7qvPzJO4e5z4nQH85J/l906kSJ4VCrqHMy+ZuyzmmmisiWlZmy8ZNCx3hgTdvEIiCKAgR
sw1vCerrU9cdRvqAbJtaPnao9kEpiMfPn2xbybkW7MFWIuVMQTeSjexpcRm8BV80QY3bjm4SLFUG
edjM4reFhheMFBvGsxiclIkU3WCK1NxZQtGZAtXquwEN7n3v0vM/n/PTlvwEyLfV4+AqI3vws6Uu
i6iM7kxjOWRygy49ulPXZrbMbMT3od33I+6V09BNGeEHwHqpSU8SDz0yX77wROSAo8r7Fa9/fA+6
QSr2viZKC/yVHkTXwCvpI9D9qZVx73b2w3Ti1klmvLutCa5QJ80UjtWBMQO2TKfcIaN7bNGsFfhc
KJEMyJfpQpGI8gK+95RV2NJB6Lkb6z0YSOfG3ctI2hMKm7U5CQvYhsM/QFBh1VkoniitDDKvUiJ6
JNxpKUo74BBsCm0DjaAHO6b50QfQKMnXlXc1vHGyIkuCrQD3AG4gZYo7qhNEVMhBGwTFJVXNjUC3
K/XQMRhLPjLXg2eCe+n8pUmYY9ckuabdwUQ9DvFPx8twPJDaNFT+csEYqMzBO+CQqZ+rXc+fLJlx
6pRp/l8TcYIEKwg8K2fSCpfVNo5jDY4p+uMhyK7kaF0GFcs7pbtDRKuZJd4exOM1qkI7PR4aQq8c
TRbrOrSHIXV4MRpWNmrcK/0e6BO0FC+C/BkdaFT+22ZtjjQppPWzOvOwkPdaIzYF/73sRjeSd52j
UYU/0qmyUqBE5r+ORixKfWP0yA16895LQ252hnKVlCSayp34Q5igOQtmN5koB56qvDKfQjXRHmwv
z8ffCe3MHWga02QIjFTL4p5uLLU014El7jjKvAjCYa5uQr/4y5N3U0pZyWN7O46nbnt9L/aQHpuK
PVE0fW8p64WNeIc8bpphKTzBFkRq/H+mY/J7N5sbEolfO+tFWxxPaqU/HkJG58SzPnt4GZSpiKZ8
M/gLuFuzcQxrzNihx/lwq6Pcpyi+g0voOJlC2LrDodVy3DjycE93OmYb73tfwzLzyCywRFdtRHWq
vIQfLhUkEY0i3lIT119j6eWLTivAWzjXnEQbzPd/uWGTQxoseuC2kvDMiDnzdEeLEoqHym2Oe5Ah
4mda7Vbze5geG+kNoO8fv2/ol13l3d6wyvpCRuSggnz2fgPc57O4LyQZM7hTuM/KnTOrL9zXFVzO
UKViD0KNzZSEJEyUl+bwfE1zQra7arxUtahusxc61VYtrBk3SpceOyGp/o6AaLyQDqUz2NexMAHV
3F8EeH7HeecK6uUtZCFnvKx6L+cg3Rkx8hOgxwXacoO7ncfbIZb2itpzkDC4ul2f3Novkp9IZma9
sGR8pjyhL6WwbuEdHG0drUUccV77MfqxpYP43ouK4tVXawgsFyXQdqNAmjlFxu+zeJI2vebW+w8C
sxA6pMsHifS2RkVKkQU+MqhLH90pHFZ72c216nhaAXA/St1887oCc0wXz7iZIYdyYS4Jn6DPHbmj
3gSOAw2hin28Dh4nJN6RUWqC5HY1wY1Q24yQzHIpJw4dKC8QsQgjjqYXQWc+CmsmjfmNBC8toBNQ
PUbyiUSvQG2TvlY3zpYlsyFvQspLvP2f1Uvijb9gkKY3VZZ4bB0In84i9cJDhdHGbn5Neypu7iOK
uZVROfoi2NmHC+Gu9Ffo5fG9HmrwgPiQ3DJx7O3FdI85fuPuEBFVSJ2KU2W6KVki0EL9prsbtRLd
nC/1sOYMVZ60UUGaoRdNbadrnKiqG+Z56dFn5rWGATghKFwJb2EUamF1rzOarGw7tGJUfdtxzJXL
I3VPWg3pv4B1aBGdvjY3ZE3+dnEU1Z44GERVIUcbESnzJ5Yg0MUY+CSj4pPCbj+c6gl9NJUpIN8H
KbsvteNtlAALJyxd2DvOuzCIPNez3O5DNMb+Fu1dBddcH896LsGJKYTqpLCTj0xdwB2dQ/tJzzCo
TSytycHLaH7NNAHynpRjRBl2mI/fPizypzVafeDZ0Oi92LI8Zl1OTLpsWQ+SAngf74aDnbXVZ+Ba
4cvJHOhWf5nAZsVsPM1THRTK65oEsGf5B8Jplb0tkUalW2A2eNjbvdALRdF2oOnIBegoyDS2MdRg
2o9QlsvTVy9GWu5IDXSsvSTz/Y5cBKlo/r0LUlT8cm47PGhwqmbGYwPxdvhPoKIGPzQ1j9nz7Rj+
mvRNXLSVSS+djyWl011v+ye0o9aaCh9lhgOVEv6Y/jKZopYG8RlWDyRAVWp//dOUze8Vq2+hfAY/
yAYaB1YmaDBXXa8kGeiSMeihPFLPY4TarVirOdjvGfWK10BVVkKECpomMicIHDknVTXydATBpO/P
xUX6JsnTosY5cAzGkPyttsXr52Vh6jYN6q0DVwZiDb9TBsu7Pt/l0Z/tc3+RL0u+I5Qf2LAxLeDu
a4sLsMS5r0uTRcOjRz9acjNFRrfb1vEzJYdM5IdyUNGdZ1ma9PE3rjVM+UL+psBaBAJ+JjCY4sh4
OLt52ff3WtJpvSbd8Wa6Ry2OFl9+NoNzIjprKm7gdoYyMek4c9u5H6pNPzysE7pWhCRyY5bK4T9o
TzoVtRvMkc8O4BvHb5z+8h4q4qUEQfwOuUvw6EYhkacMLr+vWv08PeoY4MulWadOsCxGY8Vmpa25
7uSuIlU3rwgFBNybEXR27fyVY0f0eF/PdcEYg0jbh3s5vxmE3by5HnCl2TMG32QVLqRdk5F0tLfG
a5A8KHoI1N8Rln29Z14R4LK+5zQUV7QJmPr0sQrwH96H8UWyqgY4VvxMp1RjAaNuVO1MQ/XFwnmb
JegxxWGvwQHV4ySE+Ms8mF+9sNHOoSbv2aQ5k6fHmSE70Q8IB0IZO6uG/lTS1cXOnbUIbew1vPbc
Fy0WXmlaTIUU3SxqtYp0K44K35tc6bf6o2i6Rsb8tln5QlhcJH2OHb42vrhArK40sNwRz0SM/L9Q
q45SLzyHe4i0mSt5kOg1GeXUoQgfYz7kd2iwwcxQtcjAW8Hhv5KrjsgHjKwXLCGS1EAV4Hqh+slB
pNph6FPMWBPbZoTEKr4SrOK+bb/kFXpNRqn54r+s/hAEl9uGiFykQUjRiGrne4C+IQuFgsq2uBXo
0IkVnGlpkZgU7eUZzVtsTsp3DYJRpd02fj9wOOIR2t14e4B7Sw1Ojj+3kwpnbV6t/I4KC0+M8PJX
V5o+V8XJuzuPryFTequtNSwYqm0D5GFtbvyAbgOU5VASkCWFGjj7kENt17zTa6P0Nz1botESpDyP
wTmXU1OF+TjXqAow21tsi1LcWeqd81jfZtIO8anafExfRVcaXZphAOZMpK7eCMkjyYvYi0snAF9P
Qloo+Wjc7xR5CSmIkio8VfPRBRcvpDF+uTY6VrlwUAyLJr8t+ugta48y2NVYt8U6KoqvVAG48OXT
KZvAjpYIF/dEl7baeoJr9IJhgZuS5/RtF9wr4NrViC0D3xG3Oxt+toI7tGkTFF6qAr6gZ9qwah4p
g3wBF2BWFrsD4h08sltzBGI1E/8fsaU67VeRLTqVeZmOB/j4Yn9S1BElVEugFe7JkHYy6kaah36q
8MKviRbOHTQiouX+PNTaRUZ/ERCUJxBIou1LYJQcN800zVIqbiKceNVk5IW9iW3PdkfgBa6cZUUC
WYFneQ0d6+FDEaZ+byVdop4JOiC6inxiHmohQp1LU6uSIM/PnxwUiwcdI1DuJBGBbOcWU+eymrHO
f68Yv/wVsgyrO7U4tM6sz71H1UnJZ1mCpN9SMWFdQAiJs6ccCkd32aARifgbjj9dqL+bYQr75R0C
6Af4yC+tPOPHi4/m8U+hOo4lBk9Ra9hrx+pjsWcLILcCe7uxoFy8eYcwnYwepCankAuALLge2r7K
DrKSrAIAkXDob+PCte0BJesfAqLOMkyCv+jDrUDDM2LwliTpYUdbleYUJLVsH/dP06MKptucMO2u
wfvqm1bKHCvTyEnTynoMssSPh+UDNVxMtR73bR4TCFJ98+nKZpZjjmahPc1n3rPDDuysTUlMWgpu
3sYS+j6yZo3kD+k6YAsXhnZcroJIDiXGb6E4QiajHQQWC/WIXv2rYlexGiq8yzAOk9TzcCP+k5rh
/01dHnQw0jQfrW6OYyYZjI6E4vIQ/xyhh3ldJcdE1j/QXd7S/X5WWRJqNVLGjkZF946VTXySC+aP
3tz7eVVhGbRf/bNHqugnrmqxVGjwkSYOx8kqbStr7V0cVa05T7uK6iwWQjW5KaclLVDRb2uvRi1h
/jlnz2kblUA9lVyqQWVFrRfDzZJDzq9zHmDy6R2qW5WbPQMarf6cQZ1aQek41qiKJrmrGbNJrYyY
in+8xVtly5XQ6yN9lyVUEIxblDTSyBVr/W68PJdvpeu607F7gX2yogy/DQkycAEIsaY1gwxPocfo
Y+PlD5iSAAJV6C5RbN1AaU/XYqxB0c22rPuTjiBo3zh9ZotDRuZUBOMfISNC/hZ1oXvAhVAsKUvz
yzkpflk/iLWPdHkh4hR6uHTIqzKpdJP0Ie7R6EcnBVAmYvJNmxSGoT9NGwUv6EjJ7zUNbLm2MzXh
6Wz8yb9W1ZEcam9sWpy0pLC73PuSvj6u5Cwkc/rViNYq8DRFBDJ3h/0Ty41BV9B76qsBSfTaGoqE
J0oxv9vpIndAgV8Y41TX7GGMqir4H14hL38cmXUxcbgdvKIiS6V69B1TJfhR3uE4DBBCM0SfunBl
saB5Rkh7EXSXM/Ynm5iX6QRrQAxHGDpEk5pKt6jiP5VjRHpMfTjh7X2GSll47OgH2H6ROLl+lKoH
wwIRvsK0AvnWX/LVWduvPnl4XnKRqj+Muag/kNpiQkPr5VLvzEd9+zMjKT07jGCwV1Gi9KAZs3Uf
oLzsjOjLmfza2mYYPFkdw/HXeg9vP949Vq2ojGpBttnK9BYygvJfH+3cb2M0chq3Tx/CTkO2UPo2
asEpTceH2Dbrjvy7A6ToPPwR813jf1K95yrDuiXelOablR7hHb2GUZM0EmbJZEtKvrymGVWXGxNW
QBmNjluS3uIP8Yck7ilhT26nOQPMl+ycDtlzRBQWi5uPxv4s8GcuQMpaiBiYT7CZc5GUZI/ym05z
HTC97NL0mjCkzvv1BSzLFWQBkf3QGuG+ChqYKVlj05IcTjYlqH5L12uFYvUj8Oo5D86kR1nlbI3X
WfjsDLNwUgM3+8IZmINCByaVgrR38f/MPAuy9EPVyu5SscpkO30JfUFtKNcgUikpzGIth4j0wTq4
becoaq1x4i8P+wgN10pxqUwgSUpqsEATQ0GpDK0+FnTpv1/idYAlsX+D7nCWhd+piwQAeLIZLoPZ
hX/uQM4JEHSyBlMOjrbUVsljw1Mw8U37AV2Toj6SuuJjsEqJ9r8t14GKfo9vVeFXldbb6pkobgvl
WRKAPw8UIsm7GUgtRupML/Ycf5/U1U/QbCMFBCvwj48fCBQcLB+oYfwGf1T2TbLMzLXQEzdMODDW
k0yxryAiz8Duy/nYLnRrIEJuuBWQsWWTVFTpoHqx0LN6Hw0awE3k/NMyeW90oG5xrHS8tCWrGedW
KBLB/eyrDEI+nmpsgni4vrB7M54SWxZus7XS3BHIpXE8cD2f2CnQDwUjXTZ++/r87zJD7MYRIZqZ
W33lE0nc5EP+24aNyFaYi8m2x4WHunh6fA1fydcbb0tOut7x6DSNlZKq2ZNcnVLUgMkLquNGuN0G
ARDHHMtNdnhqmBGOfg/C/42nbFKCGgC+s+qu/ecLVQQXfWohNUqdv4EYZRJdcR7LWO/xaar4Ho2a
dCRnJFSfHxLqt3NrR96kMKsFRFRFbXyG2pgyb8c2HMNZNvk2u+OEF4jSvJOof5DEukTr+yB8KuQt
sagxvJsgABgztQ7CRaJ8DQJa9KaujLicpMoYdt9gV/jiP7WjApioEvdbAQzzk+zgt5MRz61Liuv8
tb2lCaaCODcdUM+nCZzmNJIZsttM6cSRYXzo9iIyawf+CN+Kpjb57KGg2cteigg8PhuIFyWOFG3J
mUZ9m7bZE5wCrk7x5uIu0yxdDSPDmdpLOq5M/UmJOX2ORH4gxqx+jPYsdhNvzgXTY10TyNCd71x2
xbKVCqLGs9RcL+X8DYeM9TGic22L9/4H4wrGAb5/sxeZhPTrgdfGbeN8HnnVXqEulMavBsbsAvzN
MS8j/VRtnlyG1xIvuyxAu7AGwAcRL7D6OR0O10APzs/jivPcclX39hMN9Pkyg98erxxf2K4cpHqI
IjIxl8QhSAy1MaUdC+WKeG51XH9j80gy1yQsWRV//Pe9fSnAHec4i0UEuZa2Yvhg1eshdrvUCVma
APluH8cDx9i9SlaA0iXmORqnn1hAe7jUDdo2M1L7AnZPN9uqn07Wf0ARN03BPKspehwfYecsUrZy
np21FGadtdVch7pMLQVHkUcyvFkiW1kAVAnTVSQeM927wNNcaAPWHjL5Gprq5UEq8AA8bduGqt1f
OzdK+gGjpJsr/3n5Masfv8pP1hvTBPIaQBxbj7bisv6Yi8rKJwM2t5ccqz7FiKMxqO1A4ojIM6p2
h/Y5Zre+ikNh19TUKhVVOXO2SDYQwgrw6Po8yy0ZuyEVwdF3au6dkjqOHIA2rKmxFaoJCZufCp1u
R3jWnGy/FkQfdlEDH73GXWcei4OwacqB8J2i527ArB/Z59E+linQQjOlp4Mg7VMRE4MKuEpSWNb5
6OwtElIeDES+RNC5lTmci3PxRVexp0wj6/qDqA2wlMLfp+wbdLE3SaB5WOjE5x/eZo2nO7EzN3BL
31YkVHCSxzC/xkxtpghs+wtlDgV21px5F9bTK61La4dk5EeixJeZhilWzXNIOwC8SSwsEgbbS/GO
bghD5UKFRAWcOMDhXUz+A0ASD+G7Z4SYv6GeiwxjE6OVif+oNSewbTa8UGTFEH0NA8zi1kWladEq
4jv57xvlMQein8k1MME3xq3PLwYgv348t/H4Fo+QGLL9WJuybstcBhxoEbdKgW1aiL0ysjqr+kVW
Z0lkAbmUQV5UHgY84tFxyDXCdFq6jeCCO8ZiqjKiPVjEKJnXSLGiSg1XbseJP0Gk6u36CR26UCkU
cOku1vMmcZQG7CWIkIFDjED0CTp2yOJUDVe+Qih/x1KkyRjs1fbC5lOnnNOliPxwTBlzhUMiDWlY
bixpJOtFxBfhOY/hHVCLM/eHFCgzsvvs95D7hihkWmHvU7ixoPSDnrbeiWaO3YShjGkusLp5ZSK4
Ta8phdnXK5ZuSFHeE+qCjKeGjLZEDUPdB6Vdovwy07NFd3hsyi+135vFM91qRTVcebQmjVUJLqkn
vKAvgqfSW7wFGkxLCdndmcWCdJ6jNvAsZ1bJTRKM0yPF5bPG+tJVTE4Y5I5ICCalMUSsjiZm27KE
dD2yy07ZlpiwNqPkw8poXvyP1o1g006siCMTtffdY9ocSikv/SMWBbEtYhiVOUNa7Fx/DxJJegTG
Yvubrx85h6dQb9Phn6h6CJVarjx6z2naKW0ZMk1iWflf/LH3bk+g0R3FlGa9903sdeRc1aA7S3gR
3wv+86S3Gk9UJgFc/OhcWHwnRXcBJHysVbyEgvrGlkP2nqynmtpQIKeS5cDcGbQFwjuCeTt8xD3V
EZAggJtlMxTSFk8K0PddTloHUxkLeK4vM48n9eKWQBC/KoUXLT42IUpP+hVvpi6Xt9zpHXGncLdI
xp8zTDtX60HPox8aHijvc6b/4IG3m0wffmSfe3Nlb+tjj3QiHAXWmgjcp6R4njvD1AyM8Xv0gYeI
J5Dlnfthhn0sqsBZi5RJ6JD9VtOyxYxfWLB396CktP5PipPEXnfIpgxfpbCFy45DTMheiVL3PyyW
KV1MunoL7KeUYtlHC/t4qMaNUg8KXD9xlIY1sqyYu1LZai9KklVWg7T0Nl1INbjG7nomAo32i71U
ijd3jFLd0xw5zpQOrtGLsTXJXZAGavChiZzdO0ReV6F4aXzrLAQGNlYzUUq8+f0b+fQK+/mywpzJ
0wkLXAxohrPzsLf6AaHl46OqbNOge0BrafvzYx5eemUd4HYXw8gmYDuWkujvRyFP8hSD1TSWWcwq
sr1g8ISYI0S76VweDtQl+OQENFS/R0D/XIDd/oR1CDKB+mxs+BNSAg+XjB7b8BLNlPvlp0oipn3F
+KWc3PoYYgTKex9bTDBkFIoft8EyGwelOXEDnICmDI16FtlIwJINde9b2N39zO/AWFBwdPXnWWa2
YExPDQRnwtfXwrCCieYGsDGBIA16k7rpSH641cTX8gXp+KDcY0Rs6/sxPTQLcLUuwM1wFyWrtKtc
EmcohNhyibAous1CGu/qBeIAfjMHz9Tlti7LJYEh/p0LOieQ9sqThCRxmqGGIQJ4RE3dqRZelBDw
vTHYm7SW2IXKlORWbDRidzBUk16EqG1JJiV9Rx7AASag5MjFbzxlk4vYexLhyX3k+w0UZPl1QeBF
+Aq4Bq1cPBnk9zXGx5htApwCmKkUsLxP61UVALSpwEgoTjxz5637TRWbaowdgW+lhVytLLvuIDkv
V/G3UTRW8d9p4eH8JFF1gs9cvyzjbCgZ4fY2WStBaP1BbO4CW+2aT+Ds1PS6nvF5EXRfDEP7lRbL
+bybRKM7qgTyeqs7yqqdqUo2wS3pQAMQ3t7LkF1Wxm/HmiTKLYMViDW5r4CcGWWwEEGFkAW/FEme
ZyKbCIrgz2dXo70igW7oUK6zQFhS4+bE0GdAfYejlqC7JYFolRh9c5EjEg/RdUjrphZHQnGPqB70
CLjM7L/p3HvKgWQ44GN9BPGYt5G6Gq1gHpyX/r4nCuhAo+QTjbvC55zzHE/jSfa0+wLdFjGs6gLw
7lvJNkSo3H5nFbOaTQKjs5xn3eaoErZgdqiN7u8QSjIxcb6S96uhctDNGfVS9Mpj1ItecJ+9tQLN
njIR0TbRjFokSBHF+z33xWMaYnVml1BDQ+wd0zIcgBoh7qhNbAA5tPMPwrlHtEPWBYrzzSZwTd2d
K3TqU9HpVmkF/CMM6dTuiRblQPc2UbyjDMZjI5o/+fuQHlXgiw+t96V6sw3sUc6jSUGQz3XuJoWi
QeG4AYdS/Y13WMUWMk0gaMDvmxk6+N/CA6GgvySMcqOGHTcds/JSx3lP6F5kOwNiPwl2RPVXxym0
jTnxj5ctt93Obc8xdCPK5/OSthNssr63noq+d/8vaB8nBz8W2UW/rY+H2YRHnb7GK8cGeGHyS1Ur
0o4nhsFpOZBUzrtrMm2/p235uuozna235LQ4iqh7bJGHmi68rv7H1PCGZkPpE0bWOZqnRQxCa8K3
tgYrEpoqb6lJDRjHksZ1GMRyn1t0zAAaBG5/jqPr2Yj3m4gmcAjwBxj/VPcQmVr+BdV1FL8rd0oQ
dFTXsSv028iSgry1s6mbqbvRKOCMCZ/2aSlCoC3oIrqIa80YrfN2ch1LIbj1hNKApQher/gLzLpK
pc2LKgUnDK0YhhsJWkc0OiH+MCWURJDs7GQ+J6Nz61p8msT8M1aCZK1pVelWRLF5KwCeJode9OsG
WVssgC5gaV9QBzOuD86XuJWCW23S8D8JVYvctMMbjyi4akgxRMWJCeaFOJUyMu8RxfkoSk+1rMSB
fofJizLvAxV8LrohvwwdzmHoouk0aS1V6ZHGjm7OaFBt3b1umFvw/EdyzAp8LKYrX6obpuQqaRV+
hk/p1brjbYC2W+7NWaN8F++APVOFOTIYtK3bYzNidDXjJ/aJoT4yPsMDbY9/Xk4IeSNITwjLwv7y
TjaVY0rUUJ10eLrWRUcBkUZIQvbaHz30eLgJFjSUFIBwNDSjfeUbPHDpNvNQ3+Sj6IGNE9+p7g+v
vSjQn+H7G5xD4D66xbeIEd7F1WO3U//Ev3BYdo0uzNQqk5pYRum8ZUI4f1P3SYa3oXxIYyd0sESS
hCL1zY7hSBAmBTgm+p3iTyPyLnzsvwOVR/t34aLGZGXm+ApVyhkKGgf5UnNtwmra/pNseKrkI40g
VuaH3OffsCO7WT+j8enKrk4xoPHOX5SU4R8LW2FmXbJTMbdo8g8j7m59z43RAVBTUG+VCDJGA8h+
SXM8OCEEYFcsyTjo4o9fWvtOU7eeADY/yYqVBgyRQVZycuzg4HhbKOk9HM2OBLq8lVKcEHVdj9z9
PCXYGHjIAE5hxOLxm/JoQfx+rkFC1VOmIRWw+2Th45c1l55tjKHH7fW4UbzLdrr27GluPEdexyrI
VUWFJA+6qCfuG+/A6EnpvWoop6KoSQbOhxUoIDLQcOzUfWTwPX+gZr5r7TgQYTwcaIKDbDJWlE/S
pgAnswAJ+21luRlis7kRcBoYzfgkW/97LgcyNI5S86rtD+2+twSIde9h2rVVBVu/SI6UBAVXaYx/
vexKDZAVWaFMvP+ylCsFNKXI9nu2aCHp2MFDfUk2fSpfgdHEsO8bWq2xbdcQdpUK7T8nuh75LXrF
hxlV56jMi8QWveVcgAgZlbA/DBNq6EqjVuw2IgEk6Savx7MCyRBtjko30ebXh7QmFzrSOiXrfcMR
tyQ01caT080caiMj6lgcFsF+UD3vtJH2aHiuG+Kqhgg8fYxoxu8gZkNjGEnk4okflCixnJrZKdo0
YPTMXH3AnA46U4PXoQ9u8Eb0nnUDoGFLKPWtju2VGWBC4E46WeGKAt3F3vpaMRb4FE8nAQRE+u50
m0FMKE5V3KBVDeLuMRr4v6dM0rXL3oNSq2ZWOpItTAdnGcbs2PVu9bn+AqGYQXc8axFOFU6e+Ao0
8vYJdRCKqH4vSst2GDRTSp2OTYGyFj7OcNFQ5cLQad8vJW4uaLqEo4dn1RY92hA+fWqH/nYI5BFL
aWBQDQF2FrfY+vWIG8R3MRy5wLNkwth/9zsV/BlxWLoG/x0BFfrask6d6n0gaG7umV0pp0S52jBP
zsS6oPlPA/V91ppz8N057BDg3u86pTWy690cHW+fxHHcYewmnp0LbJVha4YA8/HJ9uGL2I014yzp
A5sTZOQoHSpwQzR+wJCWcTzs5MzGU98WMX7KohUcXMW6ndhhPGzfiGKloRrklMOT3m17qXCc/ged
Q/JX2P/K5lv+tV09sE2BEobvEjbu4/YqR/3I7Ixy7JsQ48qUtXpIeqTBpQOd2wQ92flLYeeTPTYt
PUMzcensN4/BAB/FCDNTCQHVzH7zObtK2AAKDasP935+3HWHTxQGeP/PVwlhJGAeYV0/xzp7YT7Z
ZGBGcp9ToxAb4jYp3fQoV2HuN1wTnzs966HzaXgWfMEeTfHhg26ROMXKZTyzoiy0RSPrLOYfqCDf
NxOzPYznScNbOIGTxYVyxdUX4PmWnxSM/U6XbcBsE8t2KMOr/D+kl0JOGOyBo3HGar8XQvTisDKJ
SZCyHNSEBBBH3tXenzn8ckSbkvtFR0DJQc5mlBEg/UAISDeH/RaWgggt9KgZ2rZzPdA8GtnTCTwo
6SY5aiEWGZ9gm1BChO/mzeoBbcF5E5S8aqEW8pggq0D6L8TqFqrP/PU9mH3rk9BD1RmrKRcki4yg
CtB+UC/h4o6sob4ucv88rtoH6Pq7U8SnniixOIu95p8ZUqEBlffPMW9hJc63Rc1Sq2ge3eZxuNdB
jSKb8qs/qXTa1v4IY2oMLg+IKYmI0t6hRoq2/6Izw5Th21oi4Rdf7woXHDYBoE+edMCBeYDEl0Fd
MATgwlviaXEgy3XLBlfOCbggJeT7vQH2UooJmbF8782zeB8LZ7pFFrQlAMN3CoBMfHaUoPYI4DWy
VfkVZd9SnEH/Y2MmFJsV/Fl5xNODbl93SVa9a1QCq8ygXQmrSgdSpRmIHevStL1hmmFXqT8Lwse+
UIAwVAl2pZHkg/7247h10Mo3OTeeWN0uwUWBVNMEcOKp0V0PvybiiqBlQLAx8IdBhBt2mBc9b6Y/
b2bQ9M3PnSdRxANXsZ3OuW/cxcw3Apmo2MBGXlv1P53lSQZWcsxIFkbMbMUrjYwPTSHMzuo1Ntoy
fXTbUWAYmxPjYdF2LwB049reKcbBWMpAaInUWB7OayISlOXPrtYb2TJHy3MhiVaAXKptwIzw7k+c
4VFu+RX0WV8qOvBm8CSCU9+30RUxnEd1XErwDtiDGuec041fCsXjG352lz0GRKnN518BLmE0KtiV
tVvJ0N7/GJN0p8N0YLU9RfTMo05cv6BsGSE2T24bpWKL3jwHC2WJwfQ8sxuqgO1a62o2EyvF1V3t
N3xnwfZ/lup+5YwyE073Ta50+mZ0c+l7+05eJYhQv9jno54GVk5Jr8Zr2QDJ/qCnb3J6/IhNczGz
bv2801b17+sZD7yvuy/d3YQwHSWViAcxnAVFQ9LJgIR1XiEBKZN3XwmS1o6lB7gofhwR4k4Mr67K
AKnyOWpbMUYKnpZQzlOUoxIybZBDJaMwKrPBtF1Qpa+pWPB0jTNYidst+9I9JJe7NSCBhOonDJ66
trfQnGkxwZdzm3Q+BL2BDCUASQ6tSsT6M1g2pr8fcc0DKR3DfDoJJdZk1bwVqwuGUESPPzMko3xC
2UXZdRpl35rdsas2Hw5HYG3N28CDSMitEiTBDTuhRH4sKaZQPFMk4nAApK0vR/gVKppFAqhq9nSB
ZqPjb53gZhkDNRkeDOsifQ6MIlBibnwkFiZyntTsVQ9qjm3Ywt+cnq+1w2OtYbrn/0n3s1vIg0JU
p7Tw/v9Y5ig/j++pEuKLErZGBORGlene+TTWx7yeqKtka+JA/Ru1K1JhduAxo57fEqL74gfD4m7c
IAqiQso2LzgAM6MQRqc/Vm0AQUaHouooMsVb2T48Fdn7iMKIit/BjQhrv2POMCjxqOjdLN7RM2xq
w4NXmfv0R9BW2scg9tVE7Jr7esIxnmnI38SZ+VNrVgTEiirypfWdTrUM5MZN72k9kNLn2bjZDiap
T3GQ7qWR6nYcwabi6X28qZFdam6RaeQ7exnHDitlIKZU9ch6jKNxuC5KP2QIFetQVcRH8FthHIY4
iy6lYWk0WBGo4+OI/RZlhJfUaGIVMvDDPvsrgubZ9wyGMhi+rska9ELQMwQHzORn2UwLnsuxC+KE
7q0hsUHfWOBYQ++8S+TfWNlGP1kuYiwFzHrLLRCgTcqOpbpWXSTMlIeWOFpInk7bExEeFJ4HzEBI
nqi09nAirVzDApDbBFguPKiqGSYGdiWl9g6T9Nx7vIizRvITZ48b8w819g9V83KaGXSYoHAK2/76
0D0tJr0jKE7eKWBxhVijhGqxMGRXaEv3WkXfIQA3HbIFO85iwUudDx0E6oWMZvhPzRiLQ/y7D2l0
GK7k0/NDw9gWw/XSOy7j3wKk5VcNthQrhU8D+dHLdoQPpi636CrtLfuyy5a08NDwIT1DHfwZdKI5
0nEhYDRhRGvfQ6xHxPW6ukeGzUEMgzQQ2fMSl6mgIDzaWOdLtuluVl8GXJIyyjmYf3Y7E2KjPplZ
RDeFKpfqHFumbZecHn7uZL8XnIqoVH6Ovwz9ygufsgcifl0651rp7IJFz3L7n4lNxbO89M92704o
e7X8suj58rqsoRfKOKf+sjm+GS/8gw5lmsHeCXtfrQ17shmLGZbMJrWhCL6vLcQtefYnubpB7EgR
PF+7gTi9uMnbReIu4D8Vo1y/LRchNBCrlVmiO3V00L5asHuvZuVkmPpvqGRqRncFx13Oxakn0EY9
F+PmwC+Tp6630lpxU8MoAcVavUFC63uoYae0PsJiLNM4GLeq1Nd0y4eHKaLy2jxrcvV6OG/EFhPJ
XF97Zjpv3Vfp4ZQPjDJN7lIeoRgCeiTKusEjzfrvzFTmKrydQ6wjcrDaL+gKfHfqil3gFk0QB9x5
Tb0H9XSD41I1PbvUmAEqa7mgcHDNIvlEGAifoSkYTb9l+UdNMjD40sH9cugbkqhCrzKFjB10/cRL
n9J5BZdY68Mn0wbLkQXpHDhyIr3aQYgiWxwia/3B2ZJt1yCfDw1XL1sy0Eo+pacQxz8CpfLVPS/p
FGCBQL82iTTNVfG4rUrWcY3GtFDplaaStMmZiGcZF43nHZmv2Nm/bplRDQ5DDDWKM4DGqSpBnitC
fWrtmv4wysIJru7irQlcVcFJYq5iZp7aGDvrHHYmHJw0MlgfS7l8Wo/Hh6MatXT1EgCorTOlqyic
BfGwtwzUQ/+ghbX5hyXkJTpDRGvC9od313WLStTqrnIeUUB8wb81ZV5QSZlAPlG0yciaa/JjH5Z4
U8J2rUi8FmiEKR1ook+XXF24NEy1F6IJnSh0JSk/7GRq7VZm5rF1QTSzGHFRdsLYo4hatH8mEeYD
B4XR+PFCD/h5uRifH1THtXGiUgfVOlhLxvr4AgZpnuFW6xhH4W6Yy0xN34dnhN8zSHa+zYQSEjRQ
tIratAT1/i3HwX2Id1nVpR+0DJUv3sWEKrCGQGDrRhrn5JB9qHRd8LYIG5w0YuNxB65S5AF5hdfd
RY+quLasigacPAnLmyPrimqq8OrzlMIC4VP8oM5WgC36E2RazyRve6nYBqH5HgROViP2SA4x7APv
UqE31fbPFZazyW+bLdqQ/z9K6IZrDGyrZqakbItordaTR/h2AYiVxxFS5cR8oWv1Q6vAq74AzltX
oYPVtXdToey9Po399MH4+v546zr+39kry28MluR3ZPwUj+O6BOmNokyx++M44mXVno76qW0pmxHX
9DDNshjulZz7S94wMIaytn96Ep8E6p8BEGiuJEQjsbn7WFIws9u+fWmw7/yqDfjcHSwpq6R/KBKS
HvTDZaDbrTWAutTv55x3sneoCvLnEC0smsHvPZ9RPpdl2jkfsi/9yoCUPmdKgGbT1TaMl/C3vyHs
HWM4PGz1BFCjbicBAjgk4BubuoDNfE29YX1RI1kCMhXO6ATjNuHnqpmEc4YsG/s9/MH4FrN+hlZr
2pOYeRF/og31HBUwC205SuPz1Gmwu7B9NRMmCamAiMd2ePkOaq+NS7fA6ThwjzgYetaKZLpC6Aty
jYFulsVvtNrqnzUKaKCCusc2H4ZUzaQnD4aT3aJ2rmcbQI1o1NHicAbd2/ldaFL/Rhho08590il7
6EWLeSrORG5CuhmZnFyxtmVyldDo+Fes3H3uQksr/nemqF6cySyKiVNSl/hOTwHGlI+Z8ta/N8E2
nbELhOXD9vSZzxUL26TiEGOGmu4ohmQumjHRuGCfhS32encRaCSsWXeDkXEEs8qKJNKRBihP2gom
dPxbv6cHIpwuSYqaZ0RFvGtfacDP28pAEQ+bvtgNcwfJsxN3Vg7z6li1gBF/J+DwsT6rmLuo69q/
LZ47DzZLd26WiYmdenkKAZ86FBLbuMzLW7uXuf3VLqdmTAIzCDUYJeMn6sw3x8jvO6+f5fI3CFVg
2elbVugPZatkp4srbfabeQq9BE/lYRmaGi1vAXQLRL91OUKnU3JXDEO7h4enbUlklhA3y6PhKdgi
d4kMsZN+VsRt3hPS1tclvQqtsL5MHmgpl9xtSWn27ZIzLcQH/iLpwax+bXo2FAh0YeiDTtSG1fr/
BAn89zgK5QIVCb9PmUb5OW3xoyg6WaotpSGIw7ucJxBURABF+jASpXyag/71thbnVEIXWE7RA0xh
GH/muRXWsIHPFN32KDZ39Wp7L8pgHYJtKOE+i3tvozJcrTnfbQ5zF7cseaP/dRl+JDJ8slw/MXab
Ww4Mqw2os0xH/+uvUil6Bpaa2471jeqxG5WA114iGG0GX6f0ifkpIakR5jfK0UHMfbW/WieY7uCV
rD337E4kOo25ueFD5gV8B6GCLBESDr5Az27GDX0Uf0CgRx4gOaKtrMzqitsteXPeRTmkJDY0FqKf
HlxBKi8wZckvsSKNN7fg0h9++iwAlS9SZ4t47o1iyds5xqdwqLZORF2TCQDshdtlgvK6wliCz7z2
X4nGO0F703BRkUtSrTNX3ktz58efOtEGdumCkg/zW29kOjwSU5sl986+4EzW7BwQ3729NgBasApT
t0wCLS3ms9Pyncb+fYCF+7OfnBqL/JrwPPZhPWd46iI90D3NLCktBwUqH4Ax4w13gVJLWyZ6CBO8
aN4hOiILqoQkXDmYybVHfJgNPxGVaDO4NUHwa88DWwy/k34TGPDLRJvuADPob56tc8q/s5lbuW61
/yJ70ADIwTo28mz/eBGqKlKHV/d+2PT8PD3q2bx8zOtDC5ZIXhzh+rTL/rauwhEOXnFjiQpl8iPe
knWfqYkzxHzrFNJFV7hiRlIgUvD6q5+ilyzyILCq5KLpTOS372L03Zh2ORmvEk2GD95tNgEbRgA5
r9stVheSOMBsM613gLMQJzuk2qOvC+UOqOkbdkNm5xtu/83r5OOIKpJf7g6Mmr+aYROtfs1a98s8
vhDC0kLSOepBolLhjKDf0i4ptovIz9UbhqwP4LCf7LxTLDnc3Y7TY1KNrAVi15lGFmrjVzU/NyXL
TrT7Kg7dkrzD6y2mC6TamBm6PAmBAib4Hv1GSJP4s5RtcfEkLZPsR+q3PqCJ5+Es1iQhp8P+KR4B
3mUUScryLzqcoRx9hKuuiw69RQ6l1iSUdin4VHvLDKBceCaAEtpK1jJYgbK6z0Fh2L0vnUkKfjB8
c51rm6cN1LAx4fGLqL+de+YJbbZmZz0Hv90fyAMmMkydDvPkYWYtHSYSZCTBrerzlnUFevpWltu4
STzGBPgaZaMRRZP27GGqGqcoJ+N34pU/08ELpT7m+CIy215tBXwFOmYp135+Jaz1zyMqiyfw6QK6
QyC2oZ27ZvWdFmOSjiCVvvIqoePNq3q8ICFqSZWORIpFMwbeFDrezid3nwh9es3rOMCFOXxqB+xg
q0M5HbPBTvxgbOvdOR93lWUuNLldIGmE+X9zMXh3P6NXSqsHvI9LtTJr4NbLwMMdTIVlSx3s2KPy
rCr9D2TK4tVg9dZfL8lmCpqUsWSDksMY5M9Eq+MrQnSUvC7NTpIw+vrKZ3zwo7mn45IA/2yQBMKp
sJgIDbICphFAKkOtOsOBlpZPqrCcGKn+VNKnJCDpKKSNQhK/jjiwmDoWmmk+2nx2EdXuyh4OSxcM
eS1EfTw6bBfqK3r+jTa4gAHRuu/LXJQHBX68YsaDMXrMcMQqGaeIkMs6QjDBtFln3KaLu6ai39d/
oYtzZStL8wdYCe7FK2dboFYp5WqHhrboa/dkPbO/v5tPuN30wWGbx/2L7vYR5UCBeW18WZQCywi6
Go8TMKKWy6/c875XpivkEtxl/lZcv+r782Umo8kmRE4LINGuh4amBC/H2Tsux3Gu3/um1fMZRKNv
5htk/sglsV56/x6USe6eBLeUBk2RG5SaRoi1crMF+P+L++ReLHF8sw0qMVeb+xLqYjIr7/lwEZhJ
f+HpEY60wlmosfEkvTL1QvMqN6XLVkhZUbCYyGKqeto9jDXOq4YLIwDh91nuvUy44kozGBL4d8jS
s7a8M7MDWwRCW+ZStwW0UfokhrE8UiI53YIaZk79XZtOCRddLMweh7FUMyefRGBPU9ukdTp0DTdf
9yTqV3DVyPzRB1ELEuPW5k08JyB/u4OGfo8z63PjbVZjhsBZpxok8+XY6Q/5BTha7JBQOlmq/s05
bP2bU929H5vrv4qHbnfAFI9Q2IGza5pU0HwgPokcqQ5tbJDcjcCSkAq6MwIaceh2evIWW+yWHrHU
VbDxIwXR4Qn2LpSr66rpD3x3Ku4lquaTAPTTqY6qHyO4FuJxH0W3vrew3EZjUg3jmmJJfb3bXjd2
W+m0BOdESxfdqxm+oTK1NZC3kKjNxpI66WKj1jEDhGOLW2249YH2WbVW8uRXRqHcsj6ML5HXv4Wh
V4T3bXV305XdPHEnMY7cmMXhfVX6oTR5ZGpjFvela3axR65i+CRPExwd7Gy7IetEhk0K00xIOBgL
Fze0XCRJYJPTxCJpFOK9f+GrMlZKbdscL+BNK9DPBPOgits5FdQxHfTrPLxBHCRZMFIQFEiQAA97
0Ye37i85nuKEuifnRObuJiDModRtQs4Ufb0EaXzx2J8hRNpgpcNoRZ5JmOQG1d13IMoX7w+VjGDL
9fN4UB/8AKW3R/1x5cGClWtuAzJUAvmO7bmCAUNFWpFR3ONQwSlQBxbY4C/XhjkKPsGjiH0QDwMr
HA9mms7uYfQBB2JIEUyrTGWmY5Zy1kzMOcM8oXbgoukE3MPW9kWCT/dVvwWkK/mvsfDubcR3iA29
c+3HPtZd+HWify8Jf9BbxCF1W5hXiRgRDFuxY6zpNaUVr4MXxfD2wzg35SqMBmkgSTGyQ/FiA4N6
Nh5CnOBKQ5zjUaJZndATcNbodIen/Y+rQMg1iB/75qt3ZEGbiLz60E9LQM2jZ5l6768GFTI8bvN2
ZVFs0WiNGEcL/ciYHzHP1MJuue47jQOEPA9ow9Gd7fCJ38V8tOMJGkk8kzIIGl/5KnkGSYgwkbI8
VjJctKC2kZdKMsNDedi3djtvw3iKEJJA3pRk8E6hpXErssAd0xZlw7xb+OnUjSPLweW9YcZGumG7
VwBYdIEGh6qZ0HZxiDhrKEd2S52kZF8xEd1QsJ41m+mU5/J0UOlvnKcARsr5rdSeMp6RkXFQiQI2
ZyV5EYJUS4rh2bFhH7QP8GVv62VvWhoyfi5sP5wwIbor6t97tA2ISiK6lVZ73mscmUP9hgQajsT+
NKOIsp6nbM5JbTw4XH/YYfUG6pbxeWsh8WCGineQ7al5HWar46PZ5vj3cq1rtZ2z8XV6u0uJSr1S
56Y92V0xM2uQdepIi2pUcMCbbtVz/NXpTmX6IkTe3JBnpFHgUvco/HlqqetzrHTnoe9GrvRcVTMm
S28gQNLby0V1uOBCFi62nVwupEofpKvNYR+LHYlc6RrK+T0BIHAWNLKi7uPdd/6fLKM6AVH7MjIH
c+m4OhHN982M+CZh7Qqcot88ZwKpl5l/wUDOhEUZFNL9Mk1zEcTKJ3yQcNQDeOWPU7Bk/Tyu6qUX
9/B6qCfLNNthRGK5+GMD3Jka8L9A5AXhR3hlr0cfz4MFUyMRJ7RqY+77FkDH3AKlpSyehJ0s+Dpl
1eMLIZsElxhJZCO+RIeHCEocSrHI1PLUvYDn7Q+JhPB+q1N2GzJ5XpeaeFbkV/8GSq3OjPYAPA8v
1ppJ4pmHBm+owYhusbscj5HMHiuhtEpsN/8i4mPINd+TxlqF7JEBeNErsc7sjqyXa0GHkby7U921
bXKdEfK7e4OSQrH6cEnxaUd7LsLlqIEVydrqigQ0gQyK+otdArwfUIxUk4stu8DnZ5njuY/QCevP
UJrPDv8fzAR1jFWzaj8AqVl8znvkMKJ0ImFnaR6n3+KjYq1mgabIR+m6YIbOaI+gtnmRSrrTP/Ek
OcSzTL6dG1Z0IOmtYfGrFYU1LikJ74zwstjlCip/QnRFyaGTomkZfMbtBsmUVMfTyYJq9CiNRc5v
a65wl0RGd+Pz/J6vL89kdKPD9h6OUUJsyAHd/UBnPhmQd1UYoGFDZaOyPhfqk5n92J1fbeaa5O2F
wajlapfqOVLMo337R0wybqdybTfFEA3TQcDiYvITE7sssb0xkX+VeAMBJBNS34EVkA0yhRTbbvjC
7Goqb5Tj1BDuK9gf/sgNinMYaoToPUomLj3MV1aOIX1sebrNf3vNR2XLSQ2XBMUmH61jfrTFOIat
ifVec5P86ghVEYZYJ4+5GmTEkX5MSI93Dk8DaC7P9JSj7F/FbBgCFOEQ8YItv++dzBfVoEuVqXtB
le0zBi0etqxpERtlZABZIbWNAM04UPIF5k06Q8ZnQIlP94M8m3sVt7OMQQOT6TusSh5PmtL99ext
gxE+Eor25zefIh51uOhSWbdK0Cvr7/zx7gDzLTt7jdDyYKyqWa1sTDUc3aDvbce9nhYhwJUmhYxG
cobwjmGzSXne1DHIUme9hmX6eCJLDZSzg8q35jUsScIZgtT3EAjTN5veEeYYSmPwjiTaXch667Sk
OLkqbID5vgA6rG0nglD9cYh77g3NXrsNjj6axHHZN8GlEbDNjeWhMS5Gi0Nl4aG+vIHBI/lrEKHf
MDCXddsuaZmjegOM8BxkUVUGMhQJ1O6uhSyq5jdwCnhQ6JL/+7IOlc8zdMY56YpYSNOah2jEBvvc
LXyvLUo7tEncq35L5sR7kgGwO//df5BUuyWnIZtl3tMB95itA+9GZlcepWEPQxPo3tUDZdVN/G40
62MrSdkWhO3tMc6ahF7VxQpZ6bFvZZUHcpeEExT6jGP63yaPkcz4FZdSKroq+MaoW8JkBAzfI8ei
7Wdwe0D652agwP8CSY4UD1VTm8f3kGPZud17t9hpe8bGGh4Q2la7hExRpRlX4vviKBMnO51kTm2x
I6l8K2hLrz0yjaEwVGZt7fO68WZtcVYeNFIaYbqXolXmsVRVkfh50KB7jHaRvUSFEQ2eKSVs7Xbc
p5kjWAchE3kKx0Mlel/GMUBoGDlkj1hfFmNi+bXYegv2tWrjzQinoloi10Whps4Jy/CpneUZ2HDs
K9U86HTKG0EgUOipPe15B9hGcQVOdfyuMurpgihSD61Qb4pvPga2OBPi/B+/rIgzuG2Tk0HsTAFa
lHGWy2qL7Uz1AVCrtY5ixS1xRe6dG/I5t0UB1ZhyT0EE0CODJpcFO5Dl8lptSzAFWXLes6Uh5UvP
j4y4nlGQCLVnHIKxjkFmE6452B5XDt0jqSVNQmBNshaCYovdAQbPZMGiQ9jXBAmEMSYgKrNPffT2
tqTma7r6dfPlzb88B/wqlftXySPVirxjOlvvIl5zbPF147v7TeLNmGkXxijrgNLIE/id1+HJDlml
a41RTUf4dxwPhtTBEG+tj9fi7I4QfuZ0RkbsUplasroVhORDOSPjqXnTC7sW0FgN2F+2D1rx7Eqt
BFNUC/pbcgcPLTcDBuO7ITodbSWlOvewi3+NLRiZWktFLhOEku6GUP81WsFxr7EdKA4UsFz4Skmo
qs3aFYDtaHlwgmv3wkxucVbT0pZ+jiC4GJ1qmmniXU88tW3aZe4P9z9oZWtIPpjV+UnJcK9dfdMA
13ig7xbP/qq9CK6usO9TaghOb0F/TsSaw+o6L5Enq9silDt2R0JkEPVCcpjzxxjO59E4693bOTUy
BP3BqyfiVE9wP41KqN23/9HqVbBBdYwHt6JsOvE+fD/7WMzCMZWfB4RkWdgzwF/iAPT4BOYDulU9
UzLrmGXrB9AOSh4oIJNpNO+T1eTjDHOa18vgaif4JpxymslAPoK6JuivaSbvUGt6T2MTeaGmwlHZ
y2kpyp0xvRUSVxRh3bLFoIdIHEhUlsEg/xAZOgaeGLMuykWlNFpANcTSUD8xtFwezCpc0tu+qTZA
Kn/fgozLqm8W8ezykl9m64+bXMooZMiuA01OaxWlnnOzLNpN2FiwgsR/45H7VGOXqe+kbGew9ptk
zN2vHiiwXApKCmyQhXlQn5OmVPhCeWnfUHrX7LRvaAJkSGx7uuF80sjvMVO3PwCPvtzb+MhGGU5j
VDvD5HF8GpORilOwuIG20g9R0/zn6tsFaDB/jJNgi672urs9BI5wsIbVZ5jh72GjuFzWjd5z8V8i
52lLyFb7nJOUsB2Vh6tv8t49Jsgbh1efSWWuWOwXgQqq45VHS0s8efOefH6bgWJdI4bbb0gdNbkC
pcFLRUWgEX1lqZfAkEpLEPYU8I8qv5WOvTfZdLJhFc2R4KNiXxllzZ1JCZ7mkSTrUDujchtIHAQw
oUFI6w2Z9jkCCb6yalaTE9kPajR32VqMeN6SvCbv6PB1roURBcIRgxzMdbgmwC0rQOWsNvNxUPDe
J38rxrEZZklGvy77/W0tsS0Cn2Le+y649C8u0QcerAtw4n1esDpKR75s69bEBzcc4UVbLiJsEVJL
3BFASMx5cL8CLCn7ai3n6GkZaREfUmM/ecOEfuWChdaNfqVY6YKx58ydW6TpqxZjWtv+RnDLqHIW
e7brqeBg3mMCUHngl3zjK6HxhU4StFw5IWSp9rELBLVuDjxhiqNluAjKdueGd9mKak7bFMdwbLz8
TchpPeCugqGuopXu+KMDQu5QB7xi44n1wEmyI+cJEZoUahhsC+bHf37EmRvXVq3/iW6x8Kb+Sppu
qcMDPTy7KznBntnxpId9sv5dduXvButoIJSqkVn2+1m+8KB130K4itmnu806a0Dwlat2ws0nUyQm
ZVePz9v/QuREZROz+Je4vKsSE+dgLFI1CDKdeAbAcSZ/8VissSolWRgO1KhL0I4mSi9q8iTIaUxP
TsTX0b3J1+YLW3xTtfe4fsBwXc/iXV61ubLx1/1SK0uguhzKBsgepCqHFKsvCw+EZ5Y5bJ0YyqzM
9CrTHSElKC2CAcb7odwGWi6XyNJVGj5ZStCTBqxmSY3Yycaza1JpR5B14QfauNURMU/lDcpbgTo9
U+pa6e+8RifdRqgNDBBo3cTZzHw3UhPp3Luem6zMXmEWUfzoL+JDx6DZlFoBu3Thtl72DoCg4wXP
G+J98qoelI7CXLxTLeuCSrN27Rbki91Xd0y9lu9lwTaTPdvEuQYaTfki9wiZg0n6VB8LvTs2bNbQ
9jKkA//oKtHwIpcwT4Foada1v2PIakwlHNPmNqrTlzBdzoQ2lGNb6go/9D3nJr5IzUoreYIcTNQk
P+Ho72MPwFeUqtA/giYsmrZkO/VI89bdDao6d013z8inTwdtlfdlfMHSS4qPu/TReenVDpxuaMJ2
hXF0APxrh2gbms/1gNJ0VFxE9YipF/oOGbqjEfr4MVijVnElCCtHEGvoczA4zRylqng8Wh5XIEuw
cdKjbf0541FEQWz5T2qlCaiDDxyuoGdeGJNE4k6krjwBftFso7YjH8Oaja7W759fJiCNkV8sUhOS
7Nygdq1zdzCgerLh+wix/pAZkN8eoh7hVzqmakRBbfUI7mzTpk/EyJ+pkKyoxIEoAhV4BPUx+Bxb
48MvW4g3DH1KnSSJgXWFUGLDsZ9BWcG4yRV3VpTgj6CVgzFHoivHj9t61YNcc8jeBdKjLyHOm192
WBy3PABTjg2Qn1tq7Lc+92/caGran8AZVsh6LR3lgVsY1sNGGcdNd3VMbUqVYkKQALL+lYy8EbyK
IBQlm1b+yVuXbHzlM1K4RQuOe5UEq0ahzobHYgcUcE0eaFRXXxOBKy3ol6q6xzYVb6oS/5oF3Kx6
D+qLXZMe/XV4aR9e0Szh8OFL+Qa2+UFjCIt3d3m9sUCw+TMEySztXicK+vJ4SBDysPM15Sg/HK9o
Qx4hfUdyGTewkPpWtwDhUHO1Lat0r9TUQWMnf8pYCYLxek78EobTvuJ8I4ZbbJ2AezMaFDXrAmDL
xL8CST3ahgt3hzsYZeuguiTENij0qQu6W2tEbUfq0HxbcTYuQ/mbTpCRGRThY/ThwVbfgH7BOZWi
7Q/YuqALDgwGLcJVhUlkxRKyqPYU6on0F2oZn/egse1zB1FynRZhqHYa+lt6AsVorMtdAADgxBB5
daIBxFpSY8Rj2tnBiHFRvWSJxWTA8JK17VGZEPvodNNsNj0Tk+Pwer4x9HsNgzPgWyraERCvM0Ys
nVJ3xfgtr076IA71Ovty79stHJ4LNV4X5Li9K2KAgjiYvDAUi/X1tyuGWfaUXYu7c5Jki9HdpUdB
gvH3EUFDb5GOlk0O21v+NgZg38JE94YvFoxIKu5uhZetUmrMSm1dCnqyBec4DjjIbLCJ8u1kHDWo
F7xL42LQ0nuBhE8GdWz1MgiWTTGj4pb7gggO+17OGx6fsFELAXue/m2enoJWsjwLmHKQZiS+sjXJ
RlOyF1nyRY91qYz0692gP4R8S4VjSgcsryceoR2PmQJtkAQbFnnfi8k8rzCir3/9H45STr7lzJMN
YydrPnL+zZMYACInQpyJi3aQrcnyk0ClSyMC1eIKTL+jPalua32Gd5U/G9kdq/jNeZmyxqXxLpTR
uHZshejHUH3310gB/LHiZbWLTwDMi436b1Zlow32YacduYUmFXK8xj7josDAABEM/yU0OBS1QCgW
a1BJlzZv1EyeJseC2dcc4n3fq+wd7PQpgTjDdfdbQTh4QW5+b8LYBttJPFw8K0xJEIakRz4hqWW1
i+eukdbO3AuEkUr9By5KnN6jMf75bmXwXKkJCOcowvcl6pOzH+XTdSaOSM5Ze5ip2/dK/TH5qql0
5VTUAANRu6EZpRfU9NuECoHXjAnCslMGLQUPfl0x2VumEw1XsVLtE6DseCxqxvcBoQ9LuyebeGHB
SSn2X+6+iVW7XstMGEZ3uuOhgIFio6dwDJ3sxaVQfQXTXsQdK8tBcSQ8/RT8bqsf9BzIhBQrY0Ep
BVIc1TlDJIiAp1CEtwd7a7S+cJapvNOmuc/nnf3JJxflVyg5Wm1BRIZVZwUCHEzIBcZSl3f20rr3
SI7ix6P75yWwn2WU/bnFq6acVjeB4KXnAK7Ke3EbZwSWXI0R9OIkneSYYQqDGCyYX28yffQqincM
qeLl80nqUSFAjDsHfXJlPItaCCv4mRsKUNoYncJLD7Odyya2jfguFs899wQdLHDsnX+XHvzLmnpH
7r0vO8Pz7NJ2pl4jusbVYg8nG+0uRY1iZQZOEd6BVwAmLt1ecS7gdBNAMpp+z2lErWDybK9qvQpM
rt0rHsRdcX6ufUdKKHhCjznifMCWfiqHzfusDW+UgNENcSPu5wAlObQ5wrZlmiCu6OOeblfPQ213
EioNctLpP3wQCp/eHfD/hg2/fUn8eFXjCJM/9bpWuD5ZzLHpeGJjsEsile9gCXUamj22pnFoFGgp
7TTARYEc7hxJqHoL1zavlHnRe1PxzS60ldv7MvlbWUAo2sC5gy6Vej9zhu5KEkiXrV6k4T79HRyK
6Q0lle4SIgFmkiCaM0IVMLK51C3S5+niXS0ANd6FL5AiFp2FFiNHBa8JjgFSuzDGt7vAtVufke1M
F8M2S5Dw9u12S5e/WES+6uJMO/aZ191O+fZE1u/3+y3+1JNXcs8643W26hgSQMWDygZ+9iDpzlj6
4s33z8HU4DvgyYUWsDw4xjAUg4C6SeXwa8GiLPUWHBkGtVIO2OtK/ZDuZgaIBcAKfzWW7Yv3cEyK
ZgKqr4zg+A1IdIS2BJQEJVS+hZ5AKkRTcc27brKvop/pkib9l0AUOMpFUML1kMDRXzVRRGdmuJFi
ahQFNOzOI8aoUlmCPVqWAafGeY2WXti1PtONjD+YESyDQB+WsCQjm8np10LnsA6GomfQr529f2yq
yeNS2fOKLPiX17E/5NxMz+OZoGAGvXD3MCAL6YxB7zGxIEf9HX42cV1ZtNQlQtyWQyfkKY260/nd
A4BpIao62ZrD6hvn+nFcLwBoswTiJwsx1p3iiKwT4cPijUQqVlBIt3BYjyLZeIJ/BqT/K+0Ttc3i
qNCwll7/KO/CSGDlIyTX0dZF3XEuDgfpthciKBIfGEXlMg+eIPuw6N/MoIEnDZ855aJWKAFe05++
cpmoGq6fQEGX0I85srNJkJH5w582ilBz5VaqkP0FqTZSPl/CFd+khL0c/Tmg4NyhuCWMnQu6xrHN
EO47SR8FRfEnBqd+aPwnMkk6I51Hk2jeJT00OOxwLqK69IhJjxieMfMrKqb4pprVRDvAQ7wN/Jxm
3pRyKdHZnYRfal3hGlp1L48x8x04YJ2nxLm7e5KIhwxXC180toaKLdHWGdraRbmSmXsR83geCc5S
eFvFgbLKn998ZcqBGyujqnomKUkvMvcN09wWxqjp35nc+SZuWVD7JQkeyrkdUdQJrsi2EZL/bh8N
UIK5qs3RqHBqwnl+bRidJJEy6vWqrgERbqF2sAvcdkcsLXv+Ciwuf2X/0oZKE6havOW0c/38/tzs
nLt9FrLYsvspjknm3kMSK4XdF46lUGMf2qHWJlBtrBEFPQ1pjp5t9qcBZsuDY2SjCR/xrYggiLg2
kW2+YvM1VTSV+vdwY5L8gWCbnrI0cL4HM9YGJ6wIM3V9BxO/954vmy9PgEs3s5znT1X2Hf9roblS
WkbLeeoMXiCz1mSkA+v8L2GwlJh95Rincfz+Dw3/gj53LlMsX/JRj7JHTHcXSKBdkmCsbtdpj0yI
v2XlJCQC9PLnda6nU+Zeq8a0HBJ2NRQNWg+S/CO8XVJoRxRFoUBRYsQkcV6K24Mm5ixM+P6bL2K8
EqZ2VFRrSHSS7UMRnnUoY6wlx1t3YsZpPQE4AphtEgIFpUEdPp34gVnB78Auu7IuBu/1UU2MXr73
m3Yc/xJKTIvYvbS+Haao4jJvueY5n5INy+tuCVuek9/J3ezgpFIOm5/QVAR4FF4b63Ke6MsrTUq0
QPEjlskHb7Yo7qPbhetNIvuaFRktACUxaHjs8MGizFl+ZwxI7B8b6vhwhV+oH5nnoA8Oo6LQfpq6
uJeSs+d+BGIvcqy356BKKX8IUokKcTg43K9IGqvgnL56rKGLSzJ6Z6X/7F3hg3LFXw64HZCY7vKV
ZlKCSJIa5XOPn8KwhZEJwnTUOhYYRQeaQO8gaCvmHiq1X76Asm70HEMQxlysFyjEiXnOabZ5SR0+
sHZOdRdYNjmrAJkafgtLPl9wqRCQSUpg3Jpmf3N+Q+c8E8zOtrsCjgW9O8IKYX1qaM4xPCypdL14
+/hfAL0FmEBFTLNTtj8SVxvRvhgffD3QFnmW9whMaWg9+nvUFDA7e9wB2w2C0jlCSrK+77bDsy1Z
6OsW7DNBKPCNrUDZ+Q6fePKRCnIUzVEU5LXHJ7VLBv4/4qyd9Kd4d8VsnQGeqkpPvyxAqrBWOp6U
QwLu8dSRRvUDNH7FudCqYYCvxYQ8+lVAYnbXBRjgM85AGBDxds+XIjk2/cbwiV4wAl2bYkKRFys6
kjXLij8RfV9k2jH2pophZPYhZTbgmtdrVrl8HvR2mnr/RjafsMTSHv1RC9wycJiV3leJg82XxZEC
cmV3Hhf4AOVaIvJrBRnXINCgBioQn5mt2P/nx0EhdlrBSdPPK+764z59eBkJ5m27s1fgv62Nk9cf
gLfYHa2X5aUcgnW4+96NoY1cgJy/gG1LT+jjNxpXThsfn1YHFJBo3Hx9IOJpU8ePG1gvr1Yk/XF4
4TX9hrWvIILJjLRTFM6N3Ra6OyUvH1SflIJB6b2c08dpyohnWGPyNHMbtUos6iWhnOfGA4SUixVZ
dFR2DByjOLU0JFLVLCMCf2AP3qldN4TfsmQUIp6zK8mZK9iluJhABLaZtrmsR2UKJTVpHZERNit2
P7/gMIR1fsrhVvXPxly/zZPwHsUI/XepGVnwdBDHsqroQ8l/4Bl4IxOdeb8fCWhYOfndIbjS3jiu
T7updphu0uvfOt36bYP5lurWQIOT/OQeklw5MUvzV2/S8HxJVkyKgUZxlD/OMkfVy3n13mEumJB+
xMnhzcuF6ivpzrpcRndccRpNeaOG2Zvb1SkbMrzz8g8E3a5GvVNCgLINw3S2Fuk8iSuoli2+gXzu
hMWVYgCNLp/303sFP8j2P0ueNlgC9matD7PXww0WwoxS+QF96bJlL4ER3W2q7aOiCsHNI4GTrEBF
bqce5/9xJd/Yy3ez/GgUmJAQGg0QAAF4/eg4WXAo15Egx8TuVKipV/Frl0eAslz2rv4n5DWhmTf0
P4wwsRqr11rg8DM2MUM/6K5gKOydmtrzw6Jg+5hLbzLdqC4RZKEmVqq65l72663Nu1TQaX7Et7Qo
X97xiBx5/tcJIkODdDEK7M73h5PGaFxnKK76NN/vth3TBnokiH0Kp7oCCun6WsRvckTxQPETST0C
Ksj67okI0Nace7tGzmYf0OAAocPZ5V4F31jN5SQ5STrD+Pk8lJnN/cXpaxyfUmyQCtaZZnqE8PxX
hjIkUO/AZgpYqwvlIbA/6uj5ARs1KzpJvSI4jrGyLS0ze7oEfWIF9tp62NfwynYGaKT+YCblUmXq
IuIcx3HFvjzXx2t1EGmBzy6kvJlcN6zsOVkmCrpgdCptjeC2hIi5aKEZbCUooNoFjI75i3MLTRhM
qZBmO1Dk5/ZyYnq177JLOL3Pgh4w8fzgXF6rtEvR098uXs8Gcr321qLdUkyrwSCR94YyH6yLQ5c4
W+Yf7IDAub/ON+/gkF0VPG+zSfzrRNivRmLQPgZzTQOpuW0w5hbCgRcP/DXjNz7iVjPnbMDH5tG1
+HRA23f3XL1FKBhQi8OxKM+NY+Ld6Bm04I7fzuFK3TA5dITT3m1tf6jxhOYUFO65xsqiHOheGRmr
SXVyUwGtgixPdnzzpvTktiGbIw5H8I/7zvoZ0vFdRZiqYkI8M2LB3sNngUlBRf+beH3ApPZ4dq7O
25688CrISZBfuzODhhY6igI7AkqiCLqt9llQlqod4AzZ88mISyY4j6lS/B8L4ZjOW+UUEMA9wqwX
HMxJOeDAMCTsFOKJcwyTapRC7DpH1jrrgLmaZo3EjLipIbay1Nu4MuMPb3ICqQ7qAZNwmNh4msq4
6du5KxstmA2toZoeGj+RCNRNwXb8bb1FGrHYKhJ37ENJNy7TqIcdd+YAQu8BpK0sxa0MTVk2jM5L
zqrmH5lweJh6TT1OeFLjmAR97POItllU8SAQAdhrQb0G0NytMSvLmL2SgTeuSIZtI8UO1AVGlY11
P+fWdnvaD2injgUHSDfMCyPK1OmFgEmDFNKoRI7JC2wzOcS/Aw9Lu6MIOi54G1iXiYypjihF2tmZ
qEiNQerAsXtxrUgMZ5P7JpgGFjfic5qUwKs5ZMe+tiFovfjyz0jLRgkwykzb1UvciN/Agjebq71G
lfUUIqALZ3I7pjFwLVEcwd730pyoPNzuY+8JyRmTMpTbzQ52bPHTHIoe5UwZrFI8U+wQOFwgtveT
YVK3E+soDCeL6VmoYfr7dPa9JKwO5GVzlUCSs6wZ4irBH95+xiBLC3702c32LJzwPKQim5o5qDW7
+auXXBtvDHCQdsO3IcqF3KFl5oyr1OzHqpYXSyUbGKj5u+0FEXaeqN0Qqf33sB35p5Ll5IujQAJI
/IDBxYrJhD3r7iAtZq2nK6QZU+i7X9NrA+xee4AV2Qc62BbGB0TitUcwHzDoCREMiwtzbaPdZpxz
mzAomU1ami7FHjSLphpfAma8E2nqN6yhorQBIwIsd9r8rVL4sTE7soSrKBKg1Q16nNl6pgESyl6a
AHWk8txUfHES0Gu/nPwvaGRQsuEU57GGGqQkFwQV8tLOfLYEC/g5RGuwvZvx05QCwGVXySevDOJE
nrSVtResFTi4jmXICXdMrjO7dLQgz1cg+abG9R5D+BQDH4x7WBFGAohNLuEgaa/ODwDxoPH/J71I
tCUkoxc8387vzlDXV4+LAuHmQrjSy0COJMe0SdfdfmhTpxMsc3aiucdTLBKfqG3H6dmFDIONTcag
8GXUjn6nhCLTR8OGU2xNXTj3cgDYuU8p87qDiQEhFev6vRHAYhFU2vaCcPq3l+DZHi9Eh7HgYVVo
3TQSyR0NNZtSvOFZkwW/12CV8I2uDamRX4Z1TE1xeO6vSiKkc/9+NnGIqGrjS0QoVkNSR6d+r3gt
26VFc80GVTapsvWTVMnhGU0AZEtYcuTKbzV49Tr2PFe5VWAOSLno98jkQQnJ8UzaNEXwLrf52E/l
iwdWBDYTgfndVWeQyO9gVO+BYLj/U2YrINyqUx/X8xHWBk01KF0RhxcN45UUjHRnYZ9L131W6jp7
l+slKw/uGXcBUeUXlp+plbqozSY4Ke98osFjTOALTFlLDsts9U4rGwQpxpwMIzPhAV5V82+LSD18
OUkZUflwMdelCvqNKm0j4H+H0sSufHdsY7upkxusUtKyIwLnorlcP78oS5lK6eEASa7DIHNfLzuU
GsspB/Ucm9ZUEFLYce+XfHmXRSk01GrXghSkzD4KT+2TwZbtRxFgBk1F1iAuQK4bOjkB6HgaL5kf
aP+YDtwZlEGe2Zv10NnNy/eJ7JswHpcKsVQDd3HL0ysEMQJsCTf574+CtjizlUFBmCYSlcW1tSBO
BijOx0MFPD9G76G9evhJ85lyBt1/fwNJzuu+TlO+Gt3FpNqNc6+73p81AGJRuS1Fx+aBInho5eew
XDzqnond2ut6vnKvsBX5sK5RIxUux4wtdUmJinI2s394BxLt9fQht42I2FD6r0U6mU/MryMBjcOn
/i4efjQy7UlGV3cofyl4NG5o02EGugCJLaGFvy5ZBTseVG0nXdoA8YkFjPMvoIajVHgBJOVnGdCZ
sPNdHjPMHIASRIELz73ETgYRMEot0g3gQ7+NYxn3V5GmkCu6nWOiUAN7jIkpMI+5D7rcPEGeJqao
Myg88taYXuhG+fqKmAQwlseAxLSXMoIuZPBr5pSn0wU8HiJngNCMTBFb3EO+IVzm6LK6syf53zqW
IUAIew3WtnLmZGn3dl4L/HmvbZQvvk7OUJJqAmuo3NfmsN0A6P07KysaQEGOZVlZw/mluBj7Pbwg
jxfkkE08U9cj/vD16CD5zSbnRBU83fSQKvddfdYpBBZpU68Kpj+HcEAYhRFezORElisDsAzLT9p1
lJkWYxO/gv8a2Gr+U61dekmyn9kASOYdoCgMT31YHyOGszLmYH4fB2GAsDmGiupeMB1j1eij80fh
YW8bIuraKK4805Loem5Na3zrAadxIDrt2XUIKtP9Pk69qtDtHwbVNKw0FoEjUA6hjWxt68eUxtMH
zvpXF4ty5VufTslRcRItqgGPvIDJDDZmIipDC3Uge5uhmOb+ztxfreJPgRHjFyUHvVP2DC5VjEBt
U9wTcvhQVdmQPvNj6v/Rz9EbGYF9UT2NT0GmmQ6gN/6CWzmBx3cUVDYDEa6T0Z71D5fxFYj+ocIv
J1JsYCv7GkRh1kbgy3rdO8/56c9OeF4IChwH95MqLXDRMAUahHR2d9KOphzaZmjgAyBZeiXtvQuW
pbPBY60lEe5lF3CiDDB93vxOqyoB3fm031oeeSBZYsOs2aoE/AuHpijQKUsFdNur1zmj3wAAx633
40ZvRH0DkRqjbcTyBVuWE3BLP0MoTx/zxrgvmbwBXby/ne232y4T/wkmIDdzA4awzep0BOe6YEiy
ADny3RbQepjtw4W8h65wHr1sSDJhMx5SgaPrMfo7YUi6Z7lFW7xC6JCn24D2Va8xMBY2cGHbVS8g
yDatFueUPYrP+dCKBVRqRVDPRe1t6knB5oNdVRKKm5y7fTpIRUOtrokhRfl4lodCG9ghYu14/xfp
uMKwdpLauIbkIzyRkSlUDWZwRtDunnrCs/OEqoeOq8ZG2Gq8aiRkMikJAOfF0b/TLhKhLwy9OH3p
N4SAvR5eF9Y0i/9xUubXCnoAwlcuyCRZlAW3KbE5yKMpZ2S3tQzykGy88dK1u5QsI54aKMuuJlwx
mC+jJwH9sv304L+a4+mFIGOhHc7rkj2jFXqH3yOQ6uySNw9doDdT9nY2KbjhEOs4SPljt7MLVgOM
aAbBTvL7R9/q7484AI13qOyBT+gkBaxZMEDC4ic0COu9FShMddajXzqBGu7V2vuPNQm7epZSgPZy
F9MsZLgom239pSlOHRNzN+ufK5BSJTtfBQpCNH7zh8vbmwASpE3qCBxhaNy6j7ec1wN96SwhI5/q
S5hlQMGJJil8EV9UJEYzlXTx28J9xBZL8qwlsAHrI4demu2SfWSjmTuhtwrkVxwO3P2L2gq9Ig1U
S2A1mjC8+/6rvbzwrHZbapM/FKPcPP/Vdk8MVyLo83VxJH5/kaugitBPCT+wjhjIn7fsiR0cH8T4
2M2SGuWUfalUMVJ6A8Q3CPDLuflGOyLmH6syGrJjok0cxb5Dq+yhJyOGt+NzBId7hZ9S6KYKtYVa
1s5R73Qp6bJa6Bie3O+b1PDcqAg3nENqliuAOK4VvXXCJeeVYNN03gwifvHGE1cliUAOTJwqq+Lu
xj0IxPTuzCZTALkbOhtzSiJgHtomZiEOhaDOs4zEi1Vkzd42NdXmyhxS+1u/zoM4M3IxIp0L4zGJ
oyTyVVbk06359xPJReEhVZR7pOlilph/7o4V1iH6ks0MeJDoHihEjtA6W6CujgKhNPlNFT1FTyk4
FSaMtKg1MOghTZMxtWB+mhOokd1YoJRLZwyjoul+3oZHUo8vd0SjySEsOWSiz5RM5HhKpYOwcpRo
ykO+bv0DkWJ3umbp5/8eaFEz7wbzmsseWoOLMTCbOz51SftMLKTs1UATxpfdTvRI4HVvR3x3Jc1R
W8seGFxenbTMio+KPxxDForjuHRxeY9W3lADdWSLryx69ovtiLaaEQrEV8CgSBfQHMjydiP6Bh6r
Tvi3rjgIUnbp9Np/Uj39sw+ZJ8DZJAqv0oED9t5Pi+t9TnqJAoIXECx6i8112wE8IH1DgVoRtKov
nszQNtWL8Fq4dK0/7d1AlrtIfLMlp1PdfyRCPSl9HM/Gn49DHJ7JmFNkeLJnhGgyEcB5EYGf1lSM
hmAgavLDc1XWHBYb4LTzJzOsTB3X5LvYG1oksD33cuKiOtypWIj0TVIjsyH8xnqmXa6gFioYFsFx
ODTZtFHh9t88iA9GCI03HiSXQWdqAAPc3fEtIMNqXUtw7JsTnsjh9E3PkyXW6fZAMjMV6GiP7A3Q
+vKDLnxJeZ59O5CGJO0XnKP/79npwBsTeqoikAWYW1w+bixIB7nzomNh8p6cQMZksZ76IznD4JKv
6MWYuffSZ6cyo4MMj2RRYls8wKPxSMJGCfeYgBjrJn836demUIz5XUcbtTD3T9RDsNAxn4A1LpQz
qZUeR7OBDca8UZSxoVSIG3i9ogBerX/jSg+RBVNpBVS8jQae+kpO6bIzXwiASIt0azFyozcDOnQi
vPUp4GA8R1Iw5KtkmSvQmoDrqd9ySVT5wn5zx9ayX5VsyKLwm+BUMYsPub1FLLGNV6hjyGvhH33S
Kj5Dq9G2vOcWWh3PNnXw985vgkrfyOLaJ6BYk5Go+H2iAr4gWWNY5xp/lqmP+rAvuKWcBzoBrojy
Jy1yvrABG+oEGptxhHBIjT/Kal9AAdN4ImOHcCX+XJ/xsxvEhsEkaXNo+4Q78uG8ReXZCdTVSjwL
ceVNm+8x1LQ7EnP83xjWHnht2QgUaIJnJT0UBR4dgEUJ2eBIAaXgaL/ph6PAjQ1rJGkshjw2/lOI
inuZdB6a633R4FcGXTBqDh/46mcPUUNHsvfZqiNepJ/zUhBAOr3NZANN6wusI4a4PnQwL/I+rO2i
Sa1W2rniAEALgpxVhEIV+pKj0jiHiwbjKiMoVgGn/Y+ELOWNv73mDBbxVaJ3w/FOnK2zayenQVhB
CBru/4d1+Pqeg4YvtVPC/Y73IEcC0rMhuBArcMveRUkJD8Kq61rJwJiTtMipKIzxiChxvEAjYwz0
C7JLUdrgPQx6EnV5kYQpjg50AXNVHbu7ErI+xwxwO3LRER/dGhzZ2Y4V79KLDVZXe1msqaQGfHuj
0WD2R+c20UIdQ7Zs2GWEjtS9C5f7wASsm1qUjZNNsGZq2YMXeIKxSLHRvK+BMjVm4oqhnYt31Q5r
qeygeimH1KAhehrymwJwqUH2S6Fre3BCSk2BZgqBvvg8IDCdKtXD6Xu6rt6L8nTqW49FtL12Gnxh
NM19m3SsF2oCyIP/b9XB37CrnQByJScvYmBf2zLK29fcHWhYu2rdJOSvydfLcz2rxB9pKejlvR7V
lfwwE1KnwEdyMFaDdK2YXk1u8UqQbcntfZnSCigacqdj3yil11uMV3daOQGSWsLM2QHXqyOldsCh
oVLLM8Q+cjCbZxs/imO+iNoSLGTaw+MA4jiAttCWQhRjiaN69YM+FXSrarF1rOfx0V1HtYtSg+om
eelpKuBAAlnBC7tCgOpHo5B3u4KQTHGh5mtHo3TKuTMU9J91QEbTfDx/RYHQD/Td8mloAh4VzopM
Ge9g4NcTaQz7DbNlCg8VGVrcggJkU1DKzx9uMFZti2/xqziSRrah62cvIt/whQt2TX8aVKqJ07mI
0Q7V0XLA+v05Lx+R1Ayah+RTy5rh1aBgvmj3EYQJFGadwRSuSjMzCchuh/CQvMUStgbsmiziNuyx
JIEdFNI/wZlruD7SWTtS5CVDzFISp8gpu7O23s8F7uWUq4uSec0F0IAKaN4bE4Nvl7inEK8WlWry
XdetqOayromZYbz3ROjr/ZTHvCC5da357AE63No9ZCIAYzhO8bAfYCJltbdykPdiJG1gKRKHRod8
uVKN4wV0tJUa4RxpFdInot54EykztZ0zEzMcVE9lCnIsEeAbQwLK14XLBCx8rPx0cpgVMfuUpbLE
WbdyB+LWEzgtguVi5417DIfFtrDHGWlCFGNG0By7lYNLjua0nnhxe5ipN5OWua/DqwwXvy+5gDW6
mMCrUi/hgbEX8PT8DrZsghxQINuqzuFK5u9zdVKn09SeECB3VBN2mTqMK4E+YMNh0fKj+KFK2Q0K
QX0XUqXznVhGcNE0p+gEy6j6fr1RFf6WDFMGuG+i4aQ2Meq1t29iVDjMQT5+zcVEJz1d65YW5TPi
VC/kYnTLfR4IxzGauaZYlJhYfM3kcB5yvhwihWB9g4eOR6uAWME7/FcsjToY2RPRU1MMEkFds5Tm
sXBUpoj32MxbTNbht/sBYjspFowYomQxNLOfas7ilzkjqmN4OlFl5Pr7DiDre5BlwjUbUpeFvxcX
B36Wkj5Po/SoqCPE1IBidmen1ZNaOZxC8DFIk9CBEQbgC3E5Vsm/jmw8hN0T9xxsBXgVduIeF8u1
eTCg8bTNXt1m3i91sQxZJu2H4N7bQtP1jElR4W9xwyx70vFiyNrNmN6l5tbh/YLQ+DZjGP0fOWRY
Jks/88mDcK5VsEKoomkavSCYtLY/xXLbb3IDTg2u4xN7YQQKBDlX8YYnZfhVaao3n3mT7uYOl8dG
Oxt3q2n9clmC7b9qvXe/7YqEgMfderRWqXE5tOOca8WodgsYiTla/jTz3FRBEk67BuoiXp5AvQ6o
86ryraypPay/7EcXFCygHzeATmmzFgONtaOqrJ+b1ljv9VTCuZOtfpgX1xgND655qVTc48/vGaYo
KAif3dtjV9O3IHVy9+Z5tSzG0KzfI6JP1HzbmyezUfB6EOpAY0SAV014aG23FWlW1UEl68xC+x4I
Bvwgx0XAxQgioSNYCoQXSoZA30DVzBbmh4VTVmVd6Fw25Qs0jok2entLCaAWr2C/+4ksdtY/dNrP
mskuvDF/QTaX53BApZSCtGuCofmj5j9vrbt6z8682X0PJTzTo59nY9kUu+JYYSrokS2EWTj5uwBs
jDMQDNn2HSr+QeTvHuzWyAtnZFMoTHCeiU4POKyj0Ib6kC3wwCTzZrnojKSw0asM8DQT/bm/CDZL
IUnn8woRZA3jfbajqKUW3Dstph7glj1P1AzF8YpZ3tdKsdEEOVxJAZAnwVwpZNQoL9Y/yEyV4aRo
8RVxsgf9sbDFCndrILwoUreD3NA1kFA+y2EtEUpSRJSEis9JNC8dYeLajsjdIOMTYBhwJpCZNYdq
zY57D8ULPFugohczk8PzOf217a3bbiOW0dndMstt1zUd/JBn+wqLgSned+sgX4zWZw9ImbN4VMmy
6r4TulgOvegfkCDKvZjG8568/kCb9uu5ia3e4LAwi9x4U3OFRDGaLX6JNduDM6TKWa5mycL5yhDW
Q7ldRvuFXdwRxy+EQvEonSzsSD8ewYXhBDF86o6JUoccxEoemUsduaVHUKdvgyZn9blZgODHwy2N
pSuoizK+3ZyL9s9cx830Y35txquu91KYZh3fqWHnGBJqSVlap4y/ccJGH1Uoy/+9no7OFYOhTDSh
ca8kC85HtS7yZ3Yve48XMvQb/BN9Ns7/uajGk4/3SUND4Lgc6muF28bHfW5Be41t80WgQVsCnhI9
yb7CYtsnMxZw++SSLBOLOu9PrsB03VsZjCrwsNFgY8y0lTOpsf3764Cl+/K5Nz14XW2k7K2bzOWX
ewJsIf8hs+6pM3sV5AbEhwbvpNfqIEwDXYijpa5l3drId0D8OL+IUIOXvRTbd3Zo4HnZwvh+98Zn
tdDulZzJ6J90ZCqz2NM7z2BcjCnp/zRn2FlkB5SSfa49I7MOFH7VI7uLnHErL4Y+vJdVxXIlX6eE
2+qJiENfDETumWT1JrIljEM3dZGzduXOIEsafxK6Xna+j10nZxDFGvNVvJdInwcdjUH1raOUuYMC
gRT/XytbSw4GgUehhIyLG8uCU4IkjDiuxNXubqr0ktdOPKSW+EUlb7vnY2lJPx4DPl2W/lZBZrro
hOIgVBgzqm0Nvwmvg6FnLItprZb/4dErYW5Ez7ySKnCfAAPP0m8Bi4ubKWQ5z2IvCrBzc8yYMyVe
AVKu7D4SW2SnI1GCjg2rpj81euFysnhiacwdVlEW+novjkVI4IaJoC2mwOk+xfKWDg5FYwkxzpsh
JAd/SX3mKaVicDY6Hyw+AymlM0bGhyflXUdSZoRUjNs8usDrHFu9v3hy8kUyzhV4qXKxWlkkUfly
rYYbsSS1T2+CsCwL9JDHw7U4KksWwkX4zfEEUR/boctWxtk5UY4idvjz4yLu18HYLaqqnOCG1yq+
wf3xemkK1WmjhvnyWw4TxcBYwiFNrTpqy0isjTu7aMc8H4CsSRHayG0pcZh57s/QuUhOxfg2gzIG
7RrVnCzrrUlikxXuSf4f2ulvgu2qsB6o+hqJtml3I10UbtssXV7+MhQIcvS2jWR3vwWHX0Iwhtuy
0cvB8uRemEA7UGJ+a12RzRl3c1josTFoHfai9PXMcIOw8KQpKBrYSfZGcVwA5pMoL7wX2QUaShdM
3JWHjL+SJf34yYfPtEwyUzGWqUTowD6jzeJ+DoKmMvlDJERHDa4BwSX98KkYm0fZbqjxRbFI0rHI
5BG7Ukg+8s0llVF9IiI7b8RDY8cyOQLNL7P27SWrJQdmvtBtc8m1be64/Iaz0nj1A0HLA5VQL23r
OjHBQi1XTyuqf4YGsa1ESUewbM7YKmMBoJ5DZ+trd21mpNl7773Wn192pfQ3JqaCoPqHme90S8+i
I2nWGTkMHT9MHrhWvIJnsdEGPsm1S6OcccvkPfZlipDP1bhDDh9Cr79ahz6GkF/AWVFPs9x52EmN
QGZBSLmD3bvHoESJ22y27vGSS1Gk1CGcVNfKKmPvoUewZnm9TBGH4B4d2A1cMwMuaOYb2SogSqOo
mi5LJY3TWcA8cSxmrvpDuBkJzzacCfENfiDeDvvs96BJ/hOMg1GKxefLmVNoOw0JwJsK3RUR3rf8
FyZg6aYc5I0OMHUSrm9aqfrcs9vReuPTidOwajaliJ5lD1JAwUJQvKQ3Li/QNWcNPMDrr63zWC5b
9+gQyDMrQCDadykwtovasVEMBp8eSiZ4pUJmSTl1gxoEYmSSm+P98Ra4ZHzfNhGzhHs+vcyFcH/G
CFjbf5bwsl+DZk4EnXjIDTv0WVZBFl2RVdnHr6laiZlvAqrFp8T90Lhq8cNcKwU5jvhnE25kkgs6
PfPqcJyEVJmPLqqEaP/GYYQmDmOPt+bCk/W0NtcoG9XK0S/1dls7mb4wfIY5tNZKuZtf4Y+NhWKM
28mpRsAvsm8kDVsrxoiKENjVftpubos+INGLRViU2sJsSuLKmAhSyO2TQ76maHX8zcCaXFqcuNPk
NFAD6jokFgSeVBtxcnp0K9i3ph48cMxF2uFi+KEPeYt4t8lG31063D0UecqwNtIi3y2AVxiSbhcY
5kx3gU4jtv9EBjw6V8FgBkMf1lcaUGSmZQe2ucAz/GUDpqUFGpu2Kkyq/mS15dIxzGP31h8LRSAz
XAlibtiPK+5v06QjpUtDcTrcHhCWdZy3FLF621PjC1Rb2nSG5UoToVX5GfTS5yQYKFt32hxA+ar2
WBq6fAlwEBd3yRn+B+i2MsIjlbFw0z/1Pt/WSI9P7xqV+aes4gROfMgymRB6XlTpT92BEG67M1z2
DARxYFaWG7mShElInmDmzFw9p5AEOy6ZyqSKFkQ4/GW2ZPA07lNyG60shK+hqoTISCXfkD8DbNlv
851hbH/iSjCetfiJnuESaPkL5ZLOUtUCKfOTCkyIG4P5uy8bMs5pESz2b7ND4Fxh/e67ew7wenx9
/0Le0IeHlFmXla47FBYx5pMUYsy31WUygGhDIFHfD9uZRCcP+mDy6PF9OineJGMjNMYTrkutGtol
gVa/xETUdHpIMUJf9g2N0xlmZoZQn+eckkLeAyaLyGSRcFTLn2yo2VFHF1oEKd+NqAL0pLAO9Abv
VxOymYHy0Vq3yDVHi/gbFUku/MzH4BDt4ySO/0UJP+UvcY5/Ts24iLegYoF50Cmiy9a5E6ssB+f+
XWqOSSvb8p1smfRxcFWZGUsX7VbZYgrfbTzJ/aSpSBb+flqJ4/Q2pxNlh4phErLR7zlbmaPDR5iQ
OYe9nETqULiqTVC9BZf4wtk2yLyPruw26Oy6Hxtt+dLtDMwRXfNfkQbS7eERyVsDQlxrjvKV1bEW
gvGFg1mFZt59Q8DVLF2rgtykrhlyq0EzgD+X3d0KnTQa76Z6VUlH1gwZ/NyPYvu0tK7B+1AG2LHl
1UrVzJwxVMFIUEBMtFQyW7wvtrA60iYeNgJj/IMMndZINxjeTOzE/4QpdTNO4RxpYHqakxWpx9ah
j5gr8CHJRoo9HbYZ/BVNrGHDBVOS5ib6qVgZS71vh8cNNK3zoNd4Xmwg21u6vA93WaxtZn91Vsqf
MhkoF6UaJSfiNRiD79YcvGLF5YQYNEPGsWu/t11r1ma6uYARrACz0nnrzUqiFxlwmMVLRFv5Pr9p
ZweSh0pWnFpYJ+PhnxvSZhxne/0FUudf7H0t+ZEaCnKh2JSPD/UOtc4ZwXlpVsPUbJMw0R2ZI/lJ
HCknL9xohlRRdfk/NkKdCUmncYQ5yE15CaOc6Elf2axEmw0AcdvW2yvNwxoWSqGbGSRBvFc/3quG
GE6mCEQlv9bpDPRtHEiOQXYZOiXwW9aLhMuJMfyhEpfSb8OnoCXom4kl3rWBzISL9ToySeM/DUem
A2qb61gp6+FR1nBU6+MdpqbeaRDKbiLdW4oVKM6C7JwMThgdH1Ptyz+RIaOvV852HSinNJVFpins
aZmKIC3QtU5i5qfPjmYX93YAvS8utmGqXYAiPBTnE279Vd59Uk2ExgnGaX9StEtfQb+xvSqGdzKv
rD4NSjnb100M91YZoRkz0DW1/UMFqqzWMQ6Sp3Lj4W7SyMVoHVB7rIcm1fQfUxJilOnDkpBCsxau
xWnni5oANRpjHDW7cbc7CUbIkcloCjs/6bGqvyO1ju5svC4rZviyE31p9hj9wl8Iv4is/sFC2w3A
ea5KBN4PImCG41loqVLA9y5bqe6Ac1SlPD93XaDDEPKOHRK9vonVlBkCUfDyF+AowPdN9CD8cAM1
nb/iYLJyyh9c1c7EE6lidQaQxsyfinXaSCLo2FdEhvzCFgqOPVKKOdW+mbMDuEBK/omPJjckt+UQ
HEkluZqrWMpSZ/bO2gLV7hNoqA+uEqDPWzMkRYLeqy18dmJkvVPhMUE6jfBhOk1doVuLvAZUWklP
UEDGGb5F/N9d7zGX1ZD9hakAcmJthYnnROM8Mhb+7c9TWh91f0YwIliEC3DlqN7ao4GMQzC2Oorx
YYg/wd6eQ1PAea0QEtLgCVIctUBKdfJ8jRqzD16hK/zGS7deX1lDWZ+5Czs1ql8kkA8Pjt8IVFeg
p4VlUsXDo9eWWGZwjxvR26dObNMnBonWF9VtWctXqU6r/RtRy+50M6S7mawNkU8O95foWfboL+rP
SihOSbg380bcAQaZKx2sE8D9WH0cmcMGVwFmqwh0Rb/evVClld5RKJxxtsi+9NVTvfCTQ72aff8j
ON3E7ryVJ3gM5tnNEZs8ST1DGsRUJ341kY6mCl6Elsj7FFq+qSIBCxbJObY7VViSc1Ss3Jw6r0QV
W01EIz/PKq7DevPlskin0CUCeiSeDz8o2nPPELojypNZAuE84xywV7czF9L16/UB0aCYFep+bY/k
c0wK8NsJ1+6KkRMu5PN41z+D1JCS37hHnoPUETKc+FwVsgw+V53ABt+0dG7sBQHcoD5SWWBut45Z
1+cqdG9oufJ2k6h6ruhf7Gf0JvrvuERdiau8Mbw1l6uEIFpusS6sdwXkNMrNcI7WtbRsGFmhA3xv
luJJ9dS5GLJw326imX+yljqL8xqGHmo3YHt6kUiV+At/WJYgtnmLEx+YGFSk0As1/TXMnoAebi43
Vz8HWnvn7HmZ49JOYfudK1nXHwYemIsI6fE7VP7UPU3gHW+CMqaN3bt3R3q+vRBu1Kg68mCLd7TQ
oBSFuG/LKS9j1fNuZvUZammUoy78VgywwPsll2YZMMnbdPXSv0gOo29ohPLJ4J2itQupXL1vup8q
tfFyshmuVTKgxpVC2PCzyXLqThYIku8emeVioMM2GLbv9xQQDPS40ofGMSc5je3XBcQGqlHoIxt9
5y8DB+lczEnj45vt1/q1Dd2Exyb2nu6ZnZ6B8GwSwSZJltg9E0icSWkFV3AcrlH2wBJZajKSFzSe
H2alg9uGimyfhGl1JQZ/hF9ZRNZySQkjHn2H0+Eysq/ZJ9u4DiZRdRDh11vp6jeBXiQdh9TuuKbW
buZQM7x6rPvf6OMArdLY7lrHK8iTwYpZW+1YMpd+oTj4SvEh2yfacSxj7WaVu7rcGIQdm+iTNgIq
fLI7zhM0NGrSRCfBXCathBOOy/JWjVEG/Zcxv/JG42SDfTPB4Q1VkkcPIHgdp/0SLuCAMENwvnT5
/QQqQwEZpYOuAWBGWIjqUd0ARQJsa0bqhw3h3PBY9P0Qikrc7Q/vQUj7S9PJQo0y7GfNJm9R1mAj
HPGTQKsxkob/nyA+NliOXY+nbpGC+5+wGIwoswJ291QbN6AHCn0zi1C+3+0VRQwtlXiBghstFj68
E5S/1A9k1bgclc50axKCTCbfuptNP0qfoLmxgZ2DDYN3nQviU1a1sBf9ogHfl7CEnZ3cTfQeLAcE
nwUZnE5gxnogCItJ1hiatIbxp5uCmwNFxLmQgtM1IZLWUiRhMLjQQnCnFmGrFX5hKM8LhoapUSk1
aWhuVu4fgKjO54VJFvnnV7lXEYX/VuZ7Xw+EGztDrNM9GaRRT2G0NAqQUwr6o8X2ee/vXOfGZibw
qh1/BKmFYkTEPHz55bbBQ54BU7RmeWw+bBnA1DS2WMPbdPkQIbKAzbDK58GQi2xzFqRzPhsu1UdN
KSCvmmXHHLVNA5JnpTMIngQNm1wWSd461zLHXe0BcF5DQ4xfnKEKBuzH6w6br75H2mDev8+VFoGm
SHac2hU3nDeTD3vNPB2yxkAKcz111c9hMFUthxTniDTbCzxEN4mUava/lC47CdGZ72dsk2wekUYI
4hBNssHcQHibcS2pmRx9gZ0OnsTqhkajrbPcTNQovbEVsttBxmYnBEFoIfqHeL0zxYJ+0iG055FD
KRU0C9CQZ8jcg1bWPOj5WoKIm6u0XGK5pcpxnqXBFcf0UQdGfx7015Zg7T4sgoNNu36dgwlNJMl4
BCmHSN47HP3t8z4wBxtn5bStjmvA25J8lPQu5sJaCf6GMSbmxFZpXWupeskb+CKf74bcwOkqouYv
5LtTaOYfyxvvfuNwMt5N3B4aij9vhm6pHN93VGQ2ctYsjeOWAwF/zl0iqm6LaLAny6tQioKqFQ+X
YU6RJcT4jWUmnALQEbkIQLZPuiFFrnq1EazW7pkUsNXqPZlW+xXmhSe6MfSQdbewqI/lCUa27Vm1
Hxom9P+MinQM7hjje2cMpI2CZAXAhlpRrUt742lN4HAXuYQA2hiR41fdWrDdw1hkXbOoOgUyKJbH
4PxmPV0O4SGSspCwu9d1GdULJgwXXL2wtoYw6TfC875RrXk7qfvcdgspNBa9jZUkJvuKUc0Gcnbj
ryKLqjuq+OLbdcQi6TeshSNU47h6Uc0K0cPT3Xw/uQ5tKoEK4E6r4LEDngUblpt5pjBqoDCCVagq
tsAyhG9c9RA6HBxapvjFBtdDYnnw8fL+itmvl0QXJfVstT6UFZ6Glltd0MNosO29jTpKH7p9nOY/
p/WckHYnIOG5LIqF4Z69Ws0oe2TvFTAbbo6Cc0lq3IWVSiCjKCsClfNQMZtwQTRUDSkSYDKgszV9
0AssTE+nZIxhx7CHhhRVeqN+vANdxh1Yka99mcHB+KC6jT55vN+ysXRqd7p2c9XUJmQtu9islwUK
0vAqRWRXqapsjBSsOTm39qiZAhCqm8a9IcRwwuE/pp3faPgkYd2ywnJjEMAGKvNFD8ryEsJURY46
FONC7cXnlYjGbmowZf9besQhodL7VdkQR4TqlaGoTnpt9Swe5tsOb0Q3acI2GVIb/ozKKZd1TCaC
iXnmzJ6b0mBTlZIfNY/swSuFX19wxkLzHTHkIJCIva+w557gpeG5eTOf3l8JUrUgn0uK8q208Zll
U9q9FGXG3Eohu1UefbasP0AbSu0FAhf6H0wg1e5LhmakAPhL+H8bJkxboCKJvE32BUfgiX0yrQQg
EzHdjzzwEm6711E6osaD3i9cGix8HzFIC+JCE6OSJL2TIX/sTEg5n2lmlPuw1gX6+s0JPttqPGVz
1uaRt1qMUIkpmvPoguJ88uWG1n6Hl3rdNhxk1RHSsJ9SPtRQPShmXWQ+3SBBnIgtifi9PZVhv128
yNIjoSfCWY6bvPoqmmRP1mAK03Lyf8ETAzqHSKWYoijEVIOJQsO2arax+jQy+69VuD+t7izsH+6k
db8v9ntoeycY4szrtNsjKgb1Gv2+13rOZVC5bsDzRGUxd03xXecYXXsDb76wi0EpYISp0Vcnyj1U
2YTZpdi9uLcuV4ypd/nu0yaHgVmqJL2AepUcsOh37/BYWx1Nkp9aMK6sb9P7z5VX8HeYEQGjqQma
hm8psTjn4NGVvyQj/wKUSiDuBvfz8PRExu/nMmW+9fbw1ww2zHKo5SB+B7owhktv75Taboa1sx/J
rESycUImaFQu7oTFkNrR8sC5ekzfLCjJSEo5OIlONAGGmPEc/0kwPQi9ktShKOZyai4xjzSvFeZA
rWa3jBtEyZriV63TyKzevMWuPAJsc6cKABSgBZ2yOq5HaO5RheC7WAzpArBBXQYPr9Dj5BV+Fs+0
YQCS1tdLADLF2eOdxfg/T4hsk5NCZgA3oEp+7wUY/Y1VSjgVQlV5zeLDjNQf8qxKh/0w4zbuiAGB
RlBN++ofEQSJnuKdn6luV+AFt7Q+HpMAN3EmdCrAotuxfzLDtQJAADDjoi21BXbi/zf+xhPf/7GY
4YQMGPggxxAIotJMHhespb/IH19/zaoWBtKzNRurUGOv+9lFwrlAzGSd/+R9G2lUOjZ9nm0GlERd
1imFo4L7Z4k2E86YC1G6etNT/GZYIQHKeCSwCVo4GVQ869mqS5xLv1EI9fQ9a1I7s7DAdunvIzfR
TNmQWZNSA01He8oqbq2W8TYhakBiuiFxD5FcE7y2OrcfTazYt8gNgUNFZOb9f/tHJo8cPbj9j+lS
wEDAryW0MeBMYytTuNbG/WSsikGdJsGdbZhIr+Bs8ZLiqyFYxDrOn8YxgoG5m++qhURiaDPmWVNt
q6NhFQhcMxBT9V18Xo7u4NXwoMJZhKFWfXkAo956t3dO2aJpkzi+LGrh7JXfres+XjSi+L4ezSog
VqGbXEtV9sfYGZF+LuijhxNwIq2+9ky0ZwklqBnsDrdqptHj4Ea4EJSQxdKXvFbkVoriorSyhYmk
p2eYiOw++xK5YEsECVPVj/MO5hsFkIjmi1Cm9L5nJ4PYIL7ibUgIGqpFcOM9DdoyNvejEoIQNiCP
O7paZTYkI6dG8By/T6nP2yTnkgW2rf3//GUTGXLAcUb5rN0S/IwAcI4gnexZUc9YufeT1eG5aiRf
UO862X2NcdODGAgVlHY+XM0o1+nfU/tC3j2ZVecba7p2HP+sMOAGBvjzs7w97/E4tCVwXy/1WYQ4
IIeE15X9F5AwOX7e/vjnED5PtZGXc/6E07MP1zyLLVVMn20XYFvKEwDwOUMeVMsB35EDP+C1PHQW
NYDxyvK8UBEBKfFiM3jqQqH3YJOvQ7FCMiGeoXSlQ489Nm8DYa0sSgSyXPIk6Gcy8WNxS8Te3pxV
+v9rUQ6r5tpz7zpeJ1m8nW93ayVJgeZAjlR0+SbUy5w+8rJJmJpa8z/C1O/wOX46P4Th1eiSkEYp
BucXARd7c4cRaQdHjoNK7y8Fg6D3BY3J8BIgozKa6qQxn3MZx7PPN5p8qPRNU6g315mT255JuHy6
a3KIWjNhWUs6WLwhQTNWb+g5e2XGe/9tfP2CqgDHW8YaRo6JtqI1IMFW+Bgr5WIFLBipYJnDFA+T
0u9Cc0adXHyCAnLludLsW+aKOxD8KNCXuZzlQOtsRU5uI9Cpm/Mx1s2b4+wU10lbJAO4LzK/0now
TXMNIhtdu7X11lEZPi9X1LF77fgHbEolrg1XNuN5EWr2pezCXCCn3NpB4l7wB9hR0M4x1myZ8FB1
V4y4yahxVfwal0f3T4DMobUTxxC5BfNGG4QQ6iCVPyz73RQRYske8+on9wxFn3vs0/y+W1Mb6MFU
zV/JLp/q9ogW1qGxssxB887RElFkg7YZUa/VtZ2sl4gKQjY6+zwTIZezbTsXc9DF2o7SrzheCbpj
45vVHL4Sm2WPuB9B/ZyOYPNQZT0du2PCdrXpWTO+TCuGS8z6ItmYnEpwasbKdFbyVcYF5QMPBIAn
daPVSttVMzvLLJlGtQkYVrRojaUllGuKLA/l9WgqGVk8yx21lHGuV1//LaL03UdBkP+CAN02Pnvb
xBtxyPxGKncAdJESuN9M95BgNgv9OwAGVdk7KJ9xq3Uv2591ktxdOLl7h7xAw6Z0LeZ1sSH7qCqF
1LOak9fo6DWBaXA6CGR82iciCaIFHqSyqJpzaj3QqFTHvPZegWLkuD72Qo+fTQT2Zi4seUIc4i4/
rJpgkjqUuCsX/nh198SXGys6co4YJVlxkW2AzI4C3LZmPC8Getuf1Uyd0p6dKHmjFsCO6ZQhIKiz
r4XrXmP+srf9az6glJJaSrdHP72ppxCMNbe/anFgsZpBhK9gNfH+tDmdU0u8Hu3GOKP3Qka70xnm
5FOwkuZFWh0xUgaTSZc/E7zUuE7H4UzcS6ETlXB/+IJKuPfAb9y+bmNv1RaOQ06jpncX4fcOKLCx
VPZZmarLIvBAOJZ2De3CK2URmLtIZGwDH1YKFJUJosOT2l+wUMiSILY8LNN22f+H8MDmi/Sl6vVF
EWFQQHpYEg22WxMCS/5whcvVgC3ks7obpEkoZoDhylHpRS/J9XjeB8nxGFGxJbbC4djkQtEi/sim
gGUqBnq+xPsawDDsqaZrB2YoSyP5HmbhTz/hCQFHGLkB8nax15B3/tbC3yV9AeZX39O5is3Mwrr/
yWdU41uDQSM1u25wMRRsCa8Uj1lGflqE48HD2vZ9rvPhJ/sYGvLmro4LJHCro3tvkcTfsUOpyppq
WB+Fwu7KqVyJYSox4yg9U6dNteUr+WZq0OdWmUMS8PhnUBwCE19UJsgHdDdZne8sIgxKo0gK2wMk
fiaVf8PmXXkO5Swf0AnOai0y1grnHVs8oM3hz7YR0Nt1TJuBfWtWUAIUR0QJ0O+TeQU/eeI0UCYw
OH2sV2RWVsda+7A29nap6BHa00I3UT5YU6PC3Tpxk/iYSa1xoQf5c2U/1dESptIGmLWwgc9Xxlna
nvVrM3U1XIenNxCbSkwoSYPQIAF1aQdLds3jO1qS25aD83lyVCv/1SPeQgeZPpsfx74NOyiRDiqE
rQyin08xSUo3s+hlhXND2xOSLjBcC6aUR+ylQ2i2oE1Ymt8p0IQx7+H7x/n8ude0Y00fwiCFqpB2
Mh11uyxCTfFFdNhPJ1jpmLrtYJeB1kAiTEIe2xEh5EgvUDivHm/StjkypKvqHPdO3C3KE9HrLJ6E
4mYEb6fFb2mHvD6odzfd/ZPNqImX+lUVrP5wsdctS3qyEdjcdolSswwR1ppu+ZxV2OEhqwbdSLuk
gjewiAfmptKu8FsJkccATMRMEtP3D4Sf0k8A4Wbs7NE77vq3RAiMjdLFoGL9XzhsP37k0yXHjcBC
EWlGLopvqAGlHsPb+RdH1BJNT2yf3+w3SrnSN4KKyzxpcyQ0PX+qEl4ET+V6ge7phWfMT+QqOwWh
P5UhIiuBf/47CzAX7HYoUIyy2IsrVdXAnrBJnCvAGEP7R1qP4sOsUNUEMwhqp1/Na+UbaLQn7ACy
VnFUodnksqgNBb7QX8/PlHRty/6SUgRBQJXG+GTMzMjdI//OG+RCKUYOmYtFYgQPX+yu50wV4SdP
Ev+TcKMo9dpBwTaL6wkeyO7sD81KHPmW4K939FfPjJ54DIh7Z9XmxFKM5uM7aKA9VHWoG009VEjL
CzIT53svzI0hfmIzA3JK86rj70q8y5fAQyQL0r7lUM3SjTA3y9T5wE9ggMWBxiNTVjM+xtNx3jLE
iuzndkNBqJ6pHGUsGEmzDpq4CBqNFZIu1EfqlQPdDDI3eZzaLs942SDYvb8PSu7AagdEJXYSSMpw
E1XFyfwW9+TfGl1pDsZL7SxLWL9HXlcjoQb1fEgwbLpVKT3XJh/uq3WUYzH7PtnH2sejSEuSZyQS
jexa8SH3xPCOt8NwOtTOhaHfoVZStFqSetburv4PUosRFCEiI+U6aE8uP+Ykm+2efhmgTbZwM5rX
ufxTDUHVINkvZf9QdkkA1G8njstehIhFo5rf8k4typnLxg3flf8ISzsjg9zyCYtMjj/t6j2MlXga
u+7Bdx7MU/9hKUZx+5LHGZx5Gh90jLWJ8JmfnIhrOqLKeN4dyTqT2cIQ1NRHTzvd+yYhgdRYWxzq
a24SFIT4wTH3QqYSFPUPSul//2TEGRcocmZavZYMtBYpY5FHoIWCctBd7cc6Kp1mKLOSVQ+VJtPe
P6yw/14OVxsdiOtcXv5M5fx/kl/wiZi2KZbZbJ3d4mL8LzEjDlzgiM2TurN5CjBTVdw+BIVL6K4m
GY+M3hZkC0Kb3YTgmhI7roEAbO9bJWjaRd8VkjVvqFPzqYT9oycxtqzSHWGXOdIBIbMgviUyAmx3
ROKlnjXJSrHEa5JrwBBjuCAfiz3RBtp6cK2N26OU++Wxw2SEfT8CxJqDkPl6TFI0QkSsOIOVIN9N
8u8GV6n9joU89LSZmrcFfE6ZXEmlkBgl3o3RpRjS4lGrWK/eRCMSWDH7Zx/YXDj5nyUVEltULRLT
t6HRYkp9sCUYnWDM3CAAhOL9RWkjm03/GEgizfy/fljZ9EdVSpCzSbTDt+65ZtpQ58yu8kL9GzIe
K1/AIxZA/8F/E94lk6Rsg/aDpaLvRgRiEbcJPPHAewHs3Wvq+bVOypidV0PAvbLbRdw7A6tivcjz
16u2yJLYZiISDPQTWhvHKahI56B62qgOIJOTT16oxT5ZaH1wPKnaCizjP9JXXfWGdDJ/LqH+QYYy
0eeHX2hwPewXVSNJ6fQvj6+guR6sj/9aIpuDde3VbTT+MRJHyn+fiAqe8z2BdNUD7XrMkbwlbrMY
UcZS641iiJC7J6Vm1Riehg9gJ6KsA11Dr4ic2Tkth4c9LlZ+AIY6Qs9HfspJWhVqQhW9XBj/Oh8C
EyXI0A/CdhUi4krLETRipP2Ug//+olRYTOLX+s3XSp4esSDiU2QwQn8BeGPkZ7TZw6oC0eWYoalg
A835Lizcsb8sHRh4pC08xXtY9vauEwfaSIxPqfICcNmSC0IjIjlzVMfVQypVt0dR7762i71vLvj/
6N0J/oLkbp1movBRWhwyFksad070Ib9HK8Or0yOnZY4x6YFYgRdLZTm9IBYG35yF1WJvw0axX9vE
XijBBc5OF5RlLr7z3WF6740eS1EQ3OLsLsefzpUO3eeWW8MlIOjcSyPZN8jao9Q/nqWoCk1Ev4Ih
LCPEYDl4cDyTc73rRMOLgapbcVnidnBVnpg2sprVQyYUqCufy62n7V8rtHxZeWVV5vzBPmHo0B50
hVhyNe+adEYzbP13nOAv3WbMi93XCPbKJ9I0QS64Yt+Utqp15C5+9yeNi9EU8qF9svAdkEyxJv0i
18kQPDxJb2qbKst8GeD5YyoN31nbimK9iRgEmpsFpSl5RiHTEYtrVwBtEaseYMYYDet/PNvGggT9
cXqVfs3pcgauWp5XvEFt7Bow+JRs5sTA9eeXrhxvn2X935yLTbfZmM/mXiNJfSBYMV848VrlY0Xx
UM6+4Lfdtp7Zy29MkGud0yi8SxICKhjxEHmWAfvgTVJStmTZETUNMNpfm7D/M/wpGZIUXkjz1Tx1
u2o9qYtBKM8hnRls2W8LCd4fQnH1KTvgrHn+m+aG0G2kjTE1PrWwIMTbWozW8Q/g0W52j/hHHGrb
Tbgrk/GNX4y7ZbOOrWUiHXtjnx6uNZV9ccuEDqtBtozAl9KV+rEAbikdfQTkmwI+qW7EfuOT9aW0
iZQRLU6vA9tMiqNGJ+FcU7VpwcJjfw2ZUWHvStjpPGfvIWK32UTU+Ms34ac/3k0n05PTp/qgzQnO
o2mfOld9J3p+IfRMBGNbSkqy32+F/C1KqbmjyJNO9JfkhcGQNjUFdKUlEMLAaWD7KxE9zkTA009F
auoFQoadgj+I84gC3oDgsWOCALdi84ASsJQSf0mK/gnhGw6rWMp3MI5CUDtz3vUGVvtCpx4UKXCX
HhX4BMeAvO0vlh0QFntSvXMAUvNFuY6rE/9TTqMx40lkvigVp8AZbIxVHTS4Jtz/t0yKEkJWnwdR
SDR2qTWhmvOjn44jsn+W1uPMHrKkmmpIB+1ZoqUSRaYymf7SaeWK1F1fRm4G8BObFiqRctQY5V8J
hPjd1zxEU/bBWlpay/zTGLZtWdWDC5p1P70hgb+VGv3gR8fPku8rjJygrvbmVK7cugP39YYEgNxH
YdpKSpdR9XMa+Af1+32t3Ju6i5QqfKuaVITuDXzhDSe9hVDtZFOn20PDZQ5Xnh1jePQyM8AptFe8
2t0EhRHp6rrbi+4297XEJEWqpaBrBUr0M1vqzEjwr7dPyejMRvVyBB3tDCPMOpJ76Jik8aVeSiu2
7i6RWPF4uGFCmb7JuULYqPn/2seXd84wKQsPvv64PjYM4PJBaX2bj6mnskzl7ldGhXpI1AMTrGgO
zBbmsbA5NW2NitHkUmwp2RpVApAd59SeX+X7DOENXdykiANlMXZmXwHhllgSbjb/QN+1MLWhRFki
+QB2tNXDsvq4Zj8DcJ8yu5G2wAqbVZ1UZ8z7zzl3flX+NGBVSxcQrvB4Y6SN2mzthja8stkcuZJY
2Aj8jDPlitK5+9bObTeSUswlyy1ZAy+HYG5b8v82PAW+ylugnvW3Lgb4G68lvBDcKR9kFHykXi0L
8kzhdzdZiGhiy3nAtp4JUyYanC+cOfPPfRqwJqjgzMhA1+zdYYwjNxpxSBmF7YwFoBaMtmWGtAMu
OOWFTcEp3EtZRcJ6ZPZDjDpsszKr8fT42SQ6+VSyccqQuHi27Gmni195gBm1MkZJmL9RAMGtfD9j
G4KUPPrjQGrUb/jmY0xF7zM38FrUuP23wU5F5a7Dl0xPhGGmBFJMI4F5xrnrb6RziJ3SABApkRmH
ZwYPRdwniFkXhwWeQSs6kkZUpwOV/R/nRv5MfhtBBa+Zk9QuFBsj71WwQB6+6kcEw2LgLc0XuyDy
nkhwnBHKDNHdH/3kuvdGAEOXud2j1m/dTCBAc3B5CbjDIyjVJKZpvMk5P+3IvnWKHoFvmQJ66M8F
A1Imo8Vn9oJlRFwDrl9Q3pUZ+GoSfxmUh+T2XSipyiwBU33Vs26Mjm2Zy7rDWTifDr9Nbvte1RA0
BNXzPwYePZrGTWX3OmjMHUzSbAaB11iKDrf4ZLyY1qn6rgnKS0KDADdKQgsxZGzVKXlEaek0h0eu
h982wxnATmQLMTlMHniBRjx35YgT1Q3gRxMX7XxbenE2503P/XTM3jZuKK4Aci3kMiQ6P3M3l8ib
Ik4bsc3Ag+e+5clst9okcFvUuKchCczglFBl70YevWecus2fjNXxJQ8XywUd71M4RLbSS8o6OfCg
Zd8z5C9CfYul+At3SJwbHOUNoCRZLQc0rpj1qHM6aPX7VChsp2FP66ULeafkplzCsGvCdJC4Eplg
AYyzfS2V0+lxIOTX2tJsDVElQnwKhlKmMFnNtQdLDyVfIMsMktdICzrIz8y+m6GKZI/feVkG6HxS
S3fIjc+cpcJRegraU1WFw0exVBApyS24p317nR7v6bvmV9nX4A4RNCJWuGft69TkjsmG+oW5M5HD
3YMqe8H60Zr4nF37hLfmMNKJ509H/PiuvVtmnBfZYbSGnQi69UyeLOXCqDGlUqQ/bI2IqWsLToim
dfMz6OHF0b47+/lIWUyk+FoYEwMUeWJxFuUpKLEkUxfBXvvbVVF4gEjBcPWprv3jihdACj4f+YtQ
s6unsj/kLyBMrPw3smcsWOqfBnijNGeSe1rfEhKyRxRRVH7j2n42m1ceS5+E4ysqpHM7M542glj/
7PXhyGiL7ATu9yPbdan821DfsJ1y29s5aqXQhHmdH3CdLy66+k29X/kcJKlNkwRi9FYUfuFfp4h8
DZaJ5QKDTsoR0ghsVpGAmbklcX49px0ArEeqElCYsx63by9kzfGMUWZG3MIEvM39ucVDWVBXdUbZ
MGJNTm2kxCia012GvKDnr+0oR7CHy9rlugzGocsJ5ZTXPazIl9N/G0wXKjCVC2CPcN7WiV0HnSId
frFKUqqD1kWEtajTHzkyW95WpMn7mm9H7mHQh3OiipQVjPp3pKUlsIH9pDuyb+DdFsAk5q66bRac
4VFrl96tL4MZ48hB/zgC+Xrjat8KNR0Pw24fJMEIwHqCJ4zFQEcjLIg7AwmYv9ZfJxoAyaxExszV
5MK03SS3uywuRmL7lD8F3+cHaUABq0ZcgzepKrWxW/37vWewcl1+0aqGmFEoXhnhuaONxqxNfjyO
giJwm1OAQE7Zxrnc3K3+pLw+ezHFrg06oBUEj+uo8EKXFpiCexYexOKDW3TJaCk/CgivOkqQkW+Q
25SD5hF8WqRNIzIgUC4WqanZvVJTmqqX0ACtuzdVEeb8D6St2w3SCkG1eIcMT15cVZmxjydjXfi2
1m3p+w8G5Fu+Ed2GRG0CConbWLNiN9gYPAsx1lfF1Z8+YG61ZyUPrlEhe+lzFSJRPbeyp2EZN0d5
7vqavhg0wiQeyWe0hMIFrSB7xDrIdQ2XM6bsbUSC3587QTRrBnV1ZB4zS/nvx0pDWUXs46E++6iJ
aMR+VHfORvL3IQtSxqLApC4oN7f3JEFrn9y97bJou9rO/ksxjr1B3nRfaMo/wFWzPKxuFerUKJl2
oumv0l2+ETKFtaHdjPc8/rdh3dNbNksgug6Wq4E7214EZJscLpwqBrl8ckXjbTa88z5HzG5P4VSI
373GQVvxztVUs9KV2LiT1vBVmVux9YEp0c7LJvdLj/VInkBEspdDonPoYAfGzGeLFjK0UWHPJYSZ
wICZQ9vPRaOyz3YA1BwcV31d5muei27XDqmlOBhiy2r7ZJ9Bwwy2ivjqM2OgOdDtn64pySwoBMnY
+Wbry3eHU8CBQ9zuutjCJJPHkDWqGtq9ebiyo+0etxmEYT9IiVpOwG2wyJ1uKpQBS6snB6XzzWX8
IGRtnXB2c/q2lK7U1KCRVt4TpZsxkzpDuNqRM2oR1Xi3bT9pakwj8pmBeXeiFiqKZ584jVR9lZCG
fUmisxMzusRNZQTj6mYajqzZvEOhD7rYtasHfGirupdWsUA11zzCOTjWg/gUXWOlS7irOZSFHb90
p6to6G9/NyLJkSn+ceMUzy55JLsY94LW6e3wGC6hP2avQcMaS8+l6QvoNkP+dJtjVEuMSTnsnDe3
ObYmQFaddIdBZVvIGbCeoZZS6EfnmGuRZqPgBNGCdw8087dzPg8vk78zdBBxSXxNCfuGk4HrVEVV
hvoz6OaRWZps7nLxlnAAh7Vb+il/AvRzeKk6LdNU5w+m0xfhG69NHfagdvKIMIQHAFPiQw5FZxzL
lfLie1nlgcoERHKSzA82TSqnU90/YZiz2HLn1LjLt24gYC/Tj1r/mnbTQ/WYaK8e+wf9mQTRk61J
esi/lEbP6REh1OvxZHWyJtMDbabtEnyNQa5DW362Mzgo3MY+2fE6FCqTYSNllQ6wslN+H37sAq6y
xNkfGzyHvgvgIK6vV3PnlWHq/pQl51C6ROLiazOcFKKSXn3qnzW6PbXKEZbKGGodhsVywiM5b8Kk
ixRo6+Xts5TdoG4UesxfJjQYvEVueOmLtepbX6CaelJt6sn9W99lCG1gmmr4XS2bsnR9Jprign1l
m1oaoTwFzDeTevfMr6kX+q4U7y11KUEtww7+QzhoS86U0NdpqsBOoUepG23Uyiqm8d2dWTpXMXUr
euDUNmxufVefKe7YN1sHeBR2oYYs9JsWpSdZK46Xz7tVAsiGFevDRedqwG5tYYrZ8EbmlMvmrW9O
R+wCgzwTKgvctaJ/vxCEi+NfEITyMczJppqbKtEy9+4JIccsveB8rOvN0q6Tk2Wn4RBOAmCvhyRp
UaHOhj/QA2pBi54Yt/6pF+diCiJGJXOIXaO6gvuKPmqXhBjSBWzNBYAKh5Z9/cbBe+w8mDl7M6sy
JQP8pe1jC3IEihHu67JEZr8nN5LYEbjE4Y4GX8V97sdYg4pbbrl6ZaCClXsBC6BONB5dceTq/5wf
lmYzli7dYWrC3TpT+ZfEE2tTY0RWJzvMBJguWdDqDe3dccCGxiFvoppIaxLOKYkfyarep1+jvCJm
avnarXkkNr2MPe/wZyQpFQ1QRXPAgFO/Y4oTlSre2UTDxoVJ8lJtHIYMBNhF+YV2GddysVSaDGpR
QePn1BFlzN/xh/9wo2IHG8YiVFhigmFPBeJHiU4T1/1TIA53UKZJIs/XN7UFPCrNxpTfGeX3YuqE
YP2xMM+LRls3xltfZkdQ8SOiH+nlT/z7rNV/rh71zTm9d//gn491buRXrMC93wZ3Hn8w3GFn8/UZ
PPjoBupY3WG65//aLRpWzvPwKwu7hcoAhbtE44mWUtN/q20JWnjtl+qbSqavJs1LwcxJVXOaCZwK
0e3pgBtKQ+uBSg6xUpyq8HzpbceoD9wmISJePmzw7Wzj1sRGiF9Y9fers4+B2M7ytFvvGABehbHA
WwAreIQrY4ITUOXqlfAflvED40GRAlFrqyZQWnJpse+xMBYxroOOOlCgholtv3eYi7SS8rBd0yzt
XQHxBJ0CGS++ve4XIUF4l7zSvkrtDjXmioOgycXqSULp2KA2yUUZGYC0K8Bv7ucpiZ/m52Xw8pIe
0FMHyogaK/ZStHRG6JE1iihX7In3Jg2NnHKjc+xCLUAVGHhs57xvXf2Liwh/+pT6fQymURl+7E2k
neQ3pE5CvD5Y+ddc5GdQED8P3xW0sKlab29acL0OfHQPrre26WGxqFsmnVDRntI4ecAY1jmuvh4U
IaQsWUUYFQqov+hFzfX88KapsuHg+v8jp0duhrCJp7OncwdQi7fPvWv5ENXJrAO9ZlwCyIQaCtvp
nSa867kSa01rudB0ZWDDD1Gsp7tpT/y/37CS/unbJnzRGme9xU1vo0eK6TOaW96LvPxs9Ut6gPcE
egPrz7XTj8NBMCdDg43gjv27/A35z08w2sdxTtCA/C77/w+gebUGRmUyAhU5iXu5GmcQUMLgtfFU
wOzQCrSdO6t3nH0MHjdqLs583pDPI11TXDZLi7edHI99Zg3Z7MAzxSfSXefBCorKWoKuvzd02wlU
ibSAfXQ/04flwVHlNjIlEJMcw46J7I6RTDPE6u7ubzZIuXpPXVBFPJb197/831eWAdCmq9KplMII
iuoCM73RrnCuDRppH7rbQMmOnYXAe0UPpJrsS/idsPqKl5T7Yu8/h/fXjHuJon3U/4/yfZltJ4hM
HaSya/O9lqWztrg8nlXMP1Kf1XxAH5ryqDWtnx7LFQ7bXdK2yczmHOW3SdiYRdAwC7va11ic/0kX
LJfv1yJ8+1+8OzQfHsk9c39ZdUGkXONBekj95eOLJZ+AW5GyQdnkXKuseEglV3TxjagMq7zkQoZa
u0w78lGfIBbMAWEe7UpcFJRehEm/1v+nbh44xC5EWu4qTbTdxy+RY7+CMXQNG4N4Sr+xkIse9+Of
EkApH6f1D+3qF1s7/Gcw/5nJePXlKCycDFI3umGfWszJUy0RE7SyIffhDaqJ161anJ3KVxbiZJFe
JBc2puRQ5S1SXae+BkIIQlZtK9+geTTAOHCz6/SIX9/W1qZz722mEFnWZG9F/y94XOrtcEOS4KLf
vjY1kyDLi10L1VKhp1jmIglfSaZFuXk5Pb68Seo60KFbY7LdPbhlZNAuCU+L/ip47pYaJ9rhIqa1
I5x6a0pu0u7Edu1WNnYSLd65NP6Q8RHXRvQEfdEmckyDlAQhoSBhPnzzWYkEzYnk+vHEAY22ARNV
0M+yilEC27LC1WCZTRY1xCKWLt3lYJ0UKxKRki7oLYCbZnQuMQBXWfwl267RbfeLLs+hnbgc3si5
UonPWmT03hcAlE4KIsJzo8CB/SUZbGMWbtMrK+D/pn1cxJmCxHgQJkU+j5eFBnblXla5mF5I5yfh
S+Aajx57CAQMIRNR8EuhSjCTE7L/C5JHrPP2cF4yUT9uBFbtVyW85VaV8vkOUu4GUAxpl8WUUO6B
tlbPu5loQXoKp1axXbswQb2UcLLFTbTAXQOYJmPJjZBsuxOh5PwO/Fss0LChNeGsqhuCIBQxgzQZ
t68pQlBKB74OCKlMusrEiiQuOLFvl6SSzzu14O5WvkEoh56oApK4Bid99v/iUOw837Qb9iTtuOzP
hyRiVepEJSvZ/Lbw8qIWoeYvjh2yNxCV5g+pqo6Rs0kr8GeRhR3FBDYu6PYabK8rFfQV0ToCn0ZJ
ebvDjfVx9WSwDKlfpTaA1ISEc32knxeYAATmxG7nS+KjWA/mrfeor9G1iQiYcZ0gH+XCugpKNHpB
MGE8hUoA7GeGvGP0VSTSgKOyY89AlGQ1DOH1FSvYnrqE0ocBc1/I8kP2kjEeG/5y/MzM7bE9vwAP
wyCilMLJ4B3L0CLJ6iv4X+DQWHHpMhoR44p0H8Kf30P0U1bIYDrB6aFpdvPB7sqtMCn+lI+gYfDJ
gjfTpnOoGJ498Q7kEntEH1N/1mv3hKpkC0iwNgchyyRtEUmZTM9DWj5sdySvS9Gcy2zz5ncY1kmQ
be97KF94NJmWsKJe5j3CN2X1bRe/dzHiRjv+jhARZz9QOA9oojmVYxIKoAPTLdSdjsFp8gKxdVuB
X6uVMNhvndf5cEMAHu7S8TLKbL6kRToLhIt/StKaUlZXHEK1JqY2sNQ81nVXSiqgojMUxLq2JkMk
W0EOU9hC25v10nOePxIKw85Mz1okiZpwEmA2U17qtEnvpBnw8DAcEQAkpK1znjC6pukh5dS1Kf5o
s1iHNrCa/xbZ2IF1iVCKeYrrcEb9XDz8ZILYZbXq0f976fc1kETrZGWw5K3c/1Z5dYccIQ0N33ib
OAQqSBVMljrATHe47rMhcmPlpM71Rxz67t3LN3pr9SiUhYlaABPXTWi+4XJvNYSECcRZ5I5K9RPk
mYbYno4XNZGmX5oaBoqt95Rx4tg/2MdR2AtPP2B+YvopAHA+SyDqrmEZDcVjDVFzz4Isj71z6FCO
8yGo+t9wt02mHHpEfa/mrbkadbZG5JjKRkrIbuKjnU+GhQV0z3jNjpmdJc8PIs7nl0UjnuMR3H9P
MuDLW8spo+uPgmJ2b+qQ0se0jO5Fmg8mfQnYV3xkb8BT7g8gDPwsCKWcjHWs2wUMvNthCmycOZs+
WrgJmGYw8hvDJY1KcpjVeHvDNkwXB6dc5kWQ+2zWwGG8HvYuDJYhPdENiiqU43iTP4KgPrBbK1M0
TQWpbFGw7w4mMsWbqXwKGa/e+LYAIYKqaKGv9I6v3EgsKjXvicNavsRvEyHsrE++nERGhw+BP0P+
kxY102gjcxxZsF5EVGKqtSGQmpZczxjTUxgVN+MuWLVztlADnah169m9/gnZfc+Hf868YR2LQ89e
AodmJhh1h05A1VqZ13Zg81iE+I1Xgg1uA3qD8YQmFvU0pDaCfkGXGOMb4e9KqzrO09LPQkV+maDm
c29Kld7+j1ApVDQ4A+0L8wAJZGLPs+D9TjboLblph+8YJVn+xu/Cpj6BvYmml9TeGLfa2Xk7bHk2
f9pKQf2syeYiXfy0PSrcxbSMCLzDy4I0sN/qJhVsRYNZu6dAVvQoqmisRjItAdxTTma67cZBllJT
NHoXy6pIQuzAUS5Fd90W9Rvu+KdGpE3pycQ8JeRp9jaad7EyYbhxipEBcLNYMjZU2nukCcf1KDV0
6mh+uPtFgc54lvBkj2CHssEJ2HpDzHTaQhrZbskvZ8N0DAHsSrmF/C33zZbXEDTqMOQ3pzNA/d4U
ICaLFeEiUv+fkLHM1L03AfZb58L4HjJ+BTvXxIUzYQQIwVI6S25qjSl+1lncqgoH7vJK4snnbHcj
CD2Tsx6TpvCU9TRD421mxwKwyjvmbAcjYEqma9EvCrl98BrqDzGUumk/McLXWF1vEAUW8MsKF11b
ZaeeY5FQP8JzcS5goqKLFd5u1Ao6m/hjIQ46SjOH0myHJ6+o9UB1MGYToqUc0mbTQcy6L3G1anPA
L2d2aKZPVhFfAGeDAa12OelzqsuHt1CtGxUj4eXfZlr2112jUrb3QhGKIbqQ/y8th3TLcVh1/Fek
NwOh3n6OPJmjG4RBi06PItgfCBMUxATlaJUgA7SVkXvJDn+8cF3nVDakbISMSmuvSNgfhQUDTymn
N1Xqg6XQeWUiBpmkX5z76c8JvEHy7wLImmVarzk/bxkxst8Y7kKe2c/3/1UvANwK3YQFvGn8Ql68
1iwMpeZkab45xq1v+hNQRRvaR0TKbgbgMuwwqM9/gckUvxHM2mgKneNBwu3tMI/zAHXteBEGs7yv
zY8G5QZeReuo+bfEdSpufCi4uY0TrgTNqlkPWamhYAtwgAeI5C+oA48v9ttOrrR9b4OXysOpzHXn
2yxmWchgtGaxEFwIjjRnWv3uztQum/1PYUjX2WejYv8c72kDrUe+Hzkbz4EcWk4c6DpxNDusAXxz
/WgfcQB2zDuszHNZZyKpM8Fb9BLjd5CJ3Ac7Tcrh+Ff19CE+2l5wC81iOK2h3rOHR12PPpGuv2rh
gKBA48ZDatlVHJp1crqz7nHF7mxuBik/+FkHZZBnZINt17DiYXhB9bhQdIp86BR7yNCaspcBJ2D0
M6AJmIs0tAHbcFi9Zr/TRIkHmlIQPG3mZAXWBcjQTLPeb6tJp8anlVjFYVRkzYVrmM6/mMHs55zx
7TptDRNQ0eO2IkBktlyvY/t+641ow5gs8HyT3BAvFhSNYtfLMJGKBNE5E3grGpMon2AsN8844mHr
YKn3tu2LMcHEx4JGlKiYEILsoBoOSq6pZi5n5Ptx9fv1mqtYf7/IXaDrXR+QDMBMAx4zX9TXBpPT
d0OVKRsms8SoisUxe/BbvKL+ng5iODc5zweJfAxEAFPSuTL5tQl2zJrArlQZu5V6my91awn2uZWm
MaQP7a/7+BCLcrt3HmUL9sbMY+pJA7YoiEXj1kcEjhYfSZU9NB3dWfsNz66ldsqdAgLOkAQDPXv6
FQS5j5uYzIq+CyGnQ65cAEW6dyRA6nIEzjPb9GiAWC3x9oYdwKkxRdubnvAoySSDw3Hd80KPs3pE
JfhoKwYOHBDhl8xLoYg7P7qoLBpM4rZJJ0ZIRtg6RiZo7YCkCw05qTQ8E43giUkdHNyBXfLbAbKA
tIfeCwixuDNI1h+HRVtM4FxjpggPP0FfzlbpW+xTRT2AegePL0nDzd9GCxKDDbwWmzu2KVuBi55X
rLZY4wjvBwy4fGHGIxGA/YMHaN1Rin2zeji5YfJeiSJ7llULZt+4k6oB+HUv+ab9Xug0vLDNHikb
mz5XfSsiJIyNmpVp/EGu8xXQYJuemqGC/MrNp7BASZMAh9k7fk/TrwaWvXx1noX+1QZZtHgY21Nx
K7Oy/7etsdsd9mfV59lG28z6e0RUNGl1CRRdNPfI0H73yvvv0rNYD+/8jb/hF0/aVh4vY3uf2hyM
CtW+jJmPtkgcy/xjUa8PbIDDFebHuUkKWhyP7MzBaO8qWxUvy3Bl3fAIjKQLMUzHcizO4//nxv8g
adlVFGW092HXnP4rGEsLRk+9BFVESd/ideuUqYZDOGUPlM0HcN3pw89hkQgs/MgKyV2dc3rMIuhg
rfM2/ZO+ZPZSYm7oMnwpZRZjcPpRUm0kZiU+tCT6sX27pbkSGmBi1jXjkZwUxHWNKnpGBjnCvmj1
jmMu9QaSpadbc9huCd80hogESg0R4NIA4cZsyuGOugak0naPVm28JN/Pi9q1+Gpxl8cz+uLgT3vo
qCwExbN85OH0u2NSdT83mPUlWYYmdAIwQivRm/28/u7Tj9+omXwdURWnJB8bungJnyd6juOBl0i6
Kgw2NBPZLGKG6KGTq8L5DLG15unls3qgDXFXD4fW+PluGjtSjKc8F5EeylhXEDgY3VFoeiYwjrln
+s6r17pm+Kth/HU3KRMLFvQdDU3hA/dntTa/zjSm9ctdh3RBMGPDAXsdyUqnrp4tp/8m4AlmtDK+
tWzxxn+ffCbL05bPvFQ7RQLa5rrFmk8ju9U+o5U81bwTscnrbyr9T/rmnlOy9nZUTAtRNg8VZdPE
5RQQj0zyAAmL+S1dO4Auedx1rJQ/5tfdRTAaCmzokd4tURzWJXkFpvQ9EgtHE/eSf8Y1LJAMtl3m
9mWfADy8RX080VkKDgjJjtifwerlu48fF3TZEnL1GqsLuC0Y6IKjqeEygoS9LD2mOC92Wg0WgILt
RWpI/HzioweFGFB3MTKJbyYZGcW5BtcuRoQvd3C1bEzexY8GUFpyqnVtOuTRCFkeVgBIHYznPU99
1YJpUqJ1lyXLTAumh6bshOnaaI1nQKmEwG7rqqIewh9Q0cZ7CeX9VGEMgkzM15XPpi4yatsTRuNT
9s2YU+srsXSMzWqtu7JrHoYIN+3JtyQmTsK09AehCthiCzvYm8FTLyiCjTVUluwQH0OEKxwc/kgD
Vv/XneU0gL7DLxqsJBWKhsbwze8T0Bs9CgZvlnklXAKaXQ/+fC/shkfeP/0UVhyGCK5fABuppppX
HQ/ufZNHE0IshZvQ60lFGV0FtJu8Q1XRMkuzrY2TdwL8Xq0gcgSCp+C+lNk4eoIZozIC8GEFNuRC
5FwlT26pu7gczD2DC07tx1slkiALrRdBgLE93YVfsMtBXGpc4CwN/jRyDv0QapWx4Tw6ogOoQxxb
XpDkk3DwucnabzxN4Vl4ypPEVMVlofDdx9NfdnoGKvlXSkobPZYU0HoVpUE3za1xggXGv8ZvPd2u
zTFeCmJ7AemyNjBIU8XWFsFkTk/d5NEJShUWmEk+BTn0erGScfuN1WMvyWGmIFHXymZ4XxypCrM0
mFjCv8TZH1/8TjAGJjTp6wvhsZefdMPHJdHIatjc/+VFVUx/lT2wznZyPODFqCL6CFZMi3deUSzZ
w4dAvvDIiETDL7qQpzEoPPUGeDFDCZvkaUHHmxEFkdc+rzcj3JIheSIwbzM1ZoRH08JjhnR7bjTu
bG+QXaavDAMn6hBJHkx2llFamyvA3mOiL8m0L0tjGyKI1gY+M+/B2YNTBhTn+aKRtyyDOPL23F9M
5MjJ7c5MWob/sk5rXi7R5eAKDV6rUJE/Hfny7SalFYG8ue7xUmjKpdsncOL5Iu2MyBtl8zSe5BnG
32bdE6MwrnqK20K70HcfQGsRcIHHYqK0F/UedoLLR1jziMp7fKsGmoZNef1DAdAoELgWHsx/28DC
nwAp7UtNQmQpnk5rjSbBbs0tru/iwEKoUbVua46kWV/lSh+Lt7uIff6isOyQQFLEITtFqwNNbx+a
YcIFfSnvpL5mZ4cQafgbe4mJ+dixk/66K+2ytN7o3OwafIoaizxmvzqTQkHFHRxxTqIh/Pn58P3Y
ZGUP0dBxVYKXmJf1pCmNfr9lk5a3QT/IHFrg/exF+rb6CM2Q/QArHZyDssaFz3QkNq6rEhcbjsce
ac8WTD8+FdDJaIU+8JyljbGqL6M1qTBvjXczR/6EjgFafrKA6vnjvnkL8qbDZx9vz3pzH4YaNJ/V
Q+eaDWH7h5fIJam7upIuVhpHjK4BC2gB1E5OIAapHf3Do8evteedt5DIhYH9Ajh6bWuXdLrto1Ds
A3W4mbrdoJFcwMVCu6Sq7sXWV3FxP3my8GqoQ88fBdHOChcs6+4EUxJFO2ahv8cOM9Ap1PL+zo80
4dwQTIESeTrlAp05LjpENGijxQd2GRtwnQJRcoNoXWMKc3O9FaWHrJQG/3Ny8LvD8NMed1wwNF4h
wU6tsfYsVV+n0yWlteKLoaUoRM6aVGn8C/pbaOJ1UTyZsu2dk12vIJQFrx3Y23EXZFCCXWRqC+pB
7mPXOjU3sMkfSzS4wB1iOytJGfL+qgt+QEJT038G5VdvFY+f9ssy7eQDrHrCo+axNOwPjCkC8Ate
nefpZ18It3bVKixmF34+dhSVaTqVftSnUV/gQmDLKszsJCtUfAlv5WIQuIZg1ux0J+qQnYE7vqOj
LdL4dfQfGdILVCHNuRXNT8DWdiDEsLp2OxkoTKL1YrC5EPN4Vv+ypUgQMCIibkuOn1H4S14tPBrC
E942OhIp17mmBAzrdFlpUyacqgXaW5aLcyVL70JxwH5zyv7u+hJ5hKahpmth4y/owM2oyBv3jCBl
fq+uNP1e8r5aLWKXstKnXSH141HGo4fsdJFEtdomCh4PwLZsZZN334EAsqll+nZXW6IqSezYqEQg
/UJDeEyEPvLqDYW1U6sVqNn7tZOaNtL6WIa/Cp3+5ZhYm7KQsNAL1ePkFDiAWHS2xp5PFLva2d7f
hvMDru5Iq2dSnBjw6Wj9V4U9Dy78XCcVPLwFpd/WPKP3ZOh4x9XEXmZznkJXhqOwEi7UDyhX4Jr3
1I1U95CZieKiO9iHK/IH2bSodVgZkuZtfdcWblnMW1NvmBRswjYvlHumnOvG/jaZa+NiKChXk+bB
6xCGt0FwOvi9t7sauizGI40DpkM9sjTI/Wk+ChjPMBDP/a5L4kOkFWCoDUc4F8ZtD2Jz3DeyITJH
gkfar69oZ+uNLjzJK6GvrfQpWtkNrdboRG4PgDPFD5MTOjI7TQzBgsMM9lj4iNOQEtIiJrvO1pnn
UGA9yWXlPOHOEYyB68sSiolz6SfowbXHBZVtVZaDgsaVdGMMWjH0SBC+RSwzaRl8/58PJHiNvP3T
roTP2A4w0j/b9Ut5FLz8nGAyka/Ifg5q7yzXOt3/y1Ub/rywQ/SG8jRzpSCOr8eCEKnsLvORgyRo
Hst1lX1rHZ99l+ftd68LoxryJ8Jq23M+OdHs3k/eUq3UgPE2movd5iBH7JgSlFHj7VxAeN6xZqpp
FksImYhbLYbusDkK7Cnh9YXmIAxnKe/DBoohqOyGD/8rI39PD3/G3CU2VBxBNb1DYSjO8sRuFY7m
tmZGiYtLp60kdrR9X387Besg2EX6WwLrH3BjLxrHI6ioIjrBZeQhqC8WiRtl2uwfpuORQw/JM1xr
XLSjBihxv4NPW0k1iNV16U3kAipif3ZdezfnraQNMxuplq8MM4JOK2ZSmiqejyNH8tKiV1aJ1Ue/
gm+BOcZit12IsoG88zttyBkd65mZ+tabGrlw5vhci2LhOkCFxP4ZGP5rRhvhQmLh9tLICyUdI6FA
kOjoaq0xv3uHRKfu+FkMq51b9anF8RmUUwCaytjd3W2NtX941/2mgw553LyCXFEKs0h9xoiiYbg+
pDbSbypXcehM4RQJvdVEBHeTvQqiWwDUbEKKNwL0s1r4GzniUg6xy9kH+BcQpp6uu1TlwkmsE46U
bjNU6KGV7VOKKunkNuUWRdIKYyQ/PtIApzDhxOqP6YubIRafO0WDuL3TBB0X2xNsJpxKnXU/+5RH
BCPDohDduQ581O/QGZJgmzT5utCNVjuVvY1PqnXEbtkRM/Q6hZ61EFUCyVUUarqKJaIInnuBKmWJ
uqgQi3c1Fn04v9AXZtv4uPk1rGHbqGRSyuSBFqZi3K2Fl02E7KlhNRdZG5frCp5KGhlalAdYPuoh
jOLeMeHx+zBauJJM1SZa5BtgPbkwHrY1F/oXpn81db5gE1YD2Md1kGUltTdtqVZrqgEpFWL0mb9r
pZHh+7XN0g8cvhUcsUkUdcNx7C7ahdfZ0on29kqNNdYAvhzasjM9mmMZ/KYgO4WiBXEA/CpAHCPp
KuwGF5biYo+CpEVMntGRDyJI/pJ1OVf0dwLfXSMcJFvpCShroXYVEigm0g1pt+ViS6H6c7YaiOV1
vPkzHhZvdIVirDpah/NkXuw9qAVEBW8IbeKjGTEjAdbrLMsFlLlBmYHoUcL7QzCSS2WoLCq15c4H
Qr32fbUG5cMZd4Aq+1iEb/hbIsyVj8j2QiT35gB492jfhfig5RodfwG90UqM3tVJbRzUAkBb1WaX
qhLvpLi7ENiVxYFP9Q4B4ezIFT7c9kcR8GVzdXBSETxgdrRSUZU5AZkJ9dpPXo1TXHLjNiL8PvlV
CflFbW6XGnzJAVUdo6CPpiaGMwg7x+pa/0bTOS2nqBmGF7eB+fblFtyn2AmDZE2f+XI4T517tUTh
88RqjF/Z9PNlfGLSpMWL1f2pJzCVfo5Wqci83GFQfNkVlQyJjWTQmBTBlpxuqgiReM5uJFCq2afA
kXo8nZ5m8kqDWhYhPJmPJRivn8mqZ6RyhlBhB5dRXRyD+Zq5GRvOwIjnlsCt0//0mwHRr1QXjSAZ
tAuQWSWLnjs48S+fkAob2DlYtsTgK65l+sMECL1zFMFkdgt9Ys28+xQ5ioOYX0JxtIn/xO68v03X
UnDs0dmySRDuVbVyvcWpvlbZw4lq5W3ZMQg+kcgxfZacfA8BtXKaEapvh9jVd+p4ZsKWPo4zEEP4
Mepc7fxWcKXQU63zitOLl2PvnJItrOssJwsMUbbyefR4hvfjaI4WjUb+rvzbuAV3CjtrFihxMyq/
2/jT1qUBmDZKFIKlLLsxcgYVFPUibipWugAz8jHlTKQK79svaCedpG/sdr6rAOzSLgBnXBia7LJw
1VZwgyGbkoubJmBiPDmQvkGjYBUR5JDz8nZSMxGcjn/FWpN6vGqbsNz+2AUf6wLqZLZHBF/uFsG1
Dn2uhsu/HBIEYTC/N3LBOkhxr4nQ2V+2p8S40ifCoIpcGAkRDVjtbj6JBLeiRthRr0m36PIFS9aa
IXZrnAg8CjNPgRC4X2aonqBAE2IoNfumRq5TL11QRp+85bUae/VHH0kNJJq2dFRSWzgfmvBVTPQW
8KOSze9L7xO8v6x64IN2SNb6QzvCpmasXUTSNB1vACqsSfsDzMolhzWnEiU/QAI6Bx+oYnmiys3w
W9gehu1uAAwxVXTmOrZMDAJTKL6rRxfQGbXR5gGIRLtUwK3t6d5y5sBqZs+5VNOhkXD8gACI44mJ
4U/4BJJVBhTaDn8gNfOe4L3tyz7IVujZ5x4yt7vMVPKlEjV6zUt4pPkjrlX1Q/Z6UhX+1x3LfSZF
0KWw6PUGhiPOEgKMMh2gSsbFXOKh0s2F7LUTKi+eUYg7HWJBajsUkR5fckNqzRgR56blGbKY/qZC
6fyEqyU2pXBngCJ4MNs0KFEszvFB6bv9UkM7b5Ax/g6dwOYBMJC6Ir7HYkxR7YSUt91bEWvH+fmj
cc8nXkntTOeVsK5yhfJf+PEwRdmLwAV7GZNcSsmjRNjnmyg78uallQlJaXXnsoTUiFgazLgLX8nS
sx7Cp0XZZUQfTRPYstz2lAGWFavqWn1Z5w4rN82w/WPnLWDsfQNhuOFw6GSiMbTrOg0VvB6jRqQy
TgNMw0m+iSO6YEW5DFbFAR+Aiffu2bTm0th4FtFwpQeS65R61ryq9xUUOOtfX8tD31h4sGYTxB13
+epCzECYNuzHFxSr6T0d6cYxbhs6foKQwngJd5hA6cD9kE11Dn9eYwWCesb8SlEFTtoLSjA2j4cc
5DzQWaPwpMOunZL1jbqQHys4srODT3ZStweR0jVzeulmVoTcWOP+ywLLHi1BKBCqoTb/J0n43/nY
HRhRnrzlyRMPj33u7Hu/W38NNE13XV/Ly1ouJ+KPd2ftKQMJlHWRDgfiSTAdQYQfMxeDzIrJHZjl
PzFtNIXtelPS42vRWs3zK8ulUr6lpLs+x84vk2JC3rI2UuyWDD9xuIsRjsZLyEWy1Qt2rfqYjt0I
aW2vybpbCSBR10lGAixYGk3r24pspKgqMVGAa107UV3Io1MMJF4rhM/CAvef58nbu7NtM1QkEd+i
bKuto8lQ/mrr3oWKD0owBJflOnTBm+DQv47o84ib9/EwFaeQF5rXc3Poov3YTxoNPTI0JQ/JLLdR
7lqIL3rv5zF5isA4QzObSkD6Pm7sR1RbetSwkL6qW5KkN8G29WnFU+eHnHnE37u7SzZzDBUvV0M1
VeMWbZZbBBI48J0sHGFjiUR/dRhzzcz/oBdPzI9Omgd0q/lV6v0btInobDM4ejtPLFOyO3yqSE8u
UCoI2kG0bz1tmvBaPfOuCX2P4pZA+PJeWMuwBpHjEIzfXO5/xvpkGf/KXIIcsyCoHcQMwkParqzJ
88Kos8OnBcPEXDSBtYuQ3hMiWDdg4xaGiZt1uV0AR+lDFQzyq3sOeZe9bvWYs3qdxwr9fHA4hpNr
j/cyyWFkU/ju3RN51hjeQhiElTguAu8RTrdONMokXHri4emZrQ/2Efb1iNEjk1bLh4FRBF7w2Jj6
2g395aehhQMRtCMBcZIR8Lo9MNemSxjK6HHv9qe6O3X7p7GQlt2wkiwUdZ7VZQGxesOod1E9tQ+W
oFzZF8XF52Dx+u1Y2QFGLFuUjWxzGdgJ2PmjREusXkEUtta1Gw8NBBZx7uODs45kZEw/6V1ujlHz
QgVl8unGrLrM1+mX5QQsH7N7PcIwgtQyz64cc2FzvjTEF2t3sI9WZN1P6rQkWLl6rAbYkR6sYfmp
0w55M6PiF1Q3E+2ZSSUUTwm+jQTzY1WLUjD512uibIHkSrm25EfLnRytoZsX/TwJz629KQY9jme9
wRcIt48Oe/lwBcQ61535mMoQWWnKPiMX81rgtoDOXOIkNrH7ij+69GxoTrzeb01D7mTDLNs5TflM
h9oBWA2sfKDmn23SdwwZmLKj+6H8g8+A68dldos5L0Gy1hQk9iMgEPSTzQmJ/xqudo7u9OA7KKac
58F9NriGT5gRsH+cfzuV0APO6ghBuvnrrx6+p29AA8Z6idwUSZhFR6a1Zn8FkT2FPEzEPd8Xf3CO
spWz6AOs/DYem+G4eL+e56Q3Ee/moB6MZFUMBrbOF0hzALwNw7sY0tWNXBwJrxJwuOTgNwe5WvpK
OORzOQYEvfzNuw09OxnCcrDT3qEx6tjER4AE3rChV403njawC4Wj1b+0aZzFsStQZwJ1CsfC28/r
WLwbf3I2kTLApIqW2aXY9OjQOfBIWwUcS2PoeYYpD04P3Et1Gllve/4ZBHPtKN2y9ok6PLJTjaY2
wzusUA1Gz6EZ7dKKVy9VTyeVckym1HmrcnNtBS+ukjvdyAtmplvwvkInOrDpliagVRsLdAQBHlkS
AxyAzKAwBd60ExfJV7dJKvwF4iXkvlTmrZCt4PgFw4jV6LXyexBGRzA1z5t+hU1hEtkJskoqm+yT
AHDazKoCYy6GLL3ZC9bZT7StB5QE3lKoPCz5a0Q0Tgw+4DJC64pHaNk0i51UNRh+ms6mbapPpsme
3ZrMz5xDUP/MrkTPDOHQB/GEGC0ZRPUEaIaFwCr8NoJLRn1gw7lc896lNsLQCkffTr6GmWvGZxOT
fSCY3ociDpxwa2kH1ipOHheJVF1rzkbr5o/3+r1wvTA1955uCCQoZyGzAeibuEboe1ftlmGATD+m
5Rf6rIzI8h5gD2fXxT/S1rm4wnlx63/VFpoGROLdQcrTvC4HllW3W8EEnz+LmeBmGNwx+FHW9aEH
zANmuop0U2lfFDlhL0nzPR9U2hrX+l5n2LKylQGEQJTjMl4W0MKaSohsvYuRE76NUn+wtoFAmfw7
tnnMIsQSh0m7Q6rqvBVY4PG9d29Vuutq06JRf0rDFz/i0QBYOUL/yC0MWXwc3IjbIuak28052bA6
Cp0l57vwGvrdgxDM0Fnsd6PozwXIrTAqP9FL8ZyJTXqADP5VlsgMwIRs5W8ZoXjMvHLXYlV5O23Y
Qax8HLCQSh2x3CZRb7Xo09sxUFW29tFhZNYpiXYkxdpCp7sICoQBtKpuXa09it5Qtqf0+nOj/LZO
MNJwwPeVLt/8JgYdQPRh/b4m7747craV4AMmn7wDHXHpJikP8DerYiIYl393+gLoS3+aKYx4R9hH
Mo7+NjN2X32ujKaYZnpLapRN6PNWy/wq0DfXWrXNhpNzxQqRbKDDUiIqIowamupvqtMChobJlUnM
2AjPDJOq3K+fiyUrLxA4pL5gqme83FxSONYvS+DAGeJP8SBrB/REi70YBUT53vs8H3ASaIfFEbWu
IoIK/1irfc0rluNTJZrWDUYFlIQj8I9d0pueF+5pkn3IyOSwwrwuA+M+ipGP8voxjpO+Zc3sd3WS
FJqhJDhiEJSDixugIrcLGpxBlMf6WSJJaN61FiExCTzKhAOZbw8hg7yiF5cIqPANJzOfv61aRk+h
WiS7f6/nmI7CB7N7lxRQXp+w1ZsARx42B99nnVyG455gkLJoa57cxGbKSM6wpc+HNGeq5xFCftQw
HSI63eQgNfne/147t1dYRMcMa29myJd989157oKIHIw8lZEll9puvjw8pDSZcPQ3/JO7ULSYxbxv
Pn4VIGHNFI+hqOa4jUH7pLrXjODSJs4tjcxUvNIRA9K8x+mBgR2HJgsRL2rxJuuiiN3v/Sgt5aSj
pXws66NtiDREiQ0WyJqo8jECkBA8vdTYJgXIZslguFs4HZiX9U1xmjfXGIotnD7zkb1Wx5y4vbAe
tOn0figvkrwccRu98TTgRNEarG841oQTF+Fhxbs7HDYFOd6V+f/1+44aAbcORgpDYqGwe0/3hOkA
GR1gWnizZgzBIakv+VP5FCfUboleExRmBh8Slu+qZOwU44bFjNXhjhQDhPoiS86nswmUsA5McIYt
iQNLUyVUlr9yH9+P34I5KV2WmHYvc2HPJeeO6UhZ7h4FQK/rPT17lY4x3rl1XE7SXhc0RieldP8k
j8ciM5BdGd/So23u2x5vxR0RTcqlmaurF9S+W8l5wJ4uOTwqtAVTe94HSO5/wKhmhyaDaXaIcw5j
pRquvlHvR2VrIyifp/3bLWQiLqzRhRy+Eu5NO4BZeCTBOLWU7ERaMiXBvXEVEEUxfZkXsJQyzwNW
bag52XQ5XzbOSq3W2fUfxaZ+tUXuqBaLSTSOOLlAiF9LiIuD5ciD175s6yozT7rW06ZFKZfL+373
AgPzFfsJaUME29E98DhFO+WV3Uk9AIoYxTqafKtHetg0f3CIQq1JhnY97/Nt91dOop6E0vA7a4jS
+Vc5GiAdaGD73xRCH1L7g6openDIKXUGX8zQFPdx+6KhW2mnfX/tZzUB0tmovjVCYEtyBkhJC5TA
4hIUfblbP6ATQJtHdJggLNJ+dmm7RQdsM7ykkZeNFck3/pTJUndTeENWmtlEnenTZKIKo7DcHI8t
Qa8P4zHuMGPemmoyESd0u0VJRUONl6+b81oykl8HIY1eAxhqJyVEZsoW+6T7ejWsf5xvXY5hPde+
mFiRTnpdZyKIGCXlAOfRICkwHdc+aSZSevrEqE4JXnv8FzTYcBtz453nWCK9cVMiaX4zBVjYs2Pu
nPpcBCjG9mflKVcaQmnFO9wCCgjOzyjbPX6qML+IcK3B9OQpTKkgC5GNBGHwWu/HYBwTWOQAd6Pl
orCdPeFN20yBahY0PDLLefggegBcMz5hCiP5cZsxv1pUnx7MCxgNyGJkTkD/mxDQ/nWuYza46+ys
Jzg64iaZ7ano25pj4CBvJUtq76yDCG14L4iI7op3DC/SXJYiL7JJ99xE5ymOSS5gDXRsMb8Gs6vq
uyLwEcB82fp6LHhQJA9OMpLR/BltOkfkH+i6DglFHzxPDj+iLqh9EN94MnhQgsekVFduOusF+L6y
fTQIkw7qexpjH5UBm+muPxxsgmqPmDZqoS6hZ7vlNRPwnRK881IHDjJtqD/yIJeZMflvXBnRZ2MX
BxmAoc9lws+WpV+XKV+YC+VJ84X+Xq76QNJeZ7cCsmscuk2kvTKqURErUjKZKwBnIVyB5C4vvGxL
6u8RkU2XaKdhGU/EPVSyxl7MnYmCWYAs+myzoUBTXgg2vRgtDU12TljuEWFHyXmec0LCmd8P0Wnd
CSfNkL+lsnusoK1FEH+JfkMKtW5Pd93ga5S8D+4IfiYxaW9OYd6A7Krv2/zsUoz6o/jHdp+I2mV6
GYsnxhdhQaM5omnthJN3qJO9LZe/J5h0Ibd7opD+K9wDJTvAiIkYLl919fNXqyczCntzZMgVWg7C
GJn6hYWp2HGEgqE6XHPYOCpX3PpTxsudhufDsalwGfSmgIsb9Uqo8ShUnLqiZ3/kbwt0ycWpJsVN
fE/gfQ70O7gsOOuS4O817cjIUJVdjzIGWuMSn9z2XND3rsNQQsn96f8hnPinYYyGk3PNENCPETIA
01UODqvD6fPgx0aevL7U1+B7CjyNYwT7EJGCT+Qy/1NuIic6W44hHeu4ZI/5RdywwBHt/8jGkYWl
8Nu5PK9oWJmIbrL0GIyTqdaWwZDe0AWjEHgnQZMZijXiDBeAM2sHop3B+qJTjMgqoEMUtNoEaoM1
ZREwBAS8ujof+Fpo3VHPbfxKV/GIA12/7dY+oNANXdCPNkldIQPKjo0f4lmJF8E+q2OMRjO519RG
ISk5lrPBAvzk85qNmP4KzfcXbyxR/HFnHGukBB9dXL5OT+OAAq/JxS+4t0DVY0cUT+fhbQZurISl
369tYG7+xe+Ok9NDv9uGUM0x/8vqB/98V1dpdksbSBM6fUvfg/qtW4/abN+4KYNoO8uxcNdX3ccL
0i+oNNEUcJiZeB6YB9kvKDtYjYMLDM8QWHve95O/LGslyIXecStUP9QzLhj8kc1tr/O3w0dNj5YV
VfINHbVPbXl2MbiC1DuWzce7LYRV/oPBxy8FuQiBu0Z7ddMIB8tMOSjt3z2kANe4THWbLS2tv4t6
BK84MC1F6QeYyfJm+V5pSiA/cvLKkULXYFoNPIsWBpjV+uiw4qIq6+HGyGzDuSh5seSDMH2iGUcw
t6bax2yQPRNjNd5VuR5p0kNTOu0G4fDPWevwofOC/ELH1r5ojeGwLIo/FmHj23RyTD6oCEj4lOq+
8syW7L/FFGjkrMPH8ISK68Tm0V+UshUR32YUQNgYV5eftRZtnq62bQpoxazTfRZDtFO5HBB3bNC+
YIyUBZlICTN+qw+Gbw7LUQuH4GOUVoHInJai1vTCsgwZSDGI9AVDhpMkvol4Qj9lg0CGVmT68D47
zglBsu78tohy9idsmchNDCbNoeKlykuPI7wd3FxZol3kYCb4pSfLtm8gAhvnpJvE6zQHq/arD01a
9lQWfsZFBaVKGs5A74vJP+jd9nMhv98sgd1IHsw2IUrmocJEd8MHTQuWPHazgsYmqFa/03thRaeJ
17UbT4I8uX4i/0Gf/wqz5TBa1eyGIQawL7vAL3xFsZxmz9XBJ5TvxRWOoZbFBomRRxxY3DaPLhPy
bzgGESCmrJA2pOHajANz281KY8rJ41+7YJiuyZHGIf59GwruN0Ep2urVCPdb71hMluR3LxXUMO4F
vQQhlAvEWDyIBv5eLaEtxm9st4NMRU/xUTqIwrxdt6pEzDlhm0UMtj4J1l1S+IsCdghopCAITF2u
FKEcV+KxHP14VKMJA6DnQ1LzfllbaxlEhK4XOATeEp9wYKzjHD4/MVq9bDbhx20OyKcgrsOLD10Q
Nn4eQdTMeQLyZBelV9upPvuvU3RbYsan9uowhaDs2YrB4p+5tx8XC8HFqRi3b/NRJe0sad2FFkTp
5ML4IYTq1jnzt3s3s9QxFDUeQiwPZ8mqANhX/21zd9tRVfqOL2SYuOGBTOw98P5vNUlze9BrJoF6
xLDqW6VH9WVAzPQRMb3+Cr/VpQvkeR5+Yog0F7hLiTleMY+mmFvPrnAZO8nmf+b2RJ4pya6biJys
hkt87C2VtG65ZQi0RqunmLJJrPnThaX5zCT/+jkCQXgwLYkVrljPdBu4NSs9vdfBSG53WPqQOMOx
saSLkvAU5oq3qa9yFtiqnEbzRaFR1XeteKDEWLykmXMfP/98imTGsZhJHRG7PUOoLVB6e3E/UBXw
gInruT2gnP3hqj6WbWj6eFbIIaJvhBuFTrns7dwrXh5ueB7ooCB+DcStWPVM1YWsxLd8dYihUmmF
JpA1u/+MlIFGZZpfyS1BXtXmPou6s4Qozs+guevlwpYscTUmzu9QAiGUdJ+/rjhczyjNZCerLlhZ
Nk1dFmn3sFChG0SiwxpfKfkrzM4weqBqIHKBqYuw+omZxH6kCAi4Xx8FvTbw8iKBN9leEH9TPkn0
jOGeNMC9FShE/WzQj87uu6XZtd+UYVjSJDrSdpft4WNL9lLDfhS/ziQb8kP2NsnJuF+UKH/0kc1u
M1w4QpyN9gzlsJu6eYaF94qgP1H+xuQ+xwCR4BlXkeJEr6krfOQzovixw8U6Dxmcc4lY0ZZoP5B5
MTD9F+uLuNPR2JB6H9l8IzIHyuXtfPxMCAnO+4FMW0CTEWA6mpNXDKS3MrUNYrkSWp8+7qazIcBB
cFscMHoWVHhFQsVFd3rDRyTYVLvA4oQDh+uVyAZIf29ZJsIGyuTpLaUkx1pfe7Q6iWQ0O7il9YCm
QPKTsQZawZpbrgJoXc6URsjgezg4MG1XQeVv1GH5qJmRyHsFFdSRkD7ybz9eH3Y4uioc3L5QXynl
36STbC7sRg0SAG+x0EG9mzeM5LWBeeAXeKshkEf0xWnfdEJu6gxbhIAJerlIC0V4Cf3GmoujQ6MC
nTu4SUMSY91zOam4ujKI8jbjewAFcgm3rMomYUZPNstEXpkEp+5t2vOkQ5rI1W7TEcPRwECzHDlu
+iYE3MstUzOROW5c0ZK5WBMwaP4C4Ky+OzmiF2YJOeoLy8z7OT7K61CbZjePUYJjSdM9bUNsj8dw
sbUxbgBFfgC3yHR9hDCBhC5C2vxHghZ/nTbT1b4DksuFuarmwdSbBElK13UNQ0u58vg1SBVavcD8
+ltZBnhmk4q9/mSrr4x6oJePeyn64b1zlUbP+PwvO22XjbDMQl/9uiKinh8Ldz6RfLv5rp+z81iz
svJj9IrwptyCzF/4QNsvZOmmBBy0YDqR5xxeYZyq2t1KhN6S897X6eCwzgxNWUtks7Z1vpE4YRHS
DaLgNrL/Hvh+QM4Zpb3079Dg4I1xswcAXZuRPV2NtvfufvNg0NWd0DtTl2xDC9jaACoQS7YGehaN
9un0AO3/Mtw4gIOexvzN7z2Jvs8jZ7mtdi0TxLNH70d1XCivw9N5DZDDFkJPNIWtumTF2f6tqtQg
CMQ04s3WMrlusYdcmCpq7Mfl3oRUjzL5TtFKicEbICBgwt8fJ3669LQNk3icTojOBnQ4q8E9w07E
eMNC6HtQDffOy/nXo0P50TVzvG8vLJV0EpMVMYg3A3fGg3szrLRixAPFHitoBAsc1JyUrwZnBEo1
g4xrtqTvzLryoJhoz5ri8uyr5bDRKXq8vlGiIfcTR8Qv6ODOB+j8wCsnPL1kcFwgAGLT+2FhnMQh
OHURhcUh7Oyhd1kwEMWQPH1SBHiU7SHrCEysKJCp9nquqCokBoGbQrPQxEx1e+xu/qnZ19+tr+ik
3peaRPa92g36YhhP7EzVbBaWUk8vlnQYO8Um5StshTr+T3AK+fFvwEQTRFxtvw4R6L3MsVZ6RhMJ
MDCF3oOk0eAXmWzQwd53TZ/01AsXOx01RnC2j5C8eJmiJVWmtAUs0FmYRQrU26NNNpbrIpO+0ukA
cRwvciUhO7DHcJUxTBKXcmUTzxoWJAPYnJo9wgzRnPlTVKWkt0OSdniVt7OuMfefEiCzwLIfq89v
TdtQPQB42zvaKgon8HDdpj+Y3p3DlRzFQqE42tCTfsP0P8t07NiQR5nAqAyme5/L0QJaVJEOPNLG
TVfDd7GQ4oSb25MdAxJouRjRygo86kOMi2jMPty5VRnbGrIafpYkACzK4OiAEC7NJUZWX825Ood+
sYV/2ghACevsyR7zP3q0a9TlMK54zB5MVQPS6A4Eez/aEffn14vV51KU2wHZQJmRUZp0ymv4KOd8
oNJmYSRx7di8WwtZH6/R5WeAzO19y2viYdeIsuwcT2JISjlUjerO/pKvz8GY8oID8HYxiSGqGPgE
zDZOS5viBao1rd8HSHCcLvekxgvTnoT+BiRtSMi5VaEuQFdybkqO3n7eZl/DMzDbKangQRTE3sXh
7Vz9mwqhalVtC9wVWHQK0lAEJ9tuvmoCQRMhAn7BkqSDu/07WWXNZYSVGRt+g2KRk4ml5JcEbG3e
Hp38rShV+DdK1ULX5iFUOKbl6Fjqv5ArztNM67+9DTqRuDEX0QKJeSbzlgfuphaFUCzYbqt3z0wb
5YLqBijJhi+fK7hgUV9vV6fyOV3sMRa/+wz1SDXDuQLhDNvP35n6m5ZAhO+wmxBYqB32snQRy0lg
1d7xBMQ8wyh2/sqFkt5VzC15U1dHJ11H3mXitGmHOSzoFTjUzCEB8r3IPjg1Ljn+cxUpId4ugoo5
olAeTf1RVsE3lypSq9zyppQbgcni2OX5NViudmG9UpMXeKY0+0X0nxhjTgTQEbOSCv345hgngGTs
C82N7WMG8w1VgSBDYMACJS3jty9iBN0OCHh8b3nmi4l2OwYT5TXA5jJlDhiJLEnegqNR1F3xoEJe
wkBWC8cDPXMLzz5VPYlm5BimIqhT7JvvjeZ0IMBlwEM9Hqqg/K5y2rQ+lGU1vZLI+IOPm89xgLm6
ZGml0SmtuUqar9r8jfYskpHCa69BgmvJ41ZHXuc7V3bb06v9qfnpWLI3LTWpnoavmV+7HQ1aHMGQ
HE6i63ptSrjM9eUCj0pSPw/yB5jGD6L7XAHsbB0WCA6d0LiEQfbCRPZ35VZzYizkhA2S8eV2Hrgc
8QBKQVg9xt4LAS471c6LQuHcHChLjC5+u7CM9vq5UlHEiSyoDtQntzQfFGJ6TfuHg7K8x/kpcjfI
NwoSnci4WsPJ2PGRY6aADR81J35Wpao1ZAgesZy483o0BUFBVO2gORP0sqKI0a1FEULmLWA2EWPb
wMdtAcNqsUt6JQbaD/doF+T/eIe0qqukzteuJ0uq+QH4NxVEoIinMMWw1xT5VhtF7sUmsifHjpp1
2AgrWpvg2HPtZ78fy01/oA2KCC4musw64B1z6baZZY3wI216PJd2rtJE/lDF5uGXzkRk85pl1mvn
qIl7sSJfKuVRSsroPnSoIrz1L6TJAOH9B5RzMgQIwP7w0Sj71INjJZoQtlyycbBj/awMQkhh+/xR
wwSrFUIcoz8Z0wdCbLr5o2GOwai7/2/peCT8k+r40AzAdbC5D+/5/X0GoOTtaJNs0Ub8SHefEIcs
3WP9VJSPzABC7ovIlFXuj3HAszZq/BW7NECTafQ8IQi8QJmB8M731ZNSREpZwh6paTbIF6febrTX
aFmULd97QwxQoflGNsiU6pdkxqupJBNlWNlmyVNGX7raUzUIvjdVmB6SttH7p2DzRre1zGY4sabh
Mvk/bjqbUy+u2chC9hUjFam2KiJrzRX2FLWSJV7hJaFBdtxxnINeIYHYos24COT0AzdRnwXCDli5
50oH3je3uJcadxjRQ+E4X2+M4oKvIvyE9t0OAs0qRbk4yppmEV1DJUDJgi+T3X+wtOWTHqinBbKb
BFKLnXKUkutGSlP56xL5oweJwjZnTAzl3n+/hSx/iLSJc1HdFIEIwFG+ebXzWjqghQZbLMAbvDPs
qzxXLRcO+KEGkFixuQiIXPXRjDcQYOEPyOzidP5sgMooSU6xrYLwLGH3I0Ed479EKg6rrk4xtKH3
OwV0mXW9a7V6bTZ6Fg+xchLDV9LG+osldH0lcMaZcZzbEhvxx5QgSUMvFuNPITU2b4s8GvVwXYLZ
nwx7m3tWQ4opEn9cJOVMck3dBqY/W8hfwK6uwCBot3NCSrcdul+DIaBv6ZtsvFBibJKbo2j0r7fF
vZxY3MzSaob0lGXjyL1rGURvJZlSX86HhWFYyLMGUiMLDO2lO6FLyOY708cx7IU4Szq5gBbq7BcE
/V1RS8/GBuf70b8UPXD5w5Bo8bcZzTNa5chKi97Dl+nSU2XMZVokX1/3AVw/CPlk+hZWNeTTmAjM
Nkqw6jhjVlCdF4YxrBR5J9ctfGrE/eHRIlrFpKNllda32sx9e6dmPhnUr7J4qrnX8lYNqtAAl1kc
Kx7OoZVIJXFtYOGxtqWan1iD6iYDJ9tYFVFtE+aQOkTqH2C86zjmdjbnFFY3NqyRl+Igl58FIxiZ
2R0LT5LXf6mgDhwiLMAwSV2xbDmck4BysmZRYl8QZ/mgLCmJTa8omTtL6ngtn3Rqxmf7IWWnOW2T
IAK3A6JJEjEPigsTZOtKqTM3IUfgTgQUtRSSb1+6wXcadJSKCJoeEULkgxf/yJ+YBTO98db0DKMI
OwxIoFg4Vz4YhbVeFX/VA7HSPEJmWlYEE65eBhT4YcHhiEYgQaowV4YBuP+d+MGWxlGMN+aoSqCh
l7uIGNjNE+nksS/YkY/dN6x7BrZOJC2QvwgBVwHNDkdnLn1kWG+6cjJN2aCrWwo527/+T3+ZE6DK
GavgWUMG9l+6CC/tq2gPZFkQEUG0a0NGiy2kr5sjcckh7koXFmXcZKUxtVEZYZXyu8RdnXkUhwxC
eQO2zmtKxJKBQoonJEe6GRkJVylWystp2qadqObqBSjlhJDBUWsFNj9msSGXw5RVmrPphu99CDoM
Gnxt5rqv9wRDmzgpGBG8qPv3IFuagcyMK3DBM6qqHssAH49IYkd2Vi3QBNeP/0LN/y06H1/1K36O
b1ZlxnBGkYBeG2vY5jglyyA2VNNvNF4ueuy0PVby1TFVzipaq4XiD5GeoH57WOunqIwvOUYUS3mY
a/05XkIoTR3dAde2PyUNgjYN5sZb34VqrcNpGhbsbqAjpTY3iNRBhZ41nRKbg4EettGdSuAci0fe
wWToEJuh9HThv+QQFp8ZMClb5w+uYNpPdPxfE9/RKthaXS6q7uVXnnb+UmSaPrhM4uN9vVWF5/JC
d1kANSufwDnghkmhKmNINMDZxjW4GdM/RsLXTStircR3aXa6bNtNApZR2X6LSpnnU0ybTpPXRiaD
Nlcst7fA5qXoQLlMLxcwkKrpyEnaCgATKne0PcrsTYXq2sKYMAOXpLPCZLAJkTBLweCAfQTvwow0
YAy63FW7y2ACuOvk9+3OTi6sMcRkEkUsycV93Xhyc6EYGaUegADE+jm21zwoAW82VeWA9kKLLc1V
SByvOwbN1+DiLccWYn9v6ygrBKBNbkXV7qudehlPcRkzy+bfGbW0E0seFWeYF6vf2I675UmDWnSx
P4qz7IOAQAEzBmvTiimbdim9UXCvwqmHYzuvmHM3WgiEiUpCSkmiBpLpIFrkAaB8AcSmo5wcIXMN
o70HPxQdPdjDhy4c1sIzwBrk7tBAdWtADobV2vvVzwpdaqp5VnHAP2BXz5fuLDZ3U33bnlqVImfO
SAOX227bY8r+YpeUr7eN0/MLWBtpmnvFO9GggIeVNsXVyOrPa0UZlcouloFULamPYvvoemMK6/EE
lqr/JQ3zjRUj36Rs/i10xRn8xAxH+I8LVWsxG8yT/K9XdXfrwSO9ID/w0xk92FDOiprZnIoozDgP
JAfZ0GWrJaWBPLQiQu+PoZfK/nbnv4aQRHqBYsTQTyd3uBtCS5SGJm6N72rp3kcSZ1OF3nlIlihN
5or8wU4JwWuDl9Tz99f9oiujbNhXkUZ8tQlau29xTggAXmS3auimOaK9YS6FUhyOD1L92zP0l7b6
kAWSoyCQv3ljs9BvHsftKlZSFDe4VpIhl0WGHMT+CbLGUbrQT+OOorq5O44u+v2JMdtqavDJMmGO
SSuQjIfCgN7zHF7JxkXkxfA91g3bOsKxCbLqpDMWlKWeRTXcFtsO3i44v25tBVN8x+u4T0hW9xso
ER64NV4vVtb/QXTfASAhzq5YaCis1aUQzre3+aIOhErV7acvb1I+hP43d60Qb62QXDk1ZdPoYC4B
hczvjoBMItp4MPwtwOu4to0narUwTVGF/Q8nwRV6BSOHTJWgxLhEH0kwsMt5FQU7bhnxbedER5Vt
7Qra3zWpsUWqW+jn40RgdAx2KykCh00UDHD6vLgenQfx2CoKvLauW9kYM8VUxST7xYO7Cuo4H/9R
KQiUVDIOIDpPReaK2oT+8O/mBN2t1ionneEtOvZeFaJ/fdi0dFJd1U41p6IjGFk5jpn09w3eTTPa
cEE9OrsO1cYpAtgASd+6CNEyNv6LTiECwv7SyR/Ag6e8OKC8avv3iZabm6KMTYMk6EAD2/IyIxqa
V8+NWreR5mfuE1TWpvW7FP25uXoOiqfAfM5nDjgMxlzWwpqH2JL7bdy8+nh7BBwYGL1Rdg8GaT07
00BnG81bLjfmeqxUf9a0ez++r8OcECSlURAMPmhemS4oKxUqcylLyBFKm47BjtIOIWZIpRrEPQhl
uJzX3h6pXN+Bh4RNcvUXHlTWZsin7xMWRKSgL0cpZJA8B5D6fLlTRqvBVktRfB0maDyzyyhBhdxd
SNOjtOB+rNPu4WYYREkuOxyw+Ln/wEZn0/h8tjYaHKZbUFhU0xfwr1FjYyL3Tzg6uRktdgYYmDWX
uWVn2xyJsplso5kR2wMCmCn2M0J91lncEh+xeBdX3ED9bcXP5Xu1hB6Vy2qRufDoy6A81U6mRF17
PeY8o1zP3MpmfthVfy26sr5mbP57ge/gmQos3drql9xkkmji4Y+s+saIPCH71nFrlfcXp/v4v/Ug
CQAZOk4Pq2p9mGlZ3jL7A4DpLOqXRTXBXfh8XOnXSi3inDT5Y5/2KMsphuQGpjocsTvwXryxZuv6
l42UVDaDMZIiAS+3NvBL68pR01a3GN/r8CIAYjlwDxfQn1G0gZTnqrM5hNTQNNNQBueH4lV1pg3M
xU0zbbByacg4XCFifN0CBJWKBh461E0cdA184lzGc5Ky21kjwTUkiFJAGj+gx7e5TEi7osBBB+kF
8ih5wiNaaRnoX47SzpDpNoEoQ0tkdpbdhCsARtKfnT1ISVAEBGlnIh3zGyC1RUL4dLcJKOsoMb9G
YJlb8npz3YGmvce2iohNvZCWLGuyV020p0nBbUaO8HckQBZVuzLj+Ixj0RZHxPhtqHCBbkU1/+s2
uvGdQCf4SrMLqmtaMRcPkf0uX2zA4ShVAQ6tYPMRQQTrWL3uGyPtr8oLDheOUyKqwWmqDP/+LAo5
YCuojhCvqjjGvfKe1plcqSoa94lsAvlldhh9T3EjI150ni4qST9+DyBFaFPU5NA4oW2Js6OpnXJF
Ts05TtnA8SQo02X7JkuCAcbWeX7YhUmrjcxGd//JHcSZJyhr7yThwEdXBA5aoWSm+z48Scd5azHd
WWQ7sXFx4C4+YR7NZgDRSlQFY5YPNxY3CKxSc2LRe+iON94w9irCd69VSMRaYQMT2Qj3AVEvpwUu
9aBDh44XGMmW6frNjNxsd/X2NSOcqYKBMLliNh8DA6RemXyNC7IoLyZMz/CDdTPa9I3V8Rqii1yo
v/UCQpRFw2RuHluv9g8hmbUoHqYqspjTkLEVU9Q6ySMr9Vd01ZxvKVDKvWRHhnUCkxWLA2uSOg3a
R7FAjec6SkSnssm6XfY0hrl7ofwwWamEmrvgN27Rl6g5Wp89O0Yy8eVtixSy79P4ttwiK30FuhaS
dl/MihQq94XjvY+WP+rziH5aaI9uc4yfHZoiK0KqcLRYV/3BiRUUZ+jsvSADlpSSsyZ9BoHPOf50
shGZKyvwMlgbR+HSU4sXM+2dVgPfbR2ALTqpjS3cyYrpmUxs8jZBhax7HMH6sfAjgTQG/SzL+jGJ
JZi+GtyQ+f4502S881VITqNszvyuyCQHfmTEtcCjSnUKZ2LTZEleRi8+/2FIPU0GM3anFsg7jxpC
0W6me4LgUqsXgyyHh5RxmsEYLojxq6wOkuS96D4fT8SNMv/bI0rQvZa0nBYDi8OnwkKceXmaImQ4
xDXb5jkF3G/gZlUKICHcjfCse+H+d+eGhD2B0rntPkYciKucp3yaTI4Fe9qvL3EfK3B/8upQxBAo
8g0oPPRxd8WTZeWSJcpbJp309FIulVfX2tEdCrC+YMKqiKkf667CTpNslLgtOLIU0tFI3gudWVEN
GreppxzkiOjydDycSpg0L4Ukv8B4Mxx/Gl/NfTRO2xtOhta77nTX9TgWR1PTKzJ49Oet4synGoyQ
98lixfF4h9eomMmZDhDcOARn0jjvmlrL2faS44r6FGNfkSxakJ0UvDJTKrb5N8CqEdKCMjBBwn0H
GTZl5G9upnfcj+7Mr4MbMU3tA/1PNnUGNbGy7SlcjvOcgBkZLK+53xfEvuPwwEKisqciq6FEO7w/
xkhbUZ969b/krQF/etf710Fh+qbdnW2khp0owB+XCPoaVMarxd92ryM0QonuJ2+DV9aJsloSH8lF
1+jAmA9V/g7ugx78lmYeGJjsIQIFR/NsQZnj6/zWLji0YbY/UZQIhIdl5CYURG5IMx6Oavq+XUqb
ArCclHOcT47ozHq93x0eOg7Obb8KY/7iv4R+ULbTscQxI1aITO2rfvB3MQPslPSa4ePKBOzDKUBs
ZHGvx4rfVyWVVoblds9rJzX6DXilcXGueGCbYOeUFuNbQspjDJOML5KqHalK/AQbsCFkllq87kyc
9+vHRi8K/kU94/5b48d1pdUE1Gt0IcaE7mM0Y2iAlKu/ZL36f0E/Qu0Q2Ah0Q33UkctyHdmI8cMy
mPsHNyBmNW4SEcPPu1OoA6D1bXZZAe8Z/1tMoRg5617Kq/eym8q8jlY36WdgTEFxjWcRguQZTWF0
NJ7Du8/qpyDtvSP0Bb5nzfZ3pQumqmLY88ZDtzwcJqYEbpnOSekOyw9srjnwguGjv5X1XBoC7Phn
DI3VNBPpqNWG45ZdLX2RVwHohLyJT+1t0QFiZtIcesUwWDU0MJWdGgzmd3qcCFYp+XyXkF6xteBS
M6DYXpe4cBMtFCYT+H7ESR9ptl3j7fzWWbt/QPiUKqoihEWvLLDJuTFTOq+K+5TYBh72Ui5wMrMF
Dgk9yOgItEevoQj7X6LSHMQOQaV2m06FERAbVefpV92cssKyxe51Of/HimcfeCilMZL23Vive1fW
HnaVqXhw/gR3j08NoC/qHnv55igF79OBD60qqx7ELzN9EfyAieZkE+hDlmcPvYyDN1YjlPpEkEip
m6kaQHqhjeuDqdh3jZ7wipmWj7feA4f86mpkXcfryd7LJD0Oa+Sr1Kqdvn1OVxxTUMyKPzKVJlDb
m+5Kv7+MTKy5pXwSVANtSUDdPQzT2YXLHqedK+d5uoI61Jn4xVhqfoFKlx5UTl3avUBP8W+sakFA
s8L1+in2ZUH7n+M3Acu5JBHc4yCSHIY1y0N1zSOZkTNgq7q2FNq9U4CRptQA+yA6sEDGbm1R/A5V
cbMxx7MIYxpqCMZucfjEb1imB3QRz3KSlBCQ6e8SmiDrJxXeISqSd5ub+eD+eKB6VsQmw74BgLCH
ZqAWWOrjGhci+8If/g0rCLaN5jmzxuAujGigQToPcwY0ilGjGyNprqOevBYTDNsxwSvCXprWBB1f
XzX0loKjVrGX94SfdPGW8d7rHPojGfkGlq/tP2PgCNrcBN7w1nG9m6RovvNMuSG4/00g63T6ldQV
xNm4etwbyYwG8slHXhBlcknj5j44XwrrQxP3yzyZYQ9HVq4Th2yUPVoNuaPbkEpZDwjrfqKdv86x
P/hr02o31pgpgM24cnZ1kyZT2IneORw6x1NsvhzV1EzvHyvjUaDrqcwEAUqy6Bi6pLt7H9sTQFqs
aX9lx1LTXp8dbHx44oofqYUXwgMWQZwZQsrvBQRxWWIW2LNm7DaCkeiulYfbJ4WPo97Z7YHs91N/
HVuJJe5C+yQGDDpPznlD0bnhyAPh6tCGsyLASLANcQNYueMAQaiTyB3n54NHXbtFdUr8RP+npVfE
DjS5QR+ObB+G6Rt4Uzsd3mcxWLzfTrdytUoQ7vVBRQO7oKjVWQEK1t8VA/czfa6l0jKYBcwEQoiV
qA0JNnkcmwH+2BpwVsoTFtssMFrNnUpyQL3ls4W9kGkdQjJfZgqrBC7xcYYrdv3VbFfR6a84HAqT
rPEAMZBzxQrB/DfoNfCKVi36EHhGKcpoC6TPaO85mDEUVwHOnMsruy7t14X3VazXOCeLJuk4w3/E
HUEiXFDWnhtySV8BWuwMNjdJAFKNMhfNYW6U4SQo7NkUeg5I8X+Yrqf35Lp+eHIzK2sr4BM4zRe/
bAIHij7zneQh+R7GBbirD7IPMHI+ym9uTZ1aH7R3Vmk3ZS5UKGoG8oyigVxYq1ICHYAko0Va4W6R
CaDTFgc+kAWWcLdFqySdVhleVqhsMLrOpXDpsBq4YLK8ZIJfG/5JYzKRLmennwlzTCSgj5C6xFkI
0F1pNSVPaQBUaMSbzrgT2ZnZgvbxFBG1qtsZyGbbrkFgwnJLYfOlj9QX/rpSlF2N6QhN9jKwQJI0
HV0x7rWdHSRTmSXFtuT6qbMMyXLF5bRru0jjFJ6Ey9j3PSPhvS1RoLlfTW2cUjH3nYkEB2kyzbk4
fGfAhBaxNeeUboMBpqQd6LkQhaBM/NAiZsMLD7GpBQwTb8CrOvpONvSihIpQ2XWCLZ1l8EHZw8iR
FbtpKYONZx8UNSVBSiqmNgpRohP4R4sF0C2yBjGSBBKySfK4GewWbAnY2lLRc8FFyjKlhSsy+9+D
Kgz7hiAMErVX4TqYN157EPdDKXrF/dY2p5ss2tK1tcf1DaQBFsw4W2BGsusYAmA8tn46Xv9B/Cps
H8oExj819a3hpT9TQQPHruIsn4J1eQxXAU1iQ/xcTQOWwfkbHbd583xzw2hViUoh6GqTO7Ld1RtD
SDowweUUxgHBT0wLXh7D23TvMrl7IZwOQPvKqnq2x9UUr3EFT8Eo4RZJF9lhqX3Ev7TcAmBh4+aS
fC/ORJtICAQl/pMZR3GgJQcPFrAlqy2wzUW69ml7guxMtze3TcNubBlGoqzWlguUuXl9HNiZXLhw
FBjXFja5p3lcmkcEDWNnnYlxySbb+ddC+8YQWH5OXflkCxNrU6N+rx68RR7ylHgl2V+WhUVbxBqJ
WiNU088F7lqSWUGYimfAhTH4pAfYX89y/R5DLVINXSpKTyQ20Qqs3RRiOqpf3nP0lTbJD9u6S2kG
w7pLoLu3iMoxwIfOeJLI46jE1SKC5HTiV9sHlOGbITLN5kxPmvqi9TA8YvhG1ksdwOj0sAsxV23I
gHUeU3MEj85CUsBkQ2QYIUeNKr57QI/x5D/+9VpvE080phStVUNRmP1ZInoVhGAix0/qYSoFlSDU
OVdSfl7IMwEOD2ozZ0Cc0EySxDC5Ltwnbe7OWxnKI5Wx5BTnBaZaSMZ264Dy9dFOr2777fDNoAni
55sJ82BEQJYcSxK8CP3JoCKSjYWgS5EfJqRNR9cefublkn2eux7UdsLV0Kcd4IBvKyQiTzR4Gn37
uBOGp2bvaSzgYxwZQYxBGVUoT5BBXxVmlT7QxuYmyKPl0zxaUO452BdcuoeKe4+0zV8aLxQ7nw4V
saD36mOobQiu/yRA/94G48elJhY1P18ZymyqbFl3viS5xLDd07xS6xSqtyMbiPo2R3UNtZIs+x8P
vr+0w9w7I0ieNIoXSRaXFE2dafEkFkGhyC1cihnlbBO09Wr1M6MOElTsPwFYCUJyT5M6Tx0wOOEN
Wc6cC/7/5IrtS7DwiHaB/dDc69bFKRsAXdYjt9D1EJjmm1GoNRIRCaGOpcJxMAGriZpLBrukF4ne
OR/kB0VTHNxUO5k05vGGlKroYB8fcei3QlOq5SNw3vk4SHFDnWuVvsyhly6k+Niu55S5B59lh+jq
t0sRBKWdoLVGx2ihFJL6mhgmsYaK/93nq29xAWgtWIt7hM9R511Oo4nqmDMT7DdEjj80gCjkeJTt
4IKvj+baycuIrbWOKqzKDQh3YnQr4xactJq8XXiZYEsJP+Y6e6p0x+E0aFRl3StwdxrmJz1hz5Y+
XJcEG2uRU8yWCwt9aPJCavWuwogzryFr44yJeFfoDVQDqe+0yWEauSMBUwUblMbvI28wUaEh7FwL
UfPsOjRJlQODaJf120hA/RAJJJf521vj4TSAeWAtV972fZcf9aRbhmqYKzc2Phq1A/5nDLmxsHxj
hCZ8XDudaxWDhg6GoDrQL3dtZbEbSnceCZp125uSIESrj8EbFMDVfdB5wvSb6KmJTdKlCYTNZaIC
7MHwUFrXF73ZhLKWHteKMX4fSaDKGxeS/wdYTNsEorTeMCFNNI1HG1ZKbubGIjdNsTF/o/UkF+GK
mCI/ROey3uutrnkuVVl/9Cwnb72Vopp/2/+7YPqX3PklS8cJbJAH+nC1sf3AKIb1097KhNrMymWc
w2SW52ZcL6M5S6QmzdtPd97HF3WWIIdialTkAZEbtocDqmN1k32e8F1QTwmn3cND4rREBy95aG6h
py1mTWr7K/8aV2ZbELA4vJLu05cd9/6b09tUnzZZ/KgsctT5UTYIf1uKBas8TzoQhPl3sjKdVRcx
ywk5NoBOQXs5AWcD/9jhkgiqdmuSJoMGw4XcYtp2/c0Eh01qXOyEoDmsE8AhCW8fcqX0nhFi3tia
oC3OurKyunh0sR78lBHJrT1IOP5zR/1X3PoWOBO9cgkSFdPdGFV8d00j9PfD5aCQFfXYLVSXx42J
vxThte0TWISfdqmJNQPSd7KGTmAlj1Srr68BihUPhALfovQfWoSU4dEBOJV8dtRgNFnyw/8G8W0b
pxE/e5LuSAcDQjiWDWnx01lJnKW9G4pHI7fFOATc0zYtyUpHeQi5/QpPmmtoB0K45wgrnTywRSJC
QpZP42C1QReI1MBg/P1oaqonmNi8dnZYd3rtmHCe0AFRc5WYjRhOrG8wiRTaMU3cn3uInkkCNAjl
SmQvM2NpfDkl/5uNzXjCj+b9Tz6WnH1Qn16f99rYG2OCTQ0fSYYx/nCaK7u+DcptE817XqHglDPr
kVSi7NRJl8rMReLT3UxodEYEBy3T8kMeb/sxlxbuEqkEySvYx3xKCKozav/b336qwzl4n2dq1uiH
ZOjOKDQTVuvVK9zibRLn9tt39L/3JvOdn5mpYe31k195gpWmBOiR1yHd8SjaN482It1ip4uwx56e
vyMF+076QaLyUwaGgOa7EWFN7IA02Gfv0zcauEh28CWKizRI6cX+cNIrmrDJnFY6TIYPheVu2swx
ZY5jGEw+KoBxxp+SqxYfgCJqKUgJtPHynko85GSrnOaLemVbe/W4lmhM4sTMbcnC989R7u3WxFBD
M9H5Zs5GSB52MSluJDPuYy7WLaDygYr6n1+wpv642iNwJf/NoYhQxeTXL0CS+PMWtTLqbn54JOio
mIVuNtl+sowqyCP3bve7QtjX2LTANC+fgZPN4mcITE6Xv3ywiCF1kMzwHKosacObdDtNzljnCFuB
yes7FGFsBQOssMW4XFqj/oRCItRNHpN6ddu7GBTpfrElDR/kKq3diliX/9dmxtkpDfZfNpZ9F/Q0
UqE0wNm3T9MOiCmwdasNFCysVyfWPWe+S+IPQnGiV5zKSW/YpClv3XXF8XqZz8+ws0SlLAaCoQC5
ovtHLRyOHjJax3M+A+jkzXePNXTeEYosMAP1x0hTeNn0W1tqApH/JqIApHbA3kKegTb3VWy27k0a
ViqzDx6nA0UQhry98GHhw3956zDFwscPI2Lmu/UF3VXozLadxmM1f3m/eEcRylNTe5xHGcZMKoPF
bpMqwLksVJp4EEVy1Ir0ZTKlk+F0zOhKBKLgs7PcQ+hHOwPmVr1VkqVtjzXu8A1+CNqoK5FGnLDv
ePipR/OWWcuOYT0p5V6rLX1LHvlqMeJwz7eeONI9iiUFk/oQSpn75DViqh91v0OOQVQtoZclGXY3
ZEaNC2uoy5NcGJVTiH4If/iWrVVo9/og+Y8HSJ2bWGTIAN+gd7LYIiOmJYHk3bGSBPW/GjDbIjE/
FHh/n8ndisUWw7fb9E3kcix/ViZy9m1FI7xEXiK/MffneQANPhVIIM6qtjZJ0TE2nixPJ3RVTgmD
dzZKKi/I9Q7LaHld0IOjzUwPvz+nLTW50B0UPD/ua+IjMKkDKlfKhb846MPfOnPpaEC7iBF5qhF/
nlzTZ9NATKb4h4YQx5o/k8fUvPbXpvcGLE4h1Tt1w4Pnr/egDN+gQ4co37W5mnnUdY1FIj5DvATx
GACiyhqgPN4hFsBARH9B0HfyGDDeGAFJ3HZoFTnV7k7BGMR4AVnzk/0/no5kQybQh+uUO0oyeyjz
cGSjXD0MylyvtZPjRHz9DCkjV+TiU13fQw7131CdWGsYSSR+MFrWuUsnC9rMXFmtkwp7pfSIJVyW
r6eVzVr7ML8queKq8fglfSfCZvkHeFAec1nAh2vaWuDiqKCdelDHc2w4d1o9/o2nPeww5ptggjlb
x1xp7rYs53TMBjdegkSQxNsauKNhx4Jky6h1mxzc8iWoPPlrcusNO2SJogg+nZSXVtwl/fxZpvKl
us24r6/NCsvSD1j7lk/hd2zIDK2zcT+LfgQb1dY0fZeMg08BDOHpuKiBA9lMnuuJ4fCZ492WACGD
Z2qdJLxE72bDFVNBnlD/TGL3KbNrcAocEa0sekaSt0BK2Ofqi0m5uS17R/3gmkfjl7fGuk80CCr/
rLcFxMQZCfskW7NES8dpYp4hAsHB7eFFSGky/RoszRnNmbnSYPeRkNuxbra5g1hN3YGFa7ors4bu
FhxoVT7L5E/1GhgIlFQ+nUHK2GKxO9RjX35fyZE/+7o924TwqziW7uKIDLhmKAeT3AHDzafxUENT
k06Ak9ja7YKyt1C3+yJ/dFBgTrHMx6el23HSiuQffPt/v8iI/uVxybJyU2S6NjWJZ+SGHphQTC9U
fN9qs4X3oMm6JS7SUbQY+sd8KPLyrN3TukAljBCznyWCmus7+NpTMEE+SAscB02V0DbvZHyU2Y/p
pgZrDx3qiEQXKDX4AaZQKmoEOeBdP9w16vL8Urhgoc/dCFaV4LLvjVosYj4pqQLJM/p5TyaIX+wY
cIxpl5mal9OS6dAxFvuFvQi9OmXoSwkUZJiTJctCL9web5qS2z0E95Ng2V0GAGZLtx86ryFwRMgB
l3G3MTaG+dI2JTxTS+8UXv73D5Nhb32l/1uRtV2pOB/R95Eo+vpryFk5sVrwjXpzsitDPkd5EE91
/Y+A0GD2IdxH9hEnSIIHHhLZ7tJnuY7cn9XWog8nVATb9JjQzqqKUSsmTYRn6VFJbkOEBcs5s1Bk
ZIa7OoSHiCd2J/bMG0kS+lT0Dgm5u8xv7CpxDXRxQgNLzyi8IQ7kQaUJzy8deDDaXbPAKN2tSkKi
DKBz33JcF6kCngzEe1B+8spjXRXCb8Hnk4qrwlL5wudU9z0kzysgqd5NYNcFpOXZwCpJ7bBB0oar
n1zyZpTfBbVpO2AtZcPeR9e0h2+XgwjnB39WxlPeTWsmOUH48KxY2IxhRnp20wViIhFJzH4zfMRA
qJ/nIaIzgatBVIWf3+SV7ezYFMmnG8X326fu7mYF99hlM+6rbtmTauMuaor1cmn59yMDZH8ddsUo
M85EaEJTAFSx3hzrdvh7HaNWrOJISxYyaIJLyIFFYUw2KeMO54/4cUZptqM3XoNtAH/8qscAGdBX
wf3bg5qbIITZK8Omuuw4LWDQlE0uxyFMglH2FlXFrDK8cZjoQrEQQKdFiIhn4MbHl/BL8nWn5Kzp
XJDE8ltg3+2svz74O7KldbV6iCjvzu5d+FmV8DLTw5JusCcy+R1zD18bHVqNPko5U1OgDlczBXBk
8UDeZKrefuc35nZrac1zbTGJ+3nnQhzAbiif7Pq+9hk0ZZebC7w2u4r8RQuTEcjOcU2D5xTrBMQt
dXM0QCfDRN+nO0ZTmM0AWzuaelHireDDSVQwSR/7L0eSK/qG36u27fcrRtIsYYIjgZYI8f6X/yvh
fI2dV7CIEq+vTrGndq7qyi2dJsh/lH92oPd4ShB/w+GI1b9k521rDuxN/+xfg6VOXRVxoPjwVuO+
YUTgk1Bp5RPTDb8X0SBOsu/jk5XO89n3KYfXN75mBTLX5inCBUpvrIyAwGIMUF50AKzHzb5/uTSn
+xDGh+MAgv9ZmdPfKlYzgZkjJqHJ/YQXakI4UaY9gnUENkidi0NPvo5626zHup7LSkWfAAdnBTe5
B2wY4RyIgVeTotRQlPywNFpqLCMcP6Hszq8TNWkQonPgLYr/7EusuzSRScTtEmxwawzX5764l9Jj
MeNBKm0RIkfUfFYMbMAUSFfgWSY+2V4GbL3yinm/cHTgL5Q4t1Kn4VBrNYB8KVY0Y167V7V9oHJm
6s/EQXGArQYVEdQHFS8gL6UgmYR/Oxuyev6vVg1oPDiKyUcVaCyhbvgpQERDj8Tvuga/o15O1CMt
fCS7b+OCBw0FkeQEQK16Neapzbzn9YtVAF1qlpZhRKrZP4aZL4GVDwNO9B7pd7zAMZPShd8pj/im
8sxGXXeZEl5oAdsgiXvqtnFEE91RYis5Ujy7dvah/bd1Dy6HvOwp21gqYBdumhIRS8YXW6jXmr7s
Fc6gxNDo0lD9JTVTHHteG74rbFXFOVTZBUYSQPGBQsmHMq+Ir+Rv0HNf3NumKyaAQMh1NJ+4CM1f
H4Yn2G91seq3H68GmKLEYBEsX1kAtfbVe2sKN6WorLCeUriRlCgExabm7THIlxjUcWvaQuZmQ0JW
cK8pdAd69uFOfuBOEw6rSXiXsU2UvlBv4pRn+W2HtU3gVGiSbTy7TR29sOiaJ6ULSERQS4znBgF4
CI/Ol8PdDcFBrU7TqLe1+NuWurFxNyPGW2OSBCP6UUcxMmU8PU8G67jqbMf9VHFGbEa1PjQedHT3
TvGfwT0lBLkO8V0VvigTAkRNXwSYmGg+wh4deecVnaCnssbDfxEFt7htZKVO83NmZzah8lTuBQkF
jP7NA3gExrBLZUXVDOTFX6CaltAWslOLqURXRanySG7v+rEbqmFjg2L2A3XWJgI8zrS1HXVw9tq7
2vHhBk88Nojj3t0fiA/Hgih5NMtugVlRQOaHF5W96v8T2b+tpl8ESCOAOJKqajZjpu2ZiLyKwAXD
V/sLhvh5ZH07AB96SHxoZ4uSDfzscNJnn1guw3OHi1zp9bhNACvBqcEH5OkDI/t0RjmdFY//iZNh
W3t2mDFAEgmrlEcdTw57CFf5KhhTz/p29dIwmQL6QvRFiVuIFVUQrccpYiGYcZNvEa1w4NXV84HN
d2ESNSNSsmKoNq9Nx4jWujQHY+sdNz4kwY8kAAHa55h2xDwvlzExKx1SM2rftFlv+1/yA185CumS
uDIxCj+IHlHPhHT063Lq9opyHRk/4As2Xhk+s5Xn0VVriVqiC3x4mUT7HE2TUvLego2uD303AQwj
6dqlw2nZP8Zfni0PN6RSrOG0+dP+Y7Ywq0oCge/K2XvrovzyDX4frey+RETLT72RBNYMZVf2pJFj
ArwUPmyHnzyPUJ5+8m9rZ+K/pXDNUVZDUFsmaxEX7P4rKj5jCJ/fMRL61OWBu1bGxbgAQUqoItDh
G+TYfMTMSd4tkXIJxHN8WnQ0x3gZ4f26EzoO/L9BRWFJnl+MO0MWEuwVgIzQ1Kot/6zlp4o5AQEt
0ONsLLInhZvnZJoeYJpAsGKO8m1mPH0dImrazE6GqRe5d7yVntCHdI9MoSskX+WA02rq6DbeJqgZ
2Jf9+9/SQqmMFw3QM2McYAJNG6hPOn0JzyQ1nYXqa+eKZiO3ygnc5X97LTIa2OAqRSqEgoqcADlp
GCnwgbu2D5URRnVz4Kx0/0qguxFuvxZw3Jjzr7et2y35ElzBGIrm98xkWu1l74uxxQIly+TgU3UW
CUado/OcCLdqDfIICEjNsa6u0yA99s5YjuBh9ZVYo+S7ns918S0YnAABFxoglqKPSR5zYJecz62G
wXMdY9epadiA/cm85w3bSXZXgf8qkkT+Rp6Z3kobaofl8GHZzpAAqfHfizFhAySYhAs3maMzUOTq
Wd/HSNF7WdQHedKJqSoKVNtIh1Sc29qEUqrB2QPhG07J21PV4Bm7oX/Q57uM8kytmRY6bKA5kCAX
iOtxaxPmeZQykBogqiELUfXzZH4nbajYGZdQW04iCj0c2DCKRx/nK3NywemP9L+IE1DQ8ScTyFFo
6dSXFJYltfyMwWxAk7lJ0QbKfvABE9ueM2caes3FUmzfeAnUQWStXqKPqtT68RMpQ/aVatkih7Gz
O2TNUx+3VxGKKc/Ompt2sYLphZXZesB+ZbXL3XeV0d5oTvigwpT30Rv0B5+rMTsz4PcHFyvEbRxT
cjVloqbYit9LvaoOKFsW003D+De2T92d02tXknSx4oMEkEHMi2/FkRLFd8JROoC72d3fm4vSz8Zr
PTxrR6i1oWuJ1YMFXs8kuY3xNEXR/mNlyyc9jb9q7+NQhU2AD8r+/X0HeqtOxn0iOVa1qOTvQ8CM
RB8bLcd5Hqp13sUbccP0lEDq/N9NGIuwyR4Ov44Dl97ldoQQqehE/NOfQNAb2EGrbn+TI+wrRz6p
p6LMHXkzB5g1DghBHIHgCmpvk6hjbDxVLgRHOG+dIU1pZfV0ZOjtJO2RmHJ6ZsUrPKSipuhbiB9k
HyhZkfP/bCm0hmvkgUExbRUl+WmnBN/zr9LIamp5A69K+ysjPzurtPQGyDKapobvtZ7lyzFZknL5
DKIL91Dnr/NvxXpFlY6izTW4sStKc00Vm6TiNfYIuDtD0a6t+swqap7sv9zQ7ZIwPHwKak1NWVHK
24/XGCEV35R0lYl76qr06Sn1N//efh1OFYZUpLOZMuP6RMY9JZmQfRF+8wUTwh0HZW9un8SaF5EN
ldVV/EgtP1rwzE/o7tqJ2c/Ad0EORouevhKvhDQhISRwQk/kH14rEq7XYbOYIfi6Rjp0PjvsNb23
X7cHQ/E88Ewno9/kaIqjBBdAqpWs1xoKN9wdMSdoMLfcekdWr6cg7GuK4T2QRUzp30NpjJWWBKxE
PMUsDK8Hf0yZYCyJ6y6o7WFoORRrazxQJX1BiMUQkFJ4VP9/G1Zmdf3uquPuhW7gVoLgXtEAnPUq
PzHfzgqMiww1ZKyCyxkISR0F+7+GfoOzfb7sKl1pZaY0ztGwwow2lmsKUFp+KXhRXw/e4g513Png
UeiVKnG0Xd3EMBioz+FDQzkBywsuPyqOamcU4jxNqgm3iPRcya2PVtIukPOC4kvuPo9aXSexc1dc
JmBjMpHwL1dKIO5VXSBdkem5RIH2CavAuLhD8+8CxuwIjAEaksx13G7Tpu3KUkmYErx/3u5+hAaa
ZA8bNOOdaZ31aNzstzWgrbeMYGXIwWF1GgqCw7vxW8CHtM/EG12RPPYB4JPYRUsTfrnd86W8XZZH
N2PxY2/7ymv5dzrRSbtuhxYrz4YwYcy64c7xcniMAaAzF0wG2ryYR7IhcHnk/Mf9oOTt4SR4uubH
6gu6RevepnmsZ1lhJiJWMl3yM9QKH2jzhmFr33TOoMgLuS0gssUv7mKvZlnT2PyZNNFcRmOWlbnk
15STGkKLtgSPYwWmKwEd3L3TG6dJiblpuxqyp59lbtL5TX3pGeUV97dWiJY6Cz3J057KZ3pgtDGM
VAQB02/iVOnDLiBwm8crfR52NHQoCtlzgGO0tRI0hIqSj2Aw4v76tUwurfW0wGkUUG9BQlH5MOMo
6paSMEiD/eYlhDlkLmw6vLGfzt3iLT2aUce2XU4aTqxj+/wMTQlUMMpP6ock+di+s2Bumg9XC/Bg
ltkccPTgZyFa5L1geEBpWn3XBXMRzFe3o7dXbll/2HG5NPelH8IfG+sBP+t2jp8SnaXCG0d34o4y
b+E00aabZbhciCRXhvmWNjvsLUA1esNYmInYsvI2sNZvqbRZELLS+CJFXVUq+8BuKiPnb5cArXfZ
ZL86lnD3k7KZQL8LEaQrO+vxo7ljcn1cdieYlY7NhQ9n37kdYdCRWCScN2+pvynkEa7ageIZox1+
bkkqtYF1aGcyQWXqxtZ9UdzAG+8KOBwekcl6olbP9lOnL8Y36cA2gs281hcZA2wY5eDRbVftn63a
QzPo1OSJB0f/WKOrTgzTj1Ff0lBkra8jwmbM+V3RjDToV7V5qiwvaKOqzFxN4u/K+Oz6NnkOg3ai
mLvhU2Re643/jiz8CQjkEt+HypbBaUvpQPYireU1yF+KserbKD5cvYjGRZrG71xblTbFD36rU4nN
8ORaYc4se6M1G0aYQ1fcPtEQyrClOW9HaHe2oDiXYXNTtKWt/nPsPdNLo3Efh9H8fVxGdgo3OVzq
URCZN7RQnVOXTEiFX+W+jbBMnvO2rXVTe7ydhWk6iU4cRpkcG9kFkfE6wT5ih5Lp7tRWgWB3Bzer
nNyY7f3WU/vd9A/3bKBFEWmv2LKNAU2ouR+WEkPp2WX7zBtvSo+4PgIrqu+nkrmXPFq2/dJnyeE6
cUBhPpinAJRrXu7aOpm5oQw5w2wqRS9Fo3fqowaZIOZqs1r8vqrt0P3rTgppN7rX4XrPsaUcjPuX
jj1OWBuE/nSca9L9rWAl984ivb3zs+my4FwoWJMWtMA9AT1zHi8d8MZp4g244SL/1U8rmHAO/Qgj
XlPOfv1MxQcxjuS7EkBQjARx0bsUhdvh8wgWimkiJZKrWwu+ngcSr+QTS8r1JTovDRsi5mzk/Kem
UDvQ/kX+mjqr5Be1EUmCtcqSQT/2ZAP73j67pjR7J9704UnQb30sEBFX0w9QG0RWnXNGZHryb6v5
+n4VvlIkR++nsZUFVE9tkO25zttrFSQzdy1O78w3aLdOU78LbJH2QG0qukBF4n/9EddKUUeAiWFq
/Aro8B8/albRhTsv1f3HpkZon8Nukk5SNbW0WNHnNZsH7tzz3Awk4ggRIIFR9VRqs5Lz14zDcGMZ
Uvw5oTLlwRFyiCXxh90PKFhD5VJ/u/E/F6WuxdpNVDCizaa2GcaZIIvbiW2fteWwC7JIojLRC6Na
nf/PcSWgiuKwLDBUKuiCu9isLPR3VDsf5eZEPQZ3gOBGbLZvUGncL3RWWyl3I/YmR2HEL/W6bs9O
6QvokxOxRerLL8u30srB/fzUB4rasPrEJKk2nl4LOAQU1+mjzyxfVZT3qznQHAy8k3kXVw6fJbrA
7W3qlrqjdsffIpVlBQBpjjx3aR/O8S94Ef0xnalzrU3+hxRZfnUOqm9/jQn32oRzehhKOuH9unUH
LC+kcztZ32MV4+ocA3qDYjMhBbaCarqTiDspYEdIJ1mCjrHD0Nwg1mDfRJeCjgu4jTFw0o/YBb9c
zGYUgpjQpMFW72egNzl+U4u2tlBr3pstclvhRYNCvDih+AoM1rtCnhU/hypBYZNnfEV5iI9Dn0mJ
Gd5EASUQduJBzZvn89eDW0cs5MV/sXcezR/I4frY5oDVLpapsKN4uGQkcd+MyPpDmzL2IR5ljvVd
kKycy26VcuedJil61XNz1V+h9yc2c9aAKx+vbj3t047Kyi9mO8MxJGS/sdaovgPAGz4mquON0Srj
AXgRgv09XVvS0OBJqWdCpvIdxZZtfDyVnlNy3eWLYAGdUFP1FyoKGHjsSQFR0vPvjqkFjgLSzGTv
b91vUMT+Q2A29EhyEZjZYE+Za9O1vwSxGSIkpb0Wt762Ie/JAmCvdrKJl2I7iomNjUpHJLM6T7Ur
w++UxGuKk7ywPw0ivRJh/hnPRH5IfgiviFLMDoUMhVvujMnqV1UZu4zG2DoVn5ynw3UOc7qp5Ym+
9UdnHoiJx62+dmpv0NAzHV+Y24cEw6wulP9mz4+xTd/QqHKbwJ5BcPne0Oyg1H+OK1dsZsYt/HEl
O5smasvwh/RxLVLHEi7i5uzJnsFzWDDJR7TTgHlbr0AQBXuRjAjnUgL+RoNWc0aMLSuHB4jv5cD/
DbR/boTGa89AtIN+dyLuotEMJxvu3n9PCBI/vmAN3ni0gEW5hx9MP4CLvhlwBVW2ePCLBbiMPIcc
PyDAP3fvyZvSdpWqycC2Mx6QUMk4sXb2ZZnvkh+HemR55v5j2iGX32lr7/vqbK89ctGJrdjowV/a
i42GRZwpF2q+unpW4jGvtcsHfMy4wIFnoUXY250QIN7MLBA+qdiPeHvmpH5FKfLhNs956DQkIV62
XbsvcMRb8Pt7/60OR+HU65CaDa95eyC25PPV23hpZdbr2nQ+5Fdan+qzIphlTa6llvbYZRkmu2Xl
v5wkKxkbDWli8ip/lCD5VNuxyxJoBsWXjOQol3omr5d00fuBA/dGQZyB+coiF9ck4OUHLN3P4mI2
E/mWIKd0BEqyTZiA6LJ+OQ7QJCXvaGFLUVVplsx90vU2DPbd/FptoxjM2UK77fA4tvdAFVE++8hK
pMZWUXccogSY3nVlOgL1u/LUNOeCXIDxg3sBn8iEv+ZP9MgImBRnxvkZv3wIR8wGmZH9NtQjsSw2
irpCsQoe5lRUqHklnEIDyMV1z7k0Zb0+u+FpIQdkbNH+H9ymM5y6s7IWq4v/vGuRWt4p1JEl089V
tuGa+SM6w82sV8wpZtnfl0F9Pf6K0DyE8bAWrxcSpXvLvr/6kjrRzTmQg31f9kuGQpOYLQpH6sKP
Kg0f4R/C/CZTPE4KHCV/GcE5LAW/tjDTo1v7ZVtLZwJt1PC89Sb/UCBngWtrgvE9HtjJD2VKA258
Nao3D8xLo10Xwzs/28HCSRSt8m5pmNa4UQjr9DXBtll6NIJ299pBMP5kjFwJIwYpxPHSAHLEHEEY
WBufGVL4GbNSvShn4ChOxL4Qs4DjSxt87Kw9dWLx+7IRYZpKd0KN+b2Fr+u/iNgnrK4je2etsOq8
Z0E6e74TbI47pwMShVUtaQlmWs07U7JO9mFDYFJGvbmDv3ietxzgMZv5Ct9/GgQXv4YxBTreDijW
VHYnYkAOaIIYMnpy8OcfE8TGeDiPq2cm1VFB6PoOgfdzoeQgZreH9OZS8TGwDuftAWGpw01DsA7d
t5Rwr3/5DbsxnOBBKYX8cE9NiXLaRSOmuR/YdDMki/+or6k+t6Mkg2Wk2lKxSXa7NDrWoQRnEtL/
5s0euQ8BuCskHj3SljL6nWFixn7bQOwrDaYTpXQ51t/cKXG8KfzTzlNYu8LlxCV3rP3TdruRExo3
ExiUCmnXFZlQiYTraIY3E0h1HJMHUlwQE4n9053PrfTC6OIaQj15CLY/DtRKnlQbtsfYAQZ9fhk6
HFcHq32QNYV9vJl7U65MuWpM+6eDU3/pRhzxr0mqK9igFl2RIO7PwUnW+PwjgWUcpc9VlZni1/Ly
vrMDOrHIANbcnoOsyldAK9F58RMtMRMM8iXcQqq5k/S1RN5TURfSKKHbMFPuOR98zwjR4y0Lz28q
Y+SltCWADmVnEs6+9ad7whVDjV2VB41o2wfEMCfZc+Tw5GAOqPMTywR3pYuubf144VwWZ4LixaEn
AFQg5GAYmYyJkMDRr8JD0lI7YweqW3v4IgHAOXKJaeLbeii0cKMGDz+Lykz2WJ3hjaUYNtEDLiFY
7t46LfsBH/bITTFcIX6mSAt25VsH8fJYisMVv7zzpRObvpSaM9LRBG2po4WmcJUdjZCESRKArX0x
k5UTBGt7kQ9V2cXeETFCB95g/uHOHfihWNyfKgHe41sSs0FQFfVn6eRiCkVMoVLST9XB/jOXamkC
1F5R9hN2IPRWwZPUjEYU1y56cQEuFRSZWZmQdAFTtHvxYYVZReYg454dqJaDja1k38sLTDe/G0Q8
Xd/+LcW+COP2ffh4MvDyfrZe++DkDxw1ONrr1455Al9outGv18P/ABXJwRjnE6/XSJZDJwy+iTdQ
X7h5Afl+eueiqMfaIWJOKjfMigrIcID5buzVbfsNbppbl7wRTgf/jZB5U51Oi/ObEU8DIELOhCdp
bOJV1PprkpySpPBWpDRFm+BeM0A9c4E1RCLPZCH50iGL6in6Z17exUp3Fqlea/oYOvDm3zBGTJ58
FPKnJcPK8WJLeZw4eQ6e17H+UX1Mp0BdHXgN6U7fpu2/Qzx973kKMuDklT7bXS6o9h/y5M3nMW3/
GQsepSxYqG1XbSRkRywteV/0+UfL5b+C21eVhHC2u8WtpOKRLkNGE+ju23A4wuU4OOMPw5zbbssR
69/amBWpNMhvHGPs92iPQFuIcmKd0LzDOyl7CJ1/4XLYzjuHMUxmW034JPYKmn92W1ZgmiNmjsJm
IHPW9gLgO+tel1OixPmHGDy3F6j6Ai5eg2JU1P0OCGz0ahTkmQbqhCPprHfv323D/3pSyZ9I9WhM
9Uk04ACJheilihg0yroSvGayyl+PNoZ6QYvRK5EZshBA1QSiD+kN4PK0bQ1Aa73xbh8CIwwOJSXA
+/aE/+5dFpdslPbWufUouCGrQnNTsQjURoZ0qKMLauMDzFyPD9C2tupMeUSt1AAZkmRTjsXVQX3N
LBU0riXdKH6FE+1OCCscxx3wwj07IpfkfNsgIzyB3Hw+yZiRidtv1qQMPIyDZtxizuMJqrdfGj+4
0Yt7suIZbSPXnYX2683T9jpQjE2NDu1T7WECszP1Q+O1K5N1sZQYj3dT9cHKSSEVePN4Da7GwHj5
FWrdpFtvKxaGY0lYPpZw5tRYyPXLztcadrKlPJ0N78UPoBN5WOYSPq5WtPT99ke1OgcisgOL/dsX
djKqFZYHLFzwaibTbUB7WJxc16hQd6SuWeM/Pqw5KrX7YcEERvk7ioxxWmE8OF91yVevIWxHm/J6
ogwggGAztsQn/0AWjWWpbVNHydCksnSFhhtuqYtOfo2hMzRCBYI+5HAsxJ2c+jPRHF0TkwL87vEs
4iIHOm+IijyldxU8DINkAiuMSHFZRbwUgdqGFdXegHD4c9Nts7dMkTmE6pOPMRGlV20XLkBQTV6K
HmlCm/Ot5VfnpkFn0RPSB2vkN2KxQRoYSWa9b2RnSaQNCZxw76mogD3EtYRj7SMkknLSG7Gt+chU
pbKslUpoiFLHhdWtTxCJsHvw/e+rwrwqL+7rrx3JeuJMXf3KwdaPL8nEfRmPqfI4kfuW/Y0m28kI
QSkSlxqM//wgCTw0SnsvUneEh88dvIOMOsAo5HKpnrZgRzT3IBUw8oYuLhTMmHC3jtStuWIMplxJ
e3Q8WPGT4dw8Iv9H4iagaWwm74IEKba/jk9va/8srxALy0eqbXksVhqNBowM6WZu9FNt7ZXcjk7J
9CVU0e9Kjo/AT9gqRcxw6X7PqcMNUb1gdgSGRaP3lA4gVwRrQcHNNUDqft+7yznK7DaR0jeUkJEx
rQWqOLW+4U8H332LAj6jzkdf+nS+lvUbYTxxKCqB4A32U8a5M5s8IQviFzoriy8kpR99A+T36o8V
TCbge/ZG+kEiX1swmTBFEUPKwJ+Q+dLc5JigoLSfSLD21YrBpaH1Ql6zMhs77DNIq95x31fIZPWK
AH8S3HrPuCDkeXOEj+viqKIZSBGOV1UrSpn0bCbctD47yUauUKbzlf4g+ONEGI350vVhTGYZ+FS8
18VsqWo3s+q6wwy56tpdcyERO4rHORdSl2hkmXjp3yemWYvXybqLjhJprIUrOEX6FHJ18f8eu0CA
MiChVdX3q0m8dPU4Jx5STpExtYfSRXPBAer6yqY/jjdwAFOgMjt/I9X6Q0XVI+Q2roZWET1G2olt
ezUtGGvFC3DxZmQqftIANB+wae58wz4KJkTj+0mTN8GaQ2q7iUtThNLljNAt8YhSf3S1iOY2AdpC
UWUS7E2KE+zSHzoP9JMc2RjGs12MgPbenkCBPXSxYRpXTQc3iH1xdsvYfoNaypCMwfAv/CZUA1qU
3btwLXEVrbwIZVwdzRMFO+9C/jyFjpOsQdGtPhix1Tw2XjL3dToF+CTuiwVrHVaFpGZgBbKYDWfT
4cUzbRMyUhd1TN0PqBHfSSy0r/aTeWeoDiuYrzM9cSYy0H6r8BRhKEwpNFI1aD/HBWLfOE+wsIlj
RR/HlVh0HHKeDP5WCThfdS5ck3bEx937f3b7yFydICZmi2x8qoXHPv/z63PPtArhbMfaNlyV0TPc
7piXGgziG1TN4652UWeNMDdjlMbHWUJ6ARVgyZvKEipzkMk9PbKh6uFFBItzG+24eEl8jEP5BhCM
zpilkDsF27v9nPQ8Ep+MzwmwJrbjm4dBYfhtmyqaLhrF5JyNe5fJWgTUCp+QXoR/cOtVUlx4xBNm
NVE8Ooldr18fNri1KY6ac91dG7KHf4B07pZCXiriXmbPGBPHbKboTcZd0N7QiYxspy8hoeZApql6
22EQIU5CX90aTRUhxF7W6F/zJ8qAOmK4lMgxg37ow4WeHowqzTR2tjlzqGIsFTX3uLm9abLa8P7b
w6IODof7F2jvLVwqr7x53benlo9uptSdoVq1rn1NCoZRTh2Grhkhts40DsGJz+PMs8e4Sr3eherD
26hFsp6oG5Bfg/YAOHi5gybXQJqT0kWJCgkCcemFYSWIJBwz/N5+tTk8yQJZ8hxWc+VW8rgWlKXC
e3u+jREQpPhn/QWEA4D3LD0xJrDlT6mr1F+QBvbvT7STApU9TfYMgnr0tj/uM7cvdKf1N+aEv/ya
E6xnNb1tgBDiMHydtiCRmLaLYYUDxf4UQkNsUo06L60EAjXDQKsJBLcy4QptKpzDR3xM6sH5G6na
BNJ2WQ1vMgPTTvo6qf26hR+5nsvgilsFjEfyPLcgxo4R6BRxKWcmyMFzpreT1uqruC0kFeonwsHS
yA1R6UEeJT+Mr/l0dtGS1wx1X80xYLXkEE/GqOPxxoNGt9EJq0HgmeXBrHKNV2qRxvmI6oqTV/1b
zeMcIWp4JPasr4MJlS3Ih9pfnW4QKrDyVtGyHsCItysCTNEumsbJZZx8ARE34bEdpJnlMOd2G6mA
tZ9mHegwboFD3aExpNKy3UabH3eEhjwqI/yU93OeJbDxb/w+c5R3QJ7z7T4JehE3eaLMiaUiW5Mu
quNq3G3d0ekIDSNilyU4HafrhTkYoI4vA0oAoQCLUQsb681u+OWFTVZBwEEAMY2jxHoidBEjZPyU
TcxQ5YtV1a7Ch5NHK0IGVqPVKoUc2+AKLVRlS5pErKYeIuzJbRwyAda8kIwFcgwaZd3K2kWXhFgs
fGyW0d3uQUJ0wTLqDb0o844bs4Rj50LrMMVy3RqXF1KTzVQXx6Pk5J6p63L3I69pSjGhdvMKFLcE
X1tGERfhL/TMW8lgj/y36t5rRM5YS06uhnHrqpg/qhJ6ZDMaD0aVWfo/xvEfsQTDi7hy096LE47F
CGe4VPLj0x4MfKvBuNf8ZVsdYVLfdvUFvmUEx10vt405ytkQDI52G0bHWt1Xvepem6OOoQZp0YJ+
LkAIxZH6eLjzfInQDRvCvEnZ98qW4goQvc6tkUnyVZyoh5eeOsOJZ8LAcOFUBfc6J+eRnLJuXWoW
Qfkwj7A0iBkc0C8aVyjNennT9CrMdKSKgtoXaLyfmkxXtu5OkciZPjJviMVPn1tYr1Fxjhne0o7Q
2Y5OKYtoDrXKSDYcFWktP03EaRCFrKgz0nqApeuH0lUXPZsg5VkDb5kLxX05IvgnxgTM5PliS6TG
fWuYlOEvUhdR65bvByiqRIKF+mgTuIJFh41M20dz0oVgxvqZACZCgG81DPHThqZZnsHC8j4d0FvV
0PTgdVSX0JoMlT9MS/qYAz7BuQBjFdebXNw+gDH/Sj7RWBoCYYGkP4/x48o6RxTYoZ05QTMzyBZH
N2/CvmKZ8VpgGuLjDBRjLEd0j0KOQAdokFxiS119fUEZbnIOzOM/EUxUrnDWsq9i3sXzmIZwMuDM
S4DkVqZMgh2qsjN2p+HsCJQbPi7bfJwT0D8UTvhUoSRJRl0TEgrfLkQ0WG/ymWwTBvc79dSqHkXt
xGWhar1abIeWSwXLuBjncDTHd7+B6647gZTXqdIl3COxfq5FS8SlNVbw7YDM1czey6cEjfzsqFXr
COdheCQGJ8qyP3UtCsR/RIN6FCqpzTcWmEHMs0GHsXioqbnSeF06OKymG5CpkuEWhIPDe1KDH/YM
dM/mB7uNJ9ScUiidvhpPSW4liYBLIwK3g9eUOqV8yazYzjQm39vEcIGR6JolHwtFVvT3iVDtif8Z
bK0E7+vNYWm7QAhKKUusAZs8Jr3W9WvJbVOb9h+73nSP4W7xnlgknZSYU8BGV3ayHCUTMCPOTzZl
e7oRfBQoFBSUHXG26Y7Kw/hI9pp90MmAuApP2psvjhI2iKC4l356nIWIk5jrrKAV0FgA7JQN4Qbt
amJC6EGg1ieBf/wJcRzkum8L+RajTcf/qNpn9mSTPZAds7MtdYCVoziFJCpS7zLAXB0scknlcxzL
fCY/F0QY8WA/ucuILx8e2nLft/kNoHIF+BIsN2w3xpHLnsQ9gTSz1345g420vOGCw4l4oVpCieCZ
4MB8x2yt618kMt+SwayOS7OImRl21UJjGtFT/Rv5EbFVPsr+Np7/Qr/D8eNOW6saf3PrzhpcP5OJ
7MbP5CLo3kuNgGfV7WFJQyxYX2hRKkwIHONdmeqXNQ7lrJxGZ2fT8PYSvWkMhHKjvMJDM5XiuI9Y
Pe9MnhYWbgxDjqpNc861ibYlfxNbbRINv/DkOEEbwf9ijUcx0TW6t80Vaqa6PSPlJXy2qaJjnF14
9qRX751sme0qeKIC0U9+ZLSZYEiwsRNd1YAspu40+UW3aNMcQLZDDmgAb63RMPUtbLXKFgpCV6Hv
ycAR2m+hIr/eUoN3i5PU4jclpBBIpYTptsO1d9RttG4WvQSKIGTKY9F/TmWc5iAu709YfoNB0XbU
fR7jKhRLeghdNQIxEVeV088WU1KGTX7h+eNhPVSgYlBgdP7Wsy5Bn2od5QAK7bDSilR4LggDUsOJ
0J8RDVNSowO5OW+4gmT6F3Apcj/gVL33ePEWIQVptEVMIwaLD2xvSgkRIMK4+zgJVW/Ocg3NcnNM
/OSrRj9YMV3p0fqcn1OgWH0VDvL3CDiCPerxq2mAw/HY6ai7biFkpFhpMB0Ugqlb5Hoo4l++sxt9
d/dNGm/zrAnLNUPwyLf+xq/MFYO8mewQIT7sEsF/j392Enr+07QxfRawo4pyA/k+jf818diGylVK
mz6LfqCuJSOe0oLb3vOP8eyYRRx4Wr6L1G/pnLkeNqh4gImiqvd/ayIKARykfrALgpSAXpXkgexK
b/qrGN3SNeWqA2zgObXox3AToVpwuVcmBskhZsVl/+R6PE/q0LkramsqgLALV4H2Ww/BZwsekHG0
ioREkNgz9L+sV9VaxqdAjeBoM2GJ33NaKi9xXxQ8DSkrIGtVnxRaqda6FFbJzwCHzYDgwE0cyOQr
YhnXfgORaHUKQpIaB++rKBido3UKoz1CJ0GXN6w7IXIpJzlTU8BgUVHvnTcXJsQDo/tO3BSFbIXn
9NmKF6yaBhjrGILult/kpx2NzOJRdwPRs7kW22R+uFv5ERwAcf9iCR1C2htBx2iCFq7Fv+WzAD7s
hCvfNL4hyIBTyOpEhHq83Vjv87XEVm3YJ6Ipryhm+5578wA+5hjHT+/vh/zMF/ym5kSmj5o9WBj6
KyBxrCECX0SAHkEg3lCVTxBezIH8mjED1zbRfXAW6X2KL6qhspjwKWEmD4TH0lZCGirnmT3zUu3O
RQETxyGQs9h+Q/3y61jJG22xb3smxkS38yRB/zAirwa3FeIxK1Hu4SMEGI+Tmvuc8I00S9Dlr8m6
3L0Ert8ovn8pCnKL+tA2o/grLy33OLtOcFCjs+zD1dtFQitimIC0IBqzjrVVwyhHRQLUTF+1waRl
b1L+LJsF2ZYelMCq11JYxryhtmqHfp5o0LJii0poBk2ehZ5G+Y1nG0jxSeiTXTkaWUPy1gsL1jNz
2z+JKQWKcmGVcE7bJLsRACevuGyvj5mZw1cUNyuIJBoYe1YAZU/F1CnjqwaA9kx7KC7FOS1EAAjB
apuXTJxiuyOjG0Sr4mEM+0b7BG9dsHpZlLQKQ59elDZ7DMhR68Je8P7BEmmQszfmxTOr9eOWH8pt
rs1H2tszUWJtCdonQ1LOCUWEwjq83BL8QgcwHrbAwCtoD17yp352T1yT1dz8SkpAxfDRvymOk65Z
T6uPDmmF8kcFUp5PG4yZNUhEMwD30ewo+KjP1Xodd/ugb7rsthrjauumHgQKjnxbSuFrYQOin9B2
TIgTN8dCBJegwhMeRC+KR7jSJGSR9KXEPDXar/wp5NUGCjpEGXVpu19N01qwMfvuvqXcC8+IMs/p
i3PqKRPgV/0jfdcYucdPisNvD+9F820gci6uHaCx+NIp7DDiQEj86XCTH3uHB5nvIphs6oosg2WV
008KAQ+7J5vM7PGshWDFMTYV2YtGAUM1dpIU7zeuP+/rOQFXCvhBGONemHG2Oks9Q2TYf0k/5Ohl
AC3FX0lpnUrQ//xBxFCxf5vKVab6Kt3S72vXmSIKae8rt4zwUXsR//+HzGRXX/wXFBDxewNpc7WS
mi20Xxitbu4OKit+v9b+vihzbxYHtlTzOrWwjo9lYu+NxL/A+80YKC0g4BmRX8TEiHTeveFfkesU
LRbNMKJHDypOSSASsXWxf9L5lawmC/Erwu7XCm3ZT9Bs5r9bOAgOkWHbePKzLf/GH5qfmCxK48yZ
aEV1evLKnYp7NZGjSpqYr2oRFeWEzSthqXGPDXTJN/WTmbfHnrFtPdet0Wtj/rrM3dGb4ui+w2N3
HzEpHZrhcwPN5IibL/SMt/f//lvX4r/CsGA00cRyGcScqDNy17LIaP65m1zzEkOLwXFeHVIRaU0c
n4ccs8LmbnHhOiLHwG30HkgluNMxZ5k1/IY0wvp3rXkucvJAeoFxf3mLqELGpco/akps9HI8WT2Z
r8KPmCoCyXpHG34dvl0wmRPVbl9b0oP4GKcvh0Fn/bowXCA776hd1Trrn0PHanOkp9OKjZAsOmDG
mJXRsfcLj21zOlp0ggDtH0eKfpdyd4BoP63YsOeNauqxlIIxXLnRfcyka0EgZTh5WuPZsdaoDgXR
khq7dWen+ccG/mLgOjRZZ6pKs0P1/LaXJFK3KUKpekNPHkYxmSUBk33AVV/sB9kP7qDj4VFrrd+U
p6vIlsZqZX/pOo/zgfPOxF7GoGy7REWp757KhpkHDpVB98O+SZHPsHMYIqnaF7HZ2e1R7+2sYDa5
b1tNDc3ZpjPIdwzaEXwSGq9bVAFVuSa1IosXxia3V4KDceGca2SJOz6G8sdH/wWbNJaselwR0b4O
9pEBkrrsAjvnrrAxnP6yyxMg6M+BXi6GMybCh/jKe1z39B8kCUg++5zaVsoS6q0w1kMZMH55kIlI
dmNOK9ZnMae1c073oF2TtdRxl186RTB5tvW3ovhpz2ONx64Ni0cz+50h0Kkdt2mXw+3QnZZmR4tE
aeFYLUAVOHQqcinL0vWg16lmpK1JGnfwxfIE43lLvUPElDeAdhaeqs9rCoJSUkSagFsYKPoERKtJ
BNr4afZ5tFxo/CQWaAW+KdF0/hnSJl/i9K7rUMr2d718zFJItP6BjujjVbKGcQSrnA38nxip6Zvb
xMj/053IK2RfLHg8jC9vutht8Eu1e1PkxFZAC15LJuJA2FAfJZWee7l8PCWthUyswmt1niAbNyWs
qVyvaMv9rorGBQgn5VWV9340wcKQcBpeWzzKrpgS5kHGp+lT8RHRtQ6WoNV+Flq8RuQsTfyWDvE/
grk/r2cq35LDoDd+TBJVz2EKbnzJxMZ/jW4WJYJVshAet2ouG4TWasuo12IM9qMr5oJGyn6SsZJB
4Rp3glcBoRXqIksQ2qrGkQ3xyKgWJyYtDeNzKaZTFpbTqvJjb+qI9HiNorfj3sffZL7nvkkuaLnS
oOWqZfqjh7wfZWV+BBKz4lNe7XOHn3g5EEnatp01YTJTE30aF7v9LqSehXJZbGeVhYWyvwQRcnxN
1Z70DEMTaIbqLQ9GKjPUu4QoGM11FpSfFB7jnDElRkMVvaSH1Nsa0Apz0B3VFwBnBvTVH7absgsH
Ks9jpfXLl9mXxd2x8SE12StuGO82DhjEUR3egNKpkc4G0oziAoJaedcKFwtpuewkNhUflNvF7S2U
GrxTbBT11PU8C6Dfw6kDWC5uBSe02429V86amah9P44S+aHiMmETXhVTCGLW9Lv0VvvVk8j7q7I4
W2VE4pR0FwLExvr3600ValILW7AkoAV04lWkOO680S7MiUFLhksQ1r8MY+0XZGHu1FEFACazCt7t
0h/tFh+kgAIxvQqHWM7AAWZ7X7d4qthxJE0FzaAobFR0opM7fjGTn3mYJ/jub2afSeVd8YqwzauK
r5wuoh1qEMAt+KP6ApzFM08vZHw2alsWYkRHmgKDhksIHtl947mplGCfRep/Lh1k27MNgD8lTxbg
wqPiwfj98mBN0Ui0q0jGAtEAKKfnV5F9j4E2G2O/DM3ld1ib5nWkN1+4tEV/wMfzR3/g3QxG8WM0
ZvQEm1yE6bjQU4seyGhxJ9pPi2JY+7rmjCbXSb83Pm8hiOMkSrfyHdVmjEQIq+/RxccSaCfP8JIQ
gCD7SqP4Vb8nODyW0iBzVIn4L7M7NR62yMCbg1JIkZnPHAVQa0jEsNb/U2Jvol4h/dU6l6TnfBdh
z50yN6S3kigC9+ObwIp/UZpqWDe5vJS8MkTyzvZiNban64WYtLGZot5bCZ0k2a//Q1wm2UDySDXH
Wsl83NAZq1honofT5Q9hUTc41rg8mpfkt+NwGefg376/PLpMkmNCJLRO0YwSQQMP4xau3vK4P+l1
hVjCeU1Db/JzhoCpMOPGLzxLCDZaEpMmN5IpukzaoHB3HZcay6cLwVuihF0YbcNevI8ULTi6S120
M2ZQub+klWyKngbW5mjI3B1FTDi3BokMlTNT26xTG7oFNj/fkSJFxgEOcKfdxffkrY8kAk01xwGy
2jsVWFyMtM18/T1OJwFa7y1NbEbYPi8ruBI0/y659JUebZqgdCDeWJsn9mTRFpLYxER4Ts/sKaU2
wnpgKbqv5k4s0e60xCvqgA59v4obG/y5We34J7nsD8LOfCPban1OfSaQqiS0J4VaeurtU/eFDkOq
/YJsq1vrFboDTBPM7W6yf29CI+Dj1QX+vRm902fYpnIawu9INqME/IXNqPhLoDFDVRgPmAjD+OQf
YpKt3m1mGE+B/PuDqqOgP5zmP6c18SlBxE3DlT8nbgGBdECZdERFhaOOaIivWeT+mqX/qj3HVa1o
PZqNLl90IkORwU4V5WPcq8nhUhPSFvvaC9rRlzTSyjL+LUoweQIwmticEm72iV6xj774SowdA1Qj
n+uJ1M4K4uVrSM1DXrOlpYxHZdygyItMUn+RsOvQNxj8BIiENqk1KapvgAKCPihwKREhMlkGd1wX
t6H3Rw24XQPGYy7PjTDRJuszHJ7P4EAiIsOxLAMFImegFntvT9kMgFiQLxKgcQ7WIJfWzBzjkIij
93dxOaReruQxwbcVLXh9W+n9IUD7b+hGA4Ill9fuX4FPFjXSwLqsZPwFD+HanHmqTs3rhg3mx5GJ
xpKalKwruejNU43yhHiMUWJ6XfdulGh97zUCs8cEseOEQ9+42MVBtfHeHJcEIG+WPyqjYN7SXAth
TxX8hvZBh66c27IfqI+7T5PSkRjsdwwp1qhsfeU5SPvIkFoSNYK4vfvMPAUQjEEHTkIrD6533Cy1
hzAqADZT8k1n+7Pb0W5TPXJDwx4sFVomkagbMUbKLpHNhVcTRaFJbN0bzV+rLs/vy8Zhd8ua3ASz
nohA3F/JSwVZxpoXgnyzdzUT+JEiPNSsoE78eHBdW7xjcuM1UUJhdYDlynW7qXKb5UbWewaOQTAm
unW/dShof1OfqN1l2BEuILwfqnKdsa8o8Foq80mYiq7IyhP6E022z9J21NHHZ3XjW8JNn0iNWAHc
llZ8GlN2KPZz1u4zu0Kd9iZRYaYArZZJH32d0goqW9rm+kEK8PovW/5hdtQVNsRh2GQkCcBpavSV
RVGS7pKh/vDlItw6VhNuzsApcfj02BSYGAWj8HxRwGm4nt6iSYt0gzfNkvQWFT9vdKjCmriR1jg0
ppqk+9voAYg/0TokVBp9rAuOF3HXBgs1baUQ4XhGa8SfhPiZIaj7UbCQgh/dv/kvv0w7FpCVC7kG
gXmYnbjyWL+3ZJrRHrx2+dkwvJ6SoaAtHAkNR4jjU443QMS3XDRXoYRLrGICXU2wn80TOEkHjA3K
voJ8JHPQ2ZOLGfytAGXc5v0Bfl4LNXrqNHA08uAYuC8iUVirosOuJZ0b6E4Esc1Esv+ZHBfXkzVz
TpZ/tLe7fe3IoJ3jEE4KY0RSuHU0qGaM9fuQBM53BhJPoxr8LMggpvQUwY2SKN2lQjHQD5B9Xmf6
r2CdUGs4D3lOAiIKjghz2HiEPKdng4yngVyf+8oQknrMpYgudgIhrmjLDtB0fysn1nUfihu1d/ie
arJkm14fkltbg41uRdBhlQB+RugnAM0C6acjCeeUSyuymqpILUjMA4iZe4/XDm0W03Bdm3jrprDX
hLkHTjjOwxQHuz4kN2RuYxD5c01pQoPQ7E4Y/Z1S2CMVoAAHIc9MwS++P11TtwM2/hZIJ0jE4Fks
2oQvJQsffjD8Izq4+XnTQ3qBC2hH5p4d+S6vcyN2w7sfJJV6etAaVll7rkHAoD4m2IHa1JCeyCBG
JZuvxgQfGzMAkoglqFsqSW98rQBXD4t1OXeX2aRpkBuw9QarjoY8LpINWGivZb/8Z9vbIlSonVE4
hg6GJkDUdd56idEUHO0rgpVDr6fgfrz6tojwmuqKpQ1brRwMCtYT/Bhh31Jya9Rx076FOtPmSR+q
lSYDZ0ml9Z56AOgr1b1FEGOxlJ/LFYydjq1IFWjgFV4mWqfSr6k02o2khgpaRhGUi4zz5JHAXNuA
pvTQ4yqzcPYLyOlC9OAk8HybwfMmFT7o6nP14sDrXhJbnda5ZRLuzpx+sAQpoMaxrPBpuoP4yzZk
vuHGi8E7ouTXCLronBjy45rtpSVBLjxTEcNMmCgu2laAG/LYmae7dd+PX0zA+9Tt8LusuBoVCi4X
hwtDznwMiNEIDvySSWYwIPUPWeVxZi6v8k9wt55s2DA/RaYaBi5TB8avTgzZhaH+vZD0L9CHLpUK
+mz2KA4Er7U2yb1sZ2shfimdfXf1q2Pd7LNV2exrwTkQovXBZEbDFgiWaI281fHM7RaxDkJ6pxpv
GimLO25pxZMjsZxT8heK/q2NbslSe6s3ZdDxR+pdEBDvns4BMwOgDbGg8HinWQrWxFmgtUSvvCvo
oU0lEc/xMBqE0mmLRKRQ8mMzWD2XE0JD7r5ET/CUs9OuzpLtaexAHL7/JJrfSOHx9Xzu8gQ7hQda
kqlBU1XLOrXQzTkRl9fUGE3jw15vuL0602PoZPgwDmOYnb1LDrnxQL9k0fzV/U69oXzJ0F0dRUf1
tP9+KLVQqYv3iBJRDbTWE63AO6FJZwMZB03Cij0TffvyCRk1GFHItKoyLO3ba41Q42UFYzHTNhCx
q7rMEfoTI1vrSpb/ecbWR1uoqNb9sQZ+Q7v7J0hLVlbrAa7iGvukFRgJVYzU2V9szkogzDFJna8i
q6OfLTjpAurv0SJQoHCrLAzgTuGfBi09AUbNaOAjFO7dGsSFOe4NKWyEEbgli8baMQJa1tdoYvjB
ojaJc/nSTpwQXkVYDZrchg1Fosi4gVapelR000Sdh/aT9ltTt0+UOBq912K2umeU1xaoG2pTSdK4
tUiUwyInKNyeD1DkvKKfMoHoxQijanTrSWDNOywl0my4ARf9YM9Hf7M8sKUsj9TV8sW69hrrlS2Q
ybUXJ+C2/LZAzFxrNEx15lr4ElRp7o4IAQceUUAKP/2G2cIdQRcRVQ0v6GR84UL3+0LSErqexOaV
UyDWKn3NrYlHWcKRC9sTdqAS12fkJY35wdfawRcjXOtYj4a3HKNtXdPYE2X3zN1UJYz298oYbqWZ
/VM3oDF9CIQiH81z0KtsnVSsKMlqUPRJBFp7rjevr4to8BoSO4AikREDFGH+vviuPiYXf9If5an2
DOua/HIlSHRzwEla6EV30e6ROIcieRXjkmfH98dFvqF5mG/j5vrsyJcb3XHCHHFQm1JxBElOXxj/
aS+VbiAXWxzY1MlwlbKAi6zFkQAdMKxlRL1SLl/rYVwR0IXLf2TZwjCKo+SAClmBd3RlkU8VEt6q
DvO0ohM9JxwsRCzLczf+GcdHz+u9ygzszYJZ0tGH9YAsYes0bac7gumkHMA4L/hoSikcE63NvQyz
d9pxzs+rbgxgDGyaT7FIcFM1FPAm29izjWhvBrcVrVDyWYaQRUgaRpu6xOZEw96Cn7ZlaHyGFSgk
QwNvI7H3IeZHhd3vPFg03jnW4sbEQ18sONMdMr/H1dXNt62vRvkjBdKVXWvU0uMjbIKbBLgzIGc8
VacZeiH5LOIqIkUchz/pJea0NqMEthCFWrfIn0VklY5MZu276qmnwzKzfd97nL8lyE/fOq7qtaZ4
V0L9V1c0zK1BLhtO8P4riPt8c0RfOLXJF0FjNwuppTjW2drJN0vjry98NvtkQd6CMmMlvGtP/7XZ
oRuMJrl+SHAiQPSXJMuvCXoNWKkU0DEhvkd+B7ikolZhOsJXgZ3dTf+HklJSkReSCcDHXL4zS3/z
BcyMTa6KltG75ms2SoS4oZEjB9WJ9gb70xs/gNl7C0imarnOCZSYINyiDz9AGZrNsJ+iQlNg4qz5
DXbWgKTXCd9SMe5teUXBZ16cFzHB62b0YmUJxqHRO5A6AKnTT85GX8yWmLYUIDDmgYIG8mnJ7X3W
MvAq4LaKKNOgx2WJ5hPOUnnvaHOOb7ac0MPP4G/r9mnN9yv5GfAGTYcWQ+ciTjVvtiXmmwrooadJ
D9ItvauuKHAiXyIpCpW5Laq2nTWUreuzugaYm4qcLJYQqfHGlPTsm3mC1q5s8vwHN7S1W4t2rweo
mvlCKaj3CKjpW3EWvboObZEZz1PpgeAowJGBnPAMqK3CbsdOVztr3IhJ9AAZy3OeDcPy9TQsp2Th
4FFt7y61iyg3OcJMiPEzyQyOdYa1b5A87ubG9Rf8fVQzP2Ee/nUlWCpTfTVP49mjlZVe3b4gl66V
X9xzGDQ8XR/AQflRsaxZfxdmmGoWdxLY3GtaGyYg5qxpqTChvJ4mwrzwachcFevk5vTIaXuPm+eR
6PhhK44FK5hH8NuCDGfavB7XUYir9Mv+fCwfHPIanf54i8Jt8iNfbTwmKOXHx8Idq+IPQEaXgW5P
s58wpTl60qwzqTWgKehfqKE09r5d2JNlo1IJSnpMhe7toSg659KF4qVbNrrf8ofAx1VjedAG90V/
huSRDa+sd/xAmW6r0kU2K5/mcehU8prWHMYqQaDDMEMJm48NFkQse51lOulY4XS23s+KS4g/xPK/
k43uf7oRbK64RDidTFmc7Xqq2KbrG61983dZaVHH5QIFRoPnPbpJuipwwKfYXkFGKJWMTbLEgDF6
hnLnbXXDkEPBGyYGyh6A5vfQ+fUPlOl+4a89SsKgfurFftg6VPV4EXgauPVCu1HryzA3/zLhb3TT
hhEQ42F2q4DY8sgkYq0SwOGE4DorAdQJuJlCeWk1/+1T67wplkgGWp8mVr6OWDEnza/803H/GMLD
4ePdXpLCAx4pNC3HntDs4R6r1L7Sihik5pfozHkZGm9vMLGfwA8KbUyoATVJavYQaAfxgbD6VSpN
kJWaBtfIMHqQoK32DNLznHlxDPl8a2d0469K/9mEW9EPkrnc3CIW9493KObmFRWl+PJURls9fedb
WerbVWdepN6nSeDXqI+nLx8O6MhtueF8flayfQUfdMYAuyuwM59sur2gzauIe0N4q5roAxnU57Fh
PEt/XfdNa47/2iQMRNEP4t0WGD60vOqlXyg8jmTYrbUYtYmJtH+N0N/7bshydPGczXxwNiucjpFe
JE9VjuEEwTMswD0VHGJGvPmpxuXORNLlZICn8zXHXHW85Fj1/b26+k6dkHlVATi8HxnM6GLx9p7E
wvqXUckiBWt/FfpGVhTXJLtJmxkacCTSUJS9o9bTimEzIBHPWkYZri3B47TDA4Rn881g6lRmoNbl
ue/n4Ysugyt9l58g9fddQMUksXto+OnQ313Nag8OawU+9XV/2btvqH86DrZC14jR71bEE74MOAij
yTBRBCM1MsSPzFKPCIMDnE7flK92YpXVEZ/ytsT6RxEOX0VeJW3+JvnFeRZmHd+z8OW4ViyqK4Ca
9jL7TbjbOKV6OHru6vlc84EbSSoPQciuk/RPq+2BKD3tgu/2n8xYTYJTcGaqFtxmw/yjwM1/asaX
TyvSXF2gvC5n435Njo+5xrY5zsTqXklQXk8ITaE7WQRPxBScixHKZpd64InWJk1jOPB/LgbNO9f9
M702MaZKsnoYsxioC6h9u9rPBTGU1FO36dNKF1vw9v9tIbnFm9Y7RJRTTTKbJzf1XeivvLY47G6W
wXGUKwkL3LuVuvSQeZr5w6zq2oTMMfhYfN6HCfIjfjf4zs7PJlfROX2PMpWqkeQtjswq4YbftmCH
yLPQMAPAAdshxNcCguf5hQFez7E+WFuoV1NHPn55ZXBTh7rtja0tQGRcPc2GbiFuqpmcw4j3T9Me
S/jnwTrpioKh/WCPGRGyghOt6oM+XJ/9maksWmv58qA3zWr7+UitedTJIwEKc+mVL+9+flcK8OpE
YM+uAEadZ6m5W0TuAGyQDrV0gemW41VqtF9abIN4WYFIMdI7ksah4sk0vhnE72x1AsfAtX2GDRBJ
cC48WMJ0wfNSp10ikTbGSJJPV/0jvsh3JujPHeUOl/c8ItZNyy0yqr5aY7ippRUAvb5KNZImsiWD
7fY+ta5RGXEsYEPVAkL174duE4OTqeoiUZQU9ngjeyx4AodTrw7niN2zY17Dr8tv/ICTlX7l6MtM
N5s89uHAEUy7RMdBBGRAUGrB5TL4lD6B4q4zaYywE4zlR+VVRbe1GPqqaeEqZ1ZIjWRvyqU02d60
q3F9pEOcFO2iZVBM8uROtvhSKIo9VXvQ834/J6eeNNJlR9O7s3kCEONOoK9YScW3g+3kvGL73GAd
KRirIfOaDci258jkW3HfT9G7A74FzckFMEyy6rPD0Kogs2yKFvOl6+tM21h6jKDRl81+zqYp9rYc
qg99ivbPMKb2ZBVHKU0907TehWzIdAEoLpNzrLhIhvKlVBwnh4usiaEeNV/MYUZetHbzWoQHypQU
OhZQV/oIeakIOsxMTLVvFRnIK8WV0EXnwXDqT9Q5p5ZP//RCi9SKaxuPJONH64tahxvyFweWu8R5
+DImIYe7aL3h0GxWCDG8bEOOXX6Dwc2jMCnb5qYt8Z6XRLMawVQ0vuD7CjtHmBDUrdeqAuNQEpTm
5DxgiyyGUd7fP34iRIf0NhU+XUHk94CZFLrP17fT5Q6pcgAWd0bpcxsdahOXhhdPKi9ZW2qH0CVE
KCS5sexRwpyyuyndgrDrVLZREQut2FqEhKZZQYgHYBDQfRhhLSDEeJbIR1MXxIexrZG38Udsr+pC
mqNWUU8eHk62QSYxBplnAjRQ+Ua2CqVmTqM12KSOEv5vJWhOs6O+XXvIzrQOiAYPSsgcgyUVt6VP
FwISouu3nf0k9JRyC++6SwV67ruZzWcGeQ0yLj8aqf1m9ZbM23F0LZC3a/yKRuSy3dCPdOSRs/zn
Y1RrmB6oPkLtMtRY1toQeMt+WsbzgXfmP7yKRNMHVB0b1sHDNw31NfwWdIDVjLXdsP8Qfj6PhdE7
u3MSG3+6Nd5SY829+WiGKNwi22c1XSMu0NQpfqmkTQKUq5PcgojbyaQN9DRXD4ZgznI7qwyk3K7T
WavQctrblPx8TFNJ44gV+GZy0jtl/1mLvb05ABm8a/1Optdmml8wkuqbjzmnCeld25VPDvf8jTo0
sqL8nosNQabLhca8JxCYON0IOh+B5lbL4LvZFJ+SxWLhNuFhbjGlAdKLPlVzqSsWviM2YZPtZcdj
ViuTkoL9ifTulw3xPQyGWBoiMzyvBNPY4BYAvKXXVxWfcTuLueRGRL2BM8HiXhqzuUD6Ef50Zq9t
tU70iZGp4B/0isLxzytO5p1tauqw0awm+9Ib6pm99UmNsYy5eiKXPj3Y5nECDnHzxZp738ry9EEK
39MIA9Ey6tVKPrYpLwLkQgDhcoyA7DIBOZVcHh4NaCnMze9tIaVeSBNOAv4i2bYBr7a+mpXKkTjq
VcsRUi+NcVwyhmKeM/+bDuwke/DV9DI+ivyXvkG5VX6rMSlrjXJxnwyl8JS6Uw4QjWw2x92rdOCL
odP5zrKzU2MEwOzdvSHiKz8M7rsdSVwsy/eO0riyqzdFnED2THdQOM6vAUzJSZCd0nPG/5CnJoZO
aP6VLVuYHdcKf7horxHAPHfasqfXkxyQEQ8TDhGcQsHD1NR1iH8NEJIBhVgN0N7LXi5mgdqB4b4U
Ej1KMzSK0jQalUy/nc9dD0aSg2mldAggZKjvPToZd7FMcf1Ovm/kVBjMREsgopvLWL0o+A8UsN4i
xcToKfErHuc5sHieeUN+xgDDSx1CkKyOQ/Ih7qC8PhLCHl2yerjeC3c3OT21iuSlpOiwwCsrbhbM
yIm/nGQLnju2cRQgghOzryDkILBCcYhPC+34bcKzFqH9QFeh6hF/ZXiwgJRKTriVk1/Yl+rExy++
qif5Gt5APuWt6oknPvQgfakpOE5iEJpadHXOFtErLViDdVDth6MKmfurN4pM/Qttm3im/5b1ZHdK
dfhbum9RbgyJBb1qRT1dGuwFoRpRBSI7yfWR2d5fcj4txWBZwyGTHz8tpHIEDMIsJlPx4MQoiuno
ocrm3llagqGDEiX2zeu7UV8eGQcxLVBrQBIHAelJRx0Jxvy85/Uq3AF3iReUTeRy3j4UCj88Eruy
OEG4gLd3e+rzj5ZRh1ET+ilKkeA6HWgPeRMdgmo6zUrGPcJ/Q+u7iuXI60v97FeUYhfoggtHPvwC
ossM6qw4Whc+MCi+lujJ9bVGdG4QwVvhQPPz5nJo0NkRm6QPoQIpoD98ZAY7SKfrRb0UptPxe2el
aJQ80pycgWpM0hVCgNeopga4SB+ZGKQhIJslSrS4R87PhCAZOo5wRSDcOLTp/vCRiysALNdbnyYv
C8i9p+PFN3SQ4UOWdeV2LWa/2M5q3xmDoZmpMiZxfqG5QYtPiPkwpvrtUq1hP6kpdaOn+YFhRbPU
rF4eRjYNFTNbY/BI7wsDO+PBThlDlrmmhajn7/Yh5iFqugUm2/vNYEOaKp12BgTqeolGA6K/LoCM
eF+uL6SODARlWwWW2vg85XIxoWarm2it73/3CmyyB4ePxE9RicOdLuFKs5fBqKFIDVK/zdEgYdgO
J/miaZ9BGXamdRu7PRnCK7CG5r+GgAwYmpxTfQejJOmwtsoqmZZ9ce9PqlVyCFwSH2TlJQVH4Ttr
KlCg2VFe3Eomqz0behZkRZTHPTMbnb1RC7arLBUQ2qIFuR/KbGcvSjZ5FpcnI6wfnTOFZD79Pgnx
YqP9SE/tDko03u1AYxuOvvdG3iJDIFTfpi7EFCRshc7kHMTOjTE34naGYG7cgQSHedfsIwmF90Dx
qb8HL5zWP5TzjMVVh8XSXtDcEcdKV91C+rfrbQ14/OWx6Kk+Lux+AZJ+l/An0HVtRBjMuSKJdwdO
ke48+VUGLG7z1Y8GmkJxjuW9nBpHWpSso4RAl4+CnYYhXl8yBroJ35+Zd8qHx9VU7bp7Dk27nIvr
wRAnZAXZMWaJ9gSbQ1eZOAjvEsOy01fgf2V0KYbFtkmH2XL89wQvrVkZyqP5U5fDP9zAcS3Rfw8l
JRK5dqGmysTMxVyn3phPgi/NZOfFoxvQGF4GYR+TwzOCp4KFOvjwj67D6mlDx9oxiTqPzK27Dw6c
G65SpceYPJGaxM56QSnNmoXwbCJZx3PSSmwS7CqRo0wGs3O51oAwMTvL0DdsR9RCMuEMhiHXitKk
g7OsbB77bexMoMUxP2A6U0uLGuKGa4PTiQpo6Opm1w1Ik9YJ1H8G3Z6RtqfaLnHu24gHEa531unf
+WXOLWh/y4fLxnoZ+Xc8xJVGmc9ccpXxlVZEIxFAm0cZW0jxoQKGIlchs9GFc+Mc06deMgD8Z5m4
ds41dOlO1XUvhmdYG7KV/7KjkKewnQL5Fu5GVGILavnHnvUMbLbLCtdAnI4zomWw7osttHw4Pdsf
ECezgiS2OuRYWxbkrJXzcygU159LJvYnIBlPDU5vU9YY1JruGQFQvKTZGafxLl1/foz3rwZh+Ga3
jIKimokv6YEDyh3dc6Daax+rdY1pUXBXSkElrUINxHIUp1KINDhPE4WFogs731z6LA1z2RgRNmox
z+1i9i29rCGDPxRpeFbkaB6Tr3YDCD/WOIbVaRm+GO0r9BePhMclqRbyE3Iw2hU/ib3Ghz5KqiC/
INjJqd5nqyly/SZTImbD0nybbC8hLgHsvjNF6PvPYp9DRWmoMnhPLhpHF6u4MdDrv6T5CEY1IA1c
UcKOsphZNAumeLsHYjJb4fvSRX5liK8fbqG5aIt+5YOS/m9sNFhB3IbapMhZ4tChs0R9nNxaDbH+
Txyu5aNSIMbnzA2AvjQDCBXtFK8fJv6USB56QrPwDn3820eE46JUtLkNNYNH8/R/i6xS0kueAt7/
wzQiwahrNbKMq4e8N3rwhdPXiLpmWQ7Eajb93cnLemE1sZ8yYR+ocVwXFMjm88c+LWYRtjVlhvdf
Rn/Fo/gsBIMZsWPJpcJ/gygPWOGfkAmmbrxOLdNxwVJcVxXq0H2l4deqB9mZCBY4fAz6v5xX7oq/
vL1stCp4M0xeaH4Xgrw7eIjmvPopr/3OW1jJu7hkzsAytnpRmDS4qSnA6iO03nQP+9hpUGMNUpsO
XDfnnDrZX1RYR72qi3B9jdxPhWF4IO1cudXDdsT86uA+hQPC7Kp/rPgd91WBdZjT4Iw8yqkKMUWE
PNKAZ2r22josdVm0kHdx+SPxMM0Wv2onPnfU1b61xjZ2YqJCuuM/jnDTh5LfaQh3ruckLTHylIki
9HLlYoa20ipGRfBCzdVzzzcryMsUv7De1U2cY2m66v7fOu4OknatiUqMJjIsgOWKIzjtTU6OBRKA
kcQutjku2lgjl2OvHjS0qpfqQuPkgT09S/aXLnq7cx/DND0UKKs/H6X4PIx3JCsHfOrEB9tPhPbc
PUmSl5oU10OHbkS7Hp8SVRdqof4zWHmGjl6nV9CcFt7Pd0do6rVNg6vbMw4G8/a5Ab07ojUj5dwl
3bd/WZsFX50f2J+ZUTJIWZMrzq2mE4oniDs2T6gKREK/0kUfoUTL7LJOwgEcHLbpwyORyDZYgj/N
Y3lsw1ruNofjLFtgO+GMCxuY+N7uk6jqVCvdhuudwMxMqcUZis4nFpbN4ZwuUUPr8bf+3aD11WXR
am74el+7L0kQT8XJyBY//cwgOhHcx/ncwwnT5/EJhzCIGLxz7EQ5FATi0nLMSzUV44dD9kdigJ1U
0GhNKyM/uuIdf1Jje69oE5sHMfZL0bmOZasHdEKdQiXln8FrlNtPKobhD8NfRsxhZ5w/apyD/uRx
8sQ+r+0XbiHXd73wmnm/Cds/FsCTygfgO2h2wCMREkY0hUDtcmofGnDZ9MqTAriOJ16U7pQzWjn5
Nggjh5HmrSMC+VRt+T8WpFZckwE8bHsJNLhM+0TAjjSsMQ8lJF4FQczutAW6U3/ejntoLcDrqWEv
6zUi4OLBHinN3McRSiXsxiGvy7Vq1ePGQnSt6yE87Tayfno+bdrGS0UZynXh9k73HMGgCQp+K+Qj
ugrE5N6HBTpw1mEEO7/VAoNW12MFlRYd7ZrmK5wGcnHQG63olcSGP+jU00HRHdp6oYxSIGj9AZsF
BLNay5HW7GhziejC0aigBEiVV6nWk3+1ELvN1SknSdBtM0DJTlOcGC9LXGJn9kyErZhDU1XPZJkZ
FH3F5oLS3sPs9ZmBtJ7+JtIURXbkZ5fAsVe5swhOwfBWW3KZigFdPgcXclbOSjSjiqvek8QcKhS5
5decfZvXN6E8w7GAHIV8wXdLVDh1vBPBEnhTl5YcacUDgSLx0RdTFyvssTEuazLudh8FAjtYBuA4
2leIC8G39s4n1XCrKWKkdIv/Hnrm6hBLkhEWmqVdCcnFojCK023nloSXKGPLftSNR1F/XUF62Oo3
JD3I1NkXeeN3nTwu4E4UhVZDVTQCjgnyFWKikW+e7HRv24QF7Vn/Nuy9AVR4vfYxHnUP/1phSsOr
fn3BFP6q3nUQ7KWzVu/lDpm1pg8EW0JOPaKHS6lOIK80dIJD0kU8zaZ9YB0XodO3iTZEezO37fek
oluyU7Wzpnt9zdGz7ZQkgGkrUhHGXCyt6p493UQKVXSnusBodN0S8PdW06qSP9YinbAKJozhTDOg
o71HlihsiN1ALtEzxC1qyu54cyyMDqxRvWuciv12+151UtF5ukAMZ8xX74W+GsbNLJWoUpyLlA+z
N4orQGwWk8kXGxtfYwfQgicqUFtsto0pTWc0ucY7EpZxQXxJRoOi/gu/QNClHXK586lM2IUpAVO1
jKpgH1Gxlhwv/4o0ow+6I2+Zd7zY7V7pYxaKZc9iMal7rv3Fdu/IyonAngE1a+30EL03oc2aYpcC
KPNxmGcymugwdR56QYhoy0sBckz+lMZ9rHQLMn7Y4ec9GQbcKVfkqgYbpn0FDMnIMam49cjzY8d+
J6Z5a1L8en6hbVk4MN64wukbuy5eDY2DG2d/VcwQ6QdyeWVQA25eq8yW5W6aLepuc1VcNpmhzeHG
8jKiqIsZ96/BIoji1tUhpQvVqcg1T5dkBubL1E3oB5HyTgxrtv/MXkwkmwZOk4tvvxrFrew/z/19
yfNf8R6mPI4Qsr9PdHYApNUEvt0YakZg7KTOofdqIWrDettx+2KCzDzSmD3QZbPvxXaMDlzL0kl9
bt7W2PNrvUOpUuocoyjLAuVEFPmy2eAYemKEZMt5OBZjKUfE46XYZUePPYncFF2JtuWBQ4RJLVyM
byEtqU26ixUUe95LoowIN4EOA8y9sZBQrhSvZF6BkfwTskKY2TbYLvHXhekrdP80DxJlKoNY7Ze2
vzhDhh8vJzpUdXIWeR1lQB5NaLu+V8wAd/ch0FQrHbiBOzLyg+zwO7V9Her6vNLwr2UmI4PlT0bJ
5vQ65p26nivC0NUQBEI8wV7Fj9j+rstrJp7hriporeBTPU2+ZmehdcimrmW+YBSQCjCl+cZTJVRv
aytkeRqVzemVj5XAlp9jUvHmzvnrF7UMkzmHwNeXTMTcCLB1OT1Mu0GEU4iYD+rTWuWfQS9EDxvr
WbGONVUU8HfduE9l+X79mraiqom2Kwd5ECH14W8olu2bMkl2g30+e4pr95DY24RxrVMY49h4WrsR
xOpSAIPwRUa3gS7lLSPiJvUu7xhE181ZlX8rVwtWTBFb9HeMSFIrmlJix8hqzWz7Q/lqXm9WKMeL
ASkJ75pgpkLZOm0LiOtYi00bf+/eltVLkwHW50CS4vJe2VfiUfhPiYhBqedQ/5Ak2o/BCoAo04D5
7N92pwDvcrKdPAnVqY9TnfvNay3W5zgCfJzdOufoYdKLvrsaWOXl47vI9DJBAe1tB5thXtcJCIla
Mqr/CHLuhrwBBZZCnnvzt6oMdWxLOZCpUZEf4D1k88nduUXAbIV3LRPdhlkW9YczKkxU2VDMtdoD
PQz11sdQWMkd/VD/trF60grdJFtax6DpAkezSpJQ7UODqVmHLUHUkr8y0y7VWA2tBjNB6+SmQgB4
3aIdl6SoX0du55SZVVb8KuiEu9JOThAFnmoUGoImunE/G8a7rkE+XWBbr/G4rYKU1m2St4n+43cm
XR7e+IvYb6T9SOcb9dNCSrddMhN8mvJ3GIZrM4FruRpVGlHm3vlB5iqjUfGkOMpviXuuVucbeawu
7p4VRfNyaxFcedwakyvpd19DboHcrauJyqkdwXPfIsDRXiOHfQh8xyNOR6+r7Q/s8Oh7JzsyqlMB
Ii9cW4sLQ+JgeZBqRcu02JdPrHp8zj+gHquD0iWIM0huirm/QH2rYbDszVWwf1tfUhZ/yzJDaHjC
90YRakUG2Syt3ZDcSWy490wDulZGZCyFBIrZerY+Ro6QogC1v/lBuygt+xVvx9qm1Vb2hvu4oP+A
B6PVxGWwqzjjUjk6hW6u2xm3JXKTS4n4y72i5S41dp4t9GGBsr4duRAImNhci1JGoZDjfzwzsxop
YyfkVE1HuN4Y3Y8Cc5UoijslXeFVUBvvf6axUyjtWaOTZWYHWFMZ/a3xQG3aCLIaRo+5e59sbGF/
GZ8NLlXHzpE9h01nyJUQ4cTUfOnqOrAWazUKDtyUCYgDadHZ0xK86vbx/m5nJdachxdSxd5sdBdN
SjbcOq8gS02hQeaPumLIZKbeI3UBToeoo1KA83ZfiKShrqXqRudOJnf7n5d9a2WY5a2PTXkRCVPP
6P3TyGxRuvP7N5SjUz+5h7zSZrv8nwNf/LNfIJcVPUa2tKliinSELqJdx3YnzMKL30dLc3ARW+xx
g6k6s5QE1PONcNi0U8W1saGE+12zZn3shD8FfuTaLL3lnfUqZPIjZNhCzUATdk6kXOatm4T9ltI2
2455jVqXeJQcivuIfRaTywE8waZLCAZJ8rK8foWGh8H75izcQOGSqkuTThzhvw2qLL2gy5Kuisr4
pbV2HwPcWKlZpfIBOaxSvwuse0xpYY1aCk+13ulNLecHizH6UwYMP24Fhh02mn4nd6Ek4Ek0CLwP
lEbVJ4fvosF4xrqEty4Jb5Yc+Hx1m/R4zu+1ClMOqRv+Y/qF8ptdtyo30V9kBOiKhszWtAR+MTgZ
bpSTidvtPa06voUFmW6WqvL55nqcLDe0/tm+0mAKT914CtEAhVbGzBPgrW82bg7iHf3E56DK+uFk
gtAN9+8ERM51pm2kUiUDBeFPaIWfDr2ntHt2BIo7hrCuWvOrfN2THsV1UGScu6Duyu1yscNDpPmD
9seYNO97GG9tLb6Bapfnu6+jXbn7TVSio0o0sYCgXdSuvHM7gMjiFILtJQafiZUjb1hW+6k9cWJG
zFg22RctXWDagkE+9fQwVwxklC4valwfd8JSWHm8d1AAZGZy9UVg2+qzdaFlkNq4kp7lT/g25KMS
orDuPI0tfTR50Z/jf4KVqxT23oAhrh3YNzZDj6Fb+YKF1LKw92aWooG4E4WEuSgGLmzqTYcE7eHs
OmS6gekp2FTuIgkLUfRfRSiCJR1o+pLIXvFBYa9Fyw7wshoXhJcIh7fo461p5KZDAE4xpML3o8fa
KV59c1kbpVqGYbL4Ev8j1NNstGYQcUxTjGj9KfOshdDUK60DF1US+0jAtL+65WgwyGDTZqv4GXE6
vj31WFuCVZc/oO3PrGyJf0yynjMCpa3QcZt0pOx9UjhonXmYMi7lMWVxWIF331s8JRR14TOWSBY7
GzPU+imcZJ8/qyxG8HVyneNGFza31pKOlxGyuVKrMYy4//ziMyepx9TRoDuSTvBbVpU0KGDtQY97
ycENZlxQHanaZ1PWS4xPlK5rOwXHuRaOMd0og7zFBIVLTIcmtG4xiE7AQWk79aI4ugjRM57zGMAE
aJZXbrwlaamwMxrbUOp3l2bxDCzLCT4u2IN30T+aKK50gkvYAza3sgEKaojQzmu7Kmln3HjSixY6
P3W5fJB5G+LQS6GKaJvO8ny+vsfg7jyhctiOuaqyIy21hRouPYBWl/oQLXK+acscPQSiRz8Pd/qF
/HQGruCSoOP9VknjY2KK1ehhdfQapwtrytNCA+cza/3EchUoWD9cXZi02mJs3w0GDSS8TVGqb3I5
Qf00AKyWF0P2z+vj4KYJTu+z3+obUUtps7o3OC6fpQsT/iOnkIo80ul4nlFaCRWKbo9iSagoTzTE
X8nuYelH9zOOHCVIRJCRqsMICYY2XyPLIrQdZVqTDNMwEOCCKCPZ6lw3R4BY61RxomAXhy23S32S
4dgGmkvT3oHkCv1XkzNauc56OYkiXCcoPyJu3p6TCnc7VWz93doLQskccwYmkKQLQvRyLD/UYU/4
9eJpk6uTODmCtFGOYYYuUtlV/Yn8fTjg0Tgb2BMsNjfOW/238xojZuPi2LfN4vMdd6o/zw+J21IP
+Xu89hM/l2JEUiEHZAlG5Jez9rakSXfV/fKa/F2Kx3GeoX/sfX5mZBAcay1xlX7HrUVJK6RRfN5L
IW2OpBTS/UgliTNvUg241+JEc2MYPzg0I0AsjfaTcjTXnk3N/ckV9DkWh/b3+w8ISnAOdeAOMbJ9
sV3ssKE+pzd9IUZ3Ef2oAQOsP9LNgxG/GxpaoNBx/yd+xuwslq8JWTeVpR0KVAWaV/8lmbY5cM2T
SKz/ZpGqmlp71i9clFLThcYWibjBjdZsIbRcQWmn14LWePLHDi8Brz4C7V/qRTUeXv+Q27Nn0A7L
IVzdwp0EHlQXtegT3roC4EdLQkngCLw6r9Djv86UWOzqVsP5KpfUoQi96OMLTOXvQbHiw1cW94rS
w9RwfhZDfz4/vnA7Zp9woRxFWukW2n99IAddoce91ku09So4qSiOQS9AGP1JJsu/PqxymprIUsNj
8SoPFBRvobLBl2/JdLug0xCXpXq6FojwwRDcwqVSi5XQZ6rvN3+dpPOOoD25HjgzL8y7yZj7zaVt
+9e6Wc7MgCjZmh2Kyv4JMMszHGPI+sToP8WanRSKDvYiBc/zYoHIJAOG3VU5uEWN4j5HpJF8MPT9
3DcGkQ0HoghHlmZuUBx3HUIR6L1A8xQ4Z/KDnjlM7s4P5bR/WNinfiPQCkCWuvpvG54HKVn9t8r3
/fbP9R+DYs2UJUnrQzVSjTN7T5s8lf8cdRv2GuWKbkAlUK4l2MLzJXy14py0GDhAFTecBXg24ku8
+UPH28ROLgFuJOG9ga553jR1R5DxVo+lB94g1WMXBqBqPk2vSt4NwkmcNh/tYk1a8pUu2I+b5SJa
K3TISXjqxbqsETiJmQAsBVl8rJO3v15NYQgs7GxrLdQ9hBF6AjzA0CkhfSnfHXu3VzHZEs0qzODV
bSRmXY/QKuCMhMZ6BGhcnTkWweJirD/AVNsxDa5maG1lS/ucQFvgUy5FvoLdGZX/5fi7gGau/xc4
t+/bYdFtLpf6C+Ezj/ZdRlNdAOd+Y9MAhFqOt18zjLid3FIqNeJnYare0gPP28F5nsZirEra5lsl
vSOBh2CdbGypg5tSjAW50FeUHhabV5qy6kZpWugu2/hR1lnwG+fkuI3aGu2VJoviNyMmXOZs8TYv
WxoiN4PUwyayELyag+uYlCSqf1WldeR6E5he3AdJp0EZXXJJNy0e08uoJRQLCu2uJJQ9Ax3+tyN5
k02LSZiST5ZKub2xYtMjrPuq13llAzQaYGiYgQhnnAeXjg1a3pbuT4+UK+PyfJbsJVIGlxtG16nx
cp8VSGU8dJCLn9b7GRBqJXqT1yzZqMhXnswwyIoAZpSycjRKt3yenguL04LHzPUCXPiX/wq0K8Rn
iDhp2vHAGGfMuiS8yNxUKKbU4y6O4TIDMyzvxfeq31vn0lhUz7gKqmWYhysVdvZ/RRpYqKuB2982
RQtUl8lOrJraWqss1HJo4Zes6Dv3+7HxiOEFuKZ/nSooGM+KR+wngwsdLE+wPWXKGhVDXRi3uc+h
DTStdT+GRboUh4GYw86FU8zi57u5awFnQe03kNyquAtLvL1z2R6MBcVM3cohzOpMBLhTDpc/lG93
AIPNsNBoTjf2GpbwY9uBc8I5G58EaJfYBslAPXMnEYzyEkPoMTVIdsZGrcuBFN5D8XVIqcwX92w8
wGuvlyJeMNXydDqx0ZAJRrNgNnNI8ZVQTPVi5+E/zGcl+tF/hCXKlujluXJ1TIgIyT73d6PQfaOO
f57GbLbQmiyxG9T0l7sllKV5eBWpPI9tY7hIut/2+/McaR7UmOSMmkBpltcCjZP8OyArofX3YXXI
gBe4RTV9GVryCGf1aGNspz9bsGYdAHnJO4Vc28Kc/3LnvQ6CQP9Mc5jr/IBnN5t+ZKJrsFRv+E7/
IVdM4847LE3kZTEhO1F4TCE+RIc+n0ZrrDBiV1VdbNH2D4MCxX1m3gncf9Tsxe4YENqQbZjkH9Og
ZsdP1zzJc9kcpRJWNUrZPB9a1/Jsv7nk95YWkEVmFgrgi+qoWH3q+xK3Uiz+3hwkEiG/IrBq+O0g
twCrlyjX6+S8FqSkdMUQZqeQouJMb7OlpJG/S1V8fzG+RjmLf7EwclBETGHtRxi1oiHn3wf60DT1
Lrj9U7OEY5gPOIMkLeYdLmEZEJsx+br5F9/tMCSl2exAYtCT++Jx1KLR7tgpW9Wx+8TmTPFK707h
77dodfekneCJgY4oaeNnWtjbnEiAN7oIa/nEVKldfIg7kJ/zehGCB+7icB0mw3iZTb9GMDlEGNry
rYH+hfrhQKeks62D2SzgGJLctS7ReBN4gkacKmXs5kI7GtD03gd8jhLSdW18ulc3CV/nh+dUGPpk
Q8q+Vo2buhTx5ZxIHdn33940Fqj6nK2L3KJm/ufN9n9rHoZb9NtRqz1k9BsXs+jjq+1V7c1Ih9sy
Mi7/S5JtlS6u667OTc1/qHmB5tmZ4fwgP7RNqWbEM5+8uxLDaUFZd1OO8wPfRJ3rsOoOAIvQ90z2
MUu22sMYk0eEoHCjvDJceDcfo5jvCmw+QcfIwqGAEns6ULGs4gSSVxYfBG44cYkxnjIqXVK3A9vg
cthLezQFDBegk0LJi+QhWXfOtQywAsugrpO4cq4burcezHr+Mw0NcTPKykC6jYPy8AsUz673wYgT
kh2NKI6pgQrS+acOmP5b8PdDq60iBamfgG3p+XJrjjKYDmP9/FoYUEe3B2p1QQnZ7Vi5hBZBuL/f
e6MhSBwX+fwnxT3YnEb2+yJDUH8HhIHrTssuCrEmzGWhv8+F0XOAuUGOHitS/ThNTxbBRkQ0a0A5
I1JRN3/15arnQ6vI8/9moVC1m10sZ9ihLAV+qcWy+bJrslXJYUQHFxv5nJBxQf1HYze0T3hkNYnS
n8RVF+g1q35hQDAlnuc2h+1uj2P193GxQrgAHfLnXwwZBqQTAPSLP/GCz/Pw9H2iJxwsJ6J6rejG
l6Op6ybrpIMc48zRm0RVGU26FO4rdxppSCHVcRBxtXg/Sc/bOBCWdJ6jzSOqhZhk4gboH/RqnSvd
kmhFBOZrcrvbUza0CkaaLcys0cb671wXYk34fWDtw4+cgoTYh19Hs+7AABz3D+NSKgKWNAl5raCw
UdJG3LM38doPCW/uJBXtbNpzLxy5IYY3kc0q/Mt9Vx/DHcU66Tmgnq197HYTI7BeQdQddH9WDa7D
5/D5Zs5NVBo6UBHRXPFWH3i5OGaD1pIBryy0c2He0rbQejMvfFzJ4TEuCaIEUxNWhW/8JL0fcc2f
Wb/Ty8jIIindG43DPEMOGJA7WlwX3joB4xN1HqfBNArLgrprYYow3lMhB/sZKLjaSxNIBzAXD5wf
4Wq8cPsGoxkx6Y+0JZqxOnzJXKSOsBstUEqcvpHQ59QPOwmmGsS4abPAYDXMOSALnsawOt9WNJ0K
aCTHyCb9qP5h/Ht27nmAqRcHqJscmhexNKuhnt1HSTn85HJHa70dWO3A3FRPW9WHNRKof3uJSGk1
q1l0+ZGPAn4NqXRdfhgi3nBa8HNOyN3Gwr1M1hdJ1keQ2PGUq0mHKpPq/PjT9NuXipCiQPEHr2zd
MIFB+mbmat52DLi92A4JqDhLR66SzlTPNt212+aN/JCuUvKYCWbApIAStiJWIE+m5fWOsgRy27KJ
HylqZY/JNU+k1uHGnFbmYs765XlMDlpzLW0bWNlxwWDzBSAFganj93eiLm9lY3bxndc6wJxYZthw
MF0kLyhJU7I8ydINPCqij5QUzqEpC/hJcD4qWIkoQ+T3yRRgHcyLMWDSM5+1CWwpyw0S/Kh+2MuH
EL1C5F1sAQEHypp33niQj6zSt5KHIXGcHXUgAehn+7g8q5cERaqTGH5F0wRfTxCyh+jUx7dJMeWm
9biE/HYdeCSMCEiuO1SMMbzF+kxi2mZY2vaOhiGcCC//ul26pbFFTIR3eQpVYTTgOA+5tjO8AYnn
Cxk7cqlW3mDiGit1Bcyq51Jdu1seVhjfZccW28ECRglkwfRzX/hKDrsp5khh+NKhOD6SEUTrnrUP
uN/zkmRz25+e2s3jyIAs2KXhidssVbb2/6TY/nUNYl7iWsVGVGGb1+JTbfMlcek7XdBwCJlnqVI1
O5hT8lVxIwUPuj9vv/exStiydsfzLEaRJzCr6iZjXTJN22+vg3amNqLShnex83HQlUaTjzDbAFaY
iz0mEnkt4xCZwnvLA4ntrpZFFq4PMFvCi35E6QMB6q1/A0T24cmedfSkyq287mjdtrwoeaehshGO
18diNvC/ikcw8+1ym6ZcncENLPQ3nW0TezkO8VdKe0XCBU6Um+KE0VefVB3IK/JT1R8S3JBKAiO7
5wE4alfeFfHUwVNFgEnMmK8N3l5IZAq7BMuUmf0pfVHBoXIcbTJ/BJzFngo5W44Hq1e0PWmDR+Kj
31UU4IdWejAHM/dUx53aJNqteMaUXqkJftaCx/cmVwxEDEcgS+bqlgBwPEtY/ZWRf1Vwztm8rOXN
qUBf29TGBRNTAhEMJfmKJn4gDoCqTL3x8PYCmh1kVpQscLVCElFDtpVfa7boLkIP3pW6nB/DFBpS
ZUS4EEQdgkhdfAKEcJftx6TVD9gyoGDGQiYKTe/IoiH4Qufz6F7ipFluFnf/4xq5PCcdYAL3Dw+T
/A3rLDa5EB3syZPP3t2smbRcZ97vNbJh1V9TPAjHtQ6vcVnFS/hFgDlSCBC6mlJ5sasT6GkOAYBx
8wWLfRxB2g+7DcJxLUbKuE8sEsN2SFCxZDJpMiQExmdMf2fQ9zRt6CrDKoJVpJWU5QsPhIn0n7Uu
TYKuu58K+DOWdfqzKty7ARz1BeJrv7UV2xG8RfBQUZpUHQo28+vaqEWEfQID1R+H7Yf1PM6XeHus
p9GIHagi92hyn5YwVH2uxxkjZmyoRi6R0LBTN5XIrcFewDCmll4f6D5AUXegR35xIzjZuU4INMkc
W2jGPqfLlWzGBvMqjd5hDb8gc1wvzM6jJHPrE4i3N7OEG7Wi0f4+OZ7G2Rspu60OxyYp831CrsPl
PGskKwZY/E1zZ/kGstjPwn04W6BFMjJty8vtoqmBnMiE5ZMKU7XUZrImOz5VaQ3vpq81iucpqGp6
v4CdFXi7KRhyUSDAiM73inlzpMgwRsVqdBRq9LMj9WTjrlg6/L4w3Gh/+XmNJNsTlxo+iqCZ30wB
ip2j7Qs6CAyOztHKSjmvK6f2DZ2MMvt/4fhOKq7CnlJoyfKv6eiPvZ7ZmQGluMrY7StdL02NiGbI
P54c3nvaSnNn5Q38YnBwE8yYldeAM8K+E/hgV/PDcWSTeqTOIVKRyfY44Fp1gAzC20tVgBK+r9Qd
Mn5I2BO10xLY661JefV6buxr8RkIKZzxfWrcdh0AcAIV0pz4NwoTupVbQFaiRns/ec9YBAoS2Wc5
NkFBpnnPTOxHn5QGiK8LHbd3hdpsYAocn4AzLEcxkMx6N3r9zRxRIXM0zQUxdAjWQXaRt+V/NTLC
ck9zKOzoK50isHWYyyICijBh6EOMjRp6Yh04HONy8+WIhfcOGvESObjxqmh0U2X/AEeyG3U54A0w
7OZWSSnAi7uFKruVSxwCoamTAKS2/Hy2XfX1hQrS6lL/MwOTllpe/T+A9VLUIMI1uaJZ8DU4VSQw
YsFI9LMndlwVoZ1KjODb2zVoZR0fRC7eqLmWjQlv4yfW1RqLs3zZ23TZ2kN0/cJ/ULpMJsM7SSCR
2Ru5AvX0WytKLqAD/LzYvIg75Q6OLSZMuEhFhgN1WegNqnB+31NUA9qc+PusaHBcG4/sk3lHrLrY
2YCabx2V1+WHGJ7EPiNUdJ4HU/f/HjB9UtDNwlmEn/9krMXkU+SDT0ljXZh15De+/IgVF9M6KUTU
Qpbb/MPcWL6XsCwzFTERBmHBOy35B3ZpTmnjl1CK5wyzOAaGToZ9UZME93ZI28Q/7Im3zkkohShw
F6TRek7vVuoXn6YrpS+W4vUaGoXenzrAp4s6ugBxoXwayWkkrfRBvXLQbfaiVeGs8SgDAUJnsGyS
ZlRqpSdtgM6dRBMATjcMFOP6hySKD2u68WXocwZrW3dzj7KHGiZ++b7k+AlcUbbt83hiGCExb2cC
2Q8S+Cgtgj9SWk19Q6hFWHSXvEaiAMm/l9CtzUQxm0QrQ9ojuly2Ko/RCbx7qLIksrAYugd+2AwS
ki4XaAovFnHV56yCXu6lLE+vOrFVeXofuFY5U0egvgwBrUkDRSQmb5uhXktOPMF41KXqRHqLJAhn
aWCZa2VG+fIEUqW7zaKDx7cc05Ui/KODcNhMGDsYS4GSXFpTgyiYGLV1oxFtmBJMcm3ijOclVWGw
E3/jgnNIaFTNQI73mt2rwoEFqXSGv/shDcdBccBvPs4GTgVzJVhs/lyNwGClKWjVg5hDiPPv8V7h
taVjDmqv+bKsm5FztxxQXiqvHTVFq2EV3Vmqmf0sTR8Nkau0kgfnmLKPe0uCFBg75koZV8Ngr5DM
BRZDUHp5fce/mqlSSkQmZBCZVnK8Cz5f6257ZuTUfcrplng2KX5795Do2Ix7u0nrxdt/Fv3QWJAm
JofbbIAwTHkHl4u3gp8ASBaxp3170nY37b83Y78uuNvgPYw6mMVY0+4zINEW9uh0nxDOxLMaTXQV
NZQBlokJkEGZt4MkR2xuzTq8loKYdtRQH0u9+D8OTu1cKLb4HFRuxNdDT/tUpd8fNg/unDxiMSqO
tmQlt4z0UWKusz3ADs10fHhrTYV6V8CwNvBPsmxZKHspI2c8KhQLnGoZGcsGQ+NiSPTVnNnuR3vM
6ur8wAN69oUs6R4BWX8BGVHu6/yHXSB3kIkNGxZtSa7UwDrOwgrYgDJuRt+/Wd5VUw3ntvAndKVC
njmvkn5bK7KpL107Ys0Gp5EoWBS4wWqN7YMeowNQ2cYHCng5+sVDxqrqSTGDu837mm0nsJFlOpz9
SzbMQYRyznptn91B3k0Bi+fwU/6fQyte0zlDHhF42LQS/rJN6cLnozqmco+mPjPEws97DcwPgVRJ
LQ1WoSgX6+4/cLwTEFqqtDUmNumJ+znU3ouDvnB7HJdD3cXob1m2In/HZtis7fv7RIQFBHuM81MG
k4lBTCDPcYbM53izTJdYv+LPoRSgyaZuLtBUx9YeSIL+FkshDQuluGKKy/3WoouJRlSutVCI46v/
n49oWSiHTf6kb+PoPhhmNE991v5YejCuJMsfPHCE9hHpJVp8aj2YP+kpM9wjXxN7eHiXgkny8yds
hUIIrDQKykG3HCoDUqBh8EOpKKs9ve9SskJOyfqYDieV78KbDyS7nzioylpMV/imoduQH2zMsi0Z
O28OQY+MtK55b/mGr+gn968RjsMrS1BeZllcLzrx6uIgBZpVvYsp9qE8rT52WgJrm5uN6KKXq4YG
7AodYkLwJdtxVnHhRV5Ykc6bHGmzIXiCgHQ/xkptRWauxiU7152fbU0ydM0aKLgyRf2vZbWdbi8I
zSwWVyjDixZYSMvFAx0EmIJnOrG6CLMpp77gHagLHKdCfJvyp6/QzZZQZ11dkI1qsPNgo86HPH5G
XCEhOig+SZv9+tBg3HSwxRrxT0w1QKjpDIZWE0klvcjRlQUxjywH//Pqwk+aIuLqMb8PRq9+cfUj
+vrNUx4mFr+ZCysDjzLYgrGMd/3S1gCFvF3lwxDiPmuwrWG3ry1VwRFNu0DBM7eSRt9p8YB/3eHZ
Dc0Cn0hzUv24EI/P3SVHGEEw/2ROUHlvUrsd1JY4oKUNTApT7obErjUts+ulO4fE752jhvR7Zyoy
fIkNoQSrM2qIgBocAgggsrjqqiCqrz+z9+0ATTXRKQklxMxoSSjhAEK0gwYIQSknWmmklLvZNvIJ
39A8E89axM+AblkJu2/QKEQAIYPpejictqGpzpyPtogRppBb1Q6y0VODYDC3C4jXTBaCIoL05UY3
Ij92tc15pVOYBIR3qqLZxBKeujye4e/rYLbYr8oyw++NrMLAAKUGXBti1BAgqZh1yGuMpDu5GS6Y
A3OG0AmLkjvn6x+eQjxbu0flaZDbvRWcTROgPQyTx5oq3Pwcc+i/LQusQipUnje8QoQdtLj3eKJt
gRRgkagqtjLAlsQ6Nsnx2YHe9PfILGEx1mw9+tqwhbJhhkj6yaeOD9lLgNso7YmXzqS0htJj60uS
zwQmrBTfUum7GPMXmLe6zDHwQtocdaHUHLohYpZkVPeews4rRLBnwPPf4LIwygXR4t+Ba2w7QZJW
owxirI1c0xTQZKYMbTLqzNPq7TBsmjDj/+Kq4GyrdDwWLQTRNqi0MkSJkaJc3uCELK6/qHmkjx+I
kwW2feXQFuiXDZrBFSKiUwJoIC+FwiJ8+bZ9O7HJKGBE5SduMnRyxDOsi5hkTBOMJgigvoma92HP
tjzN3rjaW2INzPs9Q3KMrUZsBKVkBPVoW8rswRorAWLhjcA3esIhu98ScP1n/1HlR1p/hGHuH7iY
7Slgn1nGImP8LJ7WgF+RXB0la+JRZ87veVaF+TePAHaNnX3G9yp6mqB9pQILc1Xi+SE5Sy/suQhP
U5GM+eAuPVTSCCBsWgQ33zjezBXYyVboicsickj4QKi+Po9N/xLwVQhPbIPu9LCpA8EJ76PQ/xMV
SZu94LNrFpZJAgvwRkFRibllVR1v6fe+G4ZVNKZdhWuppWeKCdpWkAk4sNrhu21nxBZ2XUBVAGhr
oLfjxn/5XNEzqE4vvLgfJbxygZkqlVv7t8QFlEe7Z9jAPUbaJ3kKBt5C6GnFJtgkUgE9rE4KY/Wk
IciayFRE7nPNNHpvlFjQTwhFcOW2fpfrcGShCciMiDuhlCq12vmQSeQQmrVdMGiA1lzQ7fb5os+R
B+49pR2l7T0ep/GUCJS2Tjyc14858NjpcsDJxpjQYNAz2w9PdMQ7s3lvKzxAUGDKYHAv4D3ry/GR
yT6NitUVx6HIwltfGIdkGWLgUGAsOdqpwSMlag0nQ60uAZ8zxeXIycy3daZ4BHcXEZ9g4rhT9of2
c8aqfHDfWQyDK5kzoGFXR/6NfXTQ+AcoL3TDKgYTElcb9bMK4Wbj/XQsZ45tH6LoZVNbUfQLGB0f
WTssxwGhp1G7g9BIstC5EwDu/ilLM/c6iYimDutn03sagFBoGeQFUFU4YNbLT3+z0AiqKO29qtKY
axcqZjaTHUbsco3jL21SbEIirQaQfiBPyI83J6W2ttwmDkvQhhgpu2tRGCNls/kyrerA+PjZQ0PY
/nqcQq8l4RkMu6vy14qbaQEiRDG3dTwsrAkdWYlLI9RvCs2Pjoikx3Bb2/Jn3DrVPYlLiLCbJ5kE
ACy3HMCwzEd5Mmt8wmwrsCtPTQdjuXVQpqV3J+YISLTs3GQcTWhKgRSU0bWD3VtrUyl9ubzJkFiW
G9yMiLk4oegAqJ/qw+0J5dTrfmKA2gfvQ9xEY2nYoXHIecQ9e8tUX61ZJjuz0qG+2kK6Jh969sgw
Bqm07sSwwjDUWyKER+6w25o+WZNnF2R9gybH/xcS8ttGQN1TpX5SWo6IJmAZf0eenCeWjK2eX/Bg
BcgdJc0w14HLsTbkvJymXPBAXidBxvb0LfRc5/AN18ixaZ/lYVbGQEMoQRqOJZ1Uk23kSRyzoe8X
lDzxYD0HTpKTUKzsb/FzMIDatbUIJM1ZiT8ScmrJ/BHnPvsk9KGM1aHBGfDAr4LMMB+vrVuAhg1+
vtAJBCTmbQZueiKndYsRfhKPsuPgrbySWSH41rQKQyWQhyIqj2maWPMAEQVVazIlL6y2M+yn796E
CVgQ9kLHSNK7ScJGVVgtgAvvL6DrTYR2v9BSewrOU26m4F+h/unxq67AyJ4RUSI2CnOX3tWOvqIT
6y2+iY8FZZvJn42vBwnZvWuNQTRC3ISk17pcttZnNRM6KyzdbC37eGDQOE2youV+yMNahk+l+049
GCX2dVGdv2bvfIr/YdqPrfqLSV0TTSYeRMlFCOLd7Y3n//r8yg20Sj7224p199dIg8xWKJ8lTW1e
YyssqFYLM64h8EL49WljhlnU31FC6m0e3LhvxjIc6+c/bsaB5fJ/TjawEfboh9jE+JsJTPuvhRsE
fr6s2gMy37vOp9ERwEF54RZPJy+sDK4AeBQsFsCZ3RC83GUAdxL0q6Q887daw9FnpmLfVxm7MOHr
d+8K1NBpFENAhcledAR21PClHTTkKRbhQ9VKmSX3IZsuipHQiD8TWlk3m+ZXFzNMuR2LBRgz/tdB
g9qtaoBIbveF8bbc8iSGKvPsrwVmmoLw4MlgRGYHtQbm3FILr969belU31dFmZ/+6UmnvisAfnq+
PyNAMYtD5LUDppg95LnjtzpSlXr0nJ4gjEK73UmjV7tfTY6GVIthPhPILmV2Gqu3EQXtzdjOYHlU
o66Yq6+tQBf9Se6R9ujbENRXmnq6r/GsagT7VifKtiS0Kr7pCl6ZzOQrNu1Jy0qA9xzdwy7AaOvQ
4Zyltm0ccZTk3BHuvTiwQSXiQydfGrDtoMhLWldj1Lntb4eiDOJoR5Ki/0LOF82K2RxX49Wv4i4F
nXeL0Qh9+et4cyqAGV391kzSJ1K/4AVGlec121t9X6Huv+h5kGEGLnlxXetiF5ZwWfAT2GjrcCTm
Hy9nMC1mQPPYUIEGwKVXsIT5vbDOFb0sg+My2QiOEmTHn01QIYTTBMIVsQFfMrRPjt1zOakiwQO8
1FhQhq5TdAU089qGnfVzKh27Vf/EBG1zvo9CMH8/ukGJ9376BJ9fuiUdrQxKfYFQcqBRiVxIJ+IS
Vy4BqpCaRl6XhuVLT14zoEwNOsQu1CZM3FBdDJlGgNAhOn5ixGvNG0HKeRLjuHdlCDpM4E1WBoYF
SC6DIrAWgfLprjm4PD8mZvmxWQWemV9TNhwXPe+5YosXMLGcr4ey9dVLPzrX9vzhJqWATenDQT6R
2++Icy3jwcSyWoehfD60n9tlQCUVh7kGHaDJ1AtcHFMXywsHr4TdDu3mxcw5+ZsJMyp0eI4M6B/F
fF0Jrecz7uh1qqK5Ry5CM4qKRHTuAxIuwbNtzID0F6evKav1Q6J8bVptYDQjYPrNsw+SU9R9V5tl
wNUujFBpKXmSxFyyWmwtUtki2VdcfOMQZJk4L492WZzkB1yrztr5oEgJW1CgI1PKf8ZRJKEIAFqd
VI7AjRBGUDCCoN8/3L+5oJsQ0SHEzwM4BE9NAmR1Soess3Z28fhiwzhuiuBw/FG/8N9YYOOTo7sD
dx2S6mHnd/M91EOQblkhJ1Z+0TU8pbmN0xcvk1clVxGA8zC2ZaQoCXxAPVzOLOUH2MSDbuEFfa5z
c63jbPQBqaN30+9r65bJJCC9HDFrpEmpf6n3QB2wVkCJsSS8NOwGl7BLCkBQF8j8ukSmPMc1ISMm
gGxl9UkodUjftOOXjZ0S9RMTRooMWnEGp/7nSXboPSBjF5gisePG5aDD+SJv78Dm5HwCJgpPHPNr
oA9nPQConvhB4gszVhQjPEHX4JkbNv63uPhpgFjP+hu6S4lVz2iL514Ui9YFN/Ryj37dmbHgTfOZ
H8BFALtAa40XJ/0vVehxGMs0WqLtNwbOGHeatY6Fg8ZcJbyHJMLDOOvTmPBQM9VGaqyZLOPlLtto
OqqgErKvGx7SciadgNmLZ/rdWd3avGIuGQqR311E6J+piJ0VY8qVIgZZVoBE4431X3D5SAQtIBwS
KfpYX9UrhdMC05hrsxM2/2kZaud9TVY3oiwSO2Kd8rjfG8s+1Xvzi57GePx9jwzdnqD9dl4axr5H
pcTCvDC3FyYU/3jmFm/6DQHjnSMG5Sx5tgsty4OwFsBFRULeMpFKMh7laaall8H3V4aH7uraYiSo
nRe34vU0z7AhzSONVSuDyMOPB9RZMjwncw5clFvFSW4VO+4KhwNxP4lYK7uTc9y3YqjXTHNDvND+
a8Fv/Ue36K+1/hJPhFGjqX9jhpx4QNL0OWvRnXzA+sBx0UFvywZ9eWoaxxtWLAEqesph94uWJtuU
Oe5AS5uf2yLOXpCpRbI9GWehKHhMdPHnKAob6sSp3PJE7zdDZ91RHX2Saa/hOPzznuaCadaxTp+b
RyJSPCN9tIE8RbEuaGDzD/shegmwy7SRlpg13jhWPei822kBAJ6J00WoF84rHeoxzqMIsOskZZU1
FMns0VzWCdgOT4IL925vaYkd7yjKPcV/eOnoirGymlnrJjCspuQrRJXKDzLxYsrpGxqk6ykxQaTi
DhpHWCyfwA6o8jnK8qSnq222oLTj71xbmumI5KDbJ9BtLQMp5jUEKBaqfRrBrOfSsnt2Ax6HtIm0
+c91xFt3AxO45RfkA8v8ZexjrFpblnRB4dcJ5OborihoU5XI6UDumAmA6lBSEhEaFUnsmQKuBwZJ
PGnl99mhYA7NM+gQOco/wlbswfxZ6ElRsulLNtJL+mH2GTaYvoz6QiEOoNW1KW2fB6TmAm4+ljrE
siore5fGS1QFORG1LmCB+q29vIqtAq3j1ognCN0ehS0d45efQBUJ1mUJPmrjakZTRPOqQ0bjfGTU
1KSsE5Q4rVEwRNsYAuR/UnLOc/hYXqlzayviS23JjASrzOy5Uew7DavyF6J8kXZtI33I3/4iVWUK
aPGPpGw1sYjLI/qT9ojSTbinGdHr6YZNsMEvjw8BWOex2PTd+5MskBZJSlZ3Cso7UN3iiBwO3li3
DObI5CXK0Iq0s+yAmIdK0JdvxodIokNOOSDAC8IBZUbXYdgY8InMXPZ8WVUK8uh+aou1kOmYftBN
6yyqFSOsg/NUWc3tBbS1sQ6RaaXuuQZg4DvSP7EmlAiA9L3V1dkXmOZjehpi/p32dwr1JK7+wyej
z13rs2rJtrJz5pxx5Ut0JAGO25hmzTAVz0GTpeF0YS0F/n8+gpAnJdG4VrrOg5ZFFSbEj5Z1iUv8
1zfMKuqFWsTKULuT9PT7hT37g9A80NdrSNWL+pYboyrfmSivkhepP9qlO7tcXzn+9Vtgb2rsxEdq
zhEqRwvV4ptJDs6eLHYdIX+alkOxcO7M7sJAwa4Hjyo50w+m4EUa7M7hWVsSDELG3jfQpCG5I2Ca
Uznm2cePit/o9sjFWb8FvGDwW1mol5aVETUCI1zqljyq3x0kghR6PGtX+Ppa04mEv4VD04lNJbfm
dYHKquXboa4JMBhU6eNjkyqJNGuGUM9+y1Xv7jJLbAqHdLVjAM1Iv9vQwPh86iwQXbIJJgwHsrFn
K2ed6jlO5Erod6VSJmeUGOMP08/XpqJG4ve2u7KXzoRudf8FPVzO4HdR9hbH5O8zD2byPUU+ttCx
xikSpgMG97eYv7u0CxzqQg52vkF4TsNryJLQmhpXXYr2EOD2JaN7FmKwJwD/HULl6Nd7Tp7I/ror
ew7CzCdn2yHwNOMa1osw/T6IPzettcN2hIAZ4pUs6Xy98jAOZBjqCXeDT8uFBNzpX2E7cfqy7Zmp
lcRIiJJ6Gvb1NhsaTI/V9JxJn/OhF1Z7vx6R3gXbkwn16MuUbbDssi04gCzCKifgvPsWXqwOAV3z
QNSKe3P2TbhZiSvGEZkEH24QY7b7lPXGYJZwywTuKY7dqBwfhr9UlYJSqe6p9EP5EFUo89zGIUQH
sITvNRwfTeBMUCOYqdcGilLWHmJQjwsyuzpNANhYVuv8SuX4FvrLnc8DpF3tyqLDtoKSxwF1iSXl
GqsWJLMWQ99Ln70OFqNSppTo5EPDRwLr3a+pDPtFIEpoW0/ZiH3u6Nc+QDcn/+MwgYbpkOH+71fo
UIeziV7MhVQwf9q89km9Y8jDq/rJtAGaTPqfDhJ6TNZCZD5bG3sQ6Wh9wlcrxCnxXB/efXDOOR6i
2ftYYGIr8dOdZ1waDgzxU2fEg1otApL5yfnlzjzcbDLNNI1KuOeEdUFEEoEiahofCs17tFv+J9xg
9DVx+9x7/z+rV0i9dZj2l1Bl4TBnMlcR4e1yfmKECFj6dUtDKNbOKWCi3/ZmADRN0+6D8QjCICzX
ZsDOPi+Oe5h/dchjpcZrBSBiRFlkVXUW/NbIYtATwawT0T11U3eDgfIign4R9F9sE6/b3ugBFahH
Sz5RqFV9d4Rxh5SMUlZ3vLIjjZr+yp5XeNQFV9lSOk2Hzhx3SbfEA1momcGi5k+Vgmez8yWn6kN2
AGKd3haii4cmY15Uoa3L7NqN9NuDvVW2Up+ChkNzruAujxhhxF/czqsrH2ISzET5JFpP27ddrw29
Fu4s0I5Zj4DshDHpRM5dMx2kklMj/k6UQKuqc1ny9g0e+g8a+xTdhg5CZ+8UbjYcW50AWFuCD6FT
EiCeyVcczCIvvvHi++egqKEXdXzLCwQjD0KoIUUYdqJufwvMF71A4ovjzy6D8oRwmHDEQu+32rfQ
JqWtdZ7pgrx+bxZPf2mg6RSSkqXWYNf5O/JjxB30ycayzahNA3vHPogL84LeGmCBykXyPVell1Qr
Uf1b8PYvwtGdQSLkprwk4pyMbP0+gI+MuK7Gs5w5FbgQ58T1mep3wJ3Kw1WPEqYJBobur5qxoE8p
v82IxWW30G2252ex70N16/kNt9WzLVwWVoVsbXdsqtjkWZfAk1Qf++nNQq4atsHeOUs6W5u/nU6A
gBTnrhfUmSXso5AKxWA9lwvOGRgdNKsZrT9CiHRYYXRHqu39AuwI0hpwnv/NNsT+qwBubQBZkxx3
PSIh9oDObvG3uNvbwZ108ydldbaG0F7KWHWxdlnR00Zkzm9RDQXOYoadEyvQH/OkdSOzPSgYZ1P0
doQvcIgQ9VNWa7bbP1lvJ7kdDSG9Ftv3KgIb+RTKhtxW/Bu9V2oHcJJJ182Vsis+grHlZLU2l03i
7msVtYMoWGcrxfd+WGwT9wyRbpEHvSMVZiL7JabWDWpw4OQfpRc7eMeOT3HoeA3O+NoOqNuO9/7Y
0KvvqoUhW8ndgrSpFCKY665ooTmGf3rE+COPH7eAoJPN5b7QsNpHz+DoXI6AnxcPX/9i8TefkKpj
52oODElfqmFwGECeVP8g/YcoIOTvhqyUHQCUIy12rCKJkxzEwYZqOR/fG4dBOF4eH6VAY2ntx4OH
V2v6DmnjjysiDb15qpY84zC2gpVAc3+BfSu/Abn2vlpws9PuhzStFxtE44capa/PlzMmQ8pfTNhA
CuO/+BFwc4i1CeKibMu5gmn+aoPtDV93H1JYBE9GNJepMTpbnBnK8951oT1EmIXxLCK9JoHHU7A2
CKi5bAsJ8bJKTX6l6+B/bLkK46RhBn+7vF92B58tFbN3ifahHaXTiKFQDkEmr6F4BsSXiyZtdobF
KFjpk8gftLga9/34i6IM2etjDdotBapaOifVFWtUWQcd8OzN/FfVtNUr+LAgzSZGxNnlwtMRY5FX
+M2qQeMuQUgdAKmqplL/84ZDolsIHLPpCR5GQm9o401wuNJQp8J29hPvB5Sjl3XCfJk920ivmu8i
FlwvfM6YXWz5libo2EyGpnhX0PgFOUbiVNTeD6rSQwzX0WPCc4ibsMPPX8GwR4PSpPvGXiK0IOB2
sqQKQ6/tFU/PoQeoi2rUuVp0S3GHh+JtyvwJMjBaNn4BUbNvRLe/WtqC4ERS+DBmSqH7zLAukj2g
6lf1ZXMMQKYF5NAT6fTCqFXbJ2O8bg+M1m2/z8VbMXQP9JgXcF9dfxd0rlWcLDWt7u14F5nm/Csy
jxXsEIcGsLQXp6d4FAfcjQzmosuYwwPJ2FpVgHKpXTtGiAFmrdiHiCjFJ+cUs9hCnrkbQqT9mTJb
XtYwk104TEVN4PuTmPEwmkSiTvB3QSZd7skzHX8hjHFo+esnf1UiM3refPTElLWdTHzI2TazKuk+
5kHa4/ja1+hM0+zjbeAbuN29wYmOmiE/UAE29SQmq1oY7rcFQ8YKOlbVFL82DZnzSnXf56Lg0McG
x3Kj9lauuZXhUhWgqxq1fxrnrQkorbGcymTTm/wCENxcvOwf/qmm2MA6qj7XY2Qb9fyHUiJJwUI9
6PCczxZMqxNcrMphU8VcDGJPVrqAvdglgYN09fc7xoNuvtTeXHy/qDgZEJujF5fY3ZwQWjAPu7cl
fHvGlHPD8Q1smZTgGrPj4DNCnyvV0ki9U8mleM1s3qPSfCXeCToUlW3DgJ9wmZOmhIODFhNvtjKo
HuqxmrN2peKgPRj/nRRGH7wsWbYomR0Na4qFshibZi7qNnLjaPrrs1Ck3fCljy8lA1wKpxftx9Yy
ecmLAf3St0XonlOgt7PWwh3NnWGM7zO8SxwuSSJJBe/BvpgbUkl5RV62yESiWn9ySayjkB01MRaw
n0L3D9earwAqGpilNbdnHOSZs+AwanTa7x7sJi8udHhv9jyoGZaFC5ZRTvBVJEqpdem7HkvnfK2E
WH7s/0q7nSi3sFyjxtPPG+C/VQZRicYIDaawRFC7qVaN5qy7TVN+FBBqOfRur+/QxdmR5DK01sD5
liP7kiuihclSqyK5QhmPojm6NpMEjXy4tZ2i/noulZ6VWfZyrdEMJ8si+LSRnUCsvtQS97PNgXUN
JDP/ECPrgjMhrjYenNScUnvtXMtJatalx89XsdGyB7bhlSfuu2BuLJAPrTDr1SvY4my0667MG/MJ
+C/WO5cDDPPslDOrg6aob/9TWx3m/KRVAzB8zh/EUC+gGP+Npnzz9c/zVl81c3NSWIa4QGxOPDns
5tJQUliyQtjQz8iV4rUSQdPzLqt0DrHVf6Aj/iUmjDhlU81nxTwdNL+ekWuSur65e/nbyE0cSZKL
99OP0DhIblRmWgIDJug9xfeWwMVVSq/cvENJcWLv1kBJFqWqBUtwxW3ZBarNh3bcXO17ivfi+NXP
GY7cH13U9yQ5UGrRIo8xVYoCs+T3IDs0gnSvP25WFoFtKElKGNlfTQXG0javD0l22RMoWmwLTn8N
pHHbOY71yJOx79cwtOh5DIRIZJUtthK4pZQGaiJcDsCAg2nzGgPU/YPA8nOdZy6bBKLkjwTdW78n
Mbl/qlVUhEECorpTu2vKIfJtwoqboNEyHvbviiLfV9oOloRgiEKJuDnRljcthllqTiOn3A1clhlg
q/vTiJUvBLYvdSEpO4U0ESvYmJ/yC6u2tfGUi/O9QmSNeSp7Z4vLjRjL1A8VZ84vKUoCl9Fdny/R
E5S7DM5G2YG3QG7WvJJH4WFC6HFoiAC8Op7qyLQk/kyo14Nn3v8pGW9MO4PXr6ImUcFjjFmD/9oT
bK0H/MqtgbmGQHWU6yq7Q5w+ax37Osjsykyk7vI2iq7xIIF94PcwfAg1O1VKoc6oocQIp9KBZL6f
quVSKb01QN52KyPuPvYO2wu8TyacTpw+bml+Q5zC0kthszQ951d7c2wkBINCQBQ3tG5+ZJ2S2rnf
O27PVtGNN2aaq0lA6hwKMbsaSEziJdw7tMUyQEwPWNTJliTpf0YGsXEcxib81UyN4uqL/AUbX7os
+4U8eDsg8S+V88/jxY7AhZ8cIRK8UNAoCDMUVluDyhB+4bFgJh3+QmvTeojU/yUZqIToLGp+VdMa
YGNHunANV6xvR/Z+gZlZlw+vgXtdWw19evG7QZaUACHumZHZPwPU6jv3hCm7N4fPl7tLoBzBlH2f
uZiw5fxTGptjIFGkFs55V1gtRvNZAdXrKNqzlOca4SvH+91EfGD1LdJrC3G8YJ9QI31er8QaVZTg
B+o6aSu4hbo9FFGs89fCjAAEC39mG9N6BR1Pwr0wfqdEfSE0+oWFmpNjuxudIReCoEt/9FA+2avK
VJ6M0FM0XsgSW9w2yJyQl1rl2uD2UfmZReyrX1su6WjhiTycNfDqI0arXzyfbaReA+ji7nV2ntKa
7xYlJx/6ERDZXsVji1hfW1SsKf/1pBtDUtl2yWR1htpa/pQ1M0kDtXUGvIFEgkrPSIzGqKqIqDT/
05zgQdH6k5VPQTJm1ak34MRJJIcI2IfYPkWLslZ9Lq0oxeOmsv1W6Ta6Fx1NFAWgJThtiGYN/V7a
FEg3bpQr5Ey8FAuc/hjX45jkQoaGfnh8nLxjjYl9l8g90CoEOaVPekBdqggFXgelXgIRLU4Z4Nbl
nl5rPnfUPuIDZrxuk/VGjAh4eIVcrpcE8MzH7mRN34z0ZQK7gzJyLa4dMgIZ6BFC9SmevQ2IHfFo
YwvZz86P3+fkYHSV0tKZwNx2eaT6y8HIDKmi4hH7zrFr4YTJeCzv9m7rIaPyYE3yZcuqeUMjZDDt
UaSRqXVMzeH/kGUdyxQJvkatHhRiWqYNqm49uwbjE5iXW5MSUi0/iH2DxmhvYhjKwFphyCJchD27
lOb+V2CKZGTPaF//svkBLYFTyjZoQ6JiVx09q6XYr5mpXZf55SlyFJoTRefteoKQOP+ax2KAc0XG
minoWH0ylGArkpH9hx/Brmocr/ibcgfqy1J0JdFmItg0qW9xm9YR0Q2u71izw4Ql11LPIA1OLZja
f9+NbLPK1smhkINXfZuQe+8Vl6i4l1Jbrna/0pRTdqczz7H9NRyEAVdCXxCoGvyF2EiYYaBZWQN+
/PM/3+GgImhCBXmcmtE9jg9pi40/b84Qbdzj2BwCK/qZMrcs7kNkGntHIkljPgsOU+6c4pre2Nw6
LyJJRPn2o4/LRHgabkV1Cs2ys926KfJm3OjHH3tcxsCUSrRjxRnJEZwBfhwlZjEZ4W6End6wGvcI
OV95assIthiyFKFPX0dbojLY3w6oC8FR46dn8eGCgKun/f1+AvSNF0l0gkDg64qRE0FNUQkkvuH2
C2Y3l7kokaaqHmhco7EfxwTCDZc+3LENR55R+OVDP6h2xLffp2xIYawz6tull3nSZvZMaZ9MWBaf
hXAfjafnrYrRHogHvRWHBQGXqrHe5fYtgLjvdHpYqCtSpCj4GyosD4+zNLAqU5+Z2buDk2+B0fZ8
2nzQ3AvMZeCAWMwEnKTHmFKyoCewM/y181W4zN0l0cG85ldMw15tkoh0M0acDWoSBL5JvttBRdwY
Pa7djiFOlHfIRdsvrMuCiYBzQcSo5CXo/vkcYrc0Uk91Ssvxil/y4HcYT4FsTpgYCH52XnGCZ7Sb
FzmwqxKpAQQxTjgK5wTc+oKjysgwoewf8To5MvAhMfY0MupyNbQ0D1zlj2TbQKK+lcAksRgyJdio
M7v+xLOHVFR9jD/1cfYvWJWm+BFTrmNdXPtNoRXmh1WTnPQhjLiESH04VbufwfIrbVw5DitxplGi
JeAFvPmelyAOjSQU6kwzeqsFzGNbqSM3u3MC2ouE1W27gSUZUuA77LMtcx6etKYz+A8uTqmMBycQ
oDHZhlVangMfb4ab7ZI/vBffzjx3wP2qftdT2QE30yL4aj8n6HTDBrhT6icpNPwEVyVlbHOHieMZ
TfN6n4P+CVnNVQQPMVoJvauf4JQab95uwMpavkjw8XqgRpbVvuesILl7xa3ZQ0j0JlobbHYmbHDX
cFQ7KGwEwt7hzOPotnOPrSIVx4+iHJTWPsnrdp3yA1Il8J8+Du6nsSXjzKU+kGJIcmjZD11bQJHg
j5LCKmi3uosUeGZZfq2h0HIKW8zqTOMEKJFAK+KkPyAtcLVloHIdyjSKef0oFWTJxzU4QpCcf+cC
muqPrR5AAv+TLX+L6cr/Uu8QcGkZ5sJAlgysWZ0Kqo2IeSOVHhMurs5dcNZOR3ktvthKZa726HSc
XvrYo4i3t0LH2IkOHOitUTbcruahE19ZheurqX+ps8lXhCYHjzJ4dpue5/DidNYGOpyO4KcEd4pl
cHwLOSJ1diEChmGFTefA82Njata7q4PdLAuKK4oLOCuix7Jt+phc1yzF0abIB8BxoGAHIhh6Wzeo
VDGR+Pa3rluXziTd4hXe53aZpI/Xqj+HoAm2mx/K4lsWZBHrYSiUmnFyOsO4SNt/2piLlqXLBdzh
3k7Klf2XEcX8jHh0Dt3JeDVzsOh6yVNfBVWao5rRKcAYCfp7HZpgelayZo3GRmYBSVuLCPUP8AMM
KZOxtJC9NK9gPjuxzQ1XfHy92jZ6TKx+g76VUkLqMZ2Kxt0rQ3FNMdUrQrnpM9hmu+183pFbXfvA
fFJ5VihB/GgR3s1DDk8XEjMPCj9BPLhPJ5LSm1ZNsODsuoaqEP4lR+liY00QiY5Fez2ONI/a4rd5
T7Ll/VdjJFdusc4urm7Q9Vcm/TwdRqkn0ta7Ecj2NYb6HcPAQW9nLFj6v4YyHj7+klKfrxqdh0J/
kUxc2dEPvpbkbOOwqCTyYSPKTdrJFnfmq3iDReoCtQJ9DI03DzpUcXHsPu0hRsTaNPhEH1odCrOv
MYUAQwLBvTdj0U68k+H63XORJnX0rKtUykwVgGrxbdVV+a5FZ3vuMYAiYlDsHWNJ2ByW++1ubkg0
VWDhCnb3SfbY4drtmIl0d/pP3eqW2tFw6hQ6NI3Y5ZqLJBVbOZ/c26PeWdlIhv2Z4cfRyVs0cEyt
f17x3RsIr2CHaFOMxFLTCIjkgwc1PlrxvyXRhVyKqcWnTGHoSYQDLoHDMLWyzt88GDxRZrdEj+9o
0ynjnLUGu7hyiSGG80L+YhUV99L5GZUWlG9WDBTE/uDav3sanI2H1/uRioUsjwlV1chUpAUyS+0n
dqOe6LTpeLwweZfYsjzzF6Cj6i0K4Fhe/GR8DGIDJTQBgeOMA3WGKbkX9Qpk/ScA5LkzO/9amLwh
xLp9LBz9jfn7NhaP0Q/fTGaXq+36+MJEU1I4JmwemQz+8360xljQdfrNXIJURIjzLIE6Cgt7Lutd
kioH3Y2F+jptQcQYBQmX/PWvnwFnQWl2kaGHqDTz7gAovNC6p7HeyGhE6jTFgJzEf01NZha8DFkv
5Wzp4g5LMLMTl71Th1wupEt4nca/sNW7ymxECPwhfo4sYIsLTNAEECoIDelscjyVWCBhtuLVL8yd
l1One19bM9I206WRUHObprsXKOZxs1Jll20hmnydS2GpGxuIcZFSoYFiT/o/9mpa0V8vxUyScStk
qdCOD/pteGUiog1Z9Ap8bi0MqG7cBC66rK30KhCNpBKUpfyvRfR6bkVchCj0SHsaoJiwsfVRqnsx
9h4dv2tIzWTZ7mUbUcFEupSwymBPsb1zbAMd8EMj2NAO8F/coBds28DrBUHhPbzan+Gk6hcEjErO
DxW15Y29m9GbxyZsN1Qh6gzwzIOxi4jf+UbBinp5S2KtJYIXgogxNi5huTx8kAzS7jq9lhQCmL9d
HJ3buxmiHz/ov2HjGoyNgSXvvuXZAZbkGQzbtwXo4k4E8sffg9Pj+ukFayWZ6Hw1I/tAAkGXIZzz
xPBave/QooTbw9VWi19rjDMWECcE+SuO6pZPHYs5ZnoFFTAoUK2nHMhf9f8+A0sccu2TjRcpZm9Q
1VWWHsmz7qRTZk/UzaSNPu+iFw6EKbcWkrBMABKl/lAk+5cLkp1KsUUYS6X4I+bE37C/ASN2U1kK
c0LBxM3i6hicTd4yNTcPHff0YkkIOVhc3KFyLjSUcgNwcY5zTh1b+exhQ0I8ga7R4wOzQ9qNVE4P
c+Yl95WWvPBDXPa6JYYXgEp//hcSA6qRGNjLR2sR++m4DtZ372Vf4t6W7htiB+aV9ZnMjq2rQxQN
ySnCKrV878LvZ6Mof60FcXLqJ0N4rUYig7UuS1FCGBbwhj/64aakAVl/tB+WxmKaVbJrPM+EAJmG
oGpuhsmL8sOjswlMuJY7MS+6lYpOGBC0E+Hn1zsHHASH6FYpKBuOoMTI57szWIFKytylZYBWwTTx
+UTtnKmLlfk//U+2Ag4jIZ9mZHYM0wlEqLlOBiXUDMqOU3kqvzmWQUKdp2Tsm8VAmjSHWpaPJ7IF
a2s2u5JDx0Mi7GQMYQILJTreJsFVVuR7U/OD3AqjCGMJSdhZ9Qg33Kml+wi4YKMC6mnCVufs4ueH
4YPn8XB9GgPJRIUV64Z0uKBJIqOS0OWsRTxHOZyiqbKVRmpYDETWquSyFpFtzrhBHsSaC/DqbAuh
q175e8g6y/cxtf5ikXurxzXv0Yp45kIY/OFzFAuC84KvPnhBrQIJ/yihDmoJO7m3U/k6hgs/IR0V
DjKQcAKBig0SRaWjjxkx8enVq2rmcWtPxsgen8Ns2KABe+h4Q4frPWS4rJ1Gf8d2HHVMWg/A/aLH
QG/4UGvdSkQNNKSQjDY4cqUHZFeiI8JO1QNJV6bOF+3sGX12sXR4l1snHZRs+rUisTb3PhWvvpku
fo8KoS44C3UCxQmSgSp1gQnjTcDSMw8lou8dStOIUsrfdPV607hNU9xNjfQ3Yxc2J1SUN/JFjBhJ
Jx1Uf5nMjMFvwShOHv4g6NSLAflag9L+u+8EpXmG0oPRQTXoIGpJm/y/2ab+Ab3Wg+sFREXxwGDS
Cq/E5Mfg23cMwEkBsH1wu0V39A06sA310HhNek4pNmUECrpT6gwR+JSxUVH8mP03KiadKggqQNMb
bivILAyoYUfSX2+KY2Mvwqs5RvB1vQZkBjsBgFwm8rPBF+SldVgJwvMQ3hUPXfz2w20S9/pyXQRA
9GxNAsvneKJ7UXatTLx1/Py1xQCkNN5IATWaWBXprZdu/ZzJ93n+mR+FNZt7sJYkyg5NjzHtiA+i
+HWSwMen2r6S74/UODClaSiThGcQoxj3VJSB2Y1Tds6mscLB+7Ff+LrM8gB93zIIdQy6/3xtCUYK
LdInXSj6I39Qoj70qOOqH7Hai2yYOP3BxXBXshgDQfAuUB+7Bs/0wtJHbEapxVo2UF30QXDHE4uH
ySHyE7e0RldJoFIeUyYZZpzMM3VOalWOXJFeX9pxQOBxvFDlZLF1Gu7rltFfAso5LR0hmVJwmeJH
UhiOzsOt3EYroa57NEJFdwgKvaJ6dpd8lPtvcrEe2MXYoze200mYx05CCiHwYJ9v6sCo8OCshpoI
OJ1Cgho0HO5pIXlZR4NzoTHwCTsQLv/ai4UUUDAKnP3vh4+aOroD1mnHLguejfgb9aakJlDkFLxG
GC3Fs9FSyk4fcQzkmBuu/Rwe9TNa9LtWksSBK63CIvEfJGderOE5CpdHL8VZQ2dz8iVAsEugcr0f
DHEEt8moJuwG7WJeMpYebaABWInEdnL/CdPzqIbVZxe5SZxXxBGsXGH3Nlok9LTuXBBGRaETqAvP
lSJO3oH98Jz5/NVkAPAbjC+g2P4s37yIR/SJx/eVa854GokrQcYROtw3WPjbAkW6lYu1HgEW0917
6jIdKXL5/5QtQ9olBqJ+50R97LRr7DpwbEVCHAu73ex/ahpWKdInaZuFMHNEHDqCbnu12LD78fOj
Oyu0zeG4JVWAqOxh1GVYlH+uwChykC7dPYqrhdtu/vi9ESk8WEzls2y43CSHzFwxeqWVhzenAg+Q
fJ5pNjsgcKKuztyFg+OOfFildQkzfz4hKpM59u0bIMpY7aKrDPwWGQy9ubyauf9DC01ueXUloq5X
pDeFL1/Ew1Ehc6Zm6nR2CY0HZMvQB30TfN8AxH0OiFrioltgh776cc2BkIZSt6MvWbrkZVHGNdsZ
kjcPBNyGfVvcKqbbC8k2TzWRhTzk6Efh+iNmC0SB2D/ODWWtwJvf8E6xPjw03L0He1p0GkrVWw+j
lMtpXX6OePeFAUJqQMJ+XxMQJufSCRcYk9mKoC63MeXLAmHFhas5OV/aZsElTyE/h0bKl1QaS0ke
4bciorYnlSZLTaJ/RPYtSLaY+t0tW1oYVehL/SXr/wsBu66B5E38kX43/CDENWdJ7WpR+GukcLzb
yllnhUmfFaZhGVbjJV+Brs9Btj1jADSzQbaLuwxC9UMKRL1ltVMGaxsgsd/ZnTo2tvj/1tH6LRPQ
Y9j8Q6Tg+VkqwRJk7KDhJ7C4jY5a86wJU19NJ2wE6H/yTt3PC0Sbhb8gdbhM5M1CSvRgulObC6Ue
F2vbhCCxzLoIZbRxirhWSFc91FgIPFue2LYVcHmO9OiquCg/h9sy4TBou5NCwHR9tiaAK/pmV0/o
ZtiRqvXYeBvuV1sLRWwJSF1r4raI4XavbibigF6U3nsfa7l6q1e8LjmFWblGapVK1g8Meg30kAfQ
Di24XyFXYrjmytC4ww+DycnYbacdbxGsG04S9Hbo4IVAeW1OXe9Fzo7OuE6aPq5Ji3fWuCwPLgn1
dK1x6jD8y+tUpgvweTHBRDGPwy03Veb92UmSCc7AR0KqUU7jRKdc9SKWHsY6WcarrdjDwo/5uUHv
3y14DB+EGQUwQ1o/V3yqg8Cx5qB1EyNZBkUxGjNKAxaYBWLeIfmbuwujsoCfQMnkamp6LdBbDZrt
8ZyFr31ns7QaEFR82R8pqFh1FMWl8IHVnnBc4oJYCHkKq8rN22tGjWR3kL6EJXyjw7cS0qpv6FEl
CiVf8pnDHZHGQ+dFU6yi8BUH4JJWodm36UY0F6ltwLMs1u/fTOSPInraX5pekwftyNtCys02c95/
ho4BP1jMi1Ns9BTKhxIm1/eGzNXdSEn8Fn4SWF3BLht2Z70ZgrCeLhPrn1L7OikEsJu25kfdGhar
nLJ5UNcRI8R3C4T1vO0ByUVYp3nq+amEFjucIaRiALYMLrGfQijMMc73kblFlC3+U+zTFDRNm1ph
pAcdonEmL+DJi7SBiPEmFxoNWifXKhBgGrVpXvc4YtjTV7VfqRzwqkmdcQ8eYsZvAmU6V8Ys8jPv
Whf49bqrxrE+GV06KfyY1wFTL6MX5Tf5rWde32QU/0El1P4+IYCB/YEx7qwNlWQIrP0VWd/0Qixi
YssEbL2b03uHoh8Sj4Fh5qRaslRrgZajKH5+GtP6eNnP3bA1xHXGJCv4Iv1kr6kQnKFaHzggVIBH
wvZpsgG3aHGXtbpLFcOg1HIyJ9hzb5GAdLjSrhVaCjXzd8h9+H90KQnFp37cMgKWqbLqJa8cfvAF
iK/S4R4ekp22BO4QTHmGsSlx9u6Gu2iywCX1Vejp+eH7LCvx1ijlIQAAYnHcL7mXW+ev93VtCODp
Ialtqg3z+QFiuWNNfnBv9DEeIjCL9d1xDbWCAU9v3hrHn7t0sISEzDqHFdOEUSkIKmNa5nKh+Uj1
2B4b4UkhKTyUXswaG3RQoknPgtbq3hviI3HE8nZIRzxYatUUO3Bn6NBSqsBJ4xzCIGaeQ9np0d3O
BrKLtfcx1J8nU+S23A3/bfx0dEdUz07l2eDrEq8SiT+zzq5qNxiav5W802KK70Mi9AVUpdPm7EAE
ySp1VDYEUFw6bO7KzMe8//SWzEcfMj9HPYgRmm7OWN8zG0u7QLEGcyznDxEMTIgH5V1Ir637K4fw
tPpxhxkn48dNza6mF+OQ+98t3poQMjdrTWxmzDDjNRAKx3g6redd0J02WTJ/f9+uJBpLYaZtG103
9YnsW7dIGpdE4UfMqSvAaswL0jLFX+jEAnk0vMluzKxdVXhn18XmUdZnKUw/FUFm6GbbeQx6VnGt
gvYHgikaCbyNP1coaqwYia+u38vJpnYbxS88qH7786Kl4jwN4XiGvqTug2Hlv5NGVYNs/oW7y7C/
wJ677SLevFRuBV3beAdsRIMzAvRO7KQ4WHiXANl0LiAOpbTol6KtBDY64hHKNQH/D0ANGpIrBIqn
6yVxSKy9aOijoG+vQr+uLNZobTrAXB6yaZriu/UENX8ZY0YMAgTV8NQHKWCo05KaYSSl5WbQH4US
HHt0uxvWqdoWVI21qw4z3MfAsEjJbme6Gm4sIAOIet+wW7d7ZMYIEEtb31/h9AHCNOxZVTGK4BoJ
8Xo023Ge0Apg4X8Nq9atl9mYUGV/0FHqkeS8Wl+wwm7Zus5h2cQTQLLmSupAFKJCgdCGadoYt94X
5O3anq6ccDr2sKFxPWjFwrT3eRVs8sz7rYH9uIulaagcFq9031F9ggCjp28zPNXZSLVsvxS7GZay
aIJ/vjP/hM0FcpyOm9Rwa2YqcRXkBLSkq0+Lkst87hkhWDgiFFZcRCPf4VUhPeiCE9km3GMtwdqR
myrqdlRd3kka3T20ErFHURmG4ZMTAjLhN1hyd1/ej6mxVl509HX6cw3V10Uph7ZWGQ0HnwXFb2q3
BYyoZ/PmSxg08OqZR5slLoSAt1yEwFMQZ4VJbzdNLFTFRtr9vTQJTgXW7wZ0ewUpD2PxJ1eCEv2m
4rrZO9Vv9tufeHoRnTeB5SrgzkkElcPutgFzQfvy9/WWtvWfS9T987ty7+THkRmz3AvN1GXc9Zl6
bcdTMRbxkrKag93UzoLWRpmbEJOHFRRAXgxsK3nBvDzmnsIta+TKQNSwRCGhkDrHK8pn88muhcma
0f3bU5Aczqf7SYu7k2KfIXiG0Jfbs7hlHWIgtkOb0X4W1xLsU1EchCvwlTpqJZ0PbW5DGIoOoADa
E22e56rXNyL5CNJXsC1Ybo5fvG0ovgDPVYDhyJRE4Soo5w6rBozjV0RwvZbqTcFgP1FrCoskpy98
XyVGpjC8PTTiXqHXssXPYunZEIjiiL7c1JBWukTCxNyexZD5VciwgCg/ZaQ8/truzwBPguChvi4H
6Wfjk+GxVix/mgBCfZHRxV1ZXG/D12gv1GN+rs8WwzhSykWd7lfzqmzZ1k5c5NwKzn1xq5Dg0/GX
Na249wYvSvsaPEf5h/xH1iye1e9vhcAlQPt6WKQidR/NEUu/xyqN0f3mwZsQmjUrHgKA3DMdLxux
KwQ7ElNpsksQi3pqOGH2mCs63kCpuf2wv7PqFiyqjHhj7uVmum68GALWGuCTc2MVTaToETkmQOzM
vbVMCZvTibqPVayND5oM2nyHQgywp0J3X8WwJEhvnJaFaNMCuGZlcRnC44Qb1sLL6QGGi5v6zb5r
lJTZIHK3gRG+oD/usWrkFibQB1vsb0xzQFYjruyrt+lffwGN3WsIr0klT1DceSfeaytTfDjhFIV3
pnXiyIlShIzuRapzuvWQWz/w68mUZX12zXlqTqF3kjNoBlCQ31btgVt+La3N7nwTmni1VGNgD4oG
olg2x5x6CrKkgj9vb2I/GIyxhHZK3QyRVA0p6v9nnBY/+S63PHgeAcrxOkugQhWJPO6qq9tXXVJH
mukkZsP9LT0D5Up478GwdKXCyZa379JLjVLeatV6jYrECRXheQL6Armd2ciOs/xhUfN2FdKEGKUt
K6x9hsnlWugUp4wJswWW69H+IP43Ce31VMgHYNCSvR5p3PGpWa0tOn9vrmViRp64YFjf1rtdJotB
Rf2vgLmMX/bLMrlD9GWGjuYJKbIDUwC0YHtA4ZzDhdQOmmKQWSG2MNFdEvgItMFDfTI3jH3QbNV0
cnU50xr5/0a5gKss1M1ZOCkNLdxSITld9GGuRw05Cv6s2/XmIrRnjTkrlgILQofSkul3BSSj2xSK
NGwPQvEnOBEGDHCDR6x7kCYe74TJboDYHGrTQKVofb8kX0ShB4l+VYiMXKPUTJfH1zRfVi/g6o9E
3OJBdm2bnDKKhzCGn+wjyGFym5XKOvHeUWmkuCq5L9LJ6As4abEybn6tWSplSTLCZAo3cva46UTD
EvTP6S0Vj13yOXm03TnPNtvC1Btp9d/x8pE2y+gz5QGhEhza5SissumCXASQ6b8J+IHGAZJE7H6j
4fa6pyu8kvq6wb9r7bMO+Mdizki8rgg2aOQAYdTjgBvy9n/vurrPD/Y69vN02mdyqRXE94nhtzNt
OiX7KA3eXM8mE/Vh0PXyFE2Y4bMsCnuv9Wbz8NUWva8D5VhVEcrOcNcocLG/NUggd8lA8hQ2zds5
M+MFdJS9izq8iXdR3q3oGmsx8Mwjrbz6Ew9aovgkwIA6cxD6+3mq966YkcpCEnqV5xF5QEeLRk8G
eiCM8Hwlr6vHnGGRlqm1jb7BCOKCSsCKfrau9DlfZDioHEY1bjFy394cgWfdSXwsIQzn6TlP5ULO
SfI2/HMCj7NRssLVBJ+Wp/0IozNwDDvfySQxm5bPmb5wA9ETGARii4fIPXpYxxXl8xRfCJMH1/9q
uRJRDXaPavZowii43xxK1W3qWVVw/M66oMAxaSBUYhiS8H7Dx3h8uFej+5c7GVcSWnP8itZxuQJF
MibqukP6aiBnyJGXIHs2VojaTu9GA1Gw1r70noOA00XHvP1k3TD2EW02Z1RU2QORaOkBOWzMQwQe
LcN72sjI1Fh+OU2VPcEMc+DSuZ5jRfkSWZnuQUbUP6Eyja4pX9zyCkbDNPDtHLrUSXSkCVMoZAg7
Y+6akXtg0mj4c4njKn5qIHvOgzX11taRWKq/jwIwxn7x23JGC3cktVYKIhEkut5x15fwzP1sBMCr
jHI2LABZ60QAuWCevuTyUWFXEFsxq6WIgzEByulNUXVIERNsMpjAqo3q8yyGujt1LAbycyKpXTB9
zlhgIaKx9mzKyvlgsHisiCMwj/v4IY7Q6Oq62Y01aTaxU+BmNfNR72At5s2f0cEgBBVy4qJOb9Lo
5JMJGIKI8dGGoIBwqMIVxpbXI5YpX8+Er+W7zvgDi58kJPW4JCnOZpvGME8K1JHXKSZmjjxBTP7/
A7n3HtcFJWSPHHFuiCiTJLSxGptKZ2rIrVeglnldj3+7eQysslFtQ4/Sck+vUuMGVYsRf2I7PWve
qBW+7C3zttKBwCTQGbp77UZPHdnE5Bi92NT1CmKwxoM4bocz6z/vfVKhfk8+ZHJ6hRLrR6/OWsCq
kNUrS0BHfjaClW4QsiFAJy1lfgVKB5Vxc2wEQ0tGRLrnA0kleX4RreYnZEssTVsGcKlJQ1xihbWS
JC2doeiVdrqGTIy3l2O0SzZsseZZ3ZZ95LCMzZllvAzUApYLVgVjh2eVXV6gctCmbMYdT5f7wgD4
l08MnZQhoduDtW5ULrVbuG6fOFbY1r+gJUWWWs5/B0BluKeNsvUaqgvS+R4TAHUPMfDkEfTK2Dqk
D4k0bskIYY7Yrw5Sc+HVzu92r7roUFZSYB4Uc3zrjMM8QYE6Bz7QwBB+I+pSX6XXt6TpOT/cDcM/
EULyoBB67yOp1yyRCfj3s9v0S8nZt6Y0WwqjoIfHt4IRJ/oRNX2L/nB8zxVTz2Z9zFqalT2T3ywz
gcfAX4IziO23SVCvWcWWApmrtwugLylyBoYxvp6kQd1ZM2TlL509rltvpIt8HuYHV00c1SUmKe4O
wLDpg9FRAEZbc3HyRJRo6VR3OGOS0iJN1gY21BrZZOPRWebACvWGd7Vf9PByc31/xZf6iWqg9XhW
71sJ/P5s6Xocf2ykbxMahXtHK5slHDWWFnYR0KIRvr7b1sS6BYM/aFoZJeq0rhzyF+0iZ50b0c6k
zTpHDIVyROei2zan9g1SxP2xEMPsioSqcnQ0iLcZ02eTJderkyqvoy0W1+Rzr3N7jJCGIoYb79E9
VayC3Xx/NSUUQGsoz9k6LajY40QbkObQu627O5MMexr+cBvX6msGphj4j43rha2AbbDJ9M1PQ7vh
jmGy/2cuH6cZrcJEa2IXL1U7MlAv9YXacvfP3IIhhp7PHKi3E1BYWp0a9VuJ9VoVQY+qlzD4DD6p
LC6bOYRspLVel3qZSENqHWR8pWYtMaDj5eA8juIs+qlQJVeunhrLLBPlw6q64miQcDfaPAn9efDL
d71cAbhaSgd6zHjMdBCwvAY2La2785yxln6nkG2wBFN9Wg8jMKdJayYU+cAOlmREWY4UudCg/EvV
bZjnrSvSf3drLzQFEfTfuyOnJWbSOWGEH93gPrXFGz2VtLHrPyTNrRDJotabftTq2cMpjjKUdV2B
BZzxVVyscsZcuTqv3IosUhnCwZ0YdYJz4F+VWKpgSyBQOSYC88z1Jf62nx7dfcWhZSiIAnfhhV/U
ih601s01kYSZnTpijVFTCzSs9tEl1vYFIhbv1aL0EWxcwioDZVURtlaqFarf3lQHZcrE2iHqCjia
PFlRwKlN5H5fbAiHCfES4fFZihS0mzBqPn9a9EzXZaezYcVhxw33hRxjqGAmhx9Qe3wTdAZNDwId
Wbw4OtcubCK4Aj0fTkNrUg1CTfLqGekRvgbakX0NYlZr0Xf9bilT4njPTzIsR02Y3I50sCsInWO5
TakT1FpmiPCmD0lI+rfqUtxxWyqiT+BCqlDMsWRvki/D6jt25ph6noGd1bccGag+OBqbLJOGRlTn
YVwjvITbHH+kOZHoJyup8+d6gJRNqGdnuaz6DDNqx6hUi14ftEaxAtFE6Ftz72Di9vhCvBVJNiAx
k5Y3RVGcoO4ehpPyTNY9kso/Ehy+jUMUc9NkZO/DIG4iVJKDLhQuiVlaa5Pylf7hT8v8c4Fb5dgH
clMjTP/EkSJoIrAmex1ZowxWbtolKNkXS4VAa6OkB5jjFGCp0D/7xITqP5g+SOsYaCI1s786Ljug
8EqoQX/H/OKRuTIbezjNQ9keSszFkIlzqHLazY4lLX1vMOKODQCGPTJu9/mgAUX14r3+oQepWbil
n3jspOM7X93uB5HKijEjS/Uno2rKIRmhOxAUlsy3H1Zfr4WKXGcyOaZEhvptBPkwLfEnsvIPo3Vo
6ramFZhSo3OjFE74w4aO/T25AB0zUonvHd3H8d4Y4cLEsqzkOwX0mWjpJwfucsDDlYRxJiiu4RWU
ZK5ZLZf3aUgV1BGuxVTHNeOzyyw+gf/se5X8Cx0kJOfu6x5xq3EbEiyGWMdUgZM38rbIuiK+LQmP
kc5jV31C0oSn6C51JMiACX5XLSCpTiV00A5Y+PQ4z390FFOgYdIF84F0m8aBRHSjZIxUsuTrbyH2
DiJXtU0iPglG7qnXkdZAzVzE+3kwo1Y0wI6NsA41muVgQXgJiRNshB7uVF86L0Klmigb0YMAR7CG
xvwpkoh7WtwgE86f2ptfK+qala7a1Oq+GSnXZA+IvIOgztpCTUpNJ+B2CDvCLAfaPsLtl2s+70bo
vi0FFZ4gA7/j9d2Q4Q539kTpezMYJOrfd2quUhCDA5hxqLI/QPLcfTSOnMNW8t0cX0mJSUXz/9Mp
RaBGo7VfBCKXc9mdAIx7CLKap6Y95cGt8vbU1y0cxpSx4lSslln+YQ4dYS67PE0jPICxBYUlEFrg
+fYnmCV/GqqcGFYPBKZeOzseez3ZFLZeh1XV8YgX3vJhXQfOImuRQ0Jl7rIbAJ9cGVOBuIZVHsX7
1W4NhvDhUXPwxZqA7UITjv4tiTm2VDXwtEl9jEXLf3227TLqr/4JNKEQXwfVDQbrJ9Wpe5yJQqOq
0GWZrTEPEON6aSmoh/slcQ7YpsFpFohJ3t0G1jqNhyepXS8A8RSEF4KxX2RyuMpQoc+isctw8MVU
tzeJQJXd+mtwLN3l0vFZoP7FehekeRLWnnh+k5Tm+4tpggEKj6gIEHlWp1i3Mr4iLVdqN7Iay56K
PGz69JiW4ta3anY+myTtnaS/rWUXh71v9euMRMuUdnLCOdcusy9mXyWjlxivY3+SSV697qm9dlGp
Nazt3B3rKvLMg2sXM7yioGE/4C570CiFDZY1DgXRkYJID3iYq+Ne0wXYyQWdAqs5uzplCZpoKIi7
tTd4ss2RbsiU750teise8osrGo8qGHQDrk9Ovhh74Gvxo2/zQeZ45Ri8/mL3LxMU3ypWPK270BP+
uhB6kvnyO+zWJQlRuBv0ObeWQXu11zrWCybc1+F4XidEYU4Uj7OYM+xACE0CKJLhSEBkdBYo/DHc
4VuJ7PS1WzWWNAVkeUu5LDeWVwg6WJrw2s7Ta9rZoPyCPne8I3ffoAM8THuwRLQ5WHO6t/rraxOR
34wUSON8cBbMYfhwebsx1JXYZ0ANqOSGCgQfSn1jHo1tNaNwuef9lGbR5vWpgoZxEq8joiYGD2ci
5h6MU6bQAd9AFCNQqLzeqeCSIkkL278i1jNTo/iisQUQAYVcFCM3E6Jvf+EB9tJX5ZIdl6X5EQvO
eMiJmGRv6DVw9cA/lSkywlpui37ipav7LU8t41XNQYunhorOHfGKPl1R4d0cnd4k5Lw7+G+RrHx7
wdm9hJVVeWLkyxfi3ssVj+We1JcsVchZGWV9CZFxe6VihDPpkUZ2E+sBD9bgB9fF3IQ8Zpo11K2d
omUuGgbV6iAY9gMv80u/Lqm/yYbsSb9S6xMN5tiwcSuQq9wIL8juW0du5Wso8tuXHBHcPphMzR5u
DjxW1018F5K7e+e4mI4wSR23rdf8PSfRoQRMCK0PkV6ljQcg9bAU9UjlmG2a/9QmBkiC6NhMiknd
ecfn6Ill11QrjC0aOTLPcTBH07zb7FzDQAmmP9OhM0qc/pX7IZwTqAcKhNp1qw583oulNbc4zWFG
r0wmbCfsSNeKrjn42J80NU/urtljhEdngqgwZGZfUoN6xOQwwpnDMwogvtGs3EZ7K8WGVeWdJayb
xwHlZwoejPAtJBiFq2vk7RZpVKMo4ZCVl9XrXtcCxs6QihfMQfSTHIjI5c0sxtYrzxoQnCF9UQps
g1f6WVqJIsBk/qFC2EprphCz7Bz59BnG1fT9FyClKWaitMSiftjReFUcr8NRTYyOFQGp43akFxsn
9PpnQZs9TqXqGLlrB3ElO0QyNSgRk+1SHAfpzparOwBS9ItweY37s3DpuUJeeDvCmcYaW9QKpeYv
qpawPls2YRch/WgeFBHi8IGtstdlvNekSnkupfLrlC/0WGcTw4Z9rAh1KCuPXQbEQPAGhgbwSFaV
Fix+kmhMfxZt1mNkqZcON/Jz2YEwmSGZl6Ld6zWggFYlr3NCPbx2pUnSK0M2G2H3mBRtfge/mDYR
5RjgojO9QB5MGRN8UjRaaK5xMrRxsyijC+ATkGnYPeo0LbHbXb8uIOfRyh/OZPCLtopLaiy1VbuC
0AfaxiWRP/pbeEWCo21WCg/IbJle6A+VHycBP1CgSRGYpftfyYh2YhnRkr72hQdXXOlfZXorMx6a
Tl6crfgvKVKb4zy1IuUSsi7TKOVfLaBnOBMrBRfEK8r25X0jIYTtNvJZerEupTVtD9Q74vYfVWuK
oSWNGs/ccCEXgmBfYjYpvl19Bh3fpf/8N2it5C9uaXHBti9scTdB8CjsJZoYGCuxbZhhXiwy/xYb
njdFv1wxX0R0ao4fcvzPIx7IoorkvttBJOnurMlcOPbHMpWfdPmTUX0GDt7HWD0I6d13P+JWykKV
wuuqiN0FLKFdL3NT2lyfsXxhnsjhoAnbog2cAskRw9oCHDINOjohMlf5O2scSaWcNZ9UVUUk5HXx
Echgok3jwBqSB/v1g5vEdUri7+lAeGCpUa8SAyEjSNSbRvHyBzSS9xaHHLXwCgpf9ISbRPT6Xi9I
Kp34eqRupYBwQgPwtYdaL7kBWKn3Nn3RKSt9Xbf3tnlOw/LESBkWFAJu32X9XEVfzw9my0uvAj+3
kq47uyHC6Pm3sI5/AJLwHh5f1nzRP/wnuGdWbELGtFEPfbAZ5gmk0KL6+w0reQHuvK4K/g4/Z8ny
dYOCx+LyUdatWD3av2A6DfiqaEe7D2K7vl/AJZxG6PYFUDZspXd0vstqMMqNrNSJsJFOcNrI2KgN
KQdhWDf29a+htV5yTzMw0gwfq7u4It2R0jwNSXfWvh2O9s0vq4sGyG43umVVtB+nOwpFbq3cTXaF
lcs3+m6In9MGWivuHonMRSZSNLpgIdH49pfv/OeqvjxYarSWPtGTmUYyZ2tIajTv+cVmja2mSavD
XD8kFxVjUGeDTy9yi49JkbLhds3g7bf43/IrwwaHOeXYbA5DdiayaVz0EB93zeeRRhfOBJ383/Xe
efcjkGmGwV/fA7Ed43EpRfM4zx782qpdgecRhAWsAEzYd7mwnzBI6hRjOe6Jy7x5erYCf0cp9MVn
Z6H7PGWAlo9GS2VdAMmtMu8yTwL63i9NiSfz9TwmeZvvWgyXvWNKH2h8TdpOQXWVuQ0Z8fKKDqOp
AqOcCtDVxc8LGTFX4ciPBeEEszlgYRT3gw0+lFG3nWZRYFvXbGholb6Z0oEE0spmpNRlGEPi12QE
wtjMsSSqdvAltbdjLdzJHFmfbuWrwA+0CUU07cA6CMBoyxQpzAvuqHeKf0c4w/ace0+OifGDHIAl
Mc65UZjodrDi5+o2qCmBihIRVqFPLcR7hb9vJ1fc7IGrjoux55MO0/eQqLCxvz2COD9gIqWgKClD
q6FhWwX55pAN7zgxRumJxxFy7vAgGHRRIjhgfsWgI4Lli6vFVehJxyUsXIisMLRDNPSUFJb/z2Yy
DxYkSu7+9pMCKq2jY0Jl5aT9WGdpela0GowiLEmPLEQOifELpPyJAhrC2dSidXMVsoZyslsmvR+q
HZub56PTDxzLOCBcPDymSHL+5EH1ErLzwzaqle14+Rb9yavMfDMo5zyCZeb6L4JUZgtlRxdyu1MP
yPIG0y9m5vXjEPj3vsSffjbih7SrLZ52LcUNGluhiM5nlpzy4lyKdYsrJokHpe28/cRPJYxhTUrt
Jw9R5RyAawO6ZtyTvygIpvT77jOZbSDP2sfnHhmpBNNfkqALosk+Z3fj/Spy4GcqBLl/qAKyifIw
Llv+3IHBudh6vW63BenKdxRG87toHLS1HuwVigXVb9STsTRbwPdLZFAhrZafx9FzV47zUvH51svQ
bPvTyqabfop4XXvyMGvT26Q5h4jLKmZt/hbh7fayJoBsY3nUXY/UO+QziUMXk5k64+ijur4gJFEy
SqVAWqfvg9JKzHcW2zlyGtcxvF22nD4qJjZQJgsDFH8NJxoL8jZqc/17fEFI52ulCH4oRDngpB2w
6nluRM75LD+I2ocFMMbV4kynjYbuZndEaE3T5n06HvxEjv0XOaC/vIBXWLyOT4SIUqPpCUBmOVSi
v0aDSafkaEpQzI9lM9bjyoEpiZ87AlHVy47ysxtRCnR4pF0Ixj629I55EkLZMRIDENP5puQC4P9A
sPcKlohKBwOF8X8Y1zQzMdFkI5Pvp+plRCJIZTYoT/acJO+2YN1JUuJwLiCvC9uSRggj0frEcKQ4
e/RanH1XWnz0KQ79OUgVtYH1/bG3j9Fd9+gsUS2ZgP3PXv+59w6rVuFCyorbj1nVODiAuaV/5aXH
CG/gzZQYr9uoGvMbYvCuRMIPhqO7Jg+xZi6++fmZT7hVoTxupJBuNjbV6nsANcXmtLksVI/VN5OC
rxdaCzU0yEa6VvGhzgEFdgaTtA90Q0in+ZIsUR3ZEG/wY8XAxv2RfDSWapg62cBWRyEUaWbEXax+
AvUMFzY4ZNoRlIOWfUTIVLIb8rACayoQDxD5ALIbUhEwDu7ldiahZTfdMvBFRm6RxEzzhbeRCvAT
M34MgWsoEuAGqX/BJ3cN7tfUaM8/d/uJ232GCtrx+H+u0EcLRKbHA8pNj8n2HHgMpJkcbBDahBxp
yygtU0iK4gV3oAXXiD2Ez2zIShdGygkuWsFrHl5rZOFNj03LeTVrTcMgg7UirweaIMpMaUW8qwlU
Hibq4x5PbR7yEQy47LjzuvD9RIt3axhpvVWZ3EmoSTHgpibe+Sw3ESpJZ2ieTXZ6gVBTGBCMPQMl
ioy6O6ezIgo5hcqQft/bzu85Gqsi5LAhfIjfUEjJtb7FbvidgsgD+ZtQTkvl7HF5UUiV7ffnHb8Z
N7f0e6bncRGxx5XpuYJUawnMu5kx9uPn1irft2S+LbKjRCsHmzRVsQ2mLwDFtAnTJ6Ro0DobmJf+
0dXPomezvOHiI9xkZeNixWRK4kjYVqAiAq4AAsB0TsL2Uri1XaD80UDbnV8TB5u5Dc9/ybOQebz9
z6QU9NTK9lOpYseTgbjlsRKu5D8InU2AtUEN/6Ed2HqA0+WPM6RLWpWDHTD+gh6jMTnOswIY/1wd
DzXgnZPlAkDf5amq3yotmhB5c5IH3WMYpvIGfdem3CybG1LfFJo697rdQ9trihC2/b437MJN7ieT
OS15duFNaSTO/V82Q2igNRhe1dYweZf3qLBqMA2mIl/kM2+CKO5alFAjxGqQW73+bY6gtN/HS6i/
r+uOd1e0t6XE13v/aMp8p9F1sJqA6LQoW+NYgh1URWR9Hn+6ugNHaej7jvxbUQDV0qe4dXQVWBQb
6zrOwoOJ9AQKhlCXA85Pm8ykwmy50KW3ORrfZfdO4eCEJzAy5JBjPivumkycIRLcEptPJLH8We0s
/C0YyL+yhXmzJJipOVU5wwC7E8fSgKk/4eAAgVkE9NdzD9vfJf8GpHH1ikGL/7VCEDI2m/28KM2x
XwualXnwMwNuoKFE9iqkHNbx+JRnDa9ThT/YZLpi0+oGIc+9Q5IY55/8uMHvoK4doDYXNcB2c5Dw
g2NpYix8X9C7zWTG4oJRqNA5KciuZ7jw1SoIzUzUwVpoleWbYUOAiiGzYDVH90iZ1nLaH8QXBGv0
ttwZ2OSYKPzJq7D2PpE+AIaInvGef6zEEsJCKFym4VLePsxUIV0rKjvUtsI17xuNGfxPro+NlqHL
155QE3abkLKgyIlsnaHsdFbPp+mkpl9g0jka6mj7FSWw8CRnFZq2lM98aXEMOp1vo5DrdOZometu
nZfBw4GU+S+owqPvZ7YWqxDY+Is9hQhAmaXf29UnQmWjAsaELxQFucZTRn3iGrFZiMRw4At/KTAm
jndncGuFPccsVYTZO2VvaH68KCoWpgVnrwmmqkt/amviSids4MmhV+WNZqzJlkj0Dnlb9ToKrGe/
Fwf2dYaqOV4gaXtCqybzjcmFde8zQUK2/wJdiIGkw6/VzT49Fd8ps8O3DaAjz7YhVNjGrDyDgdTS
QYx7PW0Fe5vqLyfClGCbxeEl9yeLJq/kuQljgFQ5lsfTrACr56qxf29aHUr58DpsqN0sZTKzrFAw
4SpbrTfwgdpJl2rlGIiXZ7oYm6cwBpxvOWf+gXco69rO1XjAY9WFytBKfIFa7reSFSXxZB79mhEo
c+2xoVr/rRYUqMnkrY6wK3XlyK3qpVLDG7C7yw+OV2nEPL4BufP3SR8hBrXnMjxgDSjkF3VcmWXO
yHzHeGRVZJ5nhP95vVN16ZeGrPlkT5afWvJSuHdqH1Pyrg7wzj6MT6WxnmR+tgyJHeyPfdDlzanN
Zf/a631a82rAWrqHamlDW3wWmebsTMZE/G15Pgphyu0iXciAZGr+Z8nTAHTybvmNv/VJbCxLD0WH
jmWcZ5ubqrO0EsOtdOeLiGY1qQ2HOSD8S+wjmobLRxRna1oVClyUdBU1A+V+xQVm9qqpvug9Z9qs
ADBV8CxgNnEgoTMB54xIIDUDYXKYDvX+Bvd/T0vQame77Mob+Yca42YNC/USrmeYJwA+XR5OoXdm
4XRCwfuD4iAx+fL2d/q6Fd/G7i7UjBJJvafOq8CH1FsSy4TgVB15YA4/9k9ff0iL3k64i/kAnXzv
tn+UbW9cOGcZvk0EINmj5UAyvLgISy1vQhQKhWUS7n/AQsgU8v5zPcClglMHw6ZIBtTF9A4/vmCg
6F/TUOHFZi9r8te0D2DNI1+Ag/M9uJMa+O66B2vWZj1bHH+G9Aw6AHYIQmAWlsS+RSUUjnfgNtjC
RokxKLm61zShS3lNU2JnpQuPp4gUny8u9jkrqDgYr167pPWf6UQP7AXPz4/4i0hdW3qr2XxkDhbP
IBCZv0EQFW+5wAL4RPwBzLlB++hXh1edUQaUpThg51I7h/FLiDq5uRfwrhSDxQcmOfO0XKRz1DaP
6vuwAYeKOhWOd/1fBDMiWOsFQuxATqwddJE9axBvEvMVctV+loy55b/A4FDKC0S4MRfsoZw/wJTA
7hfJmug9B7x8l2nMaNTIGVmEFSclrhilAk8/wCqK4EzZiGtp6/nvTeQJxlS1MumzEyiUcVl9/g/9
t/wRpbc/nzOuXIPJS4JJjqG38JoG5ud1Fog+8tOOIA7qZ/8JllV6YJZfC1LhytJeYQLXVPoVA2zw
YXUk+tHrB1BAMXA/mHE5YB1mi2nRJ7BwgUfaYEkKr+htXc+mv38TfxQ5CREGZKwqz0P9rVfsuqP2
P1RA+E+igXZnsJPkeA071INOzb1IKR7ETSwMhO9wR9CEyxDqqsREYwR21Xm0I/zH7UuoO6t7DeRy
Dpox+4SZLIIaD+uMr9uF+S0f7qTQf0/JUjN5FNlQAOTBUsBznxV7toAfXj/uwy3fe8J39vowBBox
7gSUhTmKq4fFhomGEfV0FNpLFMt19TjOtXEwJTdzm3LY+Aj+Z9mwDxP4RKNC9Etku6MYqb+BDpaT
rFhIkJpug2FMNLDgqZ8EIroirfZ+XQOZ57rwvaqmumrvBaKlnpXIbQtdQruaSTi3cqBeWzqw9VCV
dcPMhbyW6ECxUM53rDl8+POpZ32bNLuWzD5Ar6V2kSPQ4tI47KLeRju5Vc54YdNOh0Jf9pQEJasY
d+8pIB0bGX13450NWK+RCYXe1UVb+5znJPoXOGb7gcexdR4CUrhJvb7n+RdxJERqhmemw3VLEADG
XxMw4lX3qooXwRH6gQtVgIZPbAmEcze4inUlQggsJWUiRL3tV1WPHDxbYGAQ56mQM3NSGdJpBAoo
nYGOmCIOoPPAfIXfMvnjdamGeaaZc6CIQzprDL/8pvYPlONfLUy9UG+h6k8gjmuVYP7fQFEke/l5
V9PDDbPQGA665deXnurpMqiB6d5wVQ9jbXTnvccU7HEisSV7EhS+lvPY2RQoq2hux0GYdeWIuOO0
mRm3KoDlwTN3wvji3PBfZfgHjYBxLoqA9716Nm0foxvL4wZRP7ads5tNcNwnFN5VYOvrNfURuuiI
yHF7GvNbPdy8cXljxCu+6aYrp5qvHN9+Wqu03aWwmb/e7G6ZaShqeRM/oyCVyJiNfzLHfzmODTrm
MqCtRgHjSE+vp/XZWrQAFXrURoKg6/IJvYxR0LAdUtCDfYLKh4c/cQ0dqQKNwCnFHIM01PfcOSsx
Cvx3MY4HhDN0wn7/ZDuMznti3FEv6TFDtQsrakqpK7NrODES1/NZfHRt2IGAkPTJs4n1Afkq638A
JLdP7ouDWYJl6ANuVJY2qQGLo/u1zWXoS6p1hWvPQHDSFgWnsyjeecTEXgErHZmHr7FC7Z77I/Dc
rGOQbK+eyiGqJvOQvKzcAh6CW+kfFSXwPbUsc+nb+1x+5iOKpdDro7lbR9Ihu7bGrk8AI1a1DpoR
NIx4j56Gv2r7T0UT1KXSzIJk1GUl28nYCuUfZQ9zoc7RBOf53JzLqhbm2VIvfakUvVKAfWXglJ/c
paIxUNYd+19+uIlfH1gZXAYNyZrBYqP+xZ5S+YHiirlJQeq0efugjho/C2wO3Fj/dBC1tW8nAR39
CTn69FOmQfIb/Y03gj8u6X9RB58UGoA1DI6kYw2andN/ppa2EdV2925+Qy5EUpNbIk98YMXIsM24
o0Nt30eIzO+pxfv48QfoiZf94SutC2ATBnSRKPqyXUX0DgLpCSCcuNtpIHV8EjCfkNSVIS0Jp1Xe
MYzYPL6R3DjWSqCqcnK8TE0qEvBl2prTcwuDjCeXvInpaxJoRaR+BC/CU2uVdWH0YV7o0c/wgwCQ
u2Z8x4yHOmcbaKwcM+hhS7VykMWhqo9cPqgGA1LW9tZ/+/bUKmgYLiAtfU+5KWxM2mIYWmZVGJ9V
JwtyaPRyTllodOmjvOJVWJeH7tLzxBatt0mOF9G3b8+SsRk1SX/+0azVVBFSzHbAvjsfa7JJL+ZN
IninA34Ud0DDYbuwhpTHuSTCywYpMBDuJcKTToVrWhwsbcM/CAruvIxJ3Z3yIk6qbVKBXVZ9wJCi
V9BEnfHU8XfSkiTs2curf9/9BIndgTqdb9iaj7phqvq00kn6bpaFUmrr5hBKPvy2x8nn39zdacCq
2BZzZhKO6Ojj4kjMFeZ2HU+ZFrz8I3atce8NY+2Hj3PuvypGmr4aqL9ZIBP0saJMjnEAApwLlhxK
PDgta6RsjNgSJ54z1EghYSVtXY+XkzDUkgZ5Pjfaa+a6UbH3RZobR26zDc8A3naipqKOKUsUCMgQ
NsgNSWfypBCbAwoj92Y7XQy67iDgKWjDyvB8r5dd4URyCEjM/OARjfVghl+9vjdD5b0k3jGRrYQV
NOSinU45AVSJoJcA6riLs/w7ykDkGqjq4esk2RENKh7MdeSstLwNygCA35iwBXRtWW6E+2RxJFES
JNlrQ8MIou5cge2jVlipD36g+DzHdGE37xicOFA4Hf8TbEPt43cZlAx9T1e0b7jUdKVWFz8D+wN3
Zxn8uSwFedfOTKaLXU3nU3d3B1BOjKKRXhUUxrzfzLuCOp4k5uPmeAifBwWE5olLRu5/U6omDOBI
k/vK3zxUy0Xp5lhnlDmuJ/X/0Jc5mTysGpOPSPgrzpAZc1ljjZ7pjDIMtshTWhjBzOaI3HHIx2vq
zR4bexMXVVsqZaK8/qDuFWNPIcsBJNl7CReQW1MNnPDkLTsSt22xN23liPzL+Afg17RX/GxhFdcv
m9rBED0SHWO8VgY2f2qnr5mesCKrf5ToQQaFd8m1M3BlMEH4AU5P1AcbameHe5LvHXNGQTfFVV7G
vChyc0KKw1bRuzgxhvFKpOKT1e4bPaj89GqYb5VTcVVB5L+SdmenKxMZ1hPO4eP+DBAgsIQm3lAA
cnpVRIbMvvWzAvcvhcvcLaXPrzmQ7d3SAHkg05UQqT78t3WcF2C3pvkMBzSPrfAndLGNOh1OXRG8
RYyyov7we6U5XSbwO3Rn5GIukzuDXiLr2G6xRgY+DjAo9H3OpudnsnKbHuPIGOAoIloGFKKfm6ss
d31Ef8UloWWbIKndxdgTbcj1GdpJ8LVWXTO/Y/USTEUTfQYC5PCphcRhCzBZE5RvcNEkOQWL9G4v
HNBzVv5te084rDzZOfk7uKealZhcgRap69L/ggtQuZfCNPcs1tnHHahWHhjW9cXyqEiaipyjW3jY
ijztzEysuvtQtw7Ug01yMA65ynKMhff7OaY5etA33t0rwoh8HuGVkjFFKKbfFiboD9mEderrUu8q
iYRHjKA5KvAO4+wz+7JpiamJ5663AMTisN7VyOxNRSS+D4ke4DE7+EPlKw+iVCcoWBzfgCyP84G5
/1en0nEw+IW+YbwhGZgRISH2lfDWxr+miaFEE99mQSaEH0KXbMcc8kPfdL6eP/WiRxD2JyFecKsj
xf0MI6LtBlFWnnyEIKTIH8XglJAQD65dSn9yEhna6nyrFDtkjRt03RvZQhN+k1cxk/MBcLkZZlet
X29d2TKJQ00Zin88xf3tUT3ckriWpM7J5ODJzmmRLS+9ep9C4nkwbdikUWDF2LNthhGHX6bdfQHh
P/5qC8afFJxJy4/w1OVb9fYGQTeLnrPLWVoqNdDxaKN3TicXM0F7L7vCY2xIS/sZN+y0NKkBD2jx
IxsDF5sH+4XCzhanmNmz4zUNqQjr0AqHBCQgE3UjnBE43MOshFu9LtkyapQBwtYO8K3FdesblcQT
NBlBrPWekSq15qvKGbzKh0GdmjfLZG+amoVVGOlg7xuF3X1ixwKlPaYBgdemTUNlHlPQI0+2l97u
sdNFWGJAmW4fygSXPMoGeuZPwBHX2B1XHfcfOTeShHUD0Y5fWF+xIL4vOuW9EOqlGg3hpgeQ+1fA
R8eTTVhLcmee2PVDzq53XwgbxZHG6/EqO/i4JqBE5a3xs620S7CgO/6gIAdTg1+x8kvmAD3Ha83s
YX25VJpCszrSba85mvrE7mhgyeIQ8c4FM0KWmnlvsHzHQMOZQjVhMTXbBYNga2OFhlOG+DAsgymo
8Ml2JqQCFAJP1BR10A8lK77YoXr9uY/o0KhcVEoXN68fylXIdmmL/MZiGGZdbLiEkD6J/TNNIESp
GKgMcyp8WVqj5c62UU7UyXAmLgjcO2J2WUTtBl8XPtAgRrRDDy/UGP7U4uDl4Bavq9VxZWM7j/2K
6IAenA/ErthX/H/tpNe7bbzozxi41CccOnqDWc+6Oaso1WSravNZwbolmGybCbGaV+k5LLsNyEff
WlYwZNQvKqueWGPm3iXFjgsY42s+jj+rHE+mBd7harX95HL/fNrdsqEg7VSXr0mO6EW1zJlnazJk
8R7onobsW6s98YTyC4ss6W6EgR8zq9xPc76KwqUhNV40I20XEDiAEXLaKAJE9PSHHHBIdcUDfjxp
z5MmVJUaxQmjnYEYUwXF2hbG6KDj+5sWlnBkL8/q26gLq9fPklEsy8G5aZ92J1LJuwA30pOlIcK0
4b9p3fwT2V58mkVNmiMY+HXPm+F/tQjrt3JvHJmmINN7IJ7wMrS246Ua0IDCirR0zRxK/AOtFEi3
C/ubls93Aj8fjE3OEig5FIb/RE/JkpGfBaHywCN2DY+n6VdOpm/4ouER8XH3RpSSWslD/JpxmKCc
2z7W+huDDiCK8LpqWYAIbYIJtIb6aN87mkEqsYPlLCFRjg6UhCHh/OngufWzsvLEGtPDmKCui5cp
zq80+R0WfAaFJapoviMTIvV2mvte6D+YwZoyUW8nrdPCldbh/bJkfLM4t01Tbf45FMGCYg9a3Pzj
yRQSbd2jnfy9cKJIqqngFVCZzXBTr9mt5QljLFEd4exK8kz5V8uei8AJ4EH/PTENu2jVNfaLjb5g
8w7IJmcPJ7R6yfsNmU5A8MyZGGHaRCmgA4o6fP+4fXDljhAUG7UrMfPyooUv8HuxI72IF4u/B86H
677ucJdHPISrrr7sLPkLdI8wFs7wfnpdHWl01eyvboZvc/UJ/k+viHPOab9T2SQWis0nTixrF20S
1k9qrwOxB6P0TRnUfg8eTHqEcjVkNmG10Wf1RxrFXqXI/+C3RjmpdyrFQXOJ3E4Gk9yzBC+/1FnP
xiSg37ltUw4z3ZeeEEQmoVJgRRB9yIiaOOimS/gooi2XFrT9yND1HDi56tMMpE2gcMUPtpqL2QYZ
IZ6uNIUwJ/5ZxjkNO8y2BNAIUfwTk2nNmbD4bsXC2tUvfhJRXn+kLeGo0X49kRr4aR620BWpAydI
bsXNRSxETXn3rYMdSjMvss2XBUMeLDnFr8pGtVmN4LixvMFyM3vOcQFzQXo6dS0bn+MMMbZRyji6
7orZvLIfo4Ks/m1T3zXUDrWhg/dAtogdePkUpWBuQmXSiyhth3fMfrj2evUsJw7oQiRnUrdlI99c
Fadlil/LIBGPiKbPYiMvYkhiwafLqchU/CIjPVTGbS/bl+SBoIdvnUIvsx16y330mjDBEOo4j0xK
eihd1AEsgp1630lF4iB8bDz2nE9Bv+8b8QNycUeXNE0W9Wz4AXlZ8eM2sGJ8+utyKvaiM2E5GM4p
UlNitBk9YethOAZEjs+Kna0wF3OhHJ4QUxE+LXjzI4mru4dnSZKujFjRYlqQBBrR0Ka5kk7PaKQe
sZo+ygtNrcnVqdWF9fkrzQNRif/a5/nruWUS8SojeIr0SVfsEK8mBymGF9XzS0sy/tBNW6LRqH4a
Vu0PmI4/V2m4E8616pcv5sG0NoxU4VTZIbroacxV9b0E0ztmEj9yvKTxsheu//6ImodN+OjpgjRY
PfEPj02TKBoaHV4dqXTY0wTNr+cv5QCI6ZbMToKsofexNyoewlqfw94PlAEJtO3xklp4zbfNEoeR
MB4753n5suNkzkQGHd2pI0NBpm8HEKuX/fNhAIlk652/0vEFHzvm8zMx3fwwbyr7aAiVVFkoDFp+
Z/EzA51QEhCLcoBc7L8viNJp/+7qBGiKnjCbL1LLdWBIY/xetvigg+svRaW4mDOzFE1Ni/OjEGGc
chp9hI6kb1/NIG7kkl8+g16rn8+0DFUhv/hohrr2e0rOPJ3DbTeYLTdNeQAx5uEY49cn2HwuWzu0
kKbj68cvxNUZrM9i38ZU9W/wzMf6+l4ktyn5EYsJcEGpbyuSzGq/BPOcROEqOuuJNbohDjqEQ+Qv
Q2BstZrMCrwgx3iRlBPrLj5HBbEeU2PO/vwx4i3rNnjnc4SE9Z2o81bHJFmLLu0dNLRg9TzQWD65
39OIj09qE3Zr8yu1D0zbR+1yWhYx/0FBwUzYRKWQvJ7LK40bFRjGFIj9QCUU5ypGGMKMB6FTYwQI
/A3PH4QSE7qY5xXplY10LCGntnwQY3K1SuzSlRSS8tQKX5ILLdhcDUSPN5+Dogjs3vrJk4DVLimI
HNBXV8v5JEVI+LwGtfSp/25Y78rqDJekZ9vUsmCL9nNaCppj+XzljyCjObP/lL0eOmZYnNp68KOC
VWXzOA2t+LbjJ4fKpneJUmTiEXiM1X80NbFER96BkGlsxZsP6d4oKRLWO/IYVFXRdW6IX+zyQ7bS
vmdM/TthLsEQZZhbKdOsvF7W53w1tWEaEmWUnZ6B5olbKTitBhNVGyh5yZbLl0dDY9hwrTp6/o2X
cm2PdJKiJNJ8lK8McxtEuri0W19xwd+lqV0J5p75vUOckHMK4eJlOul5CrKnlR5Ur/4FYhBz5l2h
UHb+0wOA3gjQ6ttiB06jBK6luHnaDRkU+4uP9FAzxknFEP+qco92exOG5mnqTsEKmVl2HX8BSbTS
X6v9K4/JIduPOOnAolmmt4L15ESUbr3Lxam6q+0lmfhEtd4AhDlDk/Yz5H8u8H1p8X3olP/u11FE
pQkoJ6zJF3U14ixw0yH4A7K2Y2wEX0HtDHJxNG7SCAKIn5XG/ksdw2MAnN2rRYo2oXeJEdKsVb6S
YcR6PnUxypRffCZnksF2rCYRewaQpVl0W02ks4KBR3m/4It4tYyFTXGpekRvk45ZhD+30dL/pEYg
0L/iCQOUAcoY1ifu7EIVdF4NMyqS/EsImA0v04yueAzWlI+VofJkLO/PoKyOCnZW8FZqVKEi2bKd
ASwi72xQHYNe5n6S9bCjnFSzVzm+1FpNmc4Y3mNR1Fm6943V9vv5FSEu2yiHcAJw5fizdRQ51Zyv
UuoM3q624DpRjoT08Tm7kD0JKsL7OIoruz5Ne7oWuJqug/taupi7fn390thF4zjz1Nuj0NXcavjU
M46LfN8fG+eJD+DT0HyQhHqHDyTzngabHDLXs5lFFah+nySkoD+C/M2KQjvwamcL6MmfMe3xQREa
7XcRSngGpe2JgF+/CoWOI7ktBD1yqR3SyamTQFAWTgN653jyTG0m0qvdRc+E1aluDFWjHXyi96bd
MeVFmqQd4aq3A4mnF0uaEjcrvtKH0J0OZb4mAegJ5gIu7HBU/l1XRqY/EEhQZ5bgkiiojKUdwbP/
pagKgN6Y07BPjVEKAXzpEAa6IMuQmX5T4ku+3z1cTcQiipn9dABSR+1xcEXs+z7bCna3A2KwtY9C
7OasLxFmcy0zbptd2kZcD2oaKZ/cSUZGU18aPXbT5afYaTkGyvEdbghpxLgUUlX4A6Yc3dgIbLn1
l40hc6PztVznCO5475atgx4W6RqXG07DYbYTgDs+4ej9c7kt6UJQxJvsnXOq8narqMKCyPmH2bWm
JIoG7z1S/ZGKH1N757TdOK2y+yzmCiLFYdblB6lAUOsIh8sgkKutLY2nFJgtPzc/f9F+ub1NTM41
VVf59dFdUfNQQvlvWdJOjDQyYqiWAezM1LCCvuCNam1XFGKq9u8CkUZYn8UNy1BGhAUrxrso/gDl
NC+AQivoXLdmVeoo0r+fCQLTSR+3odd+z4HESzDdEvy7RbD0MCfq82xcr/Mv+YH7OjdTzD/aGPPg
lYSWneaKzSDcrp5741sLvI0kS7K9Z1FSA7Isk+VVpsLZ26YumIOpHH/mNQF4lgPHmkH6D1hjB43F
RpO1cznimG0xGUAKKKvozka/+DFgnLgR8ipjCu8O4Y1FKe1cmUGL5g0+QI0jMW1RhKNlWwTnciFk
nx89uWVivQoE7sLQXzqKpQ9OiPFEiG0fbOd2YS8rZdh2NvET0aem9UWOVYRW0zSCX7wT3GYQGqQ/
EP7+wQTQWpqvR2wbijbSLtRRZ/YxY5m7qIO2j2ckM0SnKSJa6ETZBfSZcE+1GkYQhZAm06FYa5Y0
7o7VQErdS5duVMXtGYFqoRGQ0LkbYSywNdDnEssI+WDaU9fWfHE8RVYoTKbeo0ETDTirR0Nf29H1
/Ao3pHEzCPxqIykLjqtAHYHzDHMkCRZrvfBLg30X/B9H98593yd2I7wMvhoMFIJEjyMVr3d4RUlC
ezC0+W8FLnQjD0ri0Ioql3oh4ofQOtD6n1J+tv5bJ3RSwFG8NqbjnxP8RmpKq4ycmfMREqwbQHV9
aDxzs9QBOZQXGt//sEXTMg8kxWwl7asrlcV57gT08lE88qflhte0GDeaia/cd/lLdLDwXlACIybp
mFOywVYja3C/3f5la4BP+Vzc9nHZvsYWxh7VwnmOOV9g6zxIO+3i+qm8znzE4N8Ptmo6cvaRBuMb
yHP+mvre/kvLvOkBt8UlC7Fq++TObeISriifG6+vruyzA8c6r6j0VgI0IiP78tNBNNQCqY/ml3GT
4FM0dJxgdheLgh/n1cWYBliBsA70/5KPdALYspqdf2DW3JThUzC8CGJ4zkMfk+EidF4BPJ0SPFmY
b94mwhju+8bv5xM3fyAd2KXwLTZgT9icoya4SLtnZX+hCE+VE4SMhBFtBubGa4cQuLpgLJJ7OEM4
J5SH8negsKuyUaUVAbHmFaiVGtdvIyRc3CHMskmm3vaNvdRQjPCnk72MVpKjLjmG8oHYl9oGt8FR
y0U2VMBOuY6ytFUarM1z2EmV1njiKlLB3viV0lmMGkWhSJQBV0Bo2izND9oMWyGxdtoOwcUxXxUL
I9FB9hShJBZhO9vUDNJXib9Ew7Cc48pgHR/07tWj8v7R3gcYOrs8XfkBf/SJn8SVe/GB3pjJgrXG
UCgtr6slDOcKfnRpOjoBaqe46E9PEJJEOBHfcm338+0xR3NxzF4Nsa8FdTQiA3tS7boFauDwY6zi
NVXmo7hFw/r7XRccyWJ5jehmt+G47Ebu2eWitRD7J6NL2oXuT6/rUcTjR1qkix9uy6OvWkjqTeXA
85WUeJ91jSfvoOF8v0mQ95JMRantBIkqlkgMOpfeDnuc4/L8Z4QgJQWFPYtkYcmGHvtFy+9ER832
VzTL3CgXuqZEcw7RzDyxTMWbG61wg0B3iph9uBGFGxfhdNxJc2Lj22Cf8hmaX/RIrtnMBlEriJFc
HCI+9bxGJp7xbn+spNvgjpqvz8ZS/G1/IezlU8Of45MEk3rm9mzkLYVOaJNb3zvK2sFQf2GniN82
gzH1yVba73bAltoV/dRLCheGsL8KJJaXv7CfpRIv8MOkBtKx53E6j+2tcDu5AsjDclySpBbOP+vk
+ibd7EEc6wNa2UWIdSRdXohoSZVDgfp1mOzU6xNnN8EGPDbg9zGIoOT1KFPT4nEZrsSvWvMW07Xy
iBwDWWFIzZHU4fev58GqGeqLuaEjrr6KicRtWL2XIoxThAAYQIu9PjW7vMWq2BJfYSQYH22XpA3q
lNVk5obvwJcAUl3P10Nw/oKKAd2HKz264KiPHPMgwSD+hyZtRk7qccqPInjbAi+OrXujowYRFjwa
eJZ2ze0Lsu/3HFk5+csVKtrS9YIIE4tjvLJJnLNyCg1Swdk6g3hQgJNT6/2AYB0w5DHPdsJWsrYV
qMSIPYprY9GhtUGyRRYc2PtHDeK4zk17iS5jWzlhWgpUuVuo4jZyUQLpYkywHZjxhDlpzD5ytNuQ
RH3PIRIhSydKhAAiHj9kA5prZ8W6IWP1SuGiq3DPAhPNPA26YGf0kixPqSVEr/vKKgl8+v7D3ew7
XuFTx0JrdgILAa/EYibxj9WPkbPZgnxNI6i6ffsQE9E8vGSlEQ4xNTjPp+/moD9UPr6ittcqkvcF
QHReWtepoA1QMevJQlcFLHLLiIx/9/GLKmDdH7M7Saup/fZ9n74pABbUE00mN6AZ2rUFgKULld1X
yEH8TgQ9H67DJwI2rL4L9l2r2VQC7URkmOTB0L8l+5Dc3BYP0dzfqAQNTMOR/up/+nOvkzlGP/q9
vXYMWNFyldxVN7XQo4h7Igov1AnbYX8OVOarOjjzDnVWAPb5Qtn0CaGn0MLbI19sy6BZzeFpWpaZ
asiia5EORgBTofqFncDyGGgdoruaXCJBN1+nQDzHNSoUBQ/Cr9TIPUvqZJ7bYCDJ0f5FQIcma0Fp
tPmtqhh1VUAqeRytjKeOx+7tkxt1z7eraL1G/FkZUEcsna844+afVQ3BzW/henZ29Z/AEpxZZ45Z
DB/whJa7hzdEOHjmjBde1Lraf4NiMLePxLz91/IIrhlnsHBimgHZEgl5mRtRwugHUVGPGaZVXP6r
z+OH3zdMyzBj9s3MGl2nsRhrb6JqwM+TDewVjsBtIdGPy2lxOegRbNU57oRRHM2J7ScZOGnRxDZU
f7IQY6TMrLkkZF7xXBzGlbuKPovQqUf9NLv4z/ksSPu2Iy81tagW2f4XLTsgAquKO2ss3DkRpZZP
gOx1fLcog2ZFIEpZYnjbanAKVwseyfFfPjrQljZBo+KqHgoHh0m5t5z07t6JZIZ/lG0Js7amAApl
tm/6QbWK5OvVz+rK8Iw0ZJ4qKtncNqJhJDVN+nGmxSbOZ+rfMqWdfR/bJqvgald+tqdxAzXYAlux
f96aVr7qlmtA0UrEbAAkoi2JGjT4MqoyNOzV/fw7QhveqHy9MsvKaK1zmhBEAFCcHbIeOv2T6YlB
xOvRo7Jq9zItMBhZ/nwm1AktXJFQz0o2LZ0Mm9FJ9Ymi4nQSBNIejNVSJO3FqIFyJf9NGFuwpGB3
bmcZqZ5QDBGQxGvXUUw0fwC7DsQSgBqEvFsNDtsa1EvUrhmFF+ay/kmJkILLTL2kC/2xZ1xPk20x
pKDys2sYC3GqQUehQWpgn76feMo0GkUtlf3PaXFE3/Ck+p7gySrHASyC8xM7CTl3pP/eowSwNJ1U
XgwlOrXs3ducvVdjHIHCWUBDMt+gcfQRaoeRZZ5vRe8WrJxTKXVWZ8WQ9FtJkSvqCI+7bue/PE3g
b/YRMkNyfcT5izW3Wy7jMdyz6zOxmkq96RTHoT3ic4VM+QcQrExHIsHsVeo8cLLshMlo238UEo8x
M4NdQ8quqPC7+wAh9RDw+T62UpICrDP0/vckvU3dPpNNiJT3x7mKk/CJo1iDRMCmL08OQyhqacu2
XhX6bLOtrMTeSNqcmCz1EazRLs1IGCOPKvpVNL8h7mDre3Iga7a6l4Jo3zUdBPNefTDdDvyd/Du8
IEoRRDNxREHEnkJMugqIdIUHh0VoAv8xgiVVhlOJDCBc0XtEPnAygqtZO393z0Mc3kIzj8GEILr8
ProXBtwjoTXom99c6fXNfcfvf/83pnJhc0HRO23/0ojcrmZSWpU5mffp5F1XssSxkGX1IPq0q5HE
zXuZDZNb4VoTThp5JSfPvHzVqkwNHAOpWmIz5fD1cremja2818aNTjf607BWqRqzPVBaLfCyLbIp
b8oyhemssmKrWrollQhS9ss1Fg50R7bD+Ow2TwFPpYgN2Uyy6shZw326X2HDeDsMJXQ8Gqgz0tDu
L0BAsidxkLyqCX/gT8A/YcaecgPB4y10aiY85YRFFjP5BaV+MbG3QaPy7PQXZ4TXt9j7RvzeJx+s
fIYDiWUoxzmu6jKsW8Nkx/2aIf4F/BSYT4exyXufmtCv1YLh71SEeC3rav/NGBqV0jtzHQLg6FhW
qGYtEJ1BW462acJ2zHYBYONDuCp/KyDrVOMbAQH7AGg9BQ4l43v52p57bYon7TCIKYzvOzMj9uK8
biCyrIwjTxQQPTJRfdpVMlhQ/8LDKAu5GOflPpUOYexIz3OkxJCeThkrrG5exUD3o1YnW1eQwuf5
PPS7YOmcAX7AowfSZRNTyTyLvPAKcj2sUeVvD3Tl59Ma0LZ8XwS2LgYUX8moAAzeeoyo/cYfEvlH
vq0f5kaNhpjQQ1XaN7aJNAvFu0MxMcMEH74uI0oz+RD3bvBlmqadMqAnwPNAT+gGHpnbbX556zXr
iK8GQ0bOOqTku1s0PUdzNuzXg2VWbc0idhrVTQ+zrKjmXcldS74Z8SQ+ATMuSDjHJjppCMFpSo+h
9ega4K3jLa5+VtRD6VYpSSox4Y64j5dT4Wq0+E0qDRYJI7BmlvmAnwvr9WpTUSwdw/zfzo2tZ1xb
Igj3J/3fDA5ctn9pmlFZWqpM++5OVk+9voYc7LOdT1slZqRaK2dmZjNtaBOt1IaUaQPIb8N9txpd
DCGxRvtRMDA7chtsQYlyuz7Fa/AFtdaF2tO0EzrTWwu7tzZjzsi+tBjwfaOx/WVJORogvGQ0Jklm
sobrYtMp/DP6jTb6rAsC6Vj+o+t0FSU7xAUAWmSnAgzDwnBuoWyTv2UB0IZM34srIivg2CIgdYrS
qlL/0Ph0iBiGaGwntBGMFFoMpXsK6JvLFQc+c1sIyehf3Z5eeaI4sWoKcVGgFfjjIA0DIZy3rLLW
K2ieFqCcamlcteK8vZw0uXkFJKr2nZmkWuBxzk59XTphF6PpGnHWMPZRQYuDwrFnO3c6gNWSKhjo
I7VpTOCFk5EvYl+lh3HAGyTdcjwzsu3b3C02WK0bLO4oN4vnjD1kqxImAXGWyowkojJo324hxOuw
cefKIPyPCh2Xu+sU560TGmOdpnpy8HjXpCfV0z/CwypkslAW+YvOmT0W/1aG3mTxgMyUsDb8rqBF
8iPV8OKLyCqXoqW/ywA5nMgWHiQ1mD8CMBoIMgaObguBd2FDqIwfxHvKuUM+fOGdtUO9IlW79DNB
vzchLAFhnNS9IuWO5grzC/7hsS27Kk+Mx3eZaZtk7JFxmcziWOzkdzW/P8nTsQCulseNGI18uCvd
GtYG0oja7/cacEBnYgBPooFF86D7bBJ9JJKkCVrxL0bLzXI0lowoiLtC7eCyXwKIqF/dZRMhs8KO
QKW3t951BkUj08N4tAvpKvdAHQpuWbO1wp/K1H7dJdyLcqrs7rume1YHB9UyR1wTIqpaSqCjFkeJ
vooAB5Z5BOu06vGjsze+wGZPuo9f32n7PIjp0bLq+stTNxeJs4TJkPxvR5cNQB4IOgDXd1a3BGvi
TEtJIMKs8bN6OnNvmFuuSsQP5YQXLtl0a9eOL/C2rDwlmzM3NZjyXu3AxZ7X66ZbzcElbqMOrng0
OtXQxeGc/hPcSoF1uJszY5zvL4wGGiiR3t1B6vHuZ8MKjwW3L7hX+O3LjKSshBTDY7Zv3vWeIDdJ
N9HgeMoYYJtjh68myUS92dxIuFcxtN7VGQpGl6sJmQlngdVfikIfpQD95J4UERHELDok1FAI2Wdj
qGnzDSnAlKvVe0lbQJWca/Fbf9BSo8slgQMKPQbm2ccecNYf9jEV/G2slQhbFYyvY9xvPtihkUfv
WiT1WtXhGn/jgaXoXvCniU/0FR/00vdAZopiEdoD3Hq8tqBn8+ac9gwCDC7vyfF4qeHEGsYwd6b1
4anG/vvaT6/P4AcLhyWi/F9I3zlqg8gWhU23AKLkdK+Y6v4f93cR4oyIRPplZZ8Vj5llHlg9qKWK
WUqLwxGwf1NfJlP2+jdzqaTTnLbreYvmcx/l3/C3s855eXbFXehai0H7jJN+B+j9a9yFtb1xtGxd
rCQLvj4talTsNsXkACZNmRX+gA3Q4FN0TQ3kP+QeVO7w4QFSNa7XFD00G9CniL6CCuynmvd0D/53
875e9oAfDhACQib8VXTvfD2J4aJH0xyEC5UO4H8SZjIkB2hKy2ugWx8IMHJR0992AwBlmCfzuEjA
Shy3U7bJ1PyQqmY5jfqLVwuEfTF1oZDG6YR2PvtwwUE6c6Y3yDvGnXe1KUgeEfX6PT+Ylr3aj5Lz
3MD2aKpA13yF1DHwvH1VwoGvVng4WMfr5x43rnPcDMQPWbe4TtR1hrzvlslDn4oPDeB2s0XVTwg+
bVZxODHq6fv1Lkx8g5CBmLFsZmG27Fxzd3yVq7kI+b8vMD035+Xct1xXnmU4aFOC9MqMeQ9lM3Lz
lA9INwq3vG08CUFluyQlO34qhahT/E5SAAAYmKmc8Pr11mMSptiyY3d2jPbG6W1oxTmveQCohX6q
TUogaqU2I2b2EFt/0c4SBH3WL+4lNpiL4vXFolsXSwXUcBUjM4ixvQFnyrWwwS2uZievM8riMdyt
mFx7hfpvyy3t+bkyl2jz2E/iAUytV7cTpFh7y+SbB+FjLe8ZbjDOIcY7oyq4LGvJO6pARNBuz1lv
diKV8RqhMnVboqNbdGI88xrrLDYqQOjL0g7s7LMDbqyzmbVgMbpH0JhEGsjcqmjZ/FpKSgj6u81D
kDu9S8P3TpcwWhyPOdWB2jcNRUBXQyQVHkAgoRd+AHk9XmA+2uyVXHNcTPJQZf4i2uaMSdu5Q1ha
kbYxguYpcji8pTmDY4Ftz5g+JPU2DDNs28clsYGE7SdCj94vEppnQK9YKR/QW4SEzkn6fPT4G43R
RlKeljBPDpq0y5uTNNdKoFwpmRdjig94BjpxzfdmZLzIx2QgcbDVxHNKDclhS8HFiER9JSgqzcIo
poM1FnxqsDEifA1oTSh1nuGul+z8Xlrqb+Z3RzODb0W79c58BHcaaFBLF3BUSuJ1IecI8fhk3S/w
PN5qnzv2jYmj/SW920IJl733eZf3hVaf4p2fwd2UtH0WdzIHsQfi+x8knvkvMRpCD4F5nFcKSTlW
F8X4HWkFBxARLi9/KSb0ladwdIRxf0zrwQ2ZpnIkDDV339QYHbSm8udZ+p+pSTdyRw4N6LveDDOZ
7T0ACQTEBjF1NkEhnGk87mdChnbOjtjn4tb6yAnz/GfQabuCEOXNcPZumQJrmENpXUSunWKB3VH+
h9CmRiUwvl1h//fA+cmqD1DvUMxhtZ4SK1TPMZRwHFLxXqDXc0fETcOLsPBXVFvPCG1hbaHutf2h
wcHfojDog45kY6KXOaGJGtBLaDFKeEpnRyKT+/vqR3SJsYC2fcn0NyGPvB74ZDGAsIoHPJqT4E7A
rPTqxUw2WLDEhYdZrAw0/vmN57iBJVI/rjS50d58q4+OwIjfUZg8hHIfVMCmmFbxr136wNoBMCNg
s2UCJG1bH/t1Ch3it7Amg4OhgtJSBeG2SqV+KmfuAunMt+0adwHrfRlmeyc3xgXnks9QYK+vWm0Z
RiHtIczo+CdUkojGLKManiAf84rxc/mjbgKPZrb+m6jEOkLnSVmWRvf33lHX1SqlG8M/WH12E5P1
LQT5Dz2iHoA54REoUDTVbwyAXsSm9XNTF2bqm+ETUimdZEkPYmeRwDDcx1h7ZclP2ZJgVebMyNJV
+BnAxWtEWgFSIaZ2DmdM8119Vqvb16sSH5zGuYBxmC5H98OF8bJsb/ZIbI/zGxSF6EeytfNDO2dv
jZ7pmS4vIDdfYnlO0lZrL0Zy438c74tdFR9199ERgEwfm9AIm0SxCNg+7d0jWI1oGzYQuq1n5qBT
X3N9cNC6AjBfa5Bf+G+qgba45teT+c5LZrMWl0M6xZIceqpkAiNdt04Q/kLNFOlZRjKNVc4mHloe
JKjyUYa4cmNIdphvqAlHgLU8jVVS2haHJI59nhWooJkE/ddB02JbaAeiqFbUWRpJLO+wLcgDp9C9
C0lX5cTbaUFqGVfxB9GFrBZOp4NyxuR3g/hedmQ8McB+kYBTHhq0tEeUKSEoy178TWG9TMUrczzQ
/FCI6n5jM/qC0q3ndVP/pyQPusKU219UtLZGWDoAAOloYR9at6mgxtr/FWKRDFSzZ2G2SO/sOEtB
glnKvMR6M5KqUEk/h05j1ebLTIdOIeblXV131L1Mie1+tKsdMnilVRPPjV5pz12Z3ImtqXH+yW4V
9+JIXIeRWL3eSxmmx7fEz0FUHkJlwS+hFROjP+Agv80PqJwfNE2JOWrOMbDHp+Vi+9rrr5z0K62H
cvH08JmN3yCfIMQ1rF6rFTmthHF7X8xhghygT2V8Tpl+VGBxyXsvI4kcJObNtcWKOdXWsYsAIZoQ
ZRYcXycIRcMP/LXo22clyp6WCZwTkxluGop1yRIJl5xHbmvaBa6XwaDJ1bOfvFvWMC2t5qS27WXH
2sOx6D8k2dkOQDehBeLK9oXBOFJ3RUF1F/SrUBJuJABx+qIIoXHt8bs8yjtghS0LQ50c4G98OwBt
Y67uUw1nieDv22YVeKHh4FY8vCddIKmyScpJFOs0gguWdbGKxi8j8i8mrwH4Fw6pLigArIR928YZ
FLEYBWoAcojLvHBdkwnZ4Y/oKE3I0yyULVvaHDd3GxYyQ5A53aphfJzC75h2yTkvQVcfOV1Zj2MM
LY4+l1WXZWNShG+ldhVCfP59q05X9795rdHP0znTVyadBnmHsSYHugtUajpDZFjDDfhPJwXY6lfa
USNyOXNJ2WhilVBubrZ1OjVjNLPsBdS5ngMR4khZ6FbBIi31cF6lDmPnHaEskXDj0FkqUUgIjkIh
NZ1AjEOMYQjPoJEejwYOy9TrG1gtAGtqFZNlz2mpFv4TksJLLzAgsoD2+EUDHfoY0Z1c1QZ66+31
OnG2T9QiJJtzFLxcVS9Mgj/2prl+5e437yF3K03WPvxkBt7kNjvdDVKto2jbBwi+VEKeuPQ+MvuI
GDUCIE9hsuyCgiGVr6lXsIEaMDVoEya+yYNfZDWiNo+P1utsiPaBfbClzJTE1TVqtxOcCvkSOKF5
325tKVnybkIytju0HDn/jPTLPHfmd8BRRSzhmCg/OuWJMc5X+n0QZ2KC/r5SY6mrrUJ3/5sNSj2l
DJXi7zX9uDBAteaQQwMKtpUMHzVknfBYSRc3GpPykkAIKU/x42k07UR28s6v4590KTHJDSX716PA
3MRwdaKlCcMP6zJp2IW+9iDGRgZr7v0fqFmGlfIUVu9rKpGuElLpob8vpfbNDbvmOw3NRxr/lcI2
7YPMa9UOzgD7tFuYpxG0TRp1iWNCs04TBQgHxagfuVebTdyrUzoTKWJklcPAij5vyNaOm9rRQfUw
s7gdxxTVlVstS4WtOrgizO3sWYrnzR+BRFCp5eHd2dSKwSnGXl4qh/ORQGOjySG66CJVBo2FQktO
LodYL9A2f34ko1aKj2ygwkfpjgqnBlerSvHeR94SXzH+XH1fpWOshijmzD5xkjKMIhdjv99psLp9
SCZ+4KXN+rXN20h5qJEpOCobHgVPon4MUOWCDn07XCBGz6XjQ4GqFkLLlMUPA0SynmBNmj0/11HB
uL4/lWnvV02G0U381Zz3zWuVbFA+rjCedqrWUJVZppaRBC4Voqc2AqvHtEceR7il2WcOjMiX94ov
dynLBFQVSTGr7gaOq2YMQAb2y1HQNyjsmVNs96balSgXIE/Mcj8dhTQIJxXK2qqhoPxjZeN1C0jB
dGfGhAL7RBwA+ITCvR9WYlv6pvpdH25z+b2PAKeDQGSpjkaShgMsvJwLBdpHeFpFGodip42nxp0F
2XZojUHIISnt4euYNM21XBUNbf5g9TzJMm27OrAEeYZcGbIXKPMytDQn/zN2B+8P4KTA9VZ29sSz
OYbQPEnVOjGAqpATGglfpEeFw3p6zug1WJm07aeNmRvIVplPb6cZV/HYpnYtlSjqh0m6xI25V6zm
lW9QA4Cvw73az3AU1YLePM3Pcky50lN5M522uiU5Uz2nl+o1TxkjWs9BS+mvs/uBFx7Xhb5LRGCM
CCq3oMWnAyMR9Md/Nwj1raifaxoYOPxOLOttVDEFIAgTtmce9CVpgRkTgu5BBuILF+cfDpYKYOaZ
BzOfokeXvtSQ/I4SOf1aaz3NlxehYHA2cLZ3SN9UEnrzkMnysL1CEgN1GtAjrDfqtMfizeTgFAR3
ZR2BKkKK/i9xWxg7miAqlNR+Fn0QmfmQk8icfeyYEfmH6bq3MMWMyGZtvRuKtZaDjOnWE+Vzyn4J
AY4LL7wkOYLQZvJ4C7C2F1m3Dap4IxEh+Z820oKAvfJhMGBkTlZpLV4vYRwbUEJt49Rqr7Bda/IA
YpAI5djUM1piWHC9nNT7DFyEMKAOGwDasZcGI4LABBCSjCPS1R53F8f4/8urwQF2fT72paBqsh3u
6Tt4yODkUbsqt0MqbaunYOoGQOW8DXU0jx7GosZdFgaj3MjjBYiELoZ3gJ55A710WccvCkOVLUI+
CGOJ28wcDmcVfOsRGoL2ucpBV8fx06SnEf3rB1QEiHJQoPVu+RM6x+N7WNGVMSx23frunSb6PKfH
dlicUHcbKxueMYD7Fot0A7jvzdn7//WsD5zqyqcqKrpQmsNE39d9ddHo6I495c+wxF637TBDzhTV
xtcF+Xh5kAzHQPjTzc5nRclg06GKz9vvhuE8O9UwDe7sr0oytfJBmb2R46tT7ydBXmJGWj3CK+5V
+jLlbRpT/bEXtyCGYam761BUkeb8Hvb9fiMVNTqpNv364LSADtLdPEkhDwZuu43dWT/M49DTI1aN
LfpQbxOxAQFCVvO9IjYgIULOEve+7/ayKbuRC5WNa6BobbGkILBhx69kozQYsh03eO1Ro+Ycxm+o
bwCVXf+c/8Sjrm0SFObchxMCzpROdoAey7JP3uZemNUwJfjR3BJkcvwyi/YQ2OwPUNRAmXKF7U9k
ueswYJfa2aOMl+IaIFpy5b9HzCxbcFvWCckCKgGAcAcO/TcXjG6JjHwAy6YoakGh0zchgKqybHyP
hAN0HxXuW79W7FZq0EHb7TJ8nb8QIPoNbeoxYw5ZhyYbZA9+ySwQyiIcmc0JeX5MLsAHOe9JOT4Q
xwHJ5Xu3PHaJxSo5RSS3Ygml3QnS0yIEP//lXSt/Z9f7vhe8fjvvVQyAkgSxQ0uvFyQpq3Ekiros
28QmU4+Gx9yJfAoTGptmgIc1FLrWgs1Ys9dYZiiv7jU3qZXsf0IxaS+TR7ejE76PJTL5dsRdMw7O
y4T+0p6dl8YP+2DEYDZI108ZCRTcW8dCNpkF6iHZ/U3SIvUfPGGEHLtx1YzDDYKNEKHVZs3oUckq
E9nxVj9sQ/rcIw1u3vcIfHPUH2w7r66KGnJX4+gidIXGZIXtcrLfe8CukVeJmN9bDsU5jy5vOixP
nwu6+vwytiIR/+gMg8VEGSH3cJlu516Vry1Qp4h9m5GleZ2tuaH8QQ8qjces3IMb00kbbIToyjge
dc0F7gcP/lM7/+8N0i8K2v74TntgJs+Jgdb4frSWUNm12zRlt2XeqOBdZRy/4syQrIb+Qr8LFyVK
YBUCfGTdiW5QrSFyS9MpuMwlfRt3LNTtwiiFgjk9FSsBs5kD06G324jcI6Go38sT2wi0DF/Rrt7w
LOq6l3+a601ZTHipq2EaMi5QLfOFCCsAVt74SaS2vPoSvh1DMt2ZMNurcyoTWEwcLsJfrdL2XLAv
Cy9jzyOPSwDaX3gC6758b+ON2DoBsfcXA8zoldvsm5Oy3i3CsFWbiwxY/oLK7uAW/GTn2OE6FHFX
8xgT5lYGDI2F3adj4Em5XZXIlCGi6DkC15cseAGG2HTKf25UVon/CXhjeyqz/gGRlYmC9h0LCVNI
bLitQAopr0c9D7cfvNmS7dN9anw55EZcU9TKufVWhmaq2eTQGDx0QDEM7jGEv9BbhKuPCSs/fQLs
CC8+fBVC+3HzC8ys/86W66ZsbssRPVKgtaw8fRRvnuOLImScBKUtqk6LWv+sYGntkAeIdV0Qml7+
5ymid9YOOXj+wjh7jBEXOZRFjkDGOpIY15PZQliP+HnBrzkajcvfGawQxNY7cz6up6Dft535PIXl
avlx2iZOskv/0V1CnKKuwvEU/h6mU6ykjPUK6+LJZGLOShcw0OgBJD/Coo/LmVqAdC+VVCRVvTAL
3tDRkIVvPADDduEy69CEI5beyRwfQbsxG4jn4/sE/wSEIu8g9DPEJ90UN2TLvFoHvMHJLafofNq+
cVesgwr9t5bXZHS44L0Gp/Zuwu/5pCNyphMoZf4m1TQtO5eDwF0i2EosgeqEXhHpu0phQpsHYSFH
bbdXdccP42bMFy7X3aYHGnEJ7sL6dPeVIjpIM3OqnZ6yM4s6273pl2xFddVrvuOb6AJs4c867FqQ
XYD2tT2sa+a8uyhfLyJfArREpIpqRgdN6JL9xAiElsXZCfvBdBVicZQTvXHvrB+7GXKCC4yTtvyY
hWQNCPLA9YoRJX4kCNjuVYKLPnWy8aLLoxbZBnmro8eMV1Vw898+ubwtbV6QKfAt3tnwMCfaxa6Y
fZSctAkVbf5AxbtPgO8PxxDJrVAaEqAQiFxfetgYJSLTjoRIXorn5YZirEZnkkKJApyrFrC0SVyL
Vgil8NkFm+FZHY2zSqJvhZn2kUVm+Hir8ulAGTebcmRxCJA2cyhPy5YEunJE9LxgUR1S17lFBBco
PL6c/kacn43FHNU+izCxNO2u9VQM2Ib37L9UB2S10Omyt2SWdKFDfH+bJm+0uS6jTCpvuf7oqPuA
0c2bkXIPJtrQ6wc3o/dZBFlO8ZPuxZD6BYV/G9U5BsV4vtzjPrq1DXibABt74/QlbFXqIuz8N30B
VFIFawVMk58CYJU+hGS+9yKh/j7kpC6dO3/UcnjbYB+47LCFYaMrum0t2UOwNmWOIWMZm8F+vdM9
pdBCqYZkTyIuUV6CIArjPrmKzNz8if3tRH+BnyLa5UBcnJwhTPkh2xvjP7gx94ZzPhNyBTidct4i
83DC9oVinXvZGnjt7OFk636rAi3tn73qMxCaOYpgrwLQtGMHYtQhjiXx12gl7KNEa85AAYUInbdJ
MWTqbTh7plpxoGR9+PjarHRJSivKUoqrXI8aatkbZvy/ICOF5pAnmEe8hiVyvyrIUu3GSF4YKF1N
i6yzIUkczFKpvczZGRZ1AI0wb5L/WloAjeP3JbTCS87aXqN3XS61WTRf5TUVIX45d7FJNp7wp/K7
S59qzAC8S2tR2yOfy0nSZJXDH9C93sbRLV/40FDYKUsR4Ay8uoKtqzldtBMcFONSjBPizQaXay5U
kh0TUx6IVl5YC8G0PkFsLWd3IDplWA5Ig5ogGthQRpXErb2grhz0fXvbw7okrznALwTIdnX2Bp0n
duQzFxYmw9QY/4wJoI+BnP0HvenvLZN1h9P40fs2NdpVD/4oFCkyEmNevKxq91/0pIIQ/1fo4dPR
n9hRZJtVmy+bQeMPi8zgWgvaLd9ogMXdBe92JJe7zHv1a4mWZNYYHMucVhtrAlJUdlAY/MJaWkZn
FWjInNhyD3g8A0xblCLGjDaskE6ZCnywCTFagUcGD9YpXhEqZBnH0f/h6OXFmHYS4wXjXbx9FRti
rqpy8Ma5MjoI4UhizKBp0aXqDemKJt98cTASyKoNMMEPWHGjcAcDuAahmcjIS+/nftB8/jMFZtA1
oEG74xS+Zd5HIBfKZehSzqOIQS8myatHh+aqTnEQW8qSZm7AnADAfnjMFyTtsjeIw0VCxprwMFie
FA/yGXro2tQhHNsbWdkM3VByZixvDBDZuu0h56Kp24CehEfLrf/Lx9Kwd09lwrl95TimYijdmzhR
o/3k0YsrbluEQPQJGb1h9UVrIDs0HtHjsx80PPUR6v5N5I3ctClYAJ18axqjrI/E4bQx57zxGmtJ
/hFNriLeD/4H0AJMnKEL2ov8XsPieu/nkN8fr+PVnBxizeAJrm81tETGdOJpE/1U8PZRIk8ydw5d
vMGClMJzb+lC09juN0S5wKBruSiEuTsfgK5CBW8EHgJTvovDs11XdDSQDo4VfzuIk6UnIsEXmrU2
egmYy6IpKVdMMWHOv1gyEzmajnLng3jJ5Cp5ZHc76mdaXI3g6XLAXZA9ciRU3ouG3iZUMabCNvX3
F4GKAAcCZxX1y8D/N6m05DMEWR5zKQce0Q4UE7op8rwveYiIkCPZDdOJlB48rvK9DTs1vlV22f+4
PSnVQw1hSq+M8/nYSeCehwSW5N/v/gl3xJCAFSe0gkGQDgD97ablGjioikT/a91oGXDdli0ucX/w
XwOFiLnoS1k0NBkKJAnWPIJ6WLOvkEtNvtnQHBdc6zUcgKzwubh4OzdtIQkHCeGUH0zYQ0iivdto
Is3OFt5wiUbvmxFjoXhvDeW6eeBUFHmOFatiXOpfIyqnsYkr9Lxmen3x2jp8sR4of0V+xwfIwQtH
+qjEOsvm8mHWLgrGPj+ib1kwBPJdl8bWwv1ElKH5u9Z0tumqOMe4HqTwvKltQ/KsgkRmJYu6PEzL
W5JcvUdTyujTiB4UAIAK2vg6+r6LCpHdbf0Jz+NZ+wWpTv1VdAHBs36rPGSjhoXo5hNYkbK3LOH9
DH9mg3kYC90CW7xIIZd8SB3CHGgakcZdSsoNo7ijIC+Zh04VTagwU+KSe0uV4/uOzgek6Mx89EUn
hYdp+23L6IMnp/AFZsPq8rgluP+ZWwLyJdE5IIjSOvM2sromAaCmdptWc2+cHAbXb70NqDbjFEak
yGwgrk9vYshCw+sVOjJD1yQ6oF+5FVBgkFtv42wB4Tx60MCTlBeu7j2sFN9EmaqJVZWWk/Axd4K6
Ap6QjS9us38IawOrZvogui/3guxlMN69H8BMtmrFvzmWZmhyFEEUXGw4oERve9Ov/n6x0E+CNyTr
7/MDIM4nbgPY4DzwWij3J8PmH4UIEtX5pW+qTGk0TXwzReLxH1fxFU9RUTJMu8MKJa1FEMdBho8d
pFbkzIrawF6+hSf3nlEKUV5mZzaR8rb51oI+IMaib2pS4G4YupqQMHHxHbWN0MUW1SvI6WFv5dGW
tM4JAp/6CfjMMnC5v+NzfgCBTgSNMGxzYAXBCT22Bt8yrLvzEyfJ0q68+6CF3MTv8eLZhTY8ucg7
zTlLxeSfeC3K5jnHjycWaGtcEHiEH5whNP1hfAq3M9H3wyFMN79uQAX3RrAqe49B+zrxLy9FnwRy
svDhkyPETXg+X9/KosZh4T/B37UFik+KpCS+aQgT5lo3k85ddJApeWn1zK3/9pw28FREyGRlVsfk
dG5TFQzF0pJlUGmQHkghyWc621oP6sw2bWupjTf1ythstwKqwflM3f4LkdSsytWrrgw+t2wEAM74
MPHjTDdyMSMGs0d8m6PnbQluczF7l/df9aIN4sDIZ3kyJkLETaak4ms+W2CBr44JtPf4BeKgiNno
iGNR9+WrRPRlFridIXRucIg9ZsEzq4tJcI+L8A41zfSyy8+178qncldq4NKaprpqmgOxLFyFoOrn
rt4LSO2g93e1ttXqpeYmtMvVSZ0kl90J3BDPmEkHBOf/jt1OVlf0zFttudCxNMfbLhH8srGlqNK4
w2ZPnJf3jkRZa5zRrKf+TqFZEzHZW0UDv84dux5+aFNqFTR8d3dS1M++T0t7KKujuUnt6jYDaMyj
XnFuNYvoUHDBrGQ1BBnuvGMwj1zMpSy9FXdvOb7AwnZpX/TeC9hICFMn/UKFPLZlaFTRYu7ISsmB
0HCC8G9QPLUXnOOc51tLoZXlqE1ZNhDpo0I5oWvKhOBoPhajABdyCvozsF7zongw+cogRbgcXwKk
Y/BbHMGpQFg9gAG+MLRM94NJrvQVHLBdqS7YPddFMUrYWP97/XxskSJRA6tV/eliVY7bD2oO5xgX
qMJVhGUfsYIhRT2rwKreOHLathdTf5WLoVLGp5CLVUoFMC+Cni2ujuxnhFtgNJ+TOFNuUrmq4z5k
oESi4Z18PUczUjGKDSTFc/B/RCdTDMVTvWncPnoMsW0+eN3vuf4umGGXrM+JTfU1qG8zxLVPuzqk
bU3fTx3F18XZc8L2Y3C+FE4TzNRHWXBda5fQCJBEilMT0fNFMeaJkHLY4+YgZHcBKIMlxfEc1+gK
j16qpy1a96GoFGWgqZixgMeqPqKLvuhaOFvT7Guig+yVnpTEywGY6PRz7R9FG8PZ22rXkA/caAMv
4GesV9y4E5tBP3CbXr3s82iwiaF9ayxtxNpvt1DiPR41mU39pIvsJjBSPusrF247LRVcxDhaxVvI
SR+df/NworvnxUvrl6AVyPtQ8CdojX1QL+Md7428kgFZ40r/li5ZzhvyjDZ+W3R3fL/pmPg2nop9
KAEnBT6DuAQTcHsaELvF69urfTP2XkK/f86SUPIVk464qWYF+p/ALUYkLKOUHUQltYVKYmXkFX9p
jAmjcpjHSWOdhKK+QYql3qTcKo99YlsME4XOBVLwH6ousnQ6SwvnrBJeRTImO7IIHLHFl/vZGrxn
zL2SUIuAQBAhzwSn414A/eEbSv5yXerm/IKVd+I+QYkq+Fh08DJRViH6+dy6yt/Te+jrRkEpkkqI
bzHV8zU8wnnxV5a0B0waXhHo9gmk6U/dQWxJY5l1RZoW5k+mJe1mGKVyePA1EnVRg1GkgK/Fough
pDvgMHegkGEKGIYpgDWgO3OTp+m1gAoYid2JDOX5Zbc93LiuC9xp9mrLyF0tLS7AD4Uu5iNVrPxf
+u2R20VReJ4iDiERh8QJwukEW7g+kwzP96acrHwVVlq+jdRoSax8wZFopbRy82XdD6qhqyBFL8pd
X1DVsQk26eacNDlTltA5xLzjJECeWvBGNv5J+jsT7OqjmUy7DJieeEGDYwHdKe9QPzxhLJyN9OtU
W/+4L9Tr6dDC8AS+qU+417/YA6fa7YKZ08VMD9VyUx42JJB2Cm/EmggVAzD4mSo+k2FrOYxtB8fH
d7A7oGDt2V3dNzXbkwXN2FWg2Y70IFuM4i35OJL+Vg+GEP9JGuhv2RTb+p/H3blYmoABnFeMUgjE
JsotR0w6pW8NRlCF/0w3AM0+nai7+rr+sPTYvpSPxe7w1Y4nFncciloQL0IeAPDY2K70XcM3kVkp
ZpuRhltQUr803xLoNSyXJOiIIm5kj28Rv7TD3UbDFo5kJSllHBlNuro0VGWPv86gwEr7W2zyAyrQ
oQwlwTl27zoaq9Xcc9jqRZjWT80dq+xQuXvbIYNVlXJCFMeGa5UfrkfF8/pCxHQtW0wof0wbpmfU
HLTwquOVriyJUOSCWNp/233Vj90WsDNGIOXfDNQBP9oJEF10zCEyaAFzWW81OycjEm3/m969GE8d
0fdf/+rLnDK8UDEpuaQf6DYazAImXpGHFG2ZFVtTXL59Y5JraU99C+BBt7x/NHRmlQGlMaq68x/9
vh3J9n9QFoMOYZc9KOROvzqVlmQj19ft+DZUGOnGjvF86agH+Gsb4qPdvnOinIR2E4LjMleH0THh
qq31M6+aMkr4h/Y/+9D44Z7rGQH6+QQun/cisjwcQfnOKlHYaZWZnxJz+A1ukqkrL9mzX7BDHlsf
9zYbg5vCo/6Cp/EDhZbROeBxL7CoiFYsOUJNuMZzMXyZFzBa//PPJKnWQbIKq/BL4A0P0FSsgyDL
9T5Z5L/k0bng8wmyzMc6+5ExSTNKyd/WEnHDrYyh+DyTAHOTvE/kS+kbkcqMBpGlMacTOt1J2s3E
GdAV8NxmBey7tMmw1A5VXIZPsCCGjXtYEmBpYCVWsmMxv2HvFI6BGGXYvNUEiLlyMapEP7tBVsAF
tsolxtt867q6xjQh9EaTfzf2ztfSvtXZ6O6S08J2400UCBPkq9Q20sIVncAst4Vk+8SVNjrzZxRu
0eHd3+7gTPb+138iBJUhg/0akn7zWBv5ih53fbaR6e0ZjM+jdUjekPst+Fgb+qoeUbROpM42ohFj
o7mjLEi00epfSQjh86Adgxrro4inMSXt3BcPJbdzS2vafpaqrOY3n8DFytBDUsCasUVhq9wB1XGe
uW2GXcxlSOgyig2WLsInEzFPnok8VP/4/Sx4M583wwOVq9tMZ4YoAbkwUVIWoU6luA4X5biV72wP
neEH9u34TANCkCQP8VONFcZNJX15sorGeFaxjqRA6c/P4E1pLIuukWaaQZ26AhJHNNlEPMfH98R/
e77dpUJkHpVJai5SRo9FCLtFblDVgkFeQuzTbsfn4FhtPOfWEGnepZwI2mmFwjarE+cwOEgdcuzp
nYjEk+ICpHIrLY4ADtyepoDFZ0xPK7D2dYJaYG/FtFJfjGu7Y67e0n6+o38+95y9gE2toW8nwgs0
fZ5D70Hog8ztU2KFp7Cr+HTo/YnTiOE3bgrOdZoDBAy+WfTnOnUX6jgDGKKUQF1XHP4pAdG27TkA
pQW/aCjgy6px9mQDHgmJFhn4vwAjLP12kQb+SfzhiI+buBb8JQ6C+VHfplui0VoBn2lHAQUdFHrj
uLB0Rl28Ia/CaCXCpcoZhvG1On/OK3d/IIGoecwt7xr7dm/NYUk/S1OLaDmBzasp+f8jtNW9Ug5I
vBfvhDciLXaLxAlNiExblkr1b4Mm5Erkue8CxE29md1+5woD4G4+biPilY3ZiB26FXvvszED8cie
GvYSIrE5AEzyxoC0l+rjJAD+Tk61oviRWPfgYVDbxZRd37fz5LepVdo45L4qBSPvqR0g6RjCyCi7
+ckP14OW+S/mQe8s8gAEDzvHQ+dSiKy5YiOBksHmr4Mjq4QasZPpCgYpS1LtmwEgSuEFk1d862VU
tEyNR1qwuOcfvCUS+vMRpiPg3OP68uyEI6fCAPYL1loKYZoEDbXGa2qJv7d2dFYCsdSScRhpQyZG
Ujge2yjmEZWJDgv4Wl+ry3qp53Ohpzwsa8ik/ZLGzaFj5PXbxWYDCwPmDY4Rqo69eclIDhEaQwSg
1zD/pLm0/RzR7kToK6ITNCYgjJS9lGRLBrO77Wd9EloQH6fc1OUQdufuTFqUhTK/jeXFEf9nbwY5
pF/9i0vkWji9TbdfRFI6Ml65R4D+qm2Zoh7O05fsDtRMUFZdkZw+n3vE1XsTnjH2E5WFLNsYxfDm
FzTIPP56rKYw1ewMrxNwVUZLRp5bBdmZ5teN3eefP9US+lqZ8IQW80MlXHrbR18ZCkbCyVlf9tl+
sh1btpEAMiEIYoApfrt9yVklMXIjpVIPA/l8blMFccCUzazm2e1PSoFIUgm3bKPyI+plZmhjvt/s
1KzS/5Zj1g3gx2+cFuTFfeppvRdRIpyRsUx9ZX3L/0sdKAQVBbRGC5thPAyVb70wXqldwHBY1ULh
RTwksOS/AAr7Q2A3eJFgLx7vSkudfL82K5VMthoy2gHpWTQdrBJGETl7Vxu8uECHqo7zPnvVsKxD
04b1sDBKkx20E70PlGmLlhCnb+kj1mUQTsj3f7bZOaW4LPddE4QD/h7dEj7lF0H6CUpAJBkKeNyD
bG+zLoOBnqlTtS4pq9V7HXNuuyGUO0r7MLa/eLXfbO1BV7xs+crOvlQYrdUtN7ek7ydA6pZJNvGE
+Y3/s2pCSTEssx/iYS+qJUOTCQHw2apUCRZdh86Cq3agifvXxWmjTLl9eHbVR6sv+SIvNLtzI4Rx
nWq88XbHjRrbc20PPXmfw6HUipB+qCFAphKsUd1XKYYE8PFZzCTRTPMW3BRX6jTADmMLHDyTuUJk
OcE/zPIxXrQ755UKb8eyCYdksHZkHfb++9/OXsgb1LIZNvJbWf1qbAFvxtTbdP55FilDEpPiMYkn
70CnJQRiOXemkRJkAhFsf36Uc8c2AOewhm5VeEO1hHS/yNvC9+38sFtQLDU34OHQY5w+HIdYaRdK
oqGjvYm2I+5K+YSOcQIuPeDDyCItDck2HdiZW7BdsqZNO0Sg50WidKJEjJRRiPPuteilDXH+Y8h+
1lGceRqMY8cEddmbkEBSAsO2KbLPcjgBgb3LOeP78WpDfPLlN+9k0l5ZhUkw4oHIqCSgTNeQy3Ks
JK9F71XVw/2icr4dprtgNsoo0o5fDHcmdty2evIrao6x/jjCK0OEpp4OPJqkukC1yu4MwHTvY3p2
dqhO+7Z73w2xDZ07d74tO45P7IByzD0fdBCzP5finw2gVdb6pANIL+Xk7E9fHmfyMa8XixvjjjVm
9zZ+24U8WlF5E88evHWCrtYFmaD/eiAgUFy55/E8QerNErK6HyBFkcgwqyrHpiPENf4epQ0gxamx
XoEquPIY8DpGcUsZATtTaxkf0QeBv/2R1lkyh2gMly1L92ty53M5QkYKveFCET3ph0Y1Lx46Mgta
fR4Ubj7wY1KpYwHcoA4CFw6liZ3w0aA3L13L+vbLfY+GZxpf7+D+shRITMz4EN8mEDyhPBIhjnh2
iYH8VBrCdU0Ewyr3BFDPKCUi+RP64pzRh3vf7yzC8qKxX2718JXtuutFtssZMhDB+jbIFJJccye7
3aZcYqhcPYGQt1Quh1MjuhBFZ5knlzDqwViw5v8tynvfxOvRm969puc8cjkgFvmeYMecqS1uAXVY
CBzGcXhcByc1qid7QkdO28UAn96FmZMYKPlZoSARoqCFIOtdj5S0xIehJr0ssNrIla/HiLutZLZ/
mZYrvgLswJE25nQ4cP+Y36uKcC1M1uspRX8KQdbetthNABLYg+VfCja6ldlG+FFsd64eIBbAKV/m
6BFO2mh47eg8ql1QNUXGFPfuupEPoHG5hBCPWFPaIMnipVJLYm7qkkyynOEv0usFohjnrmLbTqdM
X94IV98epPeRF1mi/Ze8v31gyN6ipFBRbMFRUx4LO7037f+PMU+EREtUMlCEl4yRWAxrBlCefX5E
RmOWWic8Cdyt2o/43QKaZnuajFP2B7r0EClH8lb0+hqpjgpCSUsu5FXgEWkTSh9cY8aqOIIw/iMV
MSZ9C3FKCKbvsZAhMyG9ot5fdnLOBDy5Zn19rArFCvlr+knWuo/I1n7Zz2PgKHJkwCcHBAnJdl9m
Y86ADyGn7cvnnp2F5+nV4v6N9NmssZyhivyV4WwRWnai1ay0DxZs6pjLRuNMyuS8m8driE9lCrZz
RkjQ0gJcCQDsYejYH+hXt6RL8QA96R5heFs3rgNtsZg6Tx5itWHNsha6LEnvDev0o9vzLr+CoTNY
oweKERRdYiD6kiYriKnazM8y+lMiF5Etmq5dItWNv0B6aTsTUXr2QMc9ym13BUj6Q7Yd8934eyxP
WUgsWg1/uIgvGG+nlLTb+e/ALvJyLciekOJImukC30yCl9rkF3xe7ObBSTZZM27d5aJ2KMvigCRi
iqo/TesZk+OArdoNWsYhI5GKcd8PeAj+ArZLtrJiGbl/NjuThSoOWYwUfH36cVoocliSQ1L4QXpw
TlZh5hGNbnTBtOxiKQfA0c2FlX+edP2iNZmnp54xROFaDhrNLPyKXJthorK1Mb9yFYdGnZaIvb8b
4lQRVIG+Mp9nSvbUjAzYpGen+mVnCPS2HWwYnFNn28Po0Obh6wAkyWBqiL2SVl0G5aApuDZ2ufTD
gW1+O1xv61GQxvUq8FSK5xGlmgqpfun4e1xo4pcCSHD81t1dl9M/KMmYe5fH6r5tGxZyNu+XrtbF
3SROeB4IVWTRyOKARIQC0U+0xmBKWUMbmFy5uAnvdWzaLIuPsDPh3DA4Hk5UVl4K+GlqiwMPZ69j
RLm7Ebucy5R50ukVlkATpmiFZlrsTYrheUkFGjjJd5gCSNr8V2UCUSwlAaMn/4bOzCqi3wuTehyi
Llw9S3mNFat4kX5aYCA1leZ0NgrScfrcR1clB++kxFOAb8n4B2K6YImptrePyFtX6Uo17QH5w9d1
ZBhCJM+mkEeR0DjoKZpHodD5T2DANkp2XPWXDDD9FnmhgK7gnqIogKxXn4J7vek2yFu4J0Ow/Kg+
54yNiXxFXp/Ph9FdVBfrsHWlky6nvDP7JPmYxccdVX9c0+8qA9thde8YdoQCzUlhcI6VcKG3fZ1m
ksg+5rARpM30DHCYLyoEkv5pBllk22rqgY4mOZwB9MJV11NsFWW9C+YNL4t+4v9bTFsRlVXe+7u0
LsZoi79ubZjm2k8FfiS4HFloyLV6SV5CbeeIUxUPwW0uTlsDx7EypwGvGIuLJVSeWQ5D1cVicfUg
j9RQbpXpFjagOZhMwFOB8yJhFLPix5QblszriSz1KQoP4TNj228GTufmacnpNlDlSOEcGUY9J4ej
XPof6FxZEi5Tsk4LKDfvs0S22AEFj1sRCSCWzud9yLjhDh3MPtaqS0Xj4mmaPVwVs/knD9MF39kz
vqhHx5jRcOcDCK5+dAgdKZ2mDy9lBmqPB0foQrRjfIlVWdqNUAdCDyxNiEml1noLVFktayLrH3PO
CRASbbUet516heJ5iaOsipH38z3SWVnCQSbJDEdWIBr0uNT+WkyyCNuvbPz9PEU0p6VYFHT+TS9t
KG6Pxc+/GWnK07g2G2224hJzGTP0QlussYebCtKxYeRwFAk9q6eP3g22FKqyFswLtBXcP/IluxHN
d60GP+cBheF3yPZ2jnac6jb32G6UU2ATfRLTFpElHQCjIGfP//6rhoTAgDGHt4pNjANy/GWEH+Ac
Srh6FgMTRjEC/9diuUbUjL12IstkzxvdhBH+8U/PQIyhgNBhDWHj+Z7kbCyYi908xhQC680292Es
Hgifr/g4mC3D3DUhLeYzmyXclk8fATQgAzRb7/vpeEiERAtPhNErbPhMzturOkMw2oLuMmguaqhD
ulLOIB61rlkVeUFuH6Sjf3IWdeRQaMrBph8+oKioQ84MbuQGXc83rRo6eyTY/SlS3YVspYM94frj
20Sv5kd7z5TtigbMkuGB4TKB2NWBtPLU/lH6HAUNqq3J0abNPcVkHQVVD4NXzAGH99FbEz7sGAI5
uclxvspgevPRANVkBylWS0Yo55qn8G+PWOUtD6vB3wwjJATdg2PQy9o7PhpjbgVm38ba31QxjJ8l
vdBwIbwqenznL77Ev92Oa+VYJBrzjxEdQilCgZ8a288cPEEBwcfTTSiJ3iu+225sS8oNjrwu9LOq
dn2xzK5kje+u5tDFMZG4kC7psiTFmG5BX2I1AVxHbULpv6H+ZXv1Im1eBt0N9mMOoVANKpxYmNFM
ZFDWPe/8wc/KMZ2OLfba6WKrCwalzTuUxbdT6OODCGZM/bveyDMRBfvVaa268XRXVtp216HXhGM/
u9svoki7gQa0EhBBDv0ABrhi4TDZO9d73m5qP3xNwjJb5xlXlr3ZOn6QcZeGkk85qvo5ZfoQ0wRc
i7g1KbcNOKM/fMl6Wsd7tseXRWvgh1HDFmAA9wZPWqORVWRDNajdiAw6JLXGZ97MMYo56OKxhhEo
WjxlKXwjx6zIPgoi32FyypW1FBdCnyBPI4WSnJMdx1IVLHHo3ZykC71kSaIj9p0fnjgfgUdwLdTH
rPZhW/V9QLq/ZvMpFU13B/6Y2sXeWuuOg6wYYPoR5g2XCVUL+n5ZRtC0TXg2XwmVK2KMIn2sU62S
NHhZJgr7uR/LO+bskgLgQ5LYspVSk5VppBsPGnHmfA7ljKPK90JvauHx2WKmbpr/nGn463VHFtVh
LezZM8dctPk6aZobxXpJEYfdUWhrO7W3dm85Qu6IdgjtWE0ghN5u9h3Hilt2Ak0Jc2vOFBCA4sDw
bd+n93u61hGnjJPV9V6OAgy3SKhr+icXTVpkTAdhaKF9TUbeSgy1yGnXgkt5FI2a3MhHtIRNAzLb
mV6dWMe+8YBpJE/pvIdntL/jLIhkicmFwwCLtipY3FpiNIohu5vSJLcbLrKrBcROQEEcFoILQNYv
m162RaKVqWKX2lyfFtFHlibllfzj7KP1BtmHut+CBtt2Tqf6NKI7FvROpjPxfCncz8Ggox2iQahQ
93P9W2WJYJxLkwo95oRhwYjMZ1tiAHYswzCpBgP7UXx0rJpPea5u5UO2b0KLsN3WH2ln0iGbbgrf
GduDzp1oef8mX4txOts2ByO0+Tp3GqlYKQs8nhqnni5JCRhmI7HqyZ1JvobUZrtMdPDcBPaB7NAx
S/2o/McQhN3IUeHxmoyx9BGtU4a7n8uJJZFysbgCRXhkd1zyNSH5OfkwTpRSJZ7816769quZh0Ar
G1TM2osfEK79jlCenbfy8xjKuSorai1yhfvEoqOj7j3AXvT1XPVdhTXOHUFbx/uVlL6cZl46YFcM
6GLpj/RvMtj3yeHaDYmD2JW1m18m5EqK7444myYtWJeLm0xCTfaMSdw0X8943drsXrJLI0Suttld
i4M8IojIr/jXmZu4yja7Bs2lLXNZiqhvOSbFQH0E/AM0lzlj4LodHTEMq7u+8ThovxD+us7Xz20h
YhHWkWvPByR9gWPZLxxi8t9DL2d0F5QcdWr69jdaeRv9eryF4LVIV4qTfYQFrDaQIg3JtlAqrSda
CkuQUVDMkfzaP1CoXnLne4GASr+g5SiKVOY/RTgAgKZGCLJ+Tx+X11xqS+j2UaPScA2NT/zlriNG
cz6N1i2RKOHU6nX+v6jyXMmcGqVIpHo3J60xccFRZ/nRWM4RpGQjOqI61VFaHAXLlvwuPaRo5u23
hhVPBf9CRbc/g53goVpNwnInea8r4dGDvJNlfD5i9jeo/RzM1C+bG0RushtMZqj6auBTrToLxiUU
IdIG1chAz6l6G7Nn16HSthVd1HgbUr6IG58WQwPzT1L/HMQXgtDPLYZjrkl0IkXuBJKVDvDcLAma
3AP7LcwOYjtFgJwjSjq/q0vMQOZZ9ZIRyempIBDXRm4ET5wjMmVsDhJLBAESOBF5eBjuXYAmwFwV
8/PyNFzFYaBS2xn+7OmePUwdrW+2q8xpuhO9+VnHL1ebvfiTO4dYQDpvrUKpBsU4Q8HYfm6fx4xw
GFNvKmNT3zo7jaWT9gi3jgUJlbUYyqd+7WJT38ThqFz0yllX1rnl+EXngp82D+mI78o0auwnnKw0
uB4Q6z+F04qZ6omlZheL3qBYZRVofWWGpM3G9IE1SmCnUjmglS7U6N9XVuGjIA+daJ+GQ625LqSn
yRWEzdR41mNih0zQUvTZ7Yjju5VmC0QYz04vNvWXXXQMonZBBmhV/o8Cs3fS+xaecLUs6fE6cdre
Z5795RX+thgFPh11IFN1C2Jflp+U93TBMgFpkOStIxKc2bc9Ysa6MjItyzumBisfqLuJRFQzdk38
Zl/XAFepKIiRNqd4mK1+7HrDaYta4kKhGlrRrA/7qvlVEf2UrqtVthzGo+uDqxe9b98ZRft68Oua
xdM21z7rnlShurmlM/5BnZX8zTEk2KwG7aVAZo8IKCaC08PATYsSvmvYE+x8J+NGiD8pDamqx6gk
Yz9RMdvE/JDN6+pkQex2et1oQbFR9xtgnGDvS5tDeDhwKs/HXBRRDNuCZJbdKZ2GfkWJ1aPslHff
i5oqZnLGog8ze92e1ENz6PIpY6KIPLeBd48Hn2HC9W+bQgemD24ZGO1KmOFJuK2CslRbnvVcrfV3
+GwpOqrIuLQp+FVGx70s9Uub4JH9KvpV1QqIEYYPD78IRZ/JqGFhTLqDAgeQd/t0IF/tEB2mnNcA
qtyHgOStajPaAArDmGzdS2eMj4pSmPhsCXCCvW+1KeUBR4QplDy/dzrpGkZbEj2cn0nOZUAhW9Py
T69wnEMA0XcXnEqGpM2jCS4qcO/rSf9V5VK4gB3Hwbl8+NHYHDXhjn4VXztvMkzIkrVKJoSxPryq
oiD4lUixC8bYtO+dsAXLcOGgXvMRguN20gTEnqIHYm6wl/7reeuxDP4lDJe1VICqkgFtOIWcyp2E
4yP1IItew3FKZugk03Mq8ewKjZB0Et/z4PC+CKO4ZWKEI1Z/Ks6450AjmWgKOkbXPyAalcW9pzkb
XmIjdSrNAYpU3v+lP6nuWVFGFlpjVayomd1UeGRZBQ/KoUOad43LrMAnLINPhBDnCZhib3ol2vdE
r4vButwIrVCBaKuKlX7NHNZCOSRwGF6ECqAU+edbFmw9Kms1WdErQGzHRRfi9Dr/pAqQeVH9LdzY
AC+rtpySn4qUGLLh37QvaktbSZlLTTqOSbv2ZowgyPw7aErjkqv9t1mlX8Tc+OC1fVZcEqLTS+R0
myVPUrH5A29kQO0aCUxaKfsVn5Micrv9zPt6wEJUw4DnInv/xvMO6vApRwMO+yNFsK/lISxquJv1
tcHJ4VO7W36rtxegdn9I0DkMUON15Slo0BBAseCYdTN0EtJQig1MhKzeTLuJd0+tnmXogp1prkht
WKYVmBF3B3OXrEgoRJClw9xfZ04HcnCvDHNTYbofcOBBfND8JyTy7yg/JtvSEDEY5eKCAzmO7uuj
LMpNxXQrgmPs3+aWuYJI+tY6wLly14e+N0f0k3CoaR0OAL/mGrPYEJSsIFO+g9wgaKVldk4vcKJR
8WDi436uz4PZV/fZTLnrZ/6BqjAKA4kIealxDjZnpfsADg6Ty3sPa3PuB7aZGn2m80YwkWC9FrW2
/wkGa2vdVcS6LG/X3YYrVHwGA2Hik3mvdqpqP9nAYm74/otWbkwPn3WzRUHEEkfqqpEgJZd2IqV7
LCZr3eXFI7KJ3p51nmJtCMCMkihDOAKf1yvS58VVE+6cWmMjiqhKLbrI+0C8r7yjpZEBZgxrrQQQ
Bm/OgHdPQ2vL5r1mwKXBqKwYVJPvhMl5eYhB3Mg0KS0NnxiHOXY5SzrpLVcTZpvoCSHtmg/HPrEl
E+YtsA3RMFu26tzyjY6g+0dWkVOHJMlvK90IyYQAaBeLQei/Xq5vA2wH159OedXxho2gC7peRQcq
rBC9DcHolOmgtZmzpK+hWiXlHQcG/Bjku1wIv6nSJwm5hn+KktOMawUtjTemNczKQmv5MgvwyZBf
nat6dOD3cy2s4DMrccYs7sbO0S0eerOgIdzg7uU44O0zDrIr98xtr8KqfAPi33nqBOGu47cvRizy
dKBsjCQuPb8S1eCKLQm+zfET5xHnBt78ebU4+Ec/PXgkLRZbbTvLyBZ8Q90L8ZkoAXAR/UOy0F8j
HK+y4ot69EVw13DbLQt5omjnJ9oGmTI/QDmiRk+ZUnQ7KsowHqh0w6BxywPPa4tCJBNZ9k1IIiYl
1WKe+HkkEAle9k/tkciWKciIdjSseKllKwOtAmmFf4yOHD08AVbqrF/iT8PagXuOzKiQw1xBqIsb
kt2QXk+vmznZBRr6ERw2o+kyAA5xHXluwvsJSIhW/jD3va9W5kF4EmrEwRETH0cRkMczsEe4ssZ9
JkxXFoNmvwj4iRBTBsKIpleqb6MQ+tCYQdWMajE/eceN3bqAs5brvYPOnf15Yil951rkQkNb61Zk
GLi/Lc3s+nE9bn7+OJsYH0XIKTrjyuXlXGlhe4m3xLA309IMqapcS92wFyKj/KsjO0wyv+7Nh71X
yFSfgLo6cpkVNV0PCdyogzeAZKzyuCcN5aG64V8coUIljHRmRQ1AcEYjET4cXl3Zm+nvznMgo0al
h2nA+8b8exN+Nsn+q5a8r2ouxN2+hptZlA2eyRqB9YzXj3jSAMwG/X7WFhReh9FyzNqXTaMf4hje
g7QbFXyTd8x4yfv9zoJpqxTG4oWPQO31TCRy4vpzsRrBqIAPus340UXRZ/gBgi15SYrYLhoHsxGS
5fdYznScLxmMonnXNfR2DRN3PKnsymmfI5n3xyGeEi6E80b2O3UhP/7aq5EsKk0uNdeEVF8x9Zvx
DiucercuGCMnVK4m6pRkA/UZAzXyZUVAFAP+LSKG3Z9xHqMWlev5DZhf46ato0OfKh8nl///786U
KdW1B/jQSO6EQezTMWyp3ob+ockPUG9kysreEIAzn9DQlX3rJ8j7pb3Ufhe0iiaDyKmg3kPoGUOE
3zAjAi6wUPrurygroVZeTx69cyBC9yeZy9ZRoa/CNrhcpVvySnoeIh89xy+jfMjJy36S0lhdStga
ficFQCuS3Yc2XPIbMGmlf8C52hYh26mJ7clMz4evPnh2TDw6+/4Z/yl7Jp6nhSAVUbjt8rkvB5NX
JvC1SeLzEmd2TsnLak32bpf5heMqkySXOqUCY9+EbMwaTyjHKlaK7L957hVAh48zW8C3VqjRYTa8
2uaT8S8YujjOjpGgg8CuRGlp7t9dIDDYH1NCVdF0Y89NdShKYaly7fvHO8qNw3muTh5euBF9TaPJ
20LDZaNJsfXP9lxLAELA+pPKG9l1MxiCmHbLjeOj7l7tt6T/jhr44BU4qY3zEEjF1MGuqcATD3cK
646R1bKTP7meFwDuVlB0HuYCYlJmxBoEZPPaLa+/cqBxh2GTj2Kg/ToRsSk7RlC+oS1eJJbScE6x
z2hzvrApAAuqTnxY35of4ZhVKpZCGKXjBxice5Uvh4169V0+0A2ajlzO+wM/15qDdgcS8ELAsX6c
9raXeV6U7PvesSxv88sGXbq4gc0LonSLD+jTh59hUotWQajs1BUDbvIS+fVMIm1lh+wqwIwPuGJ0
/FR6mfUCfR386kF66Vqxa2BkCsaQlxtTcrgnOpOjK7Qo+/zhIt2tOtSgZd1egCMDb9J2UEy9Jmms
MXquQSUElXSBi/yRSTAr0oCwwWHt6OSbl/7WV8ghZFxOKTD4T6IUYa8Dkdwgjfwm0AOuLdSBJp9A
IWJAbd82TcuVxR9bjg2KE3LPLKRAgCxDqSWGhfQ2WkXBcpX1OQS4Bah2AOnv0oThrHCOxy5UH36x
oB1cAfUmBLHd9X5yD01ZihFhxoDzz/2IkzAEU9hdaWpP4tqhgDmg53KOtwR2kWDqwTmon+Z4VvwB
2NSk9L9wYMgn4w2TSvZ0FD/HDGtnz2R9rkcnECOIBDR2Jod6JVy2pAPMj270gg52a/EsZZqje2wL
pZvxCFAfIqn2TaaaqYBvqKBZzMeSLSdlElaGm59FIG5P503rx3eI5+i5GxZckun3mrIlvhISPAg9
n7gcRUVh5QxNZuZldUZkV4ubfPTT7ZodgCi0vBhsazAoKJJBs5EPIy5ppSXe2G4Hj/lcJDLls5V4
n3aAFNeNomAPMcY3hMKIKDyfdctG3ECqPNxAS2lQxm7Z2C1HBBFYTO0EqLfHnQyiQuTSbWK/rTMc
nayq/ksN6vgRIxQr+Z5MsvwRBU66uR2WKgqGvxvB3WTZoyxj0ZfMgAH5C6apX0U1M3c4D9LyjarL
Ct6eiGW+NOJFWRhMvO5PdQgo7e8Row9i1tXMsglaVxJzUHdgoG4z3EBGdNESOD8Hwnx1OVKWSUnm
3cLj8i0O63/Oey1p6NV3bX9qKEHM7ga5dF4wXEoH5VFSnNGcFPzFkhSP1U8/XjKsKf6B0+ng3XxL
Vih8PQrWOOjaIWgb5M9Sxeqk/ysWQsnaZbB7HNLxCn58Pejw9Zjjgi05/gKrUoMc5qOr3Rq5VKiS
pZsmV2SRog/hS4hkHMdhQv8TQ4JoJ81lc49BlCn+bhNRr2QdUItE9UWHcf2dxwcHatxNxuQ/yZFU
VK9YGZ0LlV6vuXiqLrwiOMPWor2iNdERZz7kdsvQN6qeaYn3tLRdfgR3khZnffYDvIQyKGF+Jk2G
rnHi+MEodYGRs/MGu+XYCPnlh9EXFZvUeGCYzZ8GuffwY9FU5zb1S9qIqtKDXrpZztD+aZgtPqvQ
IqOHogvGgvary8+I0N1y/KICmqRCybnCbwpK8S4zbxaHsVOJEm9PgFRUOj+m6IT8wfGtaBRDsiwv
/TmOqWXttJcgISHpChbrGU5/WEfyM5TeeQmmpJKGmRvJvLZgUqA3MCl8nZB5/YlLmB0/jyme8Lyu
FPzEaM5UyCCFxiFpCzExrq++JN1G2AQZGl/rnoXP1IERd6cCCNWDrwb2PA44iwMqfzKQyUN8kJxB
ghdokBUnvhPsQ0GSBx3mo3XfFIWIk19ignSlGBh5JWuiaeAMuDm7PqJ5PUFDkJQ8c8ViZLSDyxlK
8+s9z2orpSM471L9rCFHvxjHziKWcTgiY+J4SlFMdU/SNK+UVizEoBq0+GfC6j2yG4yQBYaeJ6/i
LL8m7LEeVi1qhVmQ5cOlhK1TBNAu+icfaup+WSbcbXbPSnBMxp++mGhhZ3wmqyTaaW1uuQl4gyQC
zOq1ebzA3vnYR/EFX5nzzgR3xxtKgJvE5LttWKE3IVcTrVSggBe1dzXN7wQ4NY0dRlwQZuk2gyLr
o+2EpXupEWNHW8qiBSq6mW1mI1tuA4i3hVmb9GPVcnDigLxx7DO58sehlXXIsTYdSUh6tTCWCDca
XhMXlngcrhOzEmqDQx749EJxG7vk6uwW+OekSR7wyf2ivAhcBsL0aS9mF3uJtWzUQ3PqOP1vyJh3
uZ6dyMyeYMfXstL1wdDnwg2YlXjqlJXUfZam1V1G9kHka3LBqetiaWb6pt1bEv4xBXLacbpyqy3V
hQhP688v16K1M4YvnnCCeKRT4Pv+P6Iy2xeqxqVRvGHBQom0rcJdHd+BfNO786N/D70xtya5yAJm
AQFPLZWXyFTLIoxFFtur13aidtZS3WQGMFkijA6qPIe1zBBEuZJKAmNm1qk0qVBNjkyxia5vZIRC
idulG15TLaCyaWnq0jhRSbTKZczm5YB+FBAEygbO3J8fbFLbjhBc7bTlQ/9O5LJ8hlRSrw9UbgVe
Z3PV++22uMPbXJTzq0IY/8FdsYyCI6VdJzKcFtIeiANXNRMCbtEnzRe3p3dnQre03w2JsRzWNEXu
nXaW0PbZgXdzoi5+28w7S4l08OD9bAphDZZWoG4ukn6m+8ABi1//k5ht4VvZXgUBdN4zeg64LPxA
FpSV4/Qwnm0lXEJqjjKV+hEoHydkWRLmFR8j//vzCveDMCHASi8tdcmCEq/T7tkjI1CtlU0nsuXu
b6dnOxgDr93W9nNSzxb6GlQ8Qa6VC+hRVjzN2NqUVoDfrM7oH63w/bHgJ4t5Udf7JKsPftomNHnk
hlXZMt2bYVTYxKS88dFxdeWr74PWea7OYK6NcuG8U78UL7cOreRuegqc+GIYKcd8VvsGJw+qQA8x
zxOWgTSMMV/dqFX9M1Weq5jojeZ/aZX+y9z6pFNpUSiI1gxqGoFP5qlCTJAILVE2JfSgf1t/GoGE
MULhP3ql7Do0TQlFjJTKrbE4YWzOgMeHCyTu39QCDyAqHpgqWt6kCLk81VdP2urSJsB5yxqoRPHn
qf3BqZjYkGU31Yyt6G5DX3plGQwMfUxULAYnewTr13MjB4Xd0IMP+F12aXhENcg5QWIIbVjv6tsM
qRuqvsEPt0Ea6rDsb3RMZkJPXeZsgQSBqwWq/Zsep3sHaceRXSJi6lwTbWjGbQsppE40D25WD7wR
5mh8O3qcNVlEGmeFB5GK/VaKUYIKMl7Q8DXiH8O9BoHtS5UeUyaBYpUtteS9o8iHdMzATV9/wECB
m3Zs/ZAKqk2DqlIXTy5wp0bF3UBkWImXfvVkiPG3uXosYCyrHLle8g58+f1KCa0Y1MqwFSVAOzf0
wKm81APpyT5R0FK1OSWu+YJXyWOlCp8aT5q7pJhGyqpPwJa0vJ6pziAsvh+474sGnjg3ZoTzhxJW
1+e879XBF7PqIls3EYgrb4nN9SJj1KzdPdTsUQCupaMHqV35gvsiiRNjLTO8E785AnPNBYTQ7t3v
FISQfnHUEp5BF7DCJt/RBH9Pns5Zgf+eFDAMykmI7ibjbKBudMUcPeDcLA5eay4hEFn4ehjSWkXa
T6pF8N8LeB7MMkRgRa/3Cpz5dtFeWCNhpLh3XtiENR7YHuSF4ZMpC2542oQBykbrVd38HkAAvusC
ycsrPRbWf4vjTGSWvA+LcNfMqB0fcnZM0emQLIjZi7rd9fzEupXHQe9sf4oBCucqZDYrmK3aR0D/
1Xmu9ZU7NzwiXM7i/gllnSPDhUj6OgO9FKhcw/4MbTGM19STJM6qzXBZfNJ6Kr8KODJWHG1JWXNI
babls4zq420jv31hxSRcPoAr5uuJw72QR/DqCHLcwsH3r/iAFIBEKZZrvJ41heRY+aRF4bOhfdex
QSBhkrHwJD6RbLBPdW7faGBxG73nj4xVxlfgBG/D1ZxcLtzXXhfyVitsDgluoBm4Zp6N1GNEjecu
NmpTl4OXQZbVHA1hLHrF0L0L4M3ArPAH5vst+XVxeUatdvC+csC6RisqU0bSlq98kcbH4NkLlrux
vQoTGETZlbC5gsyP7VkevApF/IbMsKtB3zXMqU7OJLWlDq1uHV0TU2r1RMn5andnCtgTMoY7dQkm
Hgvcq2PRikiDMza9uSAQsm6MV230YM3XjCaVoXjwhgoIp5lYH3K1tR3DuEpvljRnY7PocDv0Srbu
kZZlgVOVHPgFnCeNPlneGIeCvGYMyNMNMGeJ9v3Ip7Tf66w7QGKqC70clL+efeBmK31/ZRGgUyFR
oI1JgKyoCQkUt9OYQ/9rKugWjs3AQN4Ar8xA4PO0WKA67u49AS2H8YQfB13Ge2CHnLvTjnXw2xaC
s7khqEUwne3o+zbNj7/xqe2l2dB8/4RGQOtoUFsyyP/fSxyF4pdLq7w11gKs5xnSeeSvQEFebbPW
txwM6HIRDARlZdgf+s44z+m/l6Q1sjhYJLethBWJs++7AbjrdGEK1EHTAaAz9RweWRW9KGHCaMNh
1qAGt5rmclZ0pfiMcrBOCB+9gR/dZ+P1efxKdzE+4GyQaoTWYr+NHrGFwoc9LdqA4dfyyfjQvoJ/
KKFBPvFAldOzID0lwvDLItA6i3axX8uyNSJfpmztn7ORMmYORonXxVeTGH96bajO5Ab4WXkQx6m4
5IWqWtzLSS8ATmrN0Ehp8xE+lSj3w/40JUn2Lq7TG914lXKn0uOE77q7SQfcn9o3VqiKbukmCdmI
sLL+wI5iDhVEhFg8d8RrdV1Bb3FOZBSoy4AMBusWqlg1tXMBLwCBqQBsk1TyGr55x+CtRmPtkzCQ
Mc951E5v7LJ1trsjNqk4pntESe/9NndfX5apF3KvRsFXHZaR95q3rJZqHoS70uOYjE1kySauz6MH
hFQmjOaztDQqXuGYjU9vR3c14bo6hdZWWZ37PNIU+XiVEgNFGc0wabkUGAkUHWlj3ACckiJhWH1E
rGhGrnrXjyvuTMTgz3HJlu9Vueyqbhi3+bqkMw3JrEhC4YaBPwuA+0x4gXL+xxVQV1+IA8oIrRXH
6IkOu1DC0ekwlM8YKRFlxBgLqTNIrGKmMvx1C5JGIIdXm+pEkgpv6+TXjzvqQHR9VG6FXXpNAtHi
97wlgu+aZZIyROSJhHoGgEYJ848MLY8Dyx2mW8nrPjilvTSAGTrBj4wy84ZyJqCWG3sIwS5oeV7s
ZIWaOMldfC1ASuZPePWhFEHARJxufsnPWXuyEALiHSH47vg/TXzDzjiT9b2ocx4HciHxZthgiGsn
jfiAGUoaL5yzasDLDtWXDuFnPfbt1uUg5ur3Zw8eYMxT859+2UfEg7YdT8lzqbod/N690F7S9Gat
fPWIjPmfsb6NPggrvrkNYvcwbNC6+KL4PnT5nrtIWsnJk5Sifhr0IJaVpVcgcrfYGQHaad2i7BLW
NUdP+Jz7wVm+p1+mEz40Avi3Og597rERkAfOU0S8N9xegFF0BKK8+WFzkPwDTedL2C6NYR9eroM/
8OUAeatFjVNtUgaiewyESBSVTev9uMaHd4mRvIJwxc6NWIxOzStxgCgbE0JMK73DxUK88Sv9g+ft
3oFpYzmBgQOoIbQsl+4yvdk/2MRluASbVcHUre/SBHlsOBI0gz3d51bx8EmZ0QEuqB8mXhgFV1CE
YZz4bC5EpZzrdOKcug5ARZ4Fbqaryk05W4hkuhEvz8+wuYqL6b14Z/++syB/qyF9rh89fkg+uDf6
sCSovslGtvM4Pu7U7XrD45F/L+vr7+KBKm1HhgBsaOmj0CVu3LFO2mKh2aXJxAl09l4QU6u5EH3m
NmoeE6GY16r86EXoCMEvTsRCR2F3Frm7lALY89Qc9+VIQ5mfeKKFDfA9I5KRpkoXdy6ReL35s9ns
FHKDvlctvLkkogzCBIpc+EBoCYFkse1El0g0BkELZyWHYQRXvvMo0ZsWXI3qab//sVzbLHcCdVBh
KllSzyD80UO/xnPAJ0Wy1UttRqv9vqZ9ri8V0XyaS8iwKnKP6bHqf/9odIMgRVwCKCulrjMifcqg
jlC87lo7Oja12GEfApqSD1yXlINMQoEO/RnEX8zAnr7k9JIpngBcRZdI/L0n2Rz6y9QNF4s5s4XK
ng8nozMN5bTx1EqWaSB9RHSqMwp2UwE1d5XXCmUswn5R3nR1wfAU+pj/S7wmj4LEdm5AIYkRgEIq
O3NvnX1TU9vZCyMhmuywOkRuhZu2htykWeSc8+XbzpSKWp33PDkdXOJ28Az2ylqdDzHTu094J2nz
JubAVMlKlDTKMctS2T7UKOnJsYnfhiGZqQoPTnplRolYIex2CJ25XEK53J3zlgHsONU62j6dUQNC
gAezC6stNwc63VCo80OS5nv1hS4zES/dKhZZd1W6NVZfadjGUEEnEZ6utIjQ6PDI9vvvgxsB0t1k
c/WhwHQcteNWhKhcvZe3zG3C+8iIGiVpiAW9XhXxXZmkhX9qFes8QF1O16FQC4YBjh28DL99Igph
8y7gqbEkJMtCwpDsJjEn0kB6vu+Njucx9z0vfZA2ykbd1g7elAdbzJPlaz4oZl/j8REASzxujudT
IvizDtNY93tJly/vAHZik/G2tES8sa6pU6cN18hg5dPXieMjaU0PoKtyhADvVkSCMCUqqM0g0rK6
AJBTU4awaoSFE/HnmS8JWvzCmAX2u6pznoQOoE+YxDgewqCY2h4nYXOiIOpRTJUiwXyGnmOTiOl/
+VwnSTwCKyBP2Rds6JZRu2TdvEIVeD1EUpAeK/EclVReNSAs5IeDJ2G+M+IxBEvfaePQk4fxmrix
hcCZQjPVBcoIMpgJr5zH3nkDRyc2e7YMCxqt2GNd/Sm6dD3FCfASbpLMEGh3U/9Hr2Lkq6Wuut8E
P/w6wrv1cp4XHVCYhQdOSPnejXB+lfbg7seLGAA55iyQqbfcLoIowAS1xLkPbWsGVZq7xQ1SH7hV
Rh+S/a8IFpG31WSyzE/byBIgKOT1P0aHyjZR2ofbwflz/piecrbKxGkurgnwzyYywTTxtCxEOD3U
sGtrQLXm+apmlc/jDIqSm01KRqVdSd0/yzeHr1dlV5jQKhZo8RxvYTwvq1GqPbdUGZz1zVLn68mZ
If5dxTcOltMFd2wTbfOp+2IaS1RIJhL+zH+YPnM49GvFp05Y2TPFo8MtUVb1xf6B+ffez4/hmu7H
Xphqd8sbiysQJVZxlbP2nyXWDB/mVcu+AVluamGVVhK3qToV0d1tQ+DuBUdkKjLyLKs7fNCn8w2H
QpdNuUXEpM5kfq32KgNd1PVTmELsYsBVPmU7wDxaB6fYcXmQc9p4bJj4oysoEW7b36o1whlDwdqZ
wHLd7cop9Ql2rHbC1AVZl6j7UTTiPBzJAUY+jluo594W2gncY05r644+p8Bw0jqppeatdLzLPnEq
6wXwGM+YZkjJeUbsk+hFW+ujHpc6RQZ4oElewuUL3+gwyDC1fCwTlMf0LFr6hu6OdyGHG7XPtbFE
/3SssG7HI+FVHK5QuInanBMhq7GFEA6CNH+LrmhCg+pbx/6JlFyobVR56ePv16oaCfhyiOcg3qy1
Tt7Vcrm7DvgBbPRh9QdICWWC/I9jdsERgN4yQ3i1elSVm7Va4IJ38/taTHDAMBiT4y0G4h20oVDJ
/Sjrv8UIVp2oCO5p06/qLnPgBcvfpZJFZUYHO+cG5eu5czK25ar2Xyl9YQAFPcEkaM0yc80eTJ+v
InDMWOMpwW+TgoC2EFhJzpfJ55opoDIHTyu3aopZ80oIGSHKDeJ6cBcqIiLEM7jehTMLM5p8yJ4j
C/O82iNhVArV+wYL8LP6qZTvHm/wS7PgHNMwisQPE95t53XEF6GnOgH+RMKU0DqLGKoGAkz7CHUV
MVkimUxXzngv0I43VG0yqph6yD+3neTmBj1LABMyVnrDoz0c0H2AuwVJfgIRTzJ4btgImATVxZTH
m/6tBovJMOxogXTQ4g3zltTPcVbEMNW0bAvmNbasaFD40izpBBT93iMj1XIV5IJdRmfJneCRs6GW
MeqU8BAv1pawzbw1JEit7R7enl9vdGQgsU+CaHvoeXLhVCnmsLtBbDTCgc543YEfoT58QeFuzT7M
AMn08orvTyP6Y/yxH1nPoXacnluJyRGf/GFcEl+B7iPd5Gjn2Ue8umdt/ecKd63AI0DS0mdLb3bz
+V3LhqHWgBhfa2RLOHyH81nOHPAVGfW8srubkUzxlxD3xHs4iQurGXpf0dJAlMGqwZ93uOb9vyA8
Bke3+DLAV/HcKRmW6VrTyxfuqbMrPol5GrRreGqWjxHp4N00u8soItuwsBa7/wvxMSG1ijIkNgvQ
cjGQRXKU+J6ufYndaRuRyOlMqbwL2z8YQb+uQp6Uj8tZS+9f5/twoofAU3BKRT2W4s0wEqw8S/5Z
UUKvhqki1eex+nNx0ysBIJnujRi0D9pB+86vLvPd5a7FUanK0Z+CYxjWzAWqpV8hjv9nFjVhtttZ
x6xvAAEQygJx9WeMVR3yjh7jsX55kIG4100W7op6EXYKmEjm/TeTfjj5HSVOW3OgSQ9ZuUziJr3r
a7PGX2soO2JYyCCOAk2WnOFAei/1o4BFJlOVesNYKqSIv+0+E7AKHab4T3QOryXMj4ERJOcb12y3
JGRlCpAjNb0Ozkl6OsZOrZ7CTnhtvGyPjpYpiAtvi/wgHbGtCNkwGSKwtVcoQJLvAOJYSXi/mRBz
xa3Y4xnBb+v7qSBQt9d8PemnOR2hS8UPcG73+Akjjc6kGm2irTx5cFk025X+JHqDmpS0H/5t+6fT
q+p4pPnGj0fBBQSNHkHdCPxXotSbZNUhzor+H4pYzLrXkLebzaKnolsdocxp2gz8o+qIChnRDYqH
K3CsnpEI18r2Nb2nAOxppfzYQRGZ6uBe14KWj05qVI7KR54RbBeCB8tipX97iHjiYr4TJzFcMEe7
4udr5feodKo/uyjW9Li9BoTrNWXRQptxrKgsP5nJOQ1CTTLFLoWBkDJU0ng4cVpmgllxaDtp9N3S
glCcZu1BwJU2+Q9xrqmy1qyVb4aVvVYsbcL8mo73JtZnp1JxjKKfSFUwD+Iz7raWHqebs0/OCHcK
A97+kZYRjVVXaP4/P0hozIEDaKJm9S8uEkmxdB9KPCsIL7G2wrJ2VJfN58mFOCfb66TQni/jntgM
xDbawxJRXpO42habbICNq1Zqb9e1MFWgC+Oy6BN+kYs0dlhVjCHW6Hhx/eyL9C9Z9dkrjUjNxTIT
0DxfkapZsJAZmDlAaqz6Fpzd61XHOb61+vpFsGQRywOxTybWnd4TBRIAHG9Eevs6rq6O+v3io1dq
pgYIdlRnhlyiV/MGEmZXSxy4WitaN/vBpROi7IWXvqCTiJ3ZrstG4cL1k0Q8w+9jI6OlbUa/TGp8
th3wYsJ1xZw7j6tc44l0y1XtoDNsub7boZzoX6j8KS871rnAEOhmkMg4Yxnkxh94k2Jj2O4Z0Mbh
hNv3czEaciMJ4aQ5ex57oYoGhNi1zupPkkV+vfwTtmT/ZadqLMoCedsFTPd38mG2hpi0bpNXMIs1
26U5WCsFJCp499s9ZHXXMFGfO2oA8SLArjETTPYbHrES2IQszXcj7kWJoueHIztqIQpACfd8lO0T
LtQotnFJ0k/gR4oDmmyvRvKhtAPebWOr7d0rgUGIia6zi+FPe4TGV0yWPZnxDx7XVgL1mxdySlbF
u6kaw+ZOSrEGaC1MSGTeFmwUa+kBURz6MEhUTC6jL3utCckTXoloM9noD2/2eZNLlhqb6+WDWwAU
89hwPFj37CE7kAl1exTGgO/tD8Ob77WfeP4V2wMsDtOebODUXha95bLUs+UV2tB7Ivr7WFPVn8pC
v8YbxpApD8DPYzSFh/ENEp4jzgFl3qoQ+63UvCzcGVWRlEg8l5ITQDt1DbkQ3eSKVqH+ozt5lDEr
yvGRu57CkWaRkAUET7gjnAit5agtEf2rCxLv0Hs5R3Tsd8l8xUoSvKpAE7IUaXRWDCED3yta/dWl
P4h+CHQhohsAD0jNzeTPJT6dpzE2H22KtyT1EkWWZk5Yf+KuF9Rhy6oUtZKcRpv/CtrWd+1eKOAF
ZAraVWilbv/BNtrm+paBPlJeD1/r8FNbjz6ZSCR59pwtU4BKU1KZFfuvVoQ2k7maI81j9Oos3vuC
hP1cXcyPocqx9LDl5cqDnakNAAQcd2XP+LY5/N+MYYP4q9DlKP2NxYAF7eJiVD6wC+Ppxiw9QPAQ
qIXRmL4yo25zYsL2m/7Iakj+G1YkjiQDUnqch9cdFD8dXcZw4xQ1BnRiEqHVKoyVhZHoHgTIMLah
KYDo+tdMwvI4G0gy720ss9oMRYfW3WhDkof6SKbUZds/in11Iiux+/OTdivv/Xn82qudzrUPtLRu
FQfXcjaL1CXT2c+1OVQf+xKwH6DjJ4aCLT3XAcK1PIfE9JEjlyOLYXmN/jwEh3lctzQGwwnSMESk
OE61nICsGkbhAyVyAFVyzMN+jtq6NRFGm08jmlL6t+kqO2LTlwIk4MQT7w5bKnrmVEWE4PDO2cD7
ePiBT//iz3fbgSeGeaIltUMmoDbGzKBZCFWyAQirLMlkveAmGfQ5YQLPy6g0I7/o6rLH4i8aDDI1
OHweSV/gizmuC6IVIRmXakuGMe5iJWTnkfM49tkMvcaEvelZZ/xEyPw0ZkaASCz/yGmR8Od8887s
raEDYDGMuoGMsxft9COzkf16QEfc1V8Kic8THiWrByYQAnLoMJHqKoNz+8/pEGR1ZsihrnWZBW5r
D8EgxVldqMVf+I2HTKh9wdcnQOpCon38FPQLnLcA8pDTJEbfqJlqW93wn3lwDIyMClrELtQNiOi5
XQkAjg1PPhZ51qMXw4NiyogMu94Yludtlok8KSepp9f4BpvNP+mxXNQdpv5ckGf6DzDNRdou9umu
wWfBXtXANFwAQi2pLr2xn9UeNCShHu7H3j0ZSwlMJ7gMRX6+ghRO1eCEZSSP9g7ciqBhNjGEeAK7
bsEHtmfv37zeF63OQAFC74xitnrwaUzHmBG6YREsGNUmji3zNN02VBCsff8ZC7PIOY4Hz3DJxQ9e
7SlIU1XmJquEF0rGpCA2ZsdUD6mvxpsa5harda8dmIpXRt2ArRqHAmOAxGRm5l2btcYwHwqWJKCf
5AMrzDHXXMjlKE10nspIhWXiUgPyVIL0vJzRRWJZGizxZOKZjzR4JH4yn5XtdrRJiGrKfVsdnbpu
2QXYJH/B9DPpkaRAbF/lG309w8KZNXEqDPUYZncUzKyK62x671ybeRj7mTbbwd9jgtwjAhdvKm+j
oWmi5RuVFEohnMdYOUSmHWI1NbZ9Q5342VzGBVeewidVIx6lkYCC+CG42v6YDyo3NtZdntMTjM4z
qWfaG+80joPy2KXov3AwSJLaKryBUjJ2f8G/HMvoL7l5m8217RYn8ay3XHvMBnfNYVG2euOHn8FD
RYjZUE6lqoF8yIbpQenE5B1oatJgMMlq/+bovBG+5hKy2w9+KRQsGlC5rsJbQ7oqQdWX/DyLTfiQ
NysiMbSFrcOWWPpv85b4uS+dcQnJyPYqH/3Ee9VMXP6FEbu9/Y6EyTMxup2B0DDGAgbQn910//n4
IsmoG1OKyQxJJMDARENbchWEMfj9rONEzH8mL4cEJaZ5N2MjRmXTR6E6+wb3F/4tSsYPXIxI7Fdt
Ct+Dkfh1EddvjNzFJtoMCMlcD3lqlrZlsNxrR5z3uM+EmnscCfCNC5pPjSzTDC3FeotQf9/VQCYG
ZctVmVvkk9LoO3QmTE+a4Qs4VVeOrMjd/PL+QrkJM8S1zu4rMJ9xLizO0sfwVFUZmJxOprxmTIbc
9bq8JRW7JhFhe+qAIFFVEuLblgfzJVwdOZxtxSJNKjAVbI4xOOvKjK2iVQnZ4JU56zCP1iY9GThD
68LaIVz2lkKfarSTg5h6/BrcGSlCojasChDT1TCPJ63Yu6D23a60GwcHuINJPENsprf5jCv19yyH
ks1EsWQfIBxpsRnAUzyeFHAQ0PstwQun2wAZqbaRokqfJYjL19+rLlEKWYJnAF/IQ4h8YqbXCb2w
J8c6xF51K59loZIS3PVJotcDep0Em6UKDfCrFUYjOPgtodImASxh2MZqzJSiUR/48hFlr8lvRL4+
n64FgI8fTALuKymUrEZuHEPyOooa4NeI4e+xa/z8yqXijZT4zKPyyyvB6jj2lGXYASQEHG/NsKJ8
/cUuix0plTsXDYNcZ6OVfLHcJypzP2TZl9oM42WJHtoiHHynCbY5HJ81WrjKirNtBRR/gDGnta9i
ZX9eXEFG+BtOcYw46i5SLCrD17Wt3WwidHgXKeP+b+OMhLqCOBCT70LIZcKnT5T9+xjSS2JgM32h
kiB0YB2nPffZdBdc2rGdecvUEv+oitKh76HklVXpQKmjMl+9YmJtwgrQOZtqDYRiViK5TlovHxoV
Hdsm3ptiPzPCQ2ug9+Iv0vnuyFpUmQpUiS2OJA/6Lgd1lxnbRFyKnjqLMdxCYhKZcoKaQ1Bkz2z0
GDE3XdCyH65kZn6n2LudlhH9HptE5kKHWrZIEkC7eCwzOZDchzU1Wrt8hXCTg9eTIAidBbmkNh1a
x9C0Vc6JkWaDyK34k1u5OM6BCGcb8XpzhT5igOAHNqVgPWI62+EIHq7AQQqhx1lMxBINwDsA6tNI
7oGoOQkuIahWiMnnlx1gJZhniWfX63QmHQ2FCMu73PDgmsIYKbHOONtru0Kto/dRN5KR6ix9vOn+
6ruBlPt4AI84U53RSEI/nbxQeCCP25ANC5WuVLMVcfSjZVyM2xRjAJ/fSMwQqajXNzU73LZm8mVt
t4rGoOTjR3+tk52wjfQ9vC7Xl6viHaURS6mP5HENMHAJdHzqrFFbi6/zCxg/S/g+WM08FQPPEfJ+
vNax/iMSdyfUs0Bwb9mAFMQEzJS2Yz9Ie31DDcHJQhz/QCwchwL3DwXNZ27nGPJenIB+vLYyCMLh
317vQwayOEu6juLXDWqABjJWxqqALYwDfwbKBtlR4TvNNHFjUTioEz9XJPKDweSD0NyklBKIn8d0
MeaKpDZDD3ZmjdjdQBcL+XkHEYN+yXS1WgGJCAzsZP6wHYEDRqYVLCw65Y2GQ92HihR2hFYXCyOw
r5p9MQXnbbeywCipJeC0PJi3Tv0j4v/EQyaW54ffsHkVEfmXXESrhD6y9xzRjMv3jBmMocyYsnVn
rKrJ9nWaTckqLlxywt4s4vHYAActoaq66MCT6bsG/RtZt3jrRIKNIcrLyTSqtKkqX5q7gLLcVLLV
Sdzuth1VVsYmRZiu/+pZmS9TQj0vHnY7d9AjHTvx9oWI7+KL0v5cExZTj2Yj5UI8UymsqqYY3Ezd
w2g97aUa/Qo5CGl+zt7PE6RTU1e4Vue8TuJ9NmTtUdI4LhCdeE/ECywfYX0sUiZPQ8i2f+Sa7btD
8G9UsITVtBYUZnzMkQIE+MnI+zHuz6TV7Ny8+UXCYAb7AZ0fr/gGaIMnQBRBRDJaDcmB/dQ12gSH
OEb2JqEyqZS2YJkpzxpWvvzXRPfRVZ1s+tUxPe8u8djBEuJRteFS1km6ujzMGD743HD4NNhbTWgr
gVzKXFxbWVtSCSUXguLrN+paQChD/gZ2fJWLdq9EV6FTo5vwt2Glm5JPjaQA1vNt3i9y9mr7urfO
0YbrBEcLKd+LxLn0NH6w/UofsMCmDVwvoZyoZzDwlaWaXr3q4lSeviKne9p+U62wijVYELWcrrsd
usoQWhfoAG8Dkyv+QfhZHuV/Ut4IIYQE4iHrBgR1PqsF6+/CehjCBG1b6E+kAF9xpT0SB1Ok0GFq
gxjfTqKrYI6SOK9FegcZh8sV3KRntQ05aP3/WIe48F32+BW/YjRkeLnJtLPq5+LIm0kUEplzXpUW
TXCt4lcwd0fNFm78pwqPSLTPLpcD/Y3t4ga3EFEaTh8Sb8BJIiwdQzFRDtPmiXV7Xf0jZssn/rUd
4T7kTLfmOStCvSlDTy4TzCrNPNOVeRc6SivhpUL6b6ETmX0Nv6rnrk5OEz2SuTYP5tcEMcmt8R/w
PpX6n+X/XvDlJ6VN4V5B6hEsgJhzdSgkrp/kdBMAs+24RmcU71WLngeS3XKz61R+OkEsZvQuMxTg
+axe4njlP/tfXSTRbDdhhwwCtJVmZVPrHioFcRv2aGVDeBKT+oInHyWrcgdwW6zBLixJ5eC1KGh2
jQ/EZNVUvtcjOWAoPcKr4UK8LaIY5K7sv9BL2z2IntGmN3302Ir8dcRdQKmzhyQZpI02eBZvmQ6Y
9svb3FzZykHjZrSIViKVg6Aen/A9wih/tMlLY6Z6h06yuBmWhQYYBQWv+ASvFOZ80006+e56iHbg
r4JPZ9DXzQflsXVQIBlG827aLVTAXd+DKhMuO4BAIka52erSPLMHoAjumP6i0RReQhZsPWIk2BdV
WmRw2u17IhOc+/5v8AqPQiColSvV+WowoeF0LAwtRQakBVFMglGMjW3S4cq/kpE87ASG76TjMaDw
a9O0K6JHo5QmV1Zo9gLVdecbQZ+WmFnGMveWNc2BJe2ZsWHhiD3cSH6mqf/dfxwLQnIBukgCW6Jz
rzAKWP2lpwYuxPyTyyAeSYrYJ3uYTBINekjbT5Xh4xrNhfUjnJZAXgz2J7HCETHQNlx/UIg4yMzW
B1gzLOLP7UwtVlY+WrvSQrwLBpctm650nx5j9ypy0+Glhn7q4DFAMUPXa5/fQF079erZ6nFXZNp9
34+cbH610X4pWsRt8y0vh6lD+2wMGknmGteonD8+jxgV1mDwl8yIkm7N7EiSPl+hXrKVWnYCuA/z
zJ97lpOGCWRaCbED/0qf7X3y93FxPt5OjFO5TysBaKebCeIe1rj4eXe5RFqHc1L/1s4dCQqr/FFu
eGZQPQ3VgeCQTq+OgKauvuAbqI2/m73jQlTe+btnxgYmNVtC/axR3S7MP5DQ3Zfccd9XJFYRpXlN
3qgYMv24lGsdkZteYDQ8Gk9Oy3NTvdM1I1H/aVCuyLt08fA1oehjqhd+XoY1gh4g+lewyd5lYx0r
+uImSbHKbVWZHbFHA0bKG1qLb+o4Matq5tZGXhnRNEYjmE76ByOh3WQaLpOj1q0yh9mhF6O/379t
FdXTYgoZpxpddE+5xltwJzJ5FM7MtroRbstZNDo6ytvvNNyzxdl8wMcn6mIBP7DlNuzddg9/jXpq
fyr+QWo8fO2UsG3ZjphOiSrSYEZKMCLC2IqEPq0G1CHZErjssv4c3n5AsDnS4ay10cEIo6/Tg9qB
3+Sqriv+n23j/dSxkGISUkaB5EpTM4w/icBP0wZ9ukAVm9KJxrc08u9dtK5K0F8QBO5BWpGwebfR
nQB+8yXnNWYu82VIErRNKfoEjEivnUg3QNsLueXQYpYZzKvhCs8N33wndKZpRGpdGle6GjNJqkhB
4k6EEuzykCiMdr7/3dtTHb+QSfGrTdTUmllLuvrr4Ja70Zt6poyqH/5Je6Die1dIQJsGE1xRqDfk
VxR19lykiQNWv2IcHdeYC0mcrtgmkBLU14OME9NNznI0Z8VqS7bo5UqbirRKn6zuemXW63EA5Uov
IVp84kUZlG9pNxtPazEq1y8zejre/QKMEbM5owWRp2sNky+I3+8buiNLvfSgrrTrYFC4IbBn8xWx
ffnO019cO5e+uPzA2+jQBM4X6qJdo4k9KUZzdSC1pAby/75MczRASHps3boMRU4eCHO0xrZ6yZP1
6/E3Lkvi5WMDHOBBbn6+oJl3ZqkXMRnnjYAzlwg/Jh1N6b8mhZcbJeQseIhfF0ZjEI7onmLpBnS0
4nRe4AVP8FBdUa9TQKqzqCas6njsZa4aJyA/pF3uqIxEO281EQTdWA9Jg/8YLWX8wjghmJ+D+NKZ
7cdb1waPAM4Gc/5Q/ccb8KVLSCHR9Wbsvvgfal91ggsVWqZ8DQJF25gG3bNg9h2Yqoalt/iB4Ndu
QIp97a5t8rtcITqpJkLMOIMKyqj30DpZbWK7wDC7guzVtxV0US57F3mDCBqOXnY7bokgB2/Ah0ya
5c9bcnUK/7Hzx2N7Ka+CEpVzfYsSf1o3UOXzXtjy4WZNQovdJQNawcGtnrPKJ+vY+Z1bx0v3wmCv
6OGMV2B596k5gceOtF9CV8R7thCNmHL4ra3k1HvdBWH1hNmTWwomZ14e43q6qxmeYc8aTHJCWJLb
bmb/23F7SLuY/y+CgXotQYYaFsCeMHC76KXxWde1r/0JIiy1CPyXb+8mnHGLmxUyO1rx0phgN+Hc
kqafro4v3LsRPyXdw0b3dXkbcToFLPHYaUMtJQef0f22aFowTnLvX5zOapqLvJlgNrOjWZWnrRvA
sJh4SCqgjVwXaKwd1eDLUDCpLNwu2GRbITre1ZTCGT8uyO6nifnRl27ps5XkTFLggZgvsRtp5rA6
X8ST+DBViBTN4J0HJTT4oYvtJ+xOxlNVp5hsLBpg95oCklooefHYefQcRIM3Ks7x9gN3GOUcF9xQ
ZU8zvvZg2oLHWH7pbw0MwTAPqCAXBtdhqW+0RC/1pRT6q8Y4Ma86B4QO9weqwLN21ywBs78i5Lgi
i7mQBsg2b+Dpthz4moh5NPTmTZNGCB/uASpL9pPM/S/SY2CCcusHvPZN9ZdE777dEooWQmUqIfxx
NiCNSf9rJb4EnHXmBt9RsHs78PYjMqlBk5zzKFu9BxRry7AcupOTb9hr/sKZRUR/7rff/RBjHyOM
jNxTfHcRk0/F+lgtwj2Ur1WZmvBtAK4pPlOOWEva3ZTi95jTF/65PZuMXf+oT9qko3mbpH6vVpfd
YZ2aAIegsK9OdW816A5T3Z7GLDxLfIxoG4d2NPXAQVbaiV3OpChBvN4sittkHJEKmv+qk8Cp6ef1
xKx6J/qG+ZrxBZv/UAIgKU9CDWRA/Zz+8xLSQqyt6lJDy9+3pxMO6/a3Z6xWi0/aZhNgWjT4XByX
DBJ3vyoc+4+tsHPznA+bGmnjdrPi8boKLr62vyanBo+uKNwI8Miy1hKm9T/yhJvIgyH6kDoI1m+3
5qp6WShWGR85eu5xJw1RSU34XoO0wL4WAkmt1YwcrNfFLJiOjANhK9MYm0aeFcPKBSTsA7yeXVTi
Mnxuq+r95os/jd58xf3PFDFB7ACpa2xp2MR1JbIdpVEu/Al0CObsR8CiJGgivojtBpYpX6jWTk81
EEbWVRMZKE7Ts45dQw8NyWl5gY8ZHbQz0qQc2vJ5DUwiWeu/d3Tpq082BebfYm9fqwI8sThhKsng
UcQPtZkz8ebVZi7yflAxzPeOwDv0xIxWX7g9ReqhTrJXKJBml5WT/jEw+qdsAlX642GR/9UxfULd
3spb6QcSEkNzwzdq8Ok4+cQ7ItDMQM8E924Hbmg0Oaf15NZG0m3nCGUcmyVV12wsk7b1hdrZvVui
H2nfiyhoz8gjFKizAHuYyCGqc20y6aQAC8BkgN/i0/5WSGxWB59AC0p0cI1oTUqBjLxMiXp4gOFV
YVwbO7K8iiDQksfm5UNrsiCPvh5R1cjPReecNDVMhFPGMJMGlsBjIPN3h3mgEY2uqK+e1VtP09CO
f6Eko6yAwya8rJXlCQixeNLg+3X0TWuFIPSXbHpWa7iPeNCKIRwHBzPW0AZvFi6aIIdEVPOar4U5
L3n39FEVSGviqHCIBbAx91TN8LdnM7YsJSG05UR4uKf9MDNMz5ltezMwnZCiRoDX+dbdkILgeHUs
+G2pRdFbg1QvwyBlEcxsydsOjpErZ6yFu4SzsxtAjwHl8CenoXwa5Zok9ZpCdkWwv0CIVr/FzTsW
lezgh2L9W2UxY58JLoDMAYsmW08h+4vysRKHuJTrHTeiSjYI8YMNhnr1qu9kv0yXRZRvPQJiERkD
wJoz0Fw07PW7afk/VvuL8K1ZCun92KwQZKo9khmQjZkD7cdWUApMuINdsg7kN5+hcP0Is/OFCpDF
4QJiMYwgBztDvMrkqKNdatt/LGY1Jix5RRK2+mvXze3ugRTrDKhfSunwNrN+9k69DEDawL4uRZaS
yTXeJ3y/w3TqAj4Em4gQp1iuzhTe6t4tK7K+Ynu9pApe3GI4hco5gYPeEBvyPWLNcMKKN/iQreSL
3JKTx3r+Se/kWgNN0cU5KKJ6JwBaCeRHvCotmynEZCV/y2RQCN5nQKrftddc/zlci2Okwel2IGkF
CteCrcmS4G5hU7KQgZw+n5KFaJlgdpDq11fbFjQI+GPnyuC3ZhAo7OOAxBZ1tierbFnz8r0Yh3Im
tNWd66cDlaXkyFGW/lnybyvF3BMriVgYK8zO6M8IplSrSaOm5G3xmMV6M9hnX/4raNytI0CBQFTN
mRe28rVJtMMjBO5KOTA/8JBf/Iaxb6bhbBSyOh383C3vdvVs0cXm6Bt6zrNnUKyF46HGkph8EVS7
TqMz+5oXfhRTPXsrctu6HJlnu0PzNq6O0gOh9UK6o9Fwau4/JyR0YYuP1aGcgQ3B+brWI5hAELL6
KE/9BXTT7i6j8cklZwCbVWK+nGO8HYyS1ImIbJ72WHkNm8LozEg8XkEphB40qtg2w8XUVqNMiwJH
1YA6lM6phfNzeD8F+8d83TIHZeywqKFB/RbgP/OStIMmKzUGaZvwnLByuErg+ycfm6AJEH1Zav7/
P8e7q60h5MZn+3NigvNTq0HiCj9LwPdzv322wYlqZSDadXIkLQ0fH8UEhDe18IdGKoqLJf88kG5J
Q/ewwHsS2a1X9US3Y0pH7sYEi4hi9a+TdB5SGd1xJkho/Jn0qfF8svBNVun0u8AXzshNKhS44v8H
oHQWULVqSn6/PJcIctD5J23ijueQ9Gg9qQCf4iaGy4OE18AQiwudq9rpiR9HeQcihp5sIufqTVRS
E83kfogHIy/DK+Nfn63uqp4a2VT3jvZYfh+raMXJbWpTTBMHXlGoPtPim1XRQpaDOJE6mEIaCD2V
ypU3BVms004KoTCd38Vv9BHuExkbG6UzQ4WAXxhja7P10sWb1OT8Y9KZh0Ha/lUQkypUXmxWEHjk
BtPq0l+94hQXOSOQyfLYHrR58WhxkbIslwn7hm7AJggIbUx8wGXZr7Bk424XnaFFaDo/bz0A2GZ0
WWNz//AK/Zb9gRVByAvO9FBnQI7cAmIXWlBJ0i9tBh7aN6GYoI1CNf7dlr76nsDAnYeChM0HI3yk
80nipXkHcV/F3wMyDBWuuPSP/M7SsN6nGF8VYqjfuyX9uMxdb5bfAcjp9NeQbm+axnynAU0BCWHY
DHQdzh3NrtJPsyt+C1ws6n/AtMA5KgfCBW6p9RbZa2dTbaDVqxJ1YRebKY9L6vTHnQEJnbXYCQ6S
F2hDW4iKhs1AMRH9RITzaoRjr06vEGFrEMDKLwtMU/30qotyACtrx3N/dNVLbNSu7+J7HVKqzQSH
B/iLF35KAx70/NRm7T0oXn/wSJju8hAms+UgMCLtszSdftaMVg38uFmThsYIFeeEhH01v/LBhK5q
nUm9Zk5wjBwcytEehwapT9uOVaaTRCCrls+3M7hJIw/dOg+JZh1PkYRex3ypiKFLMyHrEyA8r236
NqbUZayA18zzqiXhDTlWbaFvWXeg871Xp1DRYNHYBMlr9c8DGWRf/KI9bLF2cgJBDCNgVGt3W/wY
RSjhvYr000/5rYZgJWuTgorzbFfBULszQAInYRd8WrH4yhOl5ekq/P7pbDkdZU6DAjcV1IfoZ2p8
mxab2e7RxoadgSLQHhNHJC0Ms69kYJlmB4hOaeFnGxR3es2/hPO0zo7H92B558eVG/thqMU2XQ54
RV5yr0xSIdS74L1zoJpXKqCHUMar8qax6UCEE0xWjatmKxIbZwzbPSqCxm0J+ScxE6cZXsxe5qyV
jvkadDqRK36TR65TYUnXMzBdrrxHX/fHuo3rmp2TGZwiQYC8v9WHnUTB6TKms5kn6Fi1ENSjxeRc
Xhm0qIZvOHlC0SOpQp111BCdarCc1tIMhisjnBpGRdfiSAQmyy/PgC03jk0LotXhBTbje1FBa9Qn
/SorjkUoUL+1rIkT8wiCtdmjkgKD9/8BFxmP0hp3NiJWSkYnqt/oz3lSRYWFclirkTTeXp0ccvO8
x9luvY1IeLA75s1X3x4ankoX3SBPyhwtEnqyfb7AIHC6XuoUOKZSG+IIsyx8hrgKMs7ZQtAV6qu8
s1tqdmPoLEJDQTai3TZbnxH3pikbOvfZiqg+pBY+xg90FyPvZyxOgU+YPPtP8yB5fyjwdwsFVJW9
XUgXES08HEBBQsz17NSQy5UKUjGwOBn6SJjeXl5cYoX751g3qavjm/ChJ4XFNqnaevvy7xaZoVPN
WJeaxj5KrpKbWF/h82owNsmapoUNW6gggoU1BojrPjoBlz8oGWiT+VyplTjNuHrzX4EBE3SEbdUs
lMaBlPU796tujaKGxC6lDIfnLS/0o/tPfWWYij/KQJ/qb/d+8Tn8IQM4k95kX6q15m666QYSXiRr
lfUc83mH519nbHT5Ynu0/CS356b0ED6Gam76C0uCwBkOoiX8fqp/ArpQxZm5dWIXPMTf2UWg8Ml0
4LtD9e/e0xyqA+l9uKOC4nRq1epyJqm0D3zH8TiabzyScf9kQDhAI/YJ64V+342DeMeQt8lsznQM
txehgBaApfSuwS7Tqs3KDQH3U5emTfO8mF+WE+2hTEH2WDeYaDMRFNAy0Q6t5lzR0SQqlyPunqIV
LI/zn1yMkFGt4pQMrPLvVNiEI9T6+nWKbRwGAVttMt1gwXetPryM73KaK1QpH0/0WV9q4NOOblLF
DDBNMzUtdeWWG+ABy/+jHrPywKFNkfQZ6AyhqDvBcGp2F1OQvyz0eD9GFWOLQ9ozkYUuTnYOFCNj
ZCsI58naEx46bsTApF5gYh/YWvBYBaaI+wbtmcoyx8DvitQTqXEkOBN+4rWbVatHTHpjOchtbE3v
7YlHbPkOYL6UwlUxkgZFDamsan7G3+1r0Sr2EcGnu+WaIK8mx+TGgkmvjgS64SAbGuR6RdJvePWy
ceFAC2GaiX2WBeYEpJllnloHDIZiuEYgTl9lP+MBnWctZ/tifetcw2b9GpxepSea/N3IZeoNXsU1
PljiPvPkApvyLJKfgPOLUk53fmnGiYir4vuG9EPe64FaGPteAQig6AMVAYJVxhwKSmXip0AGooyY
3ulzqfoaV0kolUOWhCPdQePf5Pfk9S6rSTXBOrA+7y2Vl28it3sKE+GAqWKg6CqdxbFNB5DTkIgw
Z5N9NhMxPMqub0CaIZ0SLMi7DtOLImx5ylq4NvHRjDR8PUlF9simWmvz00FN4WV0ATGYW7o4ntN1
5fxm7gyd9MllWvzT461LZ91Ga1LjJPuZ4zpticIMtVmvqTV2obbRuLlJ/bO6jcDh8EUSuAnSHYlD
0Hls/cvSfWvTWx5g4NhHM1Ddg6COE6eTzOpvtSdpr4LWOQrXazBqWnls0ECLYDYwxuTf4WDKx7mZ
bpitLF6e4B9k7AQ8oYWEaj3uerqioyGeo5SGDPOi9CBHxz77F7FRvIXBPxsqaH5t5zaswFb20jmU
4C7CY/hNif/h1VJWJYX8TpYuvt8fxN1RJMUzNj9nu8IRrbFUrCLnlywISdyDPRfZMxQU4OWikfUb
sYahKrj8Rh0cY0m++oTE1HPxmKmeU8XVv5m27dc/qC5u6Db0DzxnYun8FcpHlMr1M+9jxNQZx09U
RsV0Ie1Vp/clhvfyyCyDopt1NHUQUWZkT6zjBMDgbcM9HTTaO1Sd7hAmjPe7ehe08vRZGT7kgAgx
Vrn5/uls9hJ0MextejOPhLWvDNjpmzMwVI3JC/PIaCwR9m/3I0nkF+QJ4lRNwTOcPJ3C/Y9tOGSK
2DOEkB1g7y9e9g/pgaWQi7VqaK5z0HdR0gR+YvzcMcQdMrUUg++iN7zDLzV5xWmtIMaX+Wf5HUlN
65mnDpBl1zlTQjEDpma/1ZYfqU73YGRqIhZdcATYkWi69/PXoPlSMYMp5KkKyfXs15tTr/G8TYNR
ouLkwpz/9uW+GbeuoCB1yLye7ymjVoXbhcYyZS5X5/zqR0XeGbJAmT6S6uFDf2RasMy6f6bQEkr9
UlST1FopTop+m8EGBxYiObYFxBnc7VfBncHAPv6GjjediteROd+JT6EAA/hwPFpwLpYRV7+2+Jf1
JE8IeegKH8MsLn51Tc+8Y/OMyF5x9a9d0aKTWawv/95i9Yy0bnj/jzuHm3w6sVpXofHEX3sXJF8R
YjnwPLf5BkzUb3YHO+Z+uhKFCIfN+y1/wkKBbqj1TbW7VW+4PcCLq5Nyr1dhPAaB2s/uh3mEHW/H
MsVO/YKcbx9EvJX5+cu/4GcUMpw6TkaHPzHXH48MVCaJe1Wg5Ql5Rprt+L6ocGDC9nD/QWlaqRVt
9tCdOtyEIaaYtCDw4RLsFWzAGV6O3u1C4MgnR+wo4il+6IOYem7xg/EiuX8yzhD2vNggjdemYZuc
CRtlB3XR/9K5GGE5gZHKOYSKtFDrWr+6tmXBpZwf4/5zkw/y0mxd1b+llQT8oKiHVZdrYYYdTbKo
eIyPlnUZlpDuXNAhgJN1nk9iDQIMvhDmgKlvSlZnr1jp2sdLFwQm/Z8PitSDOsue8YMbOeLxMGmz
8Rk3Nm1kndG7q4RktFibefYESU3C7n/2IR0pfR9njtf/+AhjNIZsGrUhwrIVqqc46myiEI81BAYF
pgeZ1hrWV3e15rVwKrpTl8y2qnb6/JNMD4bvJDIdJqnjjPnw7rjSGnhIKYjEu9Tt65RmH2+bUGVk
eGTNEi0Ez2oKUix7X86+11FZ1DeRefHxTW/h5bedQLXG/pEuEK/6CHcA6yIv32mt+1ncW0Jdgayt
lCUXzhEuVBE7aPAIVAX28bduwgB3FT+SlZZwVxpBITTJPcOM9ue2/DkJSOMi0RqcZugPngtaeUs7
15ao95ytpSPFi5+xUzgP7MmjEBjm+lwxHrSnAj/Y76YPvvWiN94RSt99xoxx/gZhFTI5T0FWs0E/
bp59g+xOItha5mpXMdkI5hh2qSaeE92MU/54hl9xnXlMwLxL7rXn3mxnzaqGScU1qrSCFTRFa2UW
P6Xt1Li+xKpe7ww16X216rZCxxbfXv5ug+lfpGpvP1hRAY3jr7oiPdE9/nfrf8QGTXvGwdjU7Ojx
DQ7Mvx3SUHBlRGfXbOch48HH8Pjuh2yKe2dTY9NGc00vXKcvfOvgNb76xH43g0e/yqKFsMipEb4c
fmHArcBDcr+nj3hshPwCWhwlPOFQ7fBMMI0cTSnX2h+xj5eWoH78lcK1GTgRR6mgSx4KQe7bFYUM
g3MCD9FB2rm/t5aS62qY0DHBX2RJUySk/UBOu3w3Fs0kXCnVDoN3I71PQlaEAUyGxUuY9EbYZ/Xw
BlIIOGuDMmtbJyn14tHMv8m7hsjyDAKZ5LDD/XeuLzILwU7uG+1vUAiMx+9spxbf4vxw/LEq2Tvu
Wsr0ZHw0U/8IQ84q/aBJao9Wf8XaM/MzhfIuthmXQdMIXCPBWZAwQwQPXd623sJwWAHSOyH1rAuD
0fOlaKkfWKLB7NgEbAzoMpJeCOZZmX0KbHtZ6/wbxee/9X7GlyuSnGdJg38ZwipxuZ8HkUUHJVH5
nutgfER5ESixZtvKU8SX1UVbPK0w1XrK5tuJZXi+WwUS4KrwwCd/P91AjwlTQ8yOo7U9Y3buvJJ8
YTs7abi1ggP5tMWheB4dlGpazjHjPDMeKgLhUUvq/U3ifFXaIX2heH0Kd9VbUewmcOdr54uzTk4/
SAAFxh/jxC3R1Uex7RiI6QWF59UFtNpNiwGtiWDJ+8fYFxg+YdnLZpZGNtha951A0mftL1ALcRKj
bzRulftWepTemqJc8iXOPUt9gY+OyUWE2QBZLpphcHV6PbMNsdvsdaqi3Q82DWkZwi2X2u3EQxE1
lfaLqDRd70ROFUKHDbJ0o4RU0Voc3IBpMvB3WyZ7nPpFYhbZ2WDFyRoPQgKh0li/MPLdUx9rC6f8
paxGxgiVHa4yARNy7/cMN6hQWYh5khtgBVFOXaNi27o/EG3erQR1XPaELWP/4Ul2V1SqSShi3mA3
DihDF1sQD3fTO076B0lEZpRt6QmjaLVp4v6+i50K7JoDAGb6nVbBUu+m3TZqT9L1ZH/gHEjoZQnG
W2WwnpkfXcducXvVcFCR4oWqCP7wcLc6b3ZolOMMmUCj0IzF+xqrxqFnisgJZEPLUg2eep15q7Sr
1OJnzOXCJ+QKe1Q2kETXbRN0eOFveqXuGhUJwJXEwx/8GGHWplJlsLOFZfwiPvYxKeJzYSVyx8vU
x37Ib1Nf2nsW73KYSdP+CnRZH+Jf9YVusSEa9InXN2BnwCqKLqC+cXhHpfPJQbvs94N8922+hyuQ
rZ9H60mF8/h1at4rxTKJxfC3GFTvzmHTmhEFGppd8jVOwxODrZzuEW4w+bc5ccQ65iboSoCXaMLF
AsrRW7rTk15tC9Fr/yr7rO1kYXT5/xl+VkKbqBoK0JMuAiId/hDj3feoTvlEkJBW6wD0Nml0FONQ
PH9XvkR/pskrpeR6S7roQSgJle0FeIqy0NVPb7950mFSbN0BvZmXkMnuGDq0UPtnbyGMoVM9OfgZ
OlK2Vx01mW1yEd+Hjvr8WAdl7u1hL2SXvzmSY2wVeisWNpFot7KB64/wGmdbPknT2NcKEu/OKmbk
Y5usAIJD/sj1D1E7BbrMqpoCPqDPMrFF1cyI8ZDG0AxNnkL6AU/9ze3LWlX4pS3xj1BAZYuVumq/
PkZr4RRD0Hi/FsxphMWRbxtwtEghs0WWTVBrJwycnF55FJZfMtiahQArsnuygTezoBDqFB907HmP
if4OiBAtb5KJBPtYQNfvz8tAg7NR3Oc+UeUZJK9LwOvybWfFmowym1zsb/8kN4TMKwTz76mdKNLT
/1yJMswbH0TKWy2kQYYHJ0WWRD6GHbkMGOrI9blW3f4ZJj7MqUUMRx/9HpDIWw7scDJYoNdQARAm
3HwqA+eviVw0vVFjc130CGb6WxciKJsmJjg+5YnNnTJkFkJiZakBJywgcZ1nXCGAnybUx6MXWXEV
/EAa63wAKCsK52ryXOJRrxhG/AnwZOc6OWEjLFIMYnZTCyOvCSsRPtJwvexZcOfAI0TPTY6FIAE8
NU+Rdt0LW3PSND3q8YA0Jx9FsFk3uVbkAjJ7bD7yNdKeqwMOq4fhIFz3Awrht5hXGr0FP6vaGzdT
kkyRjFZxBPjjchfyhCKvfNvucGYfHS6nceFzL3CL4QbRRos5MhcugHx2ZL70JJuBA/lAyjnc7txC
jsvzDT8t2jrK8WKX9k0sulZnQQBrNmc0WPC9Jrjyisb3MYQTmyTvzUSZ3DkRnkneOPEagNHLXGgM
AZmHnf7VaRev9x6uqc7P7a3U+Y4XCfm9zgKO+sBPJzlk8fZBZrQVjB4vfmwaUetIDD+siI675Jx+
fHFUmOC9vitF6Cl8Y8M3J/HEdRJaFczOpymkaEcLQ0ZprUacwGgsednzR9Q2IX7tz6UaoNaPakN/
6D3CwKsWwKS1mpwAJPyRXLLiKCTGMRicsB1ZZWhH7jtxPtodATbMkP9TRNIHB2hgvDdMZTmVEvx5
eHjn4BV/dcUTZ7SSR3oEHuOTo1C80w1CbKvNIdX8AkAtaB6S9K7LBvB+462RfUwVOlb6noCRcKiE
OE77YEbGxE6LlsQKyWgrowCkNXSTFNgahSYt8qD2QmDZilD+1Gj2W9MrK1zOVbJ1Z28GUBpEUo9d
MIS4idB889WSdRU1Wd9M7TveYpUI1whQbuVxZ4ED8lv8buuRFA3nhcEE3JowtzthnCo8XAHbX0N/
9f4QHoNiENliXaL5uoNAytqP4fMol5GZcqyF7gt6evLYhvmoYfdXB7LMT53HPYP12Lkntho49K65
C954/6RUrYc1/udLezKrsv4zXjpYnez4y2T57kKK7Yk0kk15TecdLkArFCm89caUfNHJhLnblYQO
0tEUuvV4vXD1qVvpjKvJIlb+RLY+4DVenC1iX1ynO3IyvFsli5qCzA9BCx2jMSOR1g5G36uupHSG
TReCIRz9V5PK8mISDKN0GcL22VJWnh7MqG6NXs3LL5kzgq4l9+7h2atX8mBDsblLTUdtSFmty+hL
ANdW7so38Ag878VDdJUhvwB3HuVvYCJ0pTuWRLaf4U48I9PnZM97pczKq0EKL9G56hAk5RtaxeOr
h52BgciK/+j6ng/fBmYYOlMZZL/rExryN1JMVpDPceSf6SEkV1MaF0yR5jVcKe7USyKiKq2HRebg
BnSaihaCTJ/2iS55LvY1GMCtXpF84t0qblz0ZJR6eQS/fRELHlxJfm2cBOYprccxVhcdc922GxAD
bXs+zAe/RT06dgyMixIvUdPA05mnIliHoM+ScrVVSWNBQ3fRLRNvQ2k1J2nOgD45uTJkPQ/F7C7y
CHz8EZ1bpGeYxSuIVLgY194BjN3RZd8iZBkuKKlnzpZT9z6WiZY4xaXtvddftNF2fFl6JY0DG3Vo
7edtPBU/iH+UNJfxrLlOpdK6T6B2Y5+P/xbD0KO3O9N+NNkeg7lcFO/aIRwWvtXI0ePvxko0L6bb
WuU6jA/kTwitYiF4NJqEolzJJcnagQ78Z8woJ1+w99qV/8Y9iEgxrgZ0IRHEmYJVbyp6tnudm8KB
OJJBstgFY+N8qjy+LvgHCZC96hUHI9U529p1BYKUNmFsM7IedZ6ECje8yc7HtnWYE6NxUVOnmK0K
dbP60bNYjF19MF6oTQxCzBsTj7ztIBEHOtrw1zyhSDAfxS6/Nxv+Kd7R35UwZ35fSJNZmx0B17z4
OzWV0Zxj7BHBznA8ijhMcN0efnblK/QCfTrG/pINr0Pa0Raof/vaIf+kF2hrXb0nGoF4rZ0xa/Dk
HLbrwazZvy7BCSE7rXT+eBguS8u01VlVwZcUtzJEVPH0nn0P8LnKB7y7WZaYZOEiK9JPY4A3aGX+
uhvN/H1LWAxsLDA5HWqkPLvihjMy++MmIts32FsHsxaLhsptoeUkve5Bu4OIHm27T54DXsXuvJo1
olRjgNIFtovW7PJekqiFO2URoNbAj4iLv6e3V8WlWMuatBTFCvAaK2BbPUmTTGy2inXlg/XINk4G
nGR6W4gt9c2u48A470RZKx0GjswWu1BFiZJAW5TFZLlvp/F8QJYVka/NFOfZDbLWY5l+x9nxIopg
5PdC1MYsYVMSS3f0jG7O8UVvzRYowVWkjLRkuK8092Y0u2j3Dm70u4eO1u5DS0SbYiCJrUFXf423
x8SL/SZl19umHIgvtTLzxiopfjNMo5wcawOuifAYsruJsZTYk48/qLIkJYVIITLY3Y1u6VNlGzAx
ZQTw/kiH8ocpQyYtYHDpXpXQCu+u5Lh87V084Tfc2Y9rDoSgw1W6JJPwow0MLb8F/JQNwChW6MxU
2uNftpQAx8DxiAzTEQEMXH87/epDXc6+qwALrPIRYDZ2rl9AAbhe6wL6Bq/o+eA9SHSvAzPI8oRU
nAs4iglXbKm3oMAkJl399hU2fv8W7MZx3AivoKLURi15dPT8lkkYTsxBMblPHFnCSrQn0FrVmTfL
uAhk960sXEV3NWlUVslU0tFwS6EKUkXtz1TRWkdFW79IVbUrJ1spgvgAXNu9UVfpvSZ1qy0ofwKJ
n7CACWNoaELBL8tMYrwMurdnB7LKTfiXf3+BBhF2CpkJ4eBWlPXIHCbhZHgdGP7L24GvBPVuLv4U
z2sH6Sb3ppxiYy1NVi+cpcPy5LTcD8YPZEQGuscZ2ja7mQ0eK0yE44Xt+MM5H5Yo5CTvQc8XJKDV
LeYeWXBqOZBAtCwQNntWxtsCmxXOkVXKS8u24aglKhuM568qnMJqGR7Yx24pNLza8EaCcHaHceom
rfNhLHjsZ2zJbVsRe54PlkopQg3xLmGL1CXWArh+ycsBi6Q7L/4YLddhGrdI3maa53kwJIwb+PB8
FJlMiFPTHKr+QzzQxg6re5n4nD/1avh2Znf3F5BgSwVlQfAYWGvGBP6IkVuYDyGlntKx4gTNlhyW
yMP8SKLkoAvImfLK2PW3NtDQhwHaQ4SXBI3MXtRKHjzFbwPDTTj4aqD9Pnpw9MtM5uK56T98cFRz
t22KI1hUUrt9K940egKBoNP2Q/9lmBdjuQ7qBoEAF+LL9LNxKSJRXN2UyI/b22bwAj1bfraIN61/
YUNnfnrCPkpOGBhTxXUnZvWmjn/7x+5tpNFCjjw8tkkLqI89xZ2Yc8CSI5bb6gy0XkxQ2MAuj5Tq
jWEEJ9QzUACMewUuVEsAxvliFOnLngpqHbkL9KJqpT3ji0wW3hupuK5jSUkCCb/su0dcHApDQp04
smM9z0lgZivPc1JXnVkrRtKaqnp/gSORFDawHRk0KrpJ8pXn4y2B0CGTbWGVTjXp/oAUbvF/1Mwt
rhazAa5iCQemU/na04UT2f8PTBoupa24maSd33knABincspLeqVDFon2yZMih7sPznNz/b6esekn
9QVjhzQo0LbqtY5SFsW2vqXygepFVbm9q0WTtA/DCyAnsXKjAs0mKRdQZQeulo5Y7IyTaHSCkUvE
uJKA1j+joIgvqWartqBx20wLXOgldCFHcM6WeN2guRuWfbCxqNrysAW+IygccuYcPpPgWQScDIdr
8f2jVvSmGRDPiFFLQp77tc6K/vX6tEz6zf2ma0JoZkFdagoqTYeyMV9IlHUf+rSL53x5TsEHuqky
z4eY7FMAQ5DhxY4LLv5gz8TQCaN2MgWnw65LeLXcf+cHyl7EElWbHmb9OjESZxItBbHgsxnj6z0a
bfC3Ctqf7a+BtcWJs4EF6wA2BKVAFgYRqBHMgFkVUaZngE93IlMl4OLiCPrAaeh9bAYDsLE46TZm
EFi7LzCdj6WXdrP+yplszKzpHUJDkqWlVDg5GQhnYSwfJlg6IYCyWgTKrmYOQ+2si/k4ggTvSbxe
hmvoL4YO6LCJzCK44szjMjbVgP9+rW0SlM7Rbp8+58ppytYG0aHOSnCP1JOylalxxLQ2mO0lLVMa
5/gAGviU4FIhUW87hHjTSGbOVMRD2OPwJuqAayiJPiWZ3PyHSC5qQzZj79mpQT1xRQFGwnTYy+Vz
njCxdyHLJK3HUvWyrz8r6QUCsCOt5/SSANdjk8E4BNoEnVFwhZ5RTjgj4uqJO+STYu0G5GaOdN82
q15pDMt8ui6S1tHkp9Fzu3XdP24nK2iqN+HK0bHwjVlCqmOWG1lfazINuL0KxlUYF0VzDudDLbLJ
07HBuDzNLbJl0/tB9DMTSD/cxLXMIZmNOils2YpKN7w1W8jljZsvrbnT34J3Twr+SjYqa27EIlUx
jZ0vKL9PibOwQqI8tWGgLEcE8HeNrEdMENROSifgs9eLfuJwUMQiiX5Ybv3RNmzFxGg+HAmG2V8c
kDdIIbrHAqIZ9SW75TcMmicb/90ILxMo+/llqfc/jOfggadtwhDf01KG6b7abmSYZ92v7/lN7jbD
hSHyw+w004AfWIUK68oGkb1IktDicdAAruQM2nCam1WNZvVVx5g56CSWzVpGQgoigQsZmzr/Cfaw
qq2KEithpy5N+3/dRiH6oL3tnMPdz+AVn+LjFAcfCRT8heCWec6I/Rri/sRBteQ0oKoyZOBPFOVs
OBtDMMhTwsSepKeM4zMg7nepxcwtZOiW7HODBgjYEE7pzgVhsFT24dUevFYoH8nFSPTamU6A7+s/
6wbn9mjVK1yx/El0+DmXf6z+DAEcplpIWZJz2Ibs8vh0jQYW/NoitUF2mJuH4R/Cfh+c2IQcLObl
rSaihVjUCp5aSVKzBA0QqWTSOx4PafS/GPno0ArurWqJEuCUveN1N0b+ABV6b2OXeRe2l0yq08N0
5mFlNNX1pMAg/UCDAYp9pzw25DJE0gepnEOHm14ANqrqdk8sIKM/p9mKD1SEGIb3cmu5k2GKP+k7
M0TofYa777VGkdBVX6NsEmeF4Q7cFA3wy3Up1Xq6NFEnovRIN7426TJUkEWw6wMcJl6rHEWpdmRj
MzLHOd5NrB9BDVT1Lyj9Vmd4zQN1w3Uafb1igayUn4+ztb4EM+WtSgOwQvV7bcdgAy+6kPx/rPqx
Eiflkyre0UsxEoDp5/zAtG4LAFashWtgyWHC88Fr5JRbCOkmZG/HcO53NnA+HI9LLRRL1siTv/SL
CgB4h7k9XOAwaUlg9grMdtDmiTZmyBd+nNQbGDQDA4FI4qrg7uda83CwWjun1VwuuV1geTljKior
NyrSB5yzceX9GrphxoDPaaURKhvlDcAxyttSP3afvEdevK0bSuclTcw0d8KeLFvwQPvcrLTjMDKn
5leIEBUkXIWlymMI/GZnDQefTN8Hi0gqokMIJ5X8AcubfwvMZdcLOw0WfVsqyroe/qvQ6Fw5vx6y
OdPel3+ppJ+EdJGEH1R/xboOsD8fHrDwGGzWHnr2+ivOR3veS1LCq0Ji81yvgCHxI1+CaayxfmVV
uZXlBzdYv/52zZAWs9GfyDsbIyVUgYUr9GhfUvbjAyWr++kR/eKgyylzbOb0BqDCit5gNZOwkOIL
hacn5OwHVkB4wsdmTNeo+RNB86BV1FR9ijSbi03M21exjBkWYFswK48l50vdrjGLEf/5mHNC0mmv
T181Og9fwsr4JEsxRorKd0QRKAmtw+KU69lKF2aggPGGIXQhNz9KWN+9qPp44jbikkEheZ6byyWK
lOSq1O05lsxZgGXGpXh6hgakHAQ/Rkx/UcE8thfNFeD+DoHHhuuwBEdO7xT4lY64u/zv+WqXePk2
F7k9FJ205aegSPWfi7a3qY9BjHUplPtesO2DG0QKI73riIN7VNMkaFE77pTVUJ7OKp91mJcguo9x
c2cS/VLGZ2LEeS89YdgKs7/3UcookcbJ1+NNWzwdfKPte4ah6MKITiXWJiJnSgP6yxzRuY+eflos
FIHriBphjpO/E/4jH8MkbK2WzzHET0OrybMS/T5t2ffwwl0e+3h8GoEJiJP3ewAqMVQEWqgavdpT
W0Zp6mukEYX4CXg4/k9JVwW6wZ6dRLuYPVK+Xw+mjOPuS93Scehc/ZK2o+tlvVWiWI6dJ00zL3eK
lBpjizMwrQ5o0AEPdRQOU3cUCNj+0k21hN5GxOxpwemti4QvAcOCX8I1J8TaEKyMfISdeK8zidGs
sF7BfwFaPlVF0ROQo4o+LHQJ4QVqX0qC1nFYxHk5srZA8Psv1i8CPpoNGPBz/Zfe0//ttSlBh8qt
8V3cV8iar3fWn2t/xSdQuwUMAJI15l4b0MWJrefqsHb5cm/B7qTncyR+Fu2VbNdYHbzygO7saTYm
ICRlS+s9uyYYwAsLx5lcFb5BsG6ozROjmFirzQJBkB09jgKF6atPNCP7x1gd9QAqHAu5whO2uDUi
m67JUBvZBoEu8uDsXmZGnOTANePmkgS0+HF1J2OVe0eCuzr+IGeNsc+URz/h2r7Sf2jEDGUgwrfE
K1T89AEROu81qCuMQZZljRCFVrfz/iQv9RCv1JMsdlICNYuqADIPcbeCFg+NGroSIU+xRvGy7dYF
HC+zOs7Av8HptCiLfsJtOcTH8/SMibPLANY0a3eFKzI3c5nd3E6/uKhPycBGZLtLFoCuVcfSkVPy
B9QsykHVW+tkJoJANad3gB9kV3eaPmStgHfrVThBZmfP0NHe6KFX/VJk7kiiM3Vqb1Y7r5gqoQ3l
QJl4+QPvnLDMRJ0LRL1rYMCgl72eJ9GB1f45d/oHJYTXQ6BNYDUKu4KnZWy5RlBPKzk5M20c7e1E
YcJI7ZJ73pUpNAe02Rc7ttmX+aIyro50pki41y4v+IA2E7kVaUK/LxG3fXxiiTNbGXrclhhnU/9T
/tmHDYjS3mAMAwZeg6hYli9aDIGHBIurnfqQsvVE2gO3LhJZ1zacHzgaolJAdGyPs8bQtpG8gLNE
rJd9ytER0FVcK8ziZg0vpR18A0M3CRDgN9I7b3fPBz83Y55dmaOuJmfyz6LZgS2cRqKg3lU06NZx
449gh/HFoCETKZPbMj/Rwcee/572Sy1KS6Oh2LEOW/e87mA+wZvRl6aa5SnkKonMm9ZCL1HqwxaZ
tAT94aFgKuzIEIDwcEt0msUBXY6SBa/4u6zVJJrblB5earnqUm3E7Jr4MebYeIFcXXSJ42/Po4Dm
5xERnTqjM1fctEaYmNFZSQx+t0FiN3fakZkbbKBNHmhhuABKyL8FV5EqFty9PmuU7oELvLrAdVPL
XvU9rS94sV6RMz/sb1xnSgkxJq5AQ+S+ynZ4l4Zm385QeNccbAZRFSanDEOlBhlmEFnkyL/Ev/kk
BO0G7qOdGIvF7zjbPOy5vG9Q/K5MEDBwEeI/ykHWlxxHO7GQ39U9eTQTaMIon0fdWu7cH74aX/5y
O19HCGWA6yVSmd2JzNtxILzZDGms/gzKkn4BhpPLfIY93wQqifltPqSpW1aE8xq+bmjmbMIxUOrs
3SCqHuTN8A3YTbWnEcA5ew4jZaMq3CnlsBwLAPrMM8cV6ZuUiaZMtWIX1RF2ROOE47iUdocEdgE9
omTXLj3oBt6+v2wsWVhG+qU4LL8VFnyrd4HK1SKG2e+bJMLJAlD8O4oxl3PqjERC35Cfcgvb0gMW
+HalwgsjP1Lm09lIdoZgyjmMXuQ/B5TK9Tm0UxXldDOFc+P/DkUJKagWxD8opzeGN9L+EzvQeYOG
XhQJ5lHFBwG439MKRDPW/ThnswdVgFYcphMqH3cWJ13yIZZomaXLAajkpfJ+zIVJjy7aKA4VwgMN
rHdstYkJGBywGtdHVlx3q47iGG+9mGSdqPR/DNxh8B01eZ/+47wCRhu8kfOsOfbucCHCUoRhTbOd
6ommuO4TytRstBj51t9oQfM0qt/dHbE5NEoKRwMt1+l8bub/OBd8TtY1JR+riS/+zbmnzQqe/bKE
rZ8cNXsCubqiZaxM5pg4JP4J4yBqbv/h9TnLuMqDyRe4/xT5YJr2vzkPKg0Md7LmXM/dcK+Wp3mn
8P/ditP5RZqqVrJUOLZ6XP0Jc0l6w7/R2RSKMHY23RfWjIJO81E8rMOnTeb9VmrqlFV6iWRUmi/O
iX7jqb/9byw8NhyB52lbHOGJPZ902E8RC/xnWetkbgigoBhBhHnFyZko5SQ8xz2ApSCzxM4sF6kE
e25UlYQQqoICX3+pDc4KfJRFvxu5b2SYMWH2Y0H+HGeRjKbA5PZkVx/tRnXNyzoyaUGZiWbXmKml
65QyGO2RGYJglti7YXyaI0jWgOo1sEADDYQNkNNrS6+Ob2Qk7r0kRqHeZriRnhrQiG8XS1naC5P4
xxvx3Y3lNUsvsYKVST8df+mj14O2C3ByVND46AGXlziEqk9++bPrCPTVJUUYRws0GVzyz8Z8Vu8R
SKGTjT2MsTbiJTb8Xsl0cHgYkX9ljbNhP88d0yINxRniMWnVgwKPRsxreIORrbkHFSdk8/IA7zVz
DI4jbA643Pqiz4ibsvqzrasJZxNZXc+xsOhtKcky9p7qNc1altWvF5zdGZKeKigrvY6sjTrmsq7h
nUcsnDAhtHSuJxf54BCH0HmS/SaIknVLpD995tykj+qvUUiC6usT6wHdZDCxkNtDC/OQyDHu5dZ4
Y6j1XnfUJFh+T2Mmz7jhFzJeWVDiAS52cdqnlZoVARIaRz/TFwJ6no7DyGSiT1Jt+/FcFuvbFJap
fghZ6Cs8rCKX21betMrai0LKSbzXk1E4D6zr49pPPv3pmuy8NozrLvwn740DHHQ2xYAh/6MrqQJ7
c2ak+KPCyoae/r06HUgesrVHcFAxBDGGh0s3aPFbfGzcIfEs0XVYPC0gsqy2LgAUWu5p4Q8p2IUQ
qusgnfdBcMR/4VYTQslEdg/I6Pyk6xgoZGUuGPj2buDTVsV6XCW1VIfwpbfTjRjeu658j2Zjy6Rl
Xqc4SXW6L0KjPKd70HPltv24+c8vPZbhnIFxQxw7XNerKlmQQ4vqlYFMyfkNUrgoKrekPxd8tfRY
jLN15vHuxwapRreiCwGsd6bBedC6i47zW6W3al3GAGNZ8k9sv5/R+uxb+vNYXIGLto1OX1Z6VELj
5PN21L2Zb4R1NVpxJU3xvfAwS72prhvLNviH3SK06JUL5FQfSFyFTV20I3P19BtfTk5R+Zp1azv3
A3o3eEpEUrXScufYY6AkaXd6F/Pznr26k2NZwL7N9aCeA9UO4PQNDlvIds6ijp53xEwnXCY/sfNI
vWmxMBUbL1WD4NB8rXvDwZZ+H0w1sQuX+SR0dZ/qrIC9zme0IEyukqt9YOpfGhylY+Jtwl8D4B6p
HvCJd1S4VUDpxDeRDTGwTTDOrZE6WJvV5fsN7C9cE0wibMQtp2INFX0/IuQJjpnUxSOJYtayktwB
N0JaU6x3WnS3omeDajurvedDSP0TuBARQWj5+nvOxMR1g8bW0aHs4q9o0MnaMFbudH9jBdNbUxUD
kTi19eOgsk3SeKksaIS16Vv3cMIsLUr9lHWZwP+PklgpGmhPH7zwmuQr7ejX/3sKE856b+o6qSsi
5m/pfKwXahMIWsz48wgFQ3hD58b7M/xRatqZqbK1OL3VMShNpDgOJzFqYwboaMqoHDlxIzbMETaY
uwyhOdtIC3+56GgKiikH8Zl/xbP8mQ+iS7sPXS9BBnveFgVEH53kyiomAlvRbSczt9Tgy2hCXxWV
8RExs6iaa3xspWtv6rvXSpnq3cpqBSSGrc6luvdMSWLQ0UgnTvbbq6h0H+bvmpHrW09tpy9euaVY
FmMYcYYLGLamOpIuVeVdCebaAImRvo5ksLBZnDTY8DyTcJNegvqILiECAK6OcBfOlIlZ4QhRLZL9
KIqHYMP0LbsJTnDUK38TJvju+graj43cedd0Okql6oLyhFoHfyw/jPk/V3a6HP+CusNIGzKqroAz
dbcH6BInWh7EwZqnIZmzZR5A4KIJbxXqQLTxlEzq6YNMhldeE5B2xV2PTDPGu32mX2cPDtiX0WNk
iUVhAXekHB7PobBJy6AK2922xfspzGA/fZzWjy1Oy2QXsgIcw2bYDdX1szN2g2h8bfX9FjTOKyi3
hWWEidYkr6LhbBHGawnHUUF0H4A/SXRREBXZOTVCHmIAxSM+jU6eZJc9KNKEo2IPsUuynDrgdS2F
disVl3n4CGnz/uh3rNW5Xa5Gjf/GyZ7d90ol9tf/EWX8lqlHs54jHZNzuHgQPE4n5Fknsfl9ImSX
+3VtqPa5gaZhR10Ibt/kaB8mDVSYsoZ6nSPbsHSJJ2Z62IjXCyzFSM+6Vl5JqnvjxppVSKxfkpoX
qZiyKHL5/Y8PWhbY6WxdMj4Qcf+CGyWoHRNp/TDs2PLjpZdbTw7snD5KZBISyIct9i/ukkciesYW
K9xEQiO5zeucIwWsxB7K5dSEpiSdlFf7JdfDBesyuX6WH63MIAXQOOxwgE+6vbj2ol8plmLLDCGa
tE+rVF54wc6etB7mfaGGcqGASmCR23iWVlcBkOUsyuFRGwhkg1VLGKUUDAQvVzbkqEO31KObZny1
qBx9JzL1fH+en4XWy9dVIjuL7tJiIqZhod9brZ2pZ5LDz5P2Sl4W3VtYb6eWEs+cR4O5Jf4iQT+L
SQ/Xxv8+5o5BQBCruUWEDQKYxOSDQn+BPIDJSQGQBwI+7WeOVnFPktmr6iYZ0mZeK9fpzNlunCYf
RKY/EuUt1eSidMzWnBVXGiVjf52z0hg9yMgr/zLjZdYTKDU8vNsQoADT2aACMG/DB0+JPY5wM5dF
pvdBtJxzM04iurbtMrjsZ0vybdoMOAdtyOl3czgFW8jD73ZbMtnDxvkYxV4RQyZYWiCp9LBPIscn
GkMZ08absrWA6JKftKPa2CfkSFtgFN5gFnT9kiuDp98+wa4yJmtbNu0Iu82kQQys2nZOjMyWvfII
JFKkolHf0trnaqAY+jm6XZE5fCZxsP1M186mu1e/Jj1qh+9cVJ2YCqe7eTl2Z76tIIObADephYrO
GL1+Y6fY3T4EVripoNMnD7ZcLFfCXlpBKMiNHgGjFz+snJGKlpFoExC7Hx/YErGI2ISKn9dZwUPU
cI+vkTgyPmkqqHf2vDQLTemEHcEuFPBjb2PuGZwxmweg4qdfotIjR4FZbXgwk7Pt/pkgP22h4yEO
IlTPaZjTwy16RoC8qKyrVDBKdSVhljpswkH8H+wvggRh/8fRdf4uMG2WO9NOweycfqVYONgCGWWR
Bigw+R44kmLiHA09/b4M7wiyWf/RjpWQuwBxKYTrd+yPkfaj04K4oWEDEVwbFeKWJ4tz86z5PHKy
7ZdKmqr65oWGxaESIw9qEiZ3tHq1M6+NRfZCsY/Afl768nbTOjoE7cJ4zoyugcUadz2kKfXLuLx4
tv6kBaB8dLHk2wFX8DdfmtSwPQc430/PLIP+79qULLNdBdYyfVa76/I60jIarm6HW09AGeufB7Wy
O2KlRISzLWCZikkA5r6e9Fqpc93xAvqOS3qwM33iOtyyaTbbTOr9dyXlJozhj2FpU3Bj9EVS91nc
I78ToDtiLnMJ4CPxjxQQ8b2JAzrPX5riLG1gsBHpchNPDP54R6EHPZP6cCaXWFgtBu5oAQKickBh
EALE4YbO0eY4jAVJCcHcxeRwMkDBLX1LHm0InxX5FDVYHYcKI9g8OVeszYifGsuhROiRWCkF0/UQ
ByPwQo6YK2XQ1rjGcHPYWEUcA6P1gZmQDUw8sQ9vDr6PtHdug59Xp1EHykn3l8LRF2axuswFIewN
jq/L9yQnJPmfvXwbiiVNzmxSn1EfZFVDgF6Xc2FjrLbd2uHTd5Q0G2c26ijn7PYMFd2Gflimro2a
AtrRxgkw8RrAjEY6n+Fuks3asMutVmJbjyli+lOQwy24GuIopRfro5M3LrCDMqx3JZJhqdkglcrQ
m8u9DHR03uoVdYmgcQPvK21Z/pzkgbhMiMlqNjFw+sKJeuufuy766Xjr6/NDoYZwZ/+Ue4bfvK4r
DCyugC20qWmxBt3mviVUpdcAxFSInV5dgpMhvlYdBeFoRUPDBchWXBHMAQhVSBfVR0WA8qBjiOrJ
G2KhtNhb3Jb8OKFwmLBN4ejZfgixPnDuBsQTtpsQXzmPeQAsjRfJR3dF7lE36/8gcZSvxW0mSsRZ
64RvIWWfSFLoW+LQNy2VNJxtHMsu98KLHt1XcAP5vPLkugpv8EX/23qsRI5Gk0Ys1qlUuEJ0jWDE
hnCAYDng/5bYlVeO50zrmnonqCzLv/K87OBYq1lVB+2IcjprmhQxVZLhSAmNZAHyMsU+BiZ2eK76
NrwAp9ets0zh/8yxWG/jzMrqK7cWlYhOoQuN4/iK/84xORmsMZcNx2z1kQLf+jaWB3IuQ+SfLOHz
uneu5gwTNT/WRWYLV0meFrJ7ynxMrJvE/jiPunUI0pZznVdqXkTFOH7JYmarSwIbR3QoYUz8uxVa
dMRzxnkSG1r+YQ0xWguL4k8bG+OgQpP2Y+82u/tvP4ZikiqHK94yjD9giUx1tFZdRvFTVsNDsdYc
cxMeuwdXt9oJhTODMy3HpVTQrrg+iaz6/BpdTV2dtoOSqJbAqPXkdlAoFZWcBBUi2mpF7QrLp915
HpxhRDUNZe9uL8t6af/vFkF1fjLTKHBsVYhtc4BDwIrgPBeSP/9pYXUxd7mpw3RfBs3cSgTx0y+K
GSqWJjX0zkdcPeDBdd0gs4ldEz4g1jHHgROb3ZIBwcOD+CpQcTJ7gi19i6D39dhI0jfnpA5OlQK1
5LMHF+TvLUFyNhfqrweIfpetSWArAfDQX8k6CUQuRP6nOjnS+gla+0jZwKXCoK1knUH5dkdpBsBp
LWbTOTg3IyGLyPcoaMzGu1IMVimQWv6vpzfYtii9rrmIsX7U+UkeUEjrfExoffHwCNmQV07QL59d
700rbBOE6GZm9KgF+KsdX1TteW79knCKfr0wlJOe5ileYe1RbpHOMdz6hGeNZXd3ABbkXkJkkBRX
oDwBvM1IT67kWSNzwVG6mOxn2Nf3KJw634HesFXUtB7LUXchpI5u1xExxFG/lue2drPkzvE+BHSz
8WiDROwqhFQES5qc6lIVWB8EMntWJJjwwmSvVntUfikbHiA0e8qoHvmCeVv7ConWokVaVpMdI3IN
TFANIbQhj6ENWhTH3TwYCjgP/SkuVIH66VzK7wTrpHMlT0Eki6MEUhk5WLZl4HdNa1Rl/qRWI2zF
MI+9dJezn5QO8O6UtXQrL8UtmwfwVYvA2UBtxpewW46nYUKzVB2XITiJxccUQ5JfrYrblwbMpEeM
GnEhyjH2OAyPoRKaQ1//dHpaDiIRMFGnSqR+FLF47Oov6Mgb9FwRQrIIqYYjjA3C46KBn/RZqy2s
l6jqCohtgCbTgH17rnZX68/t9NsFQ52zoKJbyPvtsIQ6o/M8e6/5Xmnpf6/SWGVmh25bVDZEuPmg
qXyO1SXkHyj3aPgRgS+xvJzLwNYhgBdZ3nUd4nZ9jyl59vGKETT3ivev/mvQG/Iw1K5awmDFxnxk
aEMMVLvTOJSnFCiIGXHmFQfPca6nW6CHroz7pKsr6trbO+EjmXZyEjafKleseTCHHOVld552srcR
w2OL5YkQ3/ep3rG0aZhP6ZnAePxH1iBoF2gaAH20UVFx1M52Ygz46qMWLZxhNpts8QF2n/i4f/Lv
0Xfz+9b2VW6tHUxuUfjO3g5ZMvJ5Q+KTiy5XFqUSR4XJiJ5GLvXJzDUBfrieKI5+vSbiV7C1BdUj
DrZ3sJ20TxoKLANPxD7R58z7ge7i28kH+rgi5g/DKDUc4d6dA8Gh5jU2VI3dBHa2pE5qKSzG1Til
3iPo7qCC/pRNFozODp+w6UMRzek7J2wVE8qMtlkM2sAtkAtaw91hqjylA6pxikBNXQj3SK1BKAHj
2gEdDJh2laD5Re+yYh49wOyK5OLJYj2d5y8K6HlTDUDpSdSNyQ0Ojnk31DWL5CfkbkzcYQcuw8qu
lt8k2Owi2CVRY0rhTiVFQCkN5//BoJID1Y4C0COObd73pxP0NJuBOJfbNaXAHE/n+voDEsD9m8WS
/wGv+PPMLxH0BrzUirCvStIYHsiwSpJ97L5d5RyUtOjcnuFDuwt8dCZQkdszOyVbqtdsVKU9J7O1
uo1O3LnuuHeT2RdqkxWknSYvqYqRS5zcMD8XMa1agmW24t0UIUsTw01fY1Ix+E5YHBVNkVOaVH5Q
HEMVUI12VgjDgSAxwx5COOYclImNQjbVPPfDvQ6sqGF+occ7nvAeykBsvclwEN5Tdoi4sy8znRXS
iUh9lsAN2bn5lLmyy1j/AX7vGhlfnU0VwAhEi1fdnxe1XJNRf4icj5P+VO94cXl45Cb1aXX3y/fh
14FwcEHIWNT6YS6PIZpusV/6L1S+KAFqJhfJV5/LIJCjkvdb/IcHY4735opK+GdNgTPAivuqsrT9
VLsjMP9WxUhtq600ELCcTg4VJutsymgvKxaW3u/boPZlN1Qndulb6OUHQ6hyfG+e5aiCqw+2Ilvc
ri1hhOR0NXToOlHlF2Be5HwdIrJCX++FVuHRY3fRVsz8DQvlOXCNERrPqVbgV3a5/I0eAueZbVpK
BFd7KaycfaR8AFCklOr18VKE/ZR0hs99Ja3sVudtd0gU2KqXWuYXcMIs8wakJq+wCLxcJ1PyhNw6
eR4cNvTExEC2m61H2N0cN7KVS41gwd4ZVPTOfP1CT8x8FttZA+USB+s9QFPyd+sIlcsSEGszzZRJ
V5/hp/zFI3VrGmywp9Ilkp0t1jyxyVhlvFyx9syDSvbjAJSsAuH5VsFMCxax3aE936dUGz5aQvFc
9RWBcRrElWyGYFkhTj9pR50dNL97B5j9B/1rG5MINCYvLCFXfHkWyEvAWJ+yoGTXzHOArZJrVl8C
uH2gIsOnhG8x6+gMPkYS5XzGHLzreLQ46FfbNTP0sGsd4gYQZbDHayLGUKhLgghjdJ05mIOHMxtV
n04FzW9kVDYblk9hq0ZC2bQQcTy9qFFX59wCFh4UGsLYIA/cvKdg1kKAag6p7blbL23N+v1XZaur
pDnMgvaJd8BrUNokQgseiMzm9q/5qbWO+LUtWfr3wVtni8dSXYItBiIdtt6weBu0pt3SIPGW3gU+
SEY2mB1LK+BmLulagKQD9sukyI5vvwsd60ONEebiYC4TpRxObBWL3DepAkbTN7PadIVzcZseSED/
bgc7AKLfCbjAtNDrQaRAU3EjXlFeoT3slVuzpcScLhZbDSXUVh8Xg2V78kLYq5CYBot13QszMdJX
XguutzQMqnQGCQUePqS4bJA0XF7FmBqNy82ZNkgF/KtCp3RMd8IIKGAzyatn50WEQDPe1Piuwppa
LPXK29O2H7GuEhFGA/CY4OyB8f8FJWD0+m1fwhk1xp0l3fSEKb6pCAzWw/bUOxj6p5GZ9hpxz6BL
abt0ByRq3ZVgk7q/lVEZsC8iIrWHmGZiWXeunr9lD1kSjPmSE6Xz5Va0WiUoZnsfedq1j17MMxh3
eZh9Kg4chUxpNuF16ULqAiu3C0jeyS8rIXEFEcTFmzmUQNgDqeaVqRRyzxmGdUjSa8zQDDeMM+os
/QjvFsmYLI4Ns14lfbksevmQ1TJ2AlA89p/ofzSrWCFQanQakM4KoKgpyNgGCVoRRDTR1fcXnYxd
lPVERkdRb7jtwJlJ7rKmVdk9+ys4RNHh9hc70vtJeROn/ntDrcGk0a6O2pTipg63Rh8tW4Cyuwzt
ETGwvG+ioNqVt5EiPasE4IjkQ/yaMZFEkvbkItYEK7IAG5WoXCKdD89RvIq3El/7s4TSOt9g1iOb
vUc0jhLNTI50ylKmLtRO3KpKpIALFnrDx9sCv9bgPE4AfdLVqqdaHrXq00JHL4DfMpiihh22xr7k
OhAW2dopm/Jkgnn7EMd46sinWwNtEcrq9EFh0OS0G5LFHGdF5XC+4MMjEojbTKJSSsSrEXmP/s8u
VVRgNEzdb8QHy6kidUN4Q7pXUxlzlemxEz8M5GjbYWSPIvYtJzVAZWmze+lRej3mz3KuNik2ZhuL
siMHJ4PH/ohuvIj/kznKb3Vm4QKr0q9ybs26t/wTVKKZOjFV7KL44AXfq6jr/2Ee+7aji9pTiJx3
ym8OGuFj8fypXk6084TlB8mu+UaefxEjBl7x3/RNdlfqIVOGy8r9l1PjCfdHdrccDP/+YdUnyNWx
b6kNbN2HS7vserq9eu4BBcX8O4FAUfm2WRXerppVt4ozoT8qzcMEGtSSe8SEttDDTPV2ua0pHT6d
oBqgSmFNMk7RtV54aL50B+QKKo9fjhwN65+qdMi6PekJUNMrS+9arJLMW/NvbG4fsuRm/9tjmjS2
txiVDT3DbXJCCM4NnSwTvesgYmd0PAQw9NSUU0p/HmGECo6HtZLjOZcxAzCwAU3AGNOtR70mHyC+
GxDC2dfqz8u8N/xL5cBYdAmpaa5eWGpZoGQD5SNJzlCxH2URVRAYbF29e1roGCBhTJKdpY5jMUp9
dRT9/+kmod71JjXUq9ZHMFzyQSsqHMi/SX8xk1GhGn3WySqFgrNuor1rRgEaGKSNXDP24UQnvf4Y
1BYBP3P8KRlSgqAFNcFm3mpVF4wHe8mXDZeNYdDDqXsbpxOeCOuNg092emMukoC5qq3VsZdTUEyo
nRb19Ug3zA17CaKKeTCvfhfltlLLo204rvyYKDBuaxdJut5xxSVVc2F4Aa/ZcAjpuwCQSJa1qwR9
mxePrle4qaxIOXJ0+eZUEmVCSDfImG+5qbDEcDa5+foCcSE050Y2vxdQJQIg46byg90TudfAI0E1
LgpYFOn4IM0HKzbs90DW7awXNAZLUiUKpBbfJ2fl2K0WC+R08RlbpGJV33tqOAlM46bkg+oyOUQO
14QKr5EXuEG8upI4ghSvPVnt6DUPCYXYpvl//apgtlgyM0hqvQr6J1t2EC1oleFuX/Z9xVcXrOgr
2ylVTajG7SHt+snasqZ+vKCgMq7x6MEKBEf583/PcOHA6391XuEui785JXkq69Xk6LiJYG75/TrD
sPxkoAayDARw3eDzToL4hFaqhUrG3d2CywuZ5/0GEuOWQFlgDqRFIQW/cF7edK5UqclfUH2Xd0Xu
rblJ7pvOKPox20NtAyIEyjiTdKNNghkV4q87qirnygC32orEQPxg5055Hlka3R/8Sn0etLquwVHO
8bGTGGG7E6JIqg0d0Hm9PrgaHY1QT2a5f/LWMLrgXwPLxrJ+XY4nHTsMbJ58lAo2KnqkMv1mjS7O
RtxM3b39EUqxkMqcSKAZ1dcaKYk5NOM0vwrqHHaJbZY7tzqwo8EXDHN6POgnjOW0xwtIc3THHvFE
M5KTydvjjev/ndKpOwzkv7QgTcGdexxPswLXQyZC3G3ieIfP+E1+Cxa6Nj5nghvJCdnSJD5EYyeg
3TuNy05tAjrSN6V024A7ZWrPtXp1fNNQ1HJxrr75DMaN3e2g294EX9uvBnpbprQYml+QuDHWDg77
zTstPXttKfOegYNE7O189otSS2QgtfiShXYWqdxsa+tRY1VgYAla+sbaTNJj7Rd9Y8o+fndt1BaQ
rB2BqECH/LJnYZJOhO5l1fHs29nRlIcYz+A/wg4H5OVr8rh5/ODa6XR6rkE/mLAFtMREj+RqAKjk
JQk3W3DBKrqOjdn3Ej1Mb5JtnbaPrVdJFw6cg2tEcgtyT/um5Z7gO3Bdi5vFz90+yJHlmouKoRvs
bxLvyGvsIjDqQkyPC3IVwPyWQJNnKcodpE3Zcly0ybNrP/cQJfg/I9cGPh31FrFarS6I5pACCJC0
mY+/VQENI4H0x99h/IRhoGPtheZHw2qkFX+coLu0W5G6+XVgVRqo822cERwRrGI3yDoT408yvJYE
KbCT05qglVMjcbsA/wLVCnqFrl4o6cKfIw82DtDnh5giKt8Cvjw+c8cpFl1Wh0d4IIeEW3ItFA+v
gToX/7wtpkbBHKwzsJdfuZNAQ387/xAtjCVsY9f8D5EgHTlYCg0SGstcNtKeSUefMHpW52hjVU2y
XlaPeYj1GYABUh8G1YrkUM6rVYdM3FX7F2ZOROg4K4q1hMc0WWlRdfSHWhDILIl6X5qSa2z6v8j1
sdYGIefnWvT+6G7inLA3XcRCfCphFVqoMI2L5c0QbTPZlJszacBgnWYfbLwZ/WBPPetTwqCMA0qB
3ALmdV6uEQ+Y+vnSgF0z52mcucAvHnBjMjDzACj9LFpgKXTrrpFtJwCpqdotU63lI2b5AZz/T7hv
iAo12Zam54YpeqRqTtKvu3ki36JflX90SyhEyg1/jS4vfGzt69dBWBVEwP/kQ7Ba+MOguS3VsSJ2
cjqm3thr7IbUq9uWkhmCcT5mxbiUCLFjvNFoNtTH+/Fl7RMRrUosj+38GDgwJUC6ahA23d8ZCo7T
9ZlLrUcA7kRMlEDbWcN66FuulmigFzLe+IE4qzFsZek9WVkk20i2CD8LQIEzr7f0IIax52VKzTkL
KlWl8A5p8raZmc4Wo823YKPY829mAhVTdgGjaP4F3zhdbnQgS4pDsDDbpn0Y/9x/iqakqqk6bliE
N6yABYhPRenSgmPibfkqoha+UzYzJ5DiufzoLHOwBPu9I/B32YH06mhn5JapXCyFJ9oamvNXRXPA
jZYb8IMW0YaeoPvjqF39ofezn+lRUPrcifVJzXXFoIrOI+2VfxXPfQ2jNb2kDWZcF3y3IemngCeR
LqydvOF5CDCYDPm07Hrc9gDXJ6H0Lx+ddigMJJQShQi2594aN0/CRKV0+UT6HTKh1jL/hO8JbjE0
jOOaI7MSREyCSTi53lFur3c1a2Fe191b1v3tfaacJuRFtN4fOMX5TUk93zqe+EBAPuaUK3UMgwdP
ZdbkbCSUxrcPLVOYZmd6w7RV8fqfZOoJ9Lxe/3RBpYXk4maUqwRftHjGh2f0fZuB8UgjmuS/G7xN
jMZ9+czsOBmZr7dWlGlLKb3CY/RA4dmY4LRDOsAoCMaQWtTMG5l617d5aj/AAV1vb4jV6EWqM1+s
ewK69rhiubNGsL3g7V1I0XjP0+KhgefXjBFgBnzcRvDQutvPH/QSgLGqbvz6nBuA4VuIGnSmGki1
UhdI7IyrU2pYjfSWIVb60RxWynND4LiFoEOQ4yo8cGdw1PGGpHRSqR8qzBINSF7aYSC0Vv83HvfW
wyEiXWe+PL3vsmJOYvMhg57Xn9zxmhdX0xodhdr97NVRAaecx67fQ93Z5VpQIAslAxxDvjHWodlG
PmF5/WXjaf0PanrO6bbKLOaE25DsBpj4l+Y5cSLiG7M1g1GL5aYkn5N53NvHxqAHQH5iI5tJDDym
MJXF9rYwPKaW+GgDuRLltHbqC3RqFBOqI8O62alxVK6HuH/xBXPmgz60ogl1mCfYLIbz2FdWdUj4
9g0S7FH0nUDLNp/OoRWQgk/0DHIIEK+KpsxxLEuq4Ihm9rxCaph9DRyhNUJPdZQm7iV49Yscvyzr
5RZOStVFlaQ9Zt1Lrib9FRjDYnfy9Z+mc9xiprgQlnGmqh054ZiiFrAZYMXjLg+c3ek67B3DaiE/
RdvDV1pJ8crksv6u4HgPqPDhVnigZDBhVtZDo4q+LJTdNJXGJG3nKj9aeqCqqHg7jpL0Pg3rjfwi
chmYzq68PAg1HxCjDnlcnCFa0RqGu4njzuzYPttnn53nsstQplssOj1hFq5czZ6x/av6FBx+CTBi
6Lk4xPxWDJPGn8wwHUfJG/8Nq+dcLP1DDy3n2zZX40KmZF5O0RX4mGbm9cukMxTXAMlO3gjrZzVj
VpikS0ZsQSgnw1IgCI0a67xfGpdF/7OaHWH/UieHesvAlQo7Xr7me+wb87yLZoYrZx+WZGbCBFhG
oYjoi4e5/H5GlmUkYaNyvAEBaIbe76vT1WgDjfkhfBuC2mxGqjScECTRKBmDffW0R4Htk427qKOm
+knfbIjpj+WdaI3XfBK0eeEFBi1ch/3lJCi8GHnFyE+VGHhvtdkfUT6wPMvOQHYFDzbhHu9TkZlx
qsKXuChUDZzM6LwFPln33Z2SVXermiDyVFzipvh5639mIz64sNDwPIGzBEG1/x0RKmx71OUNyMX8
EvRkU9Qqy5EkZBH03ItTwNT+uAHKO+BbEkE5Ir9f18qV7FWemeLMAcCzCZIoJAfceMWKRRM8e6hp
rmIlHpvQd+BZZDwyFpx6mEzTKFFxKP1coVBmPVCBvM29PTrsuRSq155donYB8mQH0h4S0SocjVDw
uBvew538YlmOygux9YTeoDJuf1n2uvNkjdOd4YAmCuyfzbqmzQhD8oKoEIHwZcvmfBm7sXIOALth
wEkVy2e5HZR7tY/663CfXAJYhEZbfEd3MFBIRGfVcvA7Lel+qrX9WvI8E10rfrc+focPu4tLkLX8
ICjCcIzcAsPC+P5p19phPQcH5uBnnXwnxs9fyIGieGAgMNzMh/EWdCenyZJsH2E1XVIHkRBeEvEt
AwtbsMf6d87LUOtfVP1qZXRQkS1MxXjeKkZ1sXsl8M0vOp6Mtpjnj0F2i/7NlN50W60DES0sCaK5
9zUS+ebIda7y+JqWpIPCX+rVCdzKotfmbY6WhPWnJPrpKoSXF/A6BP8kQ+JRxfMcdCmKPSCcQ/Jz
XEDgBG4qFsrMptnw86h1m1WVLp3k36QozVBNlYTSU6u750WJG33rNqIPsiqgaClW+AeIyNIqtusg
eeNKVCqF8Fp/AtaCoqkCVWATdwcYXvjJnf/zhHekNDXsrUA3iG/eRrXb0qV3MkepP0SfTLQN2N4W
mMY/hZdhWzuCVVPkYGry8WiY6m8a92AkmMQRfMHiPQxU1eYQgDDIroIxbJ6vpRgRyeFDnQOoMybr
uAT/eNKLxh8PexV/6wWVAcNdn5dgyLCTyXq/IsoXspA24bIgaJd5B2PjzcwbKk+3tm1wh9B+9I5/
8C3GQGpKnW75KGF02t/XeOT4kZbTf86inRRvaZVa/50JBfCVrjFMst6+F15XpU/qRqBJgjPtb0xH
4YgCrZKq6jjYf/e7rKgfF6w05YjP8CcQiNG/BBxp2eGDaHTD24v/5Fp4BkQewz4CIJYgcx0ZAig6
zpl+o9525PKKBHpav3hF5Nx8UU5SBMgORaZ2nZjcu2glwb6gXh5Bq4+N6npYYDIQ92X8AVmFli54
KDm0AK3iT6wuAa4Pe4QGFheLVvVQEuGlOPHsjy0nTBtPrVj6FjZ/+pMReEp78u7nFMfzOGAlanEs
cUMmP9TeYA6QuzUE4gtjYfMdi1PvpOBMYXvH9EFHVurWETJaXiSKMXUWHIteV967VxDYhSIRGnoY
zKkExiVuW4PuL0j4ADLFbGL+9qwzhRSKHvkzNv2j1lXcGUU+sPflM8DrqKCP07EFhMCS07d6RCgd
noX88tOjiqs2RmIlit7DabPxznBdhMAmtuBSVsiYAGJYFG+RN7/+/P6h86GeYOaCZVkTPnGIQyZt
kJceU1wrJDcmF6kK8yQG8gvQ9ygKFOlQgiJxBLM8UWcR+P7TZo9NxK1o6PmTRDA6wVeV3ioYaj4y
RV4WiRs2wpaMGGUx0PU+USKitKb/x6Y7eIKjcaidg6v6Y3/m2A8yMLk73A1qneazin2EwMDjRQAD
sHWGMz9R3yUat7+swGmlguUY+sdmvuMvYsNw0RQsviF7Q8HzaKOA/O7RazXdsuyXgYgyu6hRgiFd
n6u7sqeBDcGS7hgyk4DE7yVV07fz+uZVUaohU0TVdKcyH/VcRiewTCmU7/j+lVFvNPemAy1arBAH
QHTCeUGCNDBCxvxWvtsAywyakgH/BSYX9ZFCmseR1oMj4txFvQC/O+I2TM0Ph3GMJNJOKi5rkFLf
N23zDRTygu65ZMxma1ZhsvbtZhGJD6tGXP3DGyuadHg9xgf9Mk/fu2frSOCtwxvHSVJbByGfRw+e
pROXimhiW19SFA5aGnFGcjkGJUphtUwssQ3I7LKHom1srEiR9WM4d3na3fFHpDf3toLsXa+h0IzO
9aqfKAIfnZil5mKlclt2BU0FpKc1shdv6QMqZxXQ2sqXqjtU4Kdygp7RElSHhaQj3NezeUWLCZCM
eZMFp4JsxklKy2UvjzHKwQCGohcZy4E+d8/zGzMtG0qfMgnQnEP3nNgMlh1JoR06D7t5oyDjmFXB
uS9TZv/1RSVfEFYlsJydc0Xfeamfxr4axNVE2KeY3doMaMWNxeHWphADtab5NQomueTE0MKHAMdc
fTp5ewEqKVuxF9+QNph9q/2gfOoH1S8RocKSn7m+VgRm+cLfEn5Y/BK+cnecCNJ+Jeb27j0IfO8y
J53S9cnxvZjYkz3zSNROs9CQqgy+d7QBoJnGWJ74aRp10iCQWvARjFBd4GWfvlNWc2b67YYxcCq7
we7qFLs+3fHMrXHjxpOk/5iGToOXGArZQY3PpHZUZuhMOE1qiXkt8ZmmuR1/NpLeeQSI3k8GcerV
RW/hGs6p+TLN/9WB/W7u37Iiqvq3Of8Re4AoQ2BlsxmeGkaZh4P3Urn9ny0MH0Khc63rGRvE/XQe
rqFyddCB7gNYsPsTSNdCzGlPgWwksKcErmS5c07Jk2XACYPT5BqYfDjdb6FQxdF6+yNTB+RU94ox
HVpB3vungekYjWyiJ0vlvv6XyjrCMCflqLeUfdW5cOEp+Ke7Uy/ejnXUbnHKXOmmYRYyDGDA2avA
x0bk5PIwlXz50Z5f3EyGd+GrBQXbjAsCklRX+5oy+JZ6bhxbQD5OcjdSUHxLZaCIAWV+0IpJV9dk
oMtyrTmwd8kRc49Kd7KjGp38hwo+flGwGZHfXC4zmDxOtiepHMD9AKiwLrjRN9vzIcMPDcihuN3c
hBi/CAD8DGx8wQz4M/mb6eH7St0vC+esJZOFU5Gn0ape8mrePkhy2DCz5+UOjoB15pzGk/x6E5Re
OLchDXXK6qYVwcP6jkJK4/LeBcZdJF+iXQVlpDeHqotIR0qtzDASwd7suDU11rl2S03y1PFO1mKP
oEJUkAVa2ta6MICJtaHIclcMJw0nf+lhOE/dMjWiQUfmXX1Pz0h3b+UVgtCHCNODE6viO11cVA6z
g7GJE8FxnWSUc+nKUHc9r5tYAy7HCEvucJ8VNg7rZ8rSvvFwHNUYLveObZ6x2nL6pEFJE1WC6vYg
JozLSDFj0YAhgBls2i9f3nI+rW5j+KI6AuTTq27p/veegdEmk2NvBsl/Wr92BVNa/a1xaycPLdEs
SAzrBWrH71FQkGELYojazijITJtechmeVBS2Gg39JWe4314Adgq6slfvip7iGHfaeBIi5ahYmTBd
/RD4YnS9iWFItvOoVQn78os7FSdoVZ0jykGSfiHZBQdcbF77s9Duv2yNi0tXZGzNAnABzzdiGzRu
Xhu/KTL1Eic0FEnq0kARsX7Emyb6ZFAnH06xmVL0IprwG/wXECaaRgcnCJc1vBrB3vk0LiS0H6Ag
Wg+uU3meWXt8CvXi2z/TT4xFQ/4fSemfZPi+L4yHQbDj3lymm3d7j4RFUEL48Q5b7SHoH1tTqw38
6c01mYC5ExyoU5aLUOvnux6TLJD2gaqIRem2ch2JuarnbC59jAC4efAq6gcbegUZJIf4CBGwxfvv
Swqcp8RTWTrM+LS/2q8oIuvOoIl1w0+QzXdXzv/2YLTU42M5j9cFwX+3EFbIxXnV8+/IzGvuwsm8
siKi6sdrXkccktj2nmUM5g3/eGaZxKG7YvAhPWUfKrPIPTZt8Vq4kJr6tNtXws2Ejk4bUSe2n2XF
Wnv/lfPGsGSBkHF4OzoOnz7sDkASYENtJUPOhSQkALFR0ry19PxmGrrutPdAHgD4/IxV7f1XAkUD
f4h3ZFLddN+czQSyvwTOQWHcpDthA2D+GVA4oeYXFj/jXPiIeU0kQGV5++aMFVOrkt15vQXTcwzM
syulPaNsnGSxCqtiXqxgidYWX+Cl18Dl0fLvERmNVqbxG6cGjeZutNWi0mhdWX5kzRWWvbr3VCMr
ejMg3BFbZjC1DzXY4H1BM0D9WoQL1IfYFaqARGdwAsgIxCLh4PxO5mwPohwDjjcUxL/JZH3qsndP
ARped300/JOzwJ+nrf1N84wlMoBzDGRRBreb4w5bkSPNuh3QnMP8GfPUECsS534v4VMo8g9kZDCh
KGkoA+abQ+oZS85LrUXGgmzw82iYKzXxGZO2Dp/zmPFrpTRxqoyjVmze8/qlZ/LqfQrrM7fagxUw
c8QbroYCPKRffJD7w9xuj1uGuFhK4J2MC8+kZ+iq+cyf84Jw2Kj+sZKVcC4El+y78h+aPKk8NrEj
jdIrTYkHHqdJWDGfjHVg9cw9/d2r0Wvco/uf0YtUqu9Y9C4jiz2GBQQKOYiwTcZNsX0oFCKU3fUN
ZkC/vcr90GBa3JKN3v4q5Eh891PMweEzFbfgAKbXHXvOgpDCll1f0HYcWyjI30mG/ECHpE0omb7h
SJDEWBxkq3aD//JNtbGOJ2TkgwHH5acF/JdKaf7crjkVJq3jPKJOLWlY57nRZm34aCirTmNow4Wx
X8LXlSZOacPbiqAGITTaI6kOdpnW9hfwNflYHfDP8KDE3TRCi5O+P3Xx/l0jLFz48n2vyNOC2xtK
dYGPIVrxHC9+mcU08PlsSG/Gk/4Zw8+SXD+d+QBVdDgMcoIKAxo4yuMO2zKR802EqOxhWMMdCwYj
Z/86J+vI0sbUi9C+Mv5HmwLHoVRHISbMQpzwumzrgMemsbcox7TEMUFkFDLNHLlRromrZgOfa+Wg
5ajop5oVuQ/vFYW8FywL9hrrH4kJL/45vFacMdeLJWXMQdJzviKrf0v0Qwq2zHl5tcCgP41kFNtB
z7bCjkBSC0AoUT5c97UEfRlRa9vr/dnovtUvDK3v7Sbeu1Q6p7ZuCRjQIOTXrGzNfQ7Bj157X7SL
UohSjdDzDV55y+/3EsvO3AEobPC8MJFqudE62Irbtx97DqVshjRpMxJkMIIcsNHFQLNmvN9cld7z
kdD6R+TGQGVe9c69ws5yV2rTUE88hlb4iFa8ZZczWiRIW/U/Ww1YxdhwUxl6nTQ/cTG7ZHFb7dSN
N52i+bcy1C/FTaFP2A+xAGWQ5Pr2c3WF+M2V90qOlwcGv4GRG+5vFk5Jq6P+n1HNh9n7kils30kX
+Go7dFq1bsRxX6ME2H/c7hx6YUSPK6aUh9JAh1Z7p5E5h0BleOZsHYe3D7iserixsJ8diWwDTTy9
nyZ4YS04BXWpoNjJAqEan4uUdan0ypZUIgWAle1O28VWCDG3qW7DCABCuh4j6Hl75hH0ZX/CjMme
rF54o0ZCDnvxuvkv/O7qQxHmWOE4kA3EHkXJfmWUZdcmdxoSFCzKG9e+Cdv1Jkd0y5J1NdplSE3x
6ChGLOO1uR+fvXG3xTRy5OQBduwiCweLyt6FeDdVV5y5El+DAIojUD0J4qavZdmlAQMArdijnFqO
cOkWcE2OgM6/r89NDYCRg5uwFp+hECE1BEoWZzKzz7O67+5bmfNwgzNJRhlOQT4Z3J60n9onYhr0
uVeOablDOCxumGKaFvwmRtg0C4zRz3rNjE9gv5CYmL86CM0pVbn0bSKtqvLT/OLNmyiBpfV8DSrD
fTq7QmoItlCj288W400hZ3Cby0j7OzYA5Q2a5GYoD/xseqdhOfwHVbZ9qGeXGcuwK2ir6I4q6IQm
WDC+YxRGPU/Aypp3hoe5NXfR1wn0IOCRMoNynU+pw+D8l7s1WDA/R/DMBuIneDkuVpGgD0P3UkJH
9KKyy/NF3tBUvV9TwREJC85UbN6Z5SxuaTVWMMOC/iW970oQNnbPHQTNsnx5On1u2XTswip+OruE
r56HHLYYVCn7KHZKGjXbH75C4IgEMy0jD+errrKuE05PqwkE9Fj6E9+34E1BfR45ak3e+NApEG6z
sX/W8JMUM/wBiFs19cw4Yvezj3LPM72zdmPqY4zXpnuGl/iToyCScfmwErjSeEoXQEM5fKngH0oe
oIhhEDRUF3XoN9+GbMxV/PMgF/qUHKPcDZxpSZhpqfgjaMbtum8pJCNxg7dp+eGd+l/A1XeBV3Jr
YQzYAUXLf/bMYmB4GJ/xVlElKopAjYRbLyWl0GBaPJy37Yq3FHa14wq8Z6V+9ftdGVezL52Ol5UT
Ziy+0dbatK4U6jYiZHvXee95iPUs+vnE7anJEPzK/jP3yuQLH9zF2fo6baww+yvqzrwHxgsz/fZU
1DLWcedSXq12Nqa2YXfAEXuu0wxaipB5/NotCqAu1Ty5bAZgSNir09VrlE58nomdnwuYglPpyPR7
ELaqX5oWfaf0iboxteyc+HD+9ThCPYa6/PuGKavn3dBzXYJ1+wDhH4F1qjZnYMv3VbtIMu/SFWb9
zBkkR0qMTmCThd+DdicRjexUPdIwJw8O9eROp8d5M94GY9Z0dn10YqtHtgUPQnGC34HqxS/KhJcD
7fHbCTWVrrhr+BqPekNBnhhI0mwDYh3ftjLpg1HCtPC72M5Gi9rO0Sr0SHGZLMCBRo1uq3tMUAID
eOaYW/xuuEOTdkgmEz3FwqWpv/tA9UTCagibkdgLepCZU09ae4I6/3fuGbnmq2sH1XPsXdITt4+K
HmcYf2nTCRVTE5ssB8dpBa7sC029c2BUfwWpQnyDiUWX1hGmhRskNk1BhXNOVHpiRuuV2t3XYNVs
U2qJ3mwfYFU78nOxLwWAEmr89R/Km2YOo1/+7imE2ccXOynQ0RVIEqufPGsRVXfHS5lH73vnLL2p
QVsQ6eE/Gd3bqhGIb/AzrGFxHV9pfnrfvrjP7dA3wiqJtuK2Swez8KYWjK9cEDlI7janSI3G+kks
FieDFN81IRvVMrSfsKQ50aYwiCwfMhn/oIl/KqPiTusKoySff7LaQrwbcl6BMkjGptVrtx37SYiq
tWDYRZtpDPzhQblCfgdS70O/yW0IsDKg/SX/lZRaDgbzu3GcasFMj54wmxRNawQzeDyJl/5TM2nq
C2/kYzkco2dMdsHHZxLJ59TuBaUw0tQS7eDwos6rO5QanBj9aLWAxxoxPJ80N/pv5lfDRuIovorb
TRb2XcBmWY3xBJqZJf1TW/92NWYRgh+37oIzYCLAdxZyDB9GOyHShLHOw/uklWTIEPdx4y+3KH86
+2C/rtcZJ/QTpSDKS9GLnjXJz9nHJTzXb9kYld5mWFQ9DP+/1c85T3dDhuy406d4LD/ZXZSLT4FS
+18XJ/FXgSDRsKe5O0UVvzV7HWb5z0ogtQh7ZD4SMP138QJ++rQTuvq+fjZDaPu3KLU6hwAE7zKv
lLEL5lY5wtecf84zyLdwTGyRlOyCLNoyIR52xvvY/OuPNBS5f3oObyQfGpXHlGFHnUEEMYplF55t
f4Qb1yBc+R3V8OvLvfD7NPMOirl1pBAErzs8IKadMGTb44dq1AoIqxVbYpJZfJ9+8qf0ZS9x178e
IG2F7YM1nhxT/8a8/izvATf4/ZZ0gmindh3rz9iWdsZBJGPWXVdK27WosK/LiPLjPZjqcyaH/4BU
vmVR3wKFD1EPQ/eoLzDlFtVpH8DUNSGcGCrSArHIzfiJ5LnV4zdiNCsXivd8bWyt6XkqLpnbZSfG
BjeLh16ZrNHkg7+PTAy0ebCUPoJAQw5EhawC9UGAN+I2eX/dgbyIEEkVwxik/9KGziwoU2k9ZEbk
GMCpqmZt3CmJn56RjuJZiZPeukkj4ruU892OReSpo2nbeM7ybfqNQbo5+QKFIhpwAnI1VVz+qw+A
d2NjkDGN7sEmaNJIzIkzEuH3mI28RDlWFhKagA3yCWHITtS3xJV5/LBCsoaXmPQ6hNVqyMLJkK5b
BawzSMqHZVIJ+T9MN5RzAkzsHWxcQT+90JIZMT4rfykFzG/yEaekuikAZWNRGbB33xffLz7y1JAc
K74dKe1AExVxltvco8MvpUIZW0gcdEZwy1WPZ1LGJ6+Z8cS3nzNiGtn5v1ii1ZjJhXtu1PiMU8hU
dbn7nOTWqT7JAuGdvAbHtmhqeWfyU9IIdyi8byj7IuH3wHDJRuEWtPRial9q4uZkpt6WZNBAHkcl
5EJN3VJoEihTI8i2Q2pT99AzRpPlg2ZSdRnnFmFapA1m8RYmDkXbV/e1yJVpChceTKa7nNdG5kNa
rT9wqMyK0qOEj4IxcOYVrp3T3/e7NbItm/C+08RO+R4ahyKLVuqtg13Mv34+MyVSFf0TEVSoV/Cp
CzIUdGU9/PVgTUSGTEOG2jkwOvs2Sm2Y88cJTt3DbDOZCesHyG7YhVmNmVjsQtuqCQBlknJgVK62
X2FezqZJpgQEiWiPz9/Tku0FpGsumD2wB+GE5zv0zGf1euHX21ugQI4s1FVEk2Q6fF2RNCbZusL8
41z3BZ3nFlagFZqKMS/bvp/Kx28wzUv7QZKLYM/2MgG8GaAiQ3k/ITNWpjUpegqcRKyNUiWt0rTG
XbSfDeDuw6YBxNGNUXLIYZlOO4bZFp88M6VWcNYYmPLqs9gRaQ3AcveoBustMTOUqIliz2n0IC9+
EDGNSX/jjSUcNuOILdvnMKf5oMy5G1bDa65ogUbQvAB4G8qmlvJghQFn6maDzLKVZ/HufeExS6Lg
lcDtkqYmdnbhPD3xK6jO4yRlyE5RNYzzFO8IjuJLPUNI+8LEf2xk2bxip+K7zLkcab2nxEdZZNNa
JG5cJqV7JjkrIOobczK4yJ6bGGD2657qogDWc+n6RXcJtZK5o+K1O1tH8+2dzU987lbUA+s89+o2
6icpi/Z4knVOkKjTg2SLi/gU7s+iduFJs2RlyvwcmDgZmuGfmdoMf/qMae/zl92iorRYmlCpINoX
SdDDMC0yWUKb3+3fon6T+xSFnFVoMh8WvnG1QMIzGumTud1zhn74aoIDfivmlND9yUfloP4wuQ99
nVQr0521qcM+0CwkJh4+tulIh183hDk6Bkmgep6J74tjE+xryUTuhgM9qsbF73Bkio0MavNZ9jKq
1ZsruNt0jd9IGKo0bp8h80D0XqE1zUvZD6DjPmKsMY38F2LyAo7aWgJdaeJfBMyU4jfLvvPk8hVE
x7nm4keM84kz4bVHh+7IO4ocsRxcGUK/dYVovmPxFWfUi2coXYK0D3r6rwD9nFXOM3V5B1ABixA+
MRyyHzvBFtyWLShaF+eW0y5p/maVy6aFmyNZSIN3BV8rqGACaqFKPWFXD0QEhnkSkafMYoOVIp8V
s/hpXVLCbFSStXriNIhk5BdGSPM5TuB6MSHOED8YwLOrCW1yN+Q2OBYka+pfzjHYRtX/grrO1H/0
J+ujD2ej17zIrUSQ1H6CEqh9m4wGDW/7QvI6yocPoa2U7on8ALscZAKjVo1bU2praJCpxet/oWzQ
UM1sUbAA5an97+pfVro072AQpnwaD09KNH/m4iBu+ldEzwLRjq+w7YLPUH8QZ6kyL31iFcwpEcUd
3oXnNyc5GTdUfLuseLqqVUq0GDh47Gev4+37Up/2pLqOHFGYi6RZHDMSjpdQQ9eahjzLT/NE9a4T
ZG/B+IORkWzdXZ47HdrOeGdvFfs2jdbLYyJxC2Vrgkh8Hjk7v4OK4qUdBRfbWAarbR+mk2g8P1Vx
/H7OeoL0XSNnPZTZMBbJKu2LCMu5MQhBzCgwZUxy5tnNfhNfQwu42IucgfVO1fpOOAmvi/oToF6S
ean41zR9pcvVlnjx8WgzD5ilcyMI9AX8+xi0n5x0MEBq3KQMknBgCc+lxiULTT+pXSB92DOpOyd1
NVfFhPevtGoZztRf5wL3HgUlVR2cz5QYyDcpC1pWy2gQlsV3Ntk8sQXZBNC6Y+Wt8PTweiEw6W8f
QkSCvotv168jXxie71N40r18oNx39gfgVegp1xomksIgNp08bGnu3CER0eCUuCT21nfd4kLLzjk3
bWQieiN/M9rVITzlPceAQsjj0sxQYERrhpa2chMKjN0b1Pc2qLPujep1G4C871N4hV/UwcyeQQLx
MHWwSXJFYYhHrKN9V0fISm21QM9FMYP9IkA7QGdacoZast4wwWMkrz8sBWkgaq3fdnmETXDaOKGA
CEnypM8fOowgJtzIc2Q72nd5Mz7nT6xTu+ezmiWTE4JioLIPp6B9/xkjeFeLuPYCdfW/k6cTu3QK
aoLtsdu094HfHBahaSvzkG3a7kliw8Nhvn4QRwFl0cy5BJUozb+HFKRrCsvwWpm2vSUzn6DkBpUS
UhojEtBYYdGgR4chq3FvfoOFNm5hhayqDnIcQD6jBVnnQNaURX0QJxJ430+tmYqjJMhHfQep/UZH
jBRpTP69HYU3XanASknHciz696EHpMPmYvuBLq7tl0+IRcorJIQuKsyhNKHDVqjIP/XuIRzTjW5q
HA7gIH7xlhY48en6TZ/o83aSMbpTdHCvRHhKf5WiRwyZiqmCM700snc1SF0jiJw/CjCg9cQNbgHD
LRjqM5JfX6aY3xHegBhPb0Eny0Dc2DKXkciXa4x6QTqfLxMtopN1S3R/70ZIoETkCzz6I+pZGTYL
Ktm1Rn/KU5QR3rbFKp+IKGt37vKWZ/sefyLPplsA+ub2Gxv0tWbJ+jC2eFQgDynG6w2WwbHH13jM
DEhiunB/Vx9Y7P6FcAoAKEopPLe2y5OSPdOTm0PJPucT/1Mezw7fiOgAMLIf/a1YkeGEuKNDpP6p
NB0Sc1Tpag4vzU2hivt8RBLjqFymfsIVqEJBETdIN32RmDvtRlA7xmyZQsggqmBez0oklrmp4pNe
iH3KQdJCxZSGOwVNCG2A4ANKB1JTzGudVmL6eOKhx/KPzpKRKIJ7HWG3C00YYESBiJwi2zZcF0BG
4RTRKShLTZXwh9QH9JFo9qz3WT7zH38a5EG1v/k/2AaX7SNWflCPLQeEKT4eYKjavqaJ7vibBvAU
RgugiIaezfJpWW3dLasE50ydDHiC9M8XIMvvRFuiQwNlW5wF1w836xKEvtgNGu7obYKuD1CuXy20
uOrYD7SeUtHn0ZlLi775T7lIQBOJaKRtLwSvGP22nKxOX+40fLMouFj5EtQvL6xCuFxbdsoSB0R+
xXcz4HX3qegvBXIKSYiDjgqeyTLpzV9ylfLRtQQ+1K5fVWo2o3nVfhvFX0di9gBRAQlswx7NdVsW
au7qPRQ4vIv5NiiI1tNHiX4svsXXEbwN62EmXK/AMV+/peEx41ekHz1+QKBBqKCF3C7B0bcD0wvb
9bERIFdNElQSlFSOKyDNkGr770d5wM8KF7BxdS+X2SEonKXZn6ZcKnbceqF3HeOjoi/5Gfyi+lgy
fxR4m4wQA7S9ABVpSxoNwdcfDhCDxes2XgzHLsQlNboxEGGLmsDCTsRAS4DyIKIHnJKDd2ETHvHm
/5sevWHysrIKC5zI2gLjAegAKRnv/P9GkzllfKs1Kdw0awQEo/RF4LtIcs7mj/oNb3ypel+7ewdH
7s+HbdmVddeND6wMwhjOPwHI/rOLemY9evfm9uWg8dAoBD1GsLvDBpCgiKDKZUz5kauN/yS403fe
d/+RwH5DTBzCF4bHXhc80v91w/7JAIJbOSdqvquUptEyqAfVMSNz48GV7Efp9VJGncOqLs9j/sph
1CYU72M5uqDn6PGI6gvNE4zrbyU3doBNbYAy8q+Ou2tZLiEWqVK7BDHR/7Ha9q8enBZ2Gazzz3xK
Z2N7FBEvOUmm2ygKnyAWDTJJFCGpCMMgdf4Y38FoSTfx7dd+uPN2DwbWANkYqgmYU04JJUu1sZrI
+HBgtiaioJrxtqFujbUIoheOcPIZ91AsnMDb0JMhVPv+6tZeCKI6Q3MW/waykj8BHmRHvhcg51G7
ydvIEdsspGjBPBVBJts95mQO7cMTNSVAUdnoxpdz+tsQe3A9w7nSh7QZNYgGWZI6S1cCvReZVZKs
MY79sxTFgWWfvtllCfr5qzwHg0HSyvaYzkxP/H/8G/Gm+XKSbzuDQU2W26+/CjS5MTzFS4OGRVR5
mx48jXjZ9ZdKlwm/YL8HfyLm4cS7CXe/3zAlirnBHDsC80uO7NARXJitn/+1wJgGZr++4ouOgVzh
5FA/E7hjItdQadiKP0q5T9pamlzZRnAQXkq5EKD0inR/qfXjL9HHURt048qgtFyOTKY49SB+dSIY
JkaiS8sRxTvGH3Ve9La9s9B06Z0KGygIzBPQ+nV2/ExoixvKzO3CbJERYEggUr1VjVhv91jYgy9W
3PiMlcKSwUzt2eSUUVx++9yKd1xsJ8ysXh9ZzwS52yIdPZ/WMQoGaM+7mGn59G99shmx2bJS0Wvi
9HxGNino5ki/o1K7myZt4eXcpdOtcwuGhC3TeUheaHB+HudBBo/ybAsYCbZ9P2kF4MPb22zx8ggI
lV/cx/ukVb+A/rxIhn/EffINSHZyx13myCa5qhum8ckUy4HpEgDes76Vzvl1GdhX51hbdUpWYqGV
ZcPNx6Pri2rKqRxz0Jf8e3XgzGHyDifd1BPixR/Z2bJzLPvRjAOEi6LXEBYCVwPxPEPzZGgkIfX3
aT4mOkT2CMrd8+VhPC1hQM3hNT+if9HzjYHvaNPMPduF2ND9mE3f2dOp1Bt9ONNCKPMbC0s2gNAr
SHASeSC1bsVarVCsrjxI2ntOIV7RDGNx+O5WnPevA3TSD9FvLiXmIV3r1Jp1TLZ3WnAX2EYz2Une
dmx8WaHf3R0hPwE9GkWwGvb2PEmgQM7SkMb7cu3iJ46SQZDv715Mx76eF/9WNErui0cKc61jgJ41
/CGUdcEdel9S8OsDhA5FPZ7wXy49FvTDtuQO7RVoOwmFNH0PzqIoWDOaft//Us9vPoYjUpDmMg4z
ZAkY8uhejnlJ2DnJFLWW57JAeYb67qlEZcRrGkygPUT6KD/QBWomIuoJCV8lR7qIytjIbmH/L1f9
DzS7eNIzAUPgv0H4trE4Qwon4NwDQbkbl9i0wkfb9BZLCOK2wlsaLu0mNy3Z9zkBSrXKqR8eITLL
Sh/qkJylpIOP1yBb7tRsKoF3WXWvPaf+V20l4Ax3gDWGTWhVdV79YnpfzloVg9aoPR62f4jXTUwO
a0rfs39GkMTYZjMoiMWaYNK5zGYpyqmxrpvn/O8ypitEsPg/EPYD1Ud9Fn9kqjGjGDnYlLcDgMsU
hTdge2HPqEy643GsPtyd+Gp2o2qsTmNr7eV1bKA3PlKnAM21HD2BtSoKJZEaxm33BDS/ybLgkROD
LFOUavMbzn37Ms8Y7+p4qicQbH4ehkw2gISvDqIh4kFs/6GHVv8O6oe3toWp9Na1OLHIFOOY+kt3
Cu+bJNhIT745dVFC6SE0nOPGPbuLdTnKGC0M1uYHh7TJJ2c9ZZMizTUy+JPR7pRWDr8m5e+7Kfkl
1JMjYWFyjV9HOEO7cZ5O9XMxmZusqNe+8p6OcE+Mj4iKR/t1RIKbR0ldksOGNNodYZVeoGIBswgA
589DJGaGSwc3Z4gecdHQobMbo2uAPGMfqyWW2hF548g2Q1vdP3L/ypGQueHVr1ohELbELDm/rh2j
SYjiQTboht+gaXeAu+1DHYzPxoiKcVCC+Mu/kMs9ih7Bn9hhArMr6tnSZz6qLby0jz2MzTL3b1tx
9qNb+C83zluBuWk3v3flzY3E71EyiHyRcDE/d3ZIPj85jYtKxxslLW2ch+u04Cb6c5HB3StMpNSd
HddLEayihmDbY5TLth670bGLgx3eBHqKoH0C7tPTrEa/qqvbbyNIlF/9ABVnsNvGYUqPQw1XkPL/
5ii8V+zKNsemL2zWZCT9DQgUs+nhfTc9MmyOBy9nDXKvTrSUyUhx9HfmtJDs7qZ/4HWoqp54IA3N
R5VrwBLcsvv4ZeiFNAbEv1JtQOFEgiA25yNExzs8OR4W+cZhiieKDc60AnKzqeIR53K00QE63fMN
UcYOusFhhqF3slyE6DOlB2SbS4KCORL0vFtzBYz5Dl+hg1N5ZG18I1ATNHKuVKKarKowSSkrwLdg
4LbduHRwmT/bIej4Gq/VU155sBPlyqH0JwxyBMIQGHjHxd/q+sukVWWsknruEZU4pCxWc7meFWVj
pdpL3wDeBtgJERnNUmBWsz61nDwsujbuzcmjPiBKDfV4c2LyLdOMsmLYfBVccc/DHYsIEKXcfzKw
HMpaUDBItCNYOBtqFuQ/aw6kKLw2TNLis7DFnsa0h8hf2vZDlvvBFIUQ2Y9DkQoP74kfgnLO86fq
dwTXcqokbC9roUVs8F31VRApdIPGvuL925SCi7j3RK1n4k2O+U3nBAz5d229UQHHzj3wu40mzyLD
2NCMQzy+ylHoSHHlQo7xyzgHPzJabPpM/dn7l5gM9id/n3J3d03QG46j+DgOGfFo8S/8FCXWLRE1
dkspqHctedsQky+EDxugizHR3w49BxcF2h7fo36O0Mqf798v0BstPSQ0CZZVH+UBf/6zMoJ+M+1r
6FTCiiRicHLjakS1cojVbHh4Tk9Ibr+l4jbgPrMdeiHu0zOiHeY6iHroJJCFNEzeElE3dfsX1vn2
WaEyHgpmkOUN0ZoV9BH73EVe2BOjWl47550cuScbGzKS0wtY6J184XCg95MoNWlNaamGuC38Frz4
HewOwkRq8aAmUA0ThdobvhYFv9f8JA7cf2J33jhKmpqWGJVdVPCKSqm5UBeCjX0J0I0J2kFEMU5L
3w4IodjbPUS+JuZ3auLLgET0Uuqm8ZEBI773pb22RxPBuPHQ7adc+mh9Eyjjbt3xtqHYOJ6x/4bE
Ur41M1tOw6n0zPNc287x02GMcEgopqtoBwFKtEmz/ESy+rKAHTsFpJLZUPWuOH6J8VU8fOx23ywS
W3FKa6bdMbMydQ+G5CeKcBy3pN9Ro/xmYM6oZ11mcrC/FSa09Pvnaol8bQeTQ8SduPW6GErdKwHA
JOb8DC6MfYkceMSEeYBnVA8FbQ1KCJVWOsV++uVL0R0NCSooSq329eORc41b5x0x30bhYa55tWp9
JG00C4a0fPlljoaiPzivagP7MWcm1ng68e6kQsO+vS5H21vjt78/khtCBLDkebWfbON2k5yTOacZ
UMHRdovLsO8f12BLeEjXqbCuTNZ/sjo1wVp+L0DspvdmT3kf9sYRTF6exz0FqDg0fZOf1QtnGKWI
FM+7YQblqO+RfF2D066zF43gVU1ubiqUrVLM6VHXIVzezIhScSS6fkCsd6Osh74sTj5d3JXqj1cv
eob9aRnrntTYZGTLH5YobVJ8/PH54lI69Nj+1+Lwx5RJWfV6AVYlMkFFYGl7uvXu1CzLQLu5WNe6
S1Z3KO5PmpRgxsvRYOFGZr9VTnsp3Hg9/fLpDgNR6nqxpXN2SkWm7K0Dm2M3PLxTl2Ef4jjsQWFN
eGLJKUfs1p0A6S+t+ZxDV1UfW0u+LudvuQOsQvFhPR0ks61se6NrYDnd5a3sRfifXRwQtX3q8P3J
vuTy9LUNB3jR9gWauiR7v35AXuqUe7Ifb8zQZCHGi7W2ZLPeXIecwxzjMl0Rd6Z4onnAbEu3+P8E
LfJRXNvw1Z/MtK3erBnXipdOnTQOVyl3jMfwTRSqPTcSyQjBFx/WPSLy9zA8g0NbZ3snsnbggDjL
z/FLb23kJesGFnQuwPG7r7xnOF9xF9Wgf5EsugwHa8YXiRLhbPbec42T7dNGCs6zwOKnjtapVBDH
0zysKdVqEqpPeihk5+sjB8NAbSYc+yQ2qfDtwpDgERvQW6mczllGXG3kJfLrGBgGcvBdNmR/4mvi
Thnp9MVP+W5CyxAVv6iv2HcxnF+sy0Cp6Ji5NtkJ7QWSPp33gUj72vTefNx6k2XICp1NQ+rFrPmU
i6B7SNKKsdRJp6Tyv07VGV7zHOnWokL9Co72VTYZsuUaHI39vPzZJMY+tuUHzW47tpzKwjv7dFFp
0llklI1FPbOCdXStFo+awSTzVLe8d8b8U08ZVvxafv8FYbHtKIIl1yTn0C4WBKQCZbVzMr3NRh2L
cSrBEUSlJESoVgmlMJpHHqPWPyfQAQWhBri/N+hxq7+cnXwjd6lXW/YMFlGxZ2+NQBo+GR03Uep9
pF7LgYvdxedpLii0TO7YX0RmpQcjKhtt0jyaz5EKAW2Vcxaf+8uK4lld0beeMXQwhtsCeNmb9wck
RKD7rlrJgYFQ5fGWgsmcIy7UYkxdUhC2EH795OSW7rKEa1m/QjNQQ47//GNT56Twvxp42KWCjzHm
efgMT0FjME9dPC5hb5nsyo3A34ewf3xrdVp+lWkWUNA+GwK7+nBBQ4PUFyzpwZO/Q8Rv6W0U3nqE
uGcuI2jKhkEviLoOapsCFpinxamXe0XOwRkNE01qBGnrvNAfSeIm3KQ1z6gF50CgTH2pQ2Y8GRI/
s+eJXocr2+7gsWxAuV2+ZESEqF3u2QP6R81W6k56LE64epiBBymnBOk1DXhRVoldOuONVS4GRRs0
vIxjKKFDmhMn5mNp3fLi2pNWa2tONQ42vD8mjhn2R9A3cPQiY5MTn+fNZzWRGKYVKrK0O524vty7
pXZyjIIVqqERN9V2fhp+jbFeZLOu4elGcTrwFpsVZcJymiTr7EalKXbRRb+beH5rS0t//E/+lafT
7v3gsBJPLvinveGJQ2jji0W7oP4sW3wJWdch1EDaavyGcDBylE1dAa1qwzcMi1ML+9pXhxqtWbbr
0PA6nTwMwF08D3P9XHnZ4MDDQfY3VA2mcenHTI8QEuhRhT6LKyGL+0aMrQCdEGHeguGWLFgO9No4
SO2S6n716utBzOd0Jc9jaqL72G3AQGwjOSF7JuiUfx/flFagq9oNp3ZUz0PAijnfYnHJRkg5EnWV
4i4ka1p8+690zLNT6Xxxqoq1oya1xUOQl8E5AVDZsjuo8XU6znlv6dVqAAVFea7J8RiGJme+VZMa
PzXc4vHC46iur2Ci9GFIX34zEs/+dPsi7KaA4dSZpz2Cbu/WYpcMWfrDvvuP4TLJIwbT9yJwBt1W
sQj5GLIpKTkxoFp5rsbSe+nK5+qkWQ8tMrodEZcQl0BJQVYD8D4rnAAUNDkRKvT5Eu+c7Lk2tD7w
NnFcv57N16DeQz+vHO3xcWBFUguV04Lgtd/jd112/4cQeiIginRe83YufYzKOBZa7k25bgcFhtP5
kWCEeIzLaR68AGHAtJLU+5pLrc3evxiC/H/9b1j08S2caI2CPhtyPU7gdYx6SdpTuYmKJ/gFEBiV
8T6mhJ1D31CLKpdmFB6bxlimRN4+H7owgReRSckveLDo7MVUZIEb3C/W1ebSQOp7teOo4lCrzaIH
3cWFaI0FQzK2kbCGToVRi3wQSbHuhcYzyd1HD6gJundW00rLfuzLP/0gYsfi2ppKB+KM2A5AUsUf
lvRq354TGRmSFog0hpsxf5PO7JEFJH5bWLcnORqGoKgD5QTT8p41w2puo2D4cm1N8IuuzZltrJzo
TsZOv0lB/GvFnGwHs3o+Ipvz0bFkKwnLVAJeSzRuEk6OmQSXJ5M+6Sl80mAmVU3oe4aR3Nr3gC91
BePn7dyRoUF0v5gAYNOfPAOCkCtSym0AJ2q2rtWovUHYHj9zWZKqq7Efl5ku+rHG9YfOkgrGJiuc
1p8KO/p0NyWb7+DW67XY8cvneoYkqAHccqxVgND9G3ntJ+5piIsNqQgunTfAsJmCF4kwXPtlxpWr
BZmQWalPix2ohbKqX1QTvWyACkC4cOt6t9nnqAHs9RY6LQ5xQV2uQVnzzRoPsORjpEdVWudOvcim
a14fcqUE+db7z6mcKmzpVXCVtZMW8DwhNiEORLLLY2yAMW8dRUAV19ckqRP+MGEsMJPu4dQjZ7Sq
4h8vvpsg4qT4zlskmuKE1fDHG6SigMr70g7riY4rDI0vBCi9J8dYn9ep8pXsBEuuzM7xuEoxwGrT
t5u2IyaNwB/gi85rgyZb8TwFdS5Wbwu//PLjlx7xw3JeKqI1K1qfKmD5rEaAB12np79dV/IuV0ht
NYrbesQyx+NFBgWT5RTNcfrKvvoewB1HdJSgZu+z/8zU7HpagJi+ZAgrk1N9QDOlBMbxTySgYFUt
MG0CsimhzLjuJYLGZnqvz3eSPtg6D5a2aJhnlTfrzuxhPoZEuCswWVNRgzFb0gESlC7GQuQLXaPk
TRnlQY+8ebGl6GbCz+oVfKBaC+LvTyueqHKJZS25BcfBNjnLt563e4XQhqOphHFZ2SyLkQM4b5QS
1yFub96kVnLLXVCGXQax1YK/aeljzDDHRFliSmiViRnZQfcWl4gt6BtqeOjum4GAJsoDu3dz1Mfv
9AtjQCrH+H/f1hFLrMsDwRVk/pDLOmVZSRkOc7clA6tDjthcmIytKj0DNH2ASvUrKEGctEbm3Aw6
uZI/y3T0WrtVRsiva2+lMV8eRjyzcMFXAJkiYdfvpa+cIQFmasRjJvNDYD6QyAPFQ3xq8Th9MKUI
G0S/trJgBChQP6QbVDCV2E4B5Or9TOM12+TroXNCHie0c6FQo/1rKc6QqW2gjRX+HSYfGcAh+2Pq
RKHEOk6de7rv+4pcW71auTjIl95IsuEEg5UcMLKYmTi4pnkpVRlRTUHnuKK0fHN9JOgawtrY6KrO
MyF7p9nMj44IODMin1YynaMby86Tq1wUDWE54gt7ReRyyC7UhnfVWxH/mghLt4InyUPsdoNzhPn/
+hqlcmTnLJvhI92drKH/2n1kk/6zl7SktGa2eb2pEwS11sHin0riNqMAzEjI+4hbHCb+TkP33tOj
Sn44YVNF95cF9DgsJIXv4X5soJmd00AyseFBdlvKqk6Sw8dhynhsV3Nlfu5oenmdxSpJ8ndqR3Rz
8c14fZ28UTjxSAdOTZqgPG+o4gMZczmK3uhgZZo7tFEEp12KE5ry78HvJ6k4LYu0W1m5LLS4YJhN
m9lCQny6ttXFpliOmhbO5kj3CEIRR1uhb+fiRNLswtwOu3jQnv0Veoi732P59Lcd0XSgHbeUvdWF
+wZ5ft/uDLhTIg2OcDERGxPb1J3a7lEShkjyplTPycfjyaPdwOf3FXTnCm23fmLKQxXIhtgDBmx1
Tk5usoDH5t4cCXm9Z02IRtmRwsDeQwAsZvTS44KTfjjG9h0l4YwSNBM+SjcWTUdA0FpCxMKF1Yjr
2Ub7SUintQ6fJwwP2MYvotVO3uvj2PV+6L3XmcbiaiTWbEIIXIxZpnhNmmSIecOZinUpKOK2uOHm
GGfybjB7vSKodw2ffZGj9SF7C7Xn5p/j/61EZ8AZfC8Enjc+bRsQWsxQt0JNyaHF312j6aGBqjlP
vTh4nRlGRnafLFyA2TSPKfQuy8pycSYsMg6MsmC/3wbuWsTXiRuESHpnLB1xDBRoDNwK2mPN/aKv
eEdXEYviXIXuZ37NMzBMvV/eWOaWRfCVbJhB9gDwOfcpMVdsQ0b3yA/iQXkts5bOxpzvDSmZCD13
COEwj+r/Ra//ZETYC/cVAr/wBMXNDdBh24O12ibPmkm05jqohuicjT9hj++QANFsYsxA57LfOY4H
bETe0hjUQ32BshRbrbjm2WEWury2OwYNEEhwpqeRmTBFu9wYT3UfF6fOm+69NgW9P9TjZI0iDh39
jWYzXFNvJICcxdbS0qqTZdtjkVIhG1ax4npfVKH+Arz33+uT/CNP6A1wLHwUJtLLjb/4veLKfHKR
lLg7TPXjmAoJusLyLeAzsYzrpuG9k129VXwNhb4/X/R4r7qk3ERVGpITE4LiRIMdZmpWIW7VN+Zd
mUh50+gllWRRhLjBNVsWaudAEGBYT8iaFxvm0IPLG5Erm8VomZjR2cyifViKSQfovWryjF0R1370
TRvgzj1oFypP65udxHEnNs0KYjRNBghzHHd+HP0Zl3jr9h7BsBjRDyMuPIQn/vqA7zD1iwwMMUZB
IMISDzxdulNOhtnIYMIYDdnBWg8PMLW8RMLd4oez9OF5VnRWArkTtv0HOKD0l+gNUlJuQNREF2Bx
z79EDTeXwq92Q/m8rIjIMRc+UemOEoucuKoSmN24Z+k6qV1w2c23sN0Ou3R26cX2SJuUPaWWuKJQ
oYprM2UCuGnyoZV+p6MS6ITU9YRJyIpVtUJEyMQMZgl8bB/e9MTygs5s8NhFACjFlh4zBQW+Mdc4
1SHCKJZcnX5mdkhOHXzw366GVEtV09I8yG03oLaY8CJ3axyFk9n+rs3OogwFTUKBeJLfqjOfAVpJ
xud+4pOr1SF/5/0MhJhkMlQwT6fmt/+yyxyBTFxy7XezyvyXju6zznYP5kr4SOkKfy6JDuPyteB0
HCrGWFkeQcFkNfoQv2rYftopRkgeGZTvhCjkPK2B3u3HziY/xmFPGMSV3RT18XSNrZf9RK3/0ozi
SE56woojw1fKKudFW3/iQJiM+PHYDqW1zbJrgWWYduT/STbTXum/mAh1kTsGNpBq2QvIMCclp1wg
+YjD17jbGTXRk6ZuPnxNpemlWnjzDwFuZdmggCvUMwiMxZdHrxvcJn5CQqsOTQFC/g7T9wtSR/aN
wWT8y3t6eO3aq2yHeMgdZuPtdk8fv4ElTqXK8JGaxo5xcnEJM/Rfa40/fU5uQYCwWW2is8aTKRAT
L8pW5W9cZDhkgwghrD1bYKsjNNQw6z8DlFJa8W7Qcrd4eMTTv/tg/VOPFMx1RVSKyidrrTUO17zF
Mjcmbg8XcOYqzP6yYvS6XyB1e2YN4ElcDH3IeqnTUP1h2xUv3g65XyD1wTG8DoTVFRz8zFfNKHya
Gs5tPZr8IpdvAhv+Sdw81Izc2IIybXuTxT3sei6XMen7c6pbsvkFOjkbb2RkS9G8znaX4riT7eVY
+ZiG+GGEMciZsPn4c1ggQIo13bwhaLx2/5QhfegfuUO6bv+FkklbWJqPqqfP0SxNcaj5flP6x29j
1jBjd4aobpVIC8X5Zaob3eS0QEwvwHVqF4RMqaJ74Zd+KOS9bI3IpSKk1dWEOoOD0wX23c0/7VjC
dpH3gDrPorXUptM+TiudNEVZTFfnND7Taa07Cgu3ck18+3OkyKn9vm8qJow5DMXamoewmQeIilCu
RnksZdeKGRNdroI3DHLLvPOp5a3hC2S4AdG11OOFZRlXx4VllGwCK5+y/Nf5KI3Dn15YyVMbNia9
tS52RKHhKj521vuzxC9Z6+xPvwXxLKfUS6eTEHe+IXIlEgIg1QLOS3jd0FBf9jOqiT+b2QzYIr7S
26JrhJCJKIYTM0ViDSaBmJJ8mSTTXj6ZkQRXFzDmikgiArt0orYzCiLN+JfJTRfIhkXplvKLJRlS
z/TkgbNN/AYUPo4iqg3282vJ4MsgR58516J+SQwLSkaPMYLUPKwwFkgEfuuARTKn6NspFggOBH4m
NqKWL+Azp3kQQxhrWCDs7ljkAx2D6RIIXdgAnpXZCVTEQRB9l7F3xM3muGn7avaDyLklTAWfw9Wp
XrY2N9DYDEWOteAuKbyXrA9yXqjkxt5tFm1xCx0cz2coPzm/eBpKqXMPIKW1R8uxGogThjCRYciz
6zJgMG9gb27FM+D+H/AVfsKm3vhYcPhetZ0eW2MRKTMMcUJoqn3oYW6f7fWMBv6XaZE5c2c/9vxI
GG0ctPzH+UeuDGqBDPmap8j45LBqnkehbIHQKHsf1M29uGBxpbvsfC9t44Mqqc67BygV2os6Tka+
caJLPGh71ffvTASL2UI2Bh4xrcdDsgH4cmaVywDy1O9HCjvPqLlLsy8PrY0dH3tgeLFlOmlJoIFi
jjRSvUdvxc7/+ulJmMlyH4LwMmyd+dMThvr0PAruNPf0vqeBaHp8l6fpC30PkWXG9J23pPPP3X96
8KhGnWlT2HkeJV1a59K4Zt6yxiu2GMNTFKH/AjXbEwF4j+5p8ELpL71hBz/rsfQjrD5v2pWZnvuX
BeTm/rJr+9ahdj1WhTlmVbSQs6Z2cDPXGUHgcnnWmwbrP6mi2sSP+pafNXKWFFq0mKX4Tk0EuKV7
IOv0sCG+1TzgyevSKW+7DJDYFAlbV8EEygs7vHxUHnkl5heHjTFDFzgsl/EibXkMOLv0GGSbON+c
1wrEpdxd5EZRVsxza5kM7aAAxOWUCBRw3awdthHoqhEThiTiaIkc//nJ4NPMiPGekFljjP2rsH7U
XFOp7XqrWE4D3++f+MT9cVZfvbgBaXmQrmTMyNaVxge/lm4A+q9Myi3N0iSrlmDXSN0SdXJV20Id
HT6gFuUsn6Fq5/Lke2Ap3K8YPZ4SuQUx+1Wsq4a7YXXXnJTLqPNwwX108eXij75ckn+PcPoEAwrC
CfcpPCIUV+bfl0i+ya2YiMVmUicfwLeAbHEd4+hZ5RCEUl3W5Tvx/kJiptlqLH3m67RH3LyjHPJx
7MQjJrKq6ATI1Tyf4h/fM/WlO2QVLsAwUjhI3fNh51dxrI9VT/j0+F2KIpcP7cPA9eVqvPNI7Qdm
0lR0Me43094WjTZqyrHp7d9TskUcSrEckCip3n4W6Xq0V+Y0eIrwyxtkNb5WnVG8yoXO+FAZZhjt
a2UG3aM6tMiI/X/7IOrO2SvK9toA5BYX65ZrKBbxVyE9L8exn/k9k2hZdBZmEDVWshDtXHh/Dw7V
Um2Hk4Job4ZbzdS7ziTByr5ikBNxaMskJyxrB+xVR95VvEHTyM0UsYCDUwQGnHROggLLme2t1nJh
pPfOgq1xiQxVow9qzn6orGlF0O8d/FeRE6bMzoyi/Jxl2FrzYQOd7d2xAPkAp/I4UzuM5OrCMMeA
7wD3aPF9ujP3/n0kyD4zg0oL21njwGd9fiJiFSEo/VE4EzY0V9wJ5rZOu6hmlErmQyLNA53QVRBF
UGbkJ5/AdY3KugHRR6VRo42zFD5unztStLASOOL0PFKp2cu7VF5h35NJJ+Xk5bz0ILFL2phC2h5+
oj2NaFyVSFh59Gcf4dV/VB55kBCnyyJDduGZnPSX8xclW3dUFRwg7rWXIbLLs5HOSgoDA8K1mbGw
bWChvoTmx1eO5yTiS3zdaboO0aEoH6Fb/eeQ2TQyyKSkRvCaOkr4lpaAQgC4hguzr2L/G8jFd2ad
WmRWQvA91pExjfPEX853DnkugkqVXMzAxO+pvaPaHGoMxPPJdr7oOVK/xCVRW8w3ah0FCZeylgil
VZO5yH7J9lpEcFL9Agpwis/aUUlqcL4+Dg1eCETEfIxBE77CsQ8a8mgtV5M8B5wmUmqgnSZ9gi98
YButbifxnF9/yEZQNt0HLsGr3Da5vVo/E/DD8Tc6u6Eqq9qzZ8YL0R9zAqgmH39/RCoArJI7RuJO
Rg4s0xOKv/DyqCrBLC3LMEAjqGhjlsTEih1/aohvaw/AF0AiZc7XrbuL02vevXJnMCh2G+LV+X7N
7BbCGOjm7GPOCPHWx0TIrHoYgk2QrwgQsd74Ozdx30BKocSjllvzN0b8JburzaGBoGL3g7QAqGQu
Xch227piThgpz4+otcYGgh0AlDBva6f0LKanepaqbiARxaka69hhc8K9Bz1tMHYbjlZHY3jGB4E2
k2MKVObIUzUxLdCtkua2U9ZFlOmiB6PN+L4TB+ZS934A7JAtACKoZ0O9HrVijaVLut94mooM0k+L
oavMEQCna00qCMwBoapDPlMT9aXuX6P0vDshpbkQDXGEz426R/TMvKg3IvGElcydQCVCtJZk6dIA
FjjNysdVYNRmzLKp2sBQJxuGHgbtmrOBvOnk0KDF1ME2Q6cyMkvW2M4PIUULqkkoXg9udP0hQ/dc
MHBl5RkOJdqJqzNIfnIkzxbvpeRKJqYSEyW+Hph2RqD8X9a255q4yca05SI6H8ujxpVdgWUYaOVp
gNeGZ8vmJWI/vAA9MDVg5t5nZbnRtBif55Ch7WDAmfh+EHjQZzXlSrs7ST796JPVMvGrU9Gxw9wd
J2LXA7wJnjDZT97tv2H7OrPGCWCkqL5KnBMoTic6FL/GjXKEYxZ2qX9WVBA+1T3DgFS62xp25p8b
IBb19+MPHWVwRw0RVlCa8N3G3Wv8lCEJDCbEr79C1YjBopsbQ5X3TM6/NuXoDUC1ZnJGWfp4kbeb
3UdzwshX/UYFdnYkb8IhNBg7iNTHrDuOxxN2wuqC16UW5op1NK/X/efbtApdrq4Zy0wwXiVyTXLE
QyLF45a0IeEujfHFHiSsfmMVl8AMpUpqmDOkvptYvos9sOYkXq3GEGOIX0xM3dHuBkF+tF++Viuk
uzm1LR3j6FixsllFwKXwbFTJR6ENuq2wFBHkk4WHE/o+ha9TWdMBcVHTe73JEBpZQM0afeEJI4kh
gUjR4OfYAXF4naN2iajnZkEnuzhftbrCa0OZNrX+gmQrYGORKVZ/Pu9+0Yp0ep9Vb1hHawwOFeTm
uHOuaMUdfiq6pM8bvoCJfMarxl2VJmDYAth3o+p1FG1WBRuBdqZAXP5auoXPqkFyBHpbSZV8E8Pq
URNzhrdu3ef3ZKgy1JRr3KwY7TNC7gHDZ8e+b8ZJMjLePqY/Q9n/beTSeI9H9ETKhu27ItYzS/q2
/X1roIVS3ICEYhfk9PfD0tZ/lsv31vhP3hIJTQ0bSnWV4gO7d46lIuarAbflHuZDJxXExjpdSsdb
d93xVu7rJKqPLAtwY5I4lHrNG2UHzHY3CzeX8QEPvECgPLExDgiQP8+KV6fRoM/i3k3mQDn+s8Or
SZeVLZVNJ4NYrE8Lj439F9uADy73DW1SE866rNNgYF/g6Nm8D2ajZo9gJOAsvestrZEGC9H89OLu
kj08xzlJ2AGE/UYlBq2yzn21FJjgfgnYyGZsIP4//p3f1Sd7zt+RNto+cX1XZewLrcMjaM2JHYXw
/ZXOrvwTQgfYtOni2LOE5CtbyqRCDS3W5vBOeeHjeTIcPbtGYCFErZmIam275y0JKWkxG86qau6M
6Fv+kRii6PRqiTHv86xVNVRYYdpRUwlu1S9fE6ms5JG2g395lHqWRFfSHHGDu87C64EWVLwkzn6g
nEstHYkqPjTcpIGzG9bEd/VEsJjOC0vvIAztuP62/kJLrNuBlghRlc/wRsROQRjA0G5FrBvL/Sby
hjxRPl8sA53ioIXqhE+PCDFWyOfmH5HqmVW7zbi0K53VNmql/mGrjO6uELwCsQVEIZ5gWH4Iy+4a
NB+cPMgmT7RO/IxfqSAqZi363FfMG0PoTvs5PlwBFHon9u+djJjJbfiR54B3rhU+uMcX3Z9dFFGk
3fOVCD0diIFv0LQie12Un0+Zr+6qFFUzO62t0eVHWvRMjLMVoDr+KOgoMPlNZeo1VusmouDMjXWh
nWAZaWlydIKKbfGiBMtybxEdJxtMA2qiPe3ky+ofC4ef9JW3rvPpA8dD9J0OgShHLV6oCjawypRd
/eHVD/0rjLlVDUha5uJxPuodyKQmTNBJVbQ7N8AB24f3fyrPWzjV6+78yRRScu8Uvj4hHb3uHiox
2uprTQqz6XcoL9T3MKVoVw8gMKe6tFiZjNItFYnITa2XcNA+u5iT0abCUCJC8bX/tg5Mq8GNVyYW
6oemOkQSkagun4z4BqNPC2Nd+J+tmFB+A/GlwC4Or/7hkAUgiLQuXf2UCJxbnAMkKvnkuhLc4O4v
YQuauw+77bSQcFA+q4brxnghRh8JoTk/35RNedukxFTc28DzZA/2DWtWsIJX5xvLbv/jneaPoCzH
8REE7kArljw3McmBvJ6i7iS0ihMvh0BI51ORpYlOI6AxZyCV6mDclHZyA7IPs/QlecWCmFDOqbb0
G581zUHHlUsdqjgcCgZ2WcAdfGjKMPWXXQngDTfwqfL2XrpVya6fRTjbGODK0hRM4+B5LLZyxi7M
EHNprPfhth2u8fwXW/xiKkmEf6khH9Ly0iMiqyL7aGg0KCoalbVjrvqJQvYrSl28PpcDgknfbRhM
mh/lkcbL8K4V8Hsgnx5Hn4oirRFzI4kK+WNneJ9ksCYjAaaz007uavdVP+zFfXkdPU0gxmFHuE3V
13vOzXKpxJMRO+AFF21RuSdVaHhcPFWcfL+zjHEy2sGsGwVgYscDftKWSjmA7yysIJVDvN1UkxGq
2iIu7Hb6rt8O5jrDyXgnSucILTCgOoglabT48X3fDmsQM7IXmCSpNBjfMNRuXYFJGWeKgikIuU1t
2Bwxw3q0oykNTMVFbIpVuqplHvIEofkvmuhdYZ0oeW7VH/0WMpa2B0vxJ67QSJZwon+nEii6jDey
SE9n23K7IaEK/qZIs9tGBM5XzZ1+K5TcWIyh5EujZ9D+fSKlWRGm5tLmWKMCFuaEWrZwuGlVMEr+
cvpTjpg/y3SEELwApst58hSUV/5pkghSIQZePRHhlZ1zEOvClUBqIAZ5jwBRxKewQ6Z5YTP+XtUP
H3/Loj4l8K2GRB02zUICmIA93b0Al0qcdsBtV+Qe/sEQ9cwKjGAi6J9w85mmAnWczdGk9dIHERZH
li16wMVC5SBkfN/78GRePYCcN5WUN5TRNPm5uF6O4EMk+/rAYy8MFmXPHrwhjrUiULOGizKwzlpf
xSXhr7HVR8Luf0CQljosjRaX5qv+3VLR5IW42R6c/jb8Rdq+z+b2DQxR55l25Tr0gFrcB3x6NXRG
orTrSY5im9ZeUfvW0TZI1OYOVLM8UN3jjjyfCScmiUAflzoGG1ATnTX+dLL8MY0AtKzsybFPtsVo
FkpbPkU02Y648Lp9GQqD3nwwZSi0hlDrto1urbhJm20ykXp/Spvf/jx4iV/yWMhvZKxrfCRklS9S
/x8yzvNdGvqRW0D8Ebh85x5hknPQulduP9OlfXfWEbLz6YV/66X3kj8OfENW4GBT7QN8dX38KqNV
2Oyr43+nv/3hj1BZPtBx2F14HSRfjm6XAIt6o6LeNXlqjBHNwESUnrNMJdml/qFbeT/+xZzZ0iCN
A7sOUIC/BqrlspSIGfiG+dXOc/w3LGDkqSXdYk/nQzIqgMkCaK+lnKIaj1aQb1YxarUKdTgAL1vd
8a8qJDVZTtyeuoXc4hZSZOMWoqBTppurV2rI8XPpweuWMQnIouSzEyJ+zst2yO+3CO7SNndvRTME
WFHvd+vCBgErIVZcDPY85pTGSx2qZWcUaaeyrKYg9TGpbWpzvMjx2acSF+tuLBk5d1HGd/3woX6T
zmmXnHw3gcOBb3MgGa7j8WXRgUEuDqEoTcAuwYV640c123Pv/ijnA4vFdUkEvxU8ueAvahbhmDpG
LZHse2LWTMapeZB//6fkPr/ky9XapK7KEZTL0LSg5F3saV6yP9N/GXXPsr9+mrBTJcXiBNE5RPM1
2+EJFvGBxyy54xeHF0ZmNJ6RRCVzQ8XkXqMo5W75TNEnUu2ywHqDGsTGQ28FIZGruV+xjTNaDd/A
C7evqPAroerAd+zS2d6ryvr2z/hMJrvaJr1um7b/O8CkPoV0QlDdiPoIpjT6LD9RT6XujW1TyIJP
IMH7LgIWi5o4FPb86ufJ+d7UbFFElMH6tR8LYjWIuFB5hcScSXY9vrpZM6j70AE4mqrJ7opvUxJb
DCgGzFFD1LUfjQrUD3KEuZ9uYz8BaemE8dvQsKXayIMnz0K+RNlRzOFFQp7LS6rUHCFXf9xtf3DC
rpf/nTovkIhD9TYeCraprSuC2jPND3+t77cCfyQ66qkR8VLI9s+rSodeGSHF1NNLAazt41XnLF2O
BW60hTODcT53Q7l7EGwryy/rZ2bFdbbMsh5NN4z7UGVMsyhh9qYHupDOdNidu6/VWA0cmOtmfyyZ
eGZs6uCWOwRVCx/A/CD8hXxMgZno4VS9vSMLRj1pY8Lpqzo6u2MnGgDsphWLjY+Vg7+UArRrcbNY
X51o7xGGTq4l7gzZKOragYyEIU+kGcPy9OhgYMh6HYrK9kkHzYxEIMTeVG+V0CJF2E/t+vZIeH9O
tTvtiLjK0Pv/9LerLjI9gSPsLY2SIVwGgIahDSTN9xdVIc180P2BUuiL9MDBsQpk2zu1T2zWCfdq
odDPeP+JogWTkQvjiBRht4nJPenjO0tT1iOU9OgO+Cmt60sVOmW8oqDJcCcVAKcbbV+PrjBUbkIp
BQQ+c9GE7po6p42p4uC/Y13LsqI0ip/75Q98VnwAUwjsc/lZv+DFIwW0jyw6zW9upU9pBBHPPRpD
cHxH36+vy8Cc8HW1Tkh6ClBsCOXt5kCRd1s/2CZnGNJuLMiZ8L9HPWoIvon3QJnS5HvNeG4D5Bis
xeB35xpYGISXb6JiVuc4XQd+3Wd3NmcJ7W7bIgxE9JRii+nHQ36f2I40rGc3CXvx5caMQEEvhpTA
ucFL5/Viun6T98IrcRF0t8yausuktnzVNuL1PkIz42bVgiz7TcNKfh3X1WhQdyPphWENX7N5klQY
cncCeVAEzH8VnB1pXjrNc7Mh9aUmtJ1s3++M2l9LUVp7xU5txIFSS3oZiCwaUYMwdwG1EHdHSkWO
1mie5n+GBvTUXhXQVmlLOFRLmdQ481GTs5MXZSzkN4a2O+jZ9IlveQxUauoqUp4Nn099OhKmN5Gq
SwI7HJKI4QGSc7sioDCiQXaAAXhBqDQ+5BYzN6OOgBEEQh0pq8xxmVBdwyPmHCzLRZilu6BmRAxS
dQuxbM4IzVIZ6hTDX2+XUuM8kVtSbM+8VB4kUaHmZGe3Lq0GWCeFM7l5kJGgM+B6Cek2PScC5EfT
2NP87fAz2IarGhCyOhlaTuo6tNYitvKAWJukBG34w/GeXpZTBeA4aNBALckNWqf34OrX1ocdD5Sr
kySdGeUSwhcqZzhiO1ihW0O9JD4Q7NkNrcZH6kdqCFb0hdbKH+kNmfkzrge23NbLF5I/YveDe0PL
AM/PjaMgeCubGqnBCWFuPNgGoKz31nLq6OSczTFLPyNAZoGsTRt9G3yUNyXMxBzWOXn9/jTgWwHe
k2x64ZedNIStYm5x00NTVvw+AdvlBwk38A09eVbEtpykQRbi6+hpVZzHhKRzcg6TANXveWZvb8Nw
gIOnYTQfdEQQ2ZA1l60ir5MCaY2DOBBF24aMOeMvhz7G/Rz1l2ObJQp0CD4vql5ERC48lF3agMPW
N6qCgJ6CrmhjQimhFf9bItQqy5G0f5X0AbaUc8dCn3suLRkK7n+PrgSmzu6W5w7opc1UE/bs/N9J
IKUNdcbeBwG1yiV1mHuWEeanjY9xGYMkMbpo6f+U/jiwd9zp8sYQaaEZEgn60t3fxnLKbJdya+lj
0K2KlGSQIlXu+cdmnrOvvQ6Ub+V/7AzyBdH1mcwoCebIUDfuPP8C/JB1H364MzmJ82yMGYmnRzAR
1CbZEDi11o0HrYuJfkwAPaQiSF2H9d5M1MpwsVd15NnZR5MGo0pxEir0NB1VBrcQFB68CS9j2TZU
VnnymnmqOX0P0UZWbYdDL0nO3QlR5c16tFVEkV4sONQcnjdb4PgrjWksYpiVyzqSdjwfyNZqWchG
vNcHm3tTgGoGPXgIvhmxX1SUJHiuI3B1wuyyHIgLTod+4R5vtCYySz+7Pz7dg1yDtT81sUbdDzKb
+bvLHmTF4BOVhzyKTYjGjE2u1b4E4KMcyIsddcAZPTGQTy1NuJfJIgjmXwqg0V0zn8ersQfeokB+
NdszRSfDBO6c8oAjC3cYvq45XbntdkgN2/KeeFZve/jyDvHC8c301kfAqc9uaOvmMc1tSG8YVnme
4KdL5i3ldB0MDqKYOFZqQ0oyPnJIHbm2By6lxQG2krxBVu7Gnkc1+lo0YAVByZW+dTKSzjtalmc9
K+rVEltsN11XQMryr0P4UMTj9TbxEml+tgFAmaaiHPmSw6Fu/4btT1r92CfxSzYB0qwAOt375xUK
OhRK+z85Y0P7Qs3AlmkeqBYBvR69/jMcVYogCGXCILotIyAgG0ql2oio4zxYr0UfO4VcpU0b1iGQ
kMXUhDdI1QJkX3YjOxxLZSgvAKQ8d3ZQNPNCBHK1a0H05HEJ+Wj7XglmCzdOsqALvhXgRiDg78ng
glkgwql5acrFpgHbB2yrdBwPjSQ3WH/jDR++cmWCMaGckkQx7ff35To4Th3F0OwgTWRj10mdr/L+
xkCjvWDVwtZRDatTeC+zAvHa5awEOFua66gY+BTeRgWzKD44357whV354CHpvIBDcS3N+5+0atLF
179ioKLEAtaHLgaWvHlo0lNbFfYj9nKCLBBbfL3tSmPRZ5sWOjJYrA3jPhlcR2ptk17eBPdDh4Ty
3VguGkPIH4WUyHUxU/7w8G7G8MkOBjHp25Z9ntC8QxfoZX6DqssfB256hdGPn7VHoh9YMoKeeeBt
NhicImh1YaLC/q8kWCMFB2USr2pxbSdAu9w9ssTCsNgOIrYeVGgBNOmyK7/b0383VTARTNGSAxwZ
uhkMOmKL+YhpOyk1r/7N0i+U3QAiNuDA6Q51chSsB3XxS++dQ+oPW9yN6D8q4N9drlTzjUGPcrUY
cTdFSC9+0sL5Gh4uV7Ud19aoZ4OmcJUudTxIybJuMwmmtUf5PfYB/MapOxAyVALs0v6apLmYEMk8
mGtDYlLq255+1y1qg9kZyvGQSpZ7Jc/+9iv19ippcyPkmcSxJ1H0SUtRUrfwhHYh84z5kzD747gm
WeIy/ecgux9Oj8adtGApcjahC4tnK5H0tJeEtr8Aa11NPgAAbdwefTWddEa/fLeqT0zePIPMCxSO
aqYYrKonuyhkMMbtjG1nACMEuhnPA+DjhFv1Aq7mqW6g4SueQ5S65tnWjqa1AVMtV/f2gaT3UGeW
ZR5onhelLPpfywWAO/A8S+90asgIplSgWNFyKfAlpbelRqobnfZ1frzhGZtVpabddOO70vUzkSY8
uIxX4wHS2PxTyiS1AHXlLRrtOdt/ZpsziHz2ARGkBpad6o+ZGgUGD8OC3Lg2jihV+LeKf7bU65De
vGU7MY+CdBKAmstJTifhtET/wdj28m/Yw9DkPBoGaZS+7AXD+mQeVZQU2t1GX3FkxCDLsargsNr9
8CrGauUyt2O8AFO8hB4dslozVz/Q/cvupohOL1VhEjX1/0HMjf7FUlkEgILj8saE3QdvJMmd/DdY
MMbuNqySs+EqWfippl3CI9dPv8bL1dADauBMpswMSeQKpFz6QXOt8knYR5wUR8kbU5pk7/nDium7
6XqbqkBf5YQgKVx5eO2IBWZhjvlE8I15XNVyVtxRJEB+klel24VepG7uhDGbrP0BPuLqZopA3sVp
Ftc3t+cNMFm4mKV1QDviJbOcTBmolo2akbf49yRWE9a5ROoUUwji4iqM6S2nfWAw8BvFb0oyS0RX
UA0JXeqp6HOyxz6rWffRYi9Kkdx0rGhAUSInYl086D4Y6h9rkxpZ2/4lazhjmqcEPH/mobAOsbOG
Q8I3aPAGK0tCzhT0NmvcvSTvVsGosuiiDSjJx2HV6+kVIhQ11m2+IsGF/KfxlZyhR+El9LW16FYk
H0tojhbdYgsBnFeVJfg33vsi/H3C8tDveGYumV4rrDRh2WZPKtLqJiVICuKulU1GXnYqt3B8ysNH
hWztJQJ1b5cZWUrTIIAlc17/r0W+pEBaU2zE5TN2oUFg3bFhOrO64pTE9e2OW7cn5zQeN94rFBxO
COBk42WYb5uXHuYGfHiKJ2fgG56l321yQtaHzpJnKBcv/rcsXHWjSXiMlGv4kfo4hzxfrTbD9cgJ
DTCfRa0OLWKsLC4GEUboW27KoxgEAvw3sQYLtsrR+ibDtUvRK7qqibnrUv7UaLwxQBPqYZO2iABp
NL6uD9As1gMLcrHp4DtYillKqMOsQA6F9ot+PWrzYqZ6kQId4+FOHRYdvWV9ZUBYsRiuBp/axzVH
hyLijqbpatvwHRVVGJHIMTunLQSARYR5+6X/A165O/YbEx5mmU3gb6Bu0MEgSRoJFjzGh2D9L/9C
lPTUoe0OfvU1KRZndTafFvL2+PFgdL9qHdHPQuQPXgkRsYsoAjtN7lqubiDvttioO2bbUXqrGPJa
TNOucegsvx3nkO8Qe+WpvZuIwV0V5ic+SwYJjJ7ABmAynJoXtlWRyUtyvHwQbhczfCw3QlEmfiND
gIxI5e1THru8JXXtLJ746Iyu69vyAT7oBuW5VPIxKSmjRLoS+tfICeQHy5xDLCsUqMzplJPuLPl1
lYlyRcDJ+3BvQtBD/0tx7qEuMRqdqSoAM4cWX5uEqDt8K75Qfn6YvLjTPGhsowVufLLhEJJ6Vk1F
RulAM0vV1WW2dmBmWgLen2rJxQnGx6RIeC/12TBzgpqNzI9iVNbAPszL7ceCdVEvPVD/6yCRtZ/8
nz4P0PPMVSw9iJLTvZIcu3Y3xfC35sO3TlIVbKwm2JialSkO7L/nwM1kj0DFOQ8B8nrblciMyGTw
pGnzRn1vuS7qmyCH5NJPSf9tToUdrFH786i4EnyeQ67voC+B4z/PAxeUMZO4RDRstdeJIgyx6H7Y
fHrTYyOsKrjm99ZU3uTcXGSca76blRLcgS8ZDX69hcxTP3jU4siG/oo4S1HT7PiflyaLPdk5mzAC
oEnSe2tjccwi5I7dLq9ugyPK4dlKbnzKEK+pHH/xo1TvNWu+yF9Hd95/A51tLbummAmOQxs1dz+A
NquU+5NTYhbA4V5FCmylxDaAPswRgTkw6JbFbBmBR1CNiXGDs1FsYyZabZQAY7IsgHImfFixnXUf
Wt2vuWf7IcoDgPcuNpx/L0hRRrCmLJXgLFwrlHKTkQmpCuG4bv85KPfQB0uEVAWauGmCW3aKJyej
zIrbVH9M1IvMce6c6TIyau4R6i9r6nRUL7WU6+jXeGLs76cFVGaD5lX4mu524/X81kQIUZPEozt8
/bg9sP4Xn+1Yuv7Ttz/BCvSC4s9Q8zg/hnTQ5DkVihy3lM2lki3fjb/M65Z9KqhjZS9Zt0Ia1iJP
yc2bOzSm5BPzs/NXv4MaUaX15AHz36HaOVfQPt78ll79wfRcTifIvfXLNNiSO0AzGkt5DI79aRiL
6ty6klOVdMqgDJMoB5xQLE77EqJZ7iBuqMi2E+JSC77KB9aVu1nCszTmgvPpyK82l7Qpo5n+vais
PTJG4AtScZz4Tp6wt+9l0/4B6bofC2IZKMUc+q/sPKVN5L7NNU31GEchOqgOQ9ahILg7FE9e7WT/
p/6zWpUEZ8mEL01oOBEHCwZuZcDuDbbm4IL6lCT0JYBtIiYHoCOoiPCe1QwgHIT0qu5efjvD37Y1
KWKVGOZEEpnurv0ytJ3S/XYasXXeZ06V1S1MC5C/7v68bst7wEeFVYfclwDmU4AtS/hJpW/IVgPV
Bi9a48Z39y4PaV2eC4wGLNDz0ZJUeFC8ERifHGC2Keay+x7OrtorvturRCiyWFWipIwxl7anXjlS
rzidTmJnhcJtD8zSnfrmD1PD+loMp9FEZOSbNt/zyjYUJ88gprCTIFE0ihuszQRcti8UAA+WtrNU
cu2sY0mRcU2QA3BlNpjF61HEtk3zkebqpIC3IDGNXKPROfP5v7D8rrIzeAp4mMtUNgt1Kg7EGsGC
UdjgGPZdtHZWu5qv7ixgySqrsBz4JRRp42z7kfKaPIbcKbIXX/rKaYJ3GGuXqADLUnMek5driFVR
gE6rlhdg0o6B6vzGnJdjuHNeRp0fvhuyf3aMM+tMlNCNXcKFOLGk36o7ep6XocufBxlZFk8ADjje
yrKBkFXuWfC58mWDYwbH8ovuYX//tE68+InajuQ3etdoCu3VOyUQTp7IQaetK2B6ndWIa5uGqg1/
bSLrZFJFWJzFVg3HRcGXVtTAV7TmsDcbHoYPQMTvHW5qCek60jIJdyfoc38ZZY3/amsE2X3aFqxW
NRtPAKWnHJigMY6ttnj2eC+2lW/lPuu8xuh04DHFU2ev2o90sLuvM2TKbVxFSeGN4mzMcINQGZoS
dUEDjANpf8nNRKi9Q55q9gNNNfzAotWs2Q4tFp9SnfDcOut/mmUpxGhx2KVMG2JKTGujE1XjfJLC
TtIlKvdzaie+4SZAVdLsFgXhrclmWggWnMNRR0VYr9b7W8W79NcNS4gKUqk1b6eoAfkxMcBJKeYa
qh98omlhQKr+p2DWcMsCAat6UxS61D6DDkT/T+OOIHwLE75f1goVvxyhZHsXtN5RauNq55Ej2iov
YRQ2RiyEt8uY2C3sHikfT5IG+9URsfM81abQfkdcDZpApVzOzOownvYjHxNQliLL+aCAuwwKIBFF
PAiQgbj4OxY8infOCPPO3pzJL8zVR/KeYxqEeTO654pCrywRH+EzYVqyStqBZ0+uKLg9zk6/z1hQ
RLBliUV6PUhNtS+nWTze9pfqrjNs9mLg65oh2iteEi2LA6DJBz4vh6ar1P0VOUzbNWHPsS6Rd8sV
GYk7x+liZkV7jONQdFf8UYdKzicq8okACyRVg5g9mzyBtLjX4fZmPqI+Hx6GXb0IIwvoh06mbfOy
Y8j8KVMMPcp1GnXW6M7ts19ExgITyCG6T3BtIHi0xkEPfnC15GJF3dET9QcEssC5QDp+U1pRe0yl
tFoZczgslEKQ9laQQ8ZIjAgvWBK44ySWjuIUW6Gmv/TuBayE9jVLWPPvSYVs6jp3mc6cDuPS22jp
JmjZpg3eSW1Vdt8ylP8ipE5Jh0Tc0lN7Mp+q9pXfL2uhXetV4WoYQqCy9pTD5UHIUfX09JuxYqIW
7K9xpBKoceikveDGQ10+VVDOy8g0hGoecojHPHORlMuOkVikJUULc58jARsU/iXrA0un8t6sHAl8
j8UxsguTBsVrOQU1bl1WwGz+8ycu5CmZo9YMu/oIWgQbgZnFARx3JtEoY6BbcfdEvpF8khdzdO5l
a2X95P0p9jJOFf3Npvbbj2F/DG96VeO7ez23oG1EO+cpoUKL0syCZG2Zz29+7lhlLC7kSVtQE7w9
JN4nOcFnd5RBrMBHy0hLSgrJ4989oiFYIhtkM79Y1phWBfrLTmuYT0C0xFjFI/VQER8dM3/GQ+OV
FAjV6swPmN/LDV0jDCQ2OD1F1nes8MN4Jg2K3iM1OKKcv5gv5+BMDEh44FVT5tNKEEuglljDYCC7
3GhK2daT1ywePD1p31eoj7w59+ASPAHtsnLmZCAWw4NuE9FrpaSrDMxQc/FUrTnnRqQzO4F/Vvjb
Jeziav1RrA0VQnbiKPN1PLlFia3BePhlKu5yflHFGRj39b+Hor8aKMSSE3hJ4ZBbka9ngQMGYmLq
GW2mDVv/jH9g5y0zb8EiAoKz5q3h4epUQFS6C9jweyjCwDtJ8Grt95fPJQeBFZiiG9UGQCHN63PD
yfC4WeuzWfpaCh13sGwswMnyJkUW50SV/IUvXuevNNyekw8+uguNCdpaHcqK/5zAdgRPZRB4oxvO
CnonZXqjTymLmQDhyMyFx6dZ+VHaqSlOz4tq0eqaxGx2ALESTvDfSw2NOGQLqAi5snyH8UlDD2gd
iMdwA+LywDpN+Mvugl8GfIYu82jCI4YWo1G8fFscjRdFxG3CSoOxyW+WKpuKu+5tIpPCV1zfqUKC
FI5q8XEloG4M5wPohz6z1v1wUHGgTMnNhY5CxmD+2CIPDeAEEvbe4MryiRZU+IOIK2XH1AEVZjzW
1QRL0iRYebzkUzC+RlhumPmaEdIUZIpjnJkQakYOMFrTR/4GQhB4wR2hhg/UaUwF4PQ/xCDjzvDa
sg500rY4Pa3hW0f+hb4g65fv6FQzZKTVt9eDHFdBzzKC4IBDpwGrpRWSWoJ8hnqTsgIHxV2QmNBt
LemzWLocI1Zql1bJJuJbL1XkP0USYGNabO7AyKVbWBe9YGsFzUXAhyG/NDBHpmINx3ewiv6dFTsK
XtkWvABF9/86zB11973XNOubwg0/jmgYfIHUjDXZcKBTdHHsa9+aVNcl6rLyZcXtSUwVl70DAqUY
I5iOlauAxK662Kfh1UmrJL559rWR6YFIJnyILES1PDKfK7ps5oz2FI2dUUieHoP/PFRlH5UjnjPn
fGdMmJqf42JdiukJSSv2HpBgKC+x5JA+Jj1Emq9AVrsiYiw6PFAsmBgfUs5vU5nR7NBXVIXasX3/
FF9Eqvfg3YL++CNh6ZSrZwemLh0ZGtFCJvMw3k0UJzRHdRRe+Rlfvp3JSz/KmPuPbvTCl80dhK7t
w3DDxJlj+fn3LYZt54sHlz8wzGYbIA0FQS9X2u6OySP9y376Bfa8DXlolbLd8+132xntyJ4hqQCV
/XPdhGPEpNDDxBrYhDJCX/52l5pramTPvjNOn9+Qu2Kd+n80vFgreQWbE6Kdg/CcweJXKGDs7Zlt
IwA+0LulaAmr+NmA+NdwTVwMw1XLEC12BcM92ewoNRQvnnkDHv+refzVo4zJReZdtnZ3AMa2EhYh
0rqpKb066TTSTuAJIf0BE6GAwqFe4rB06A5oq3SsDsdePD2w+ISLoUhqhH1ct5TLMbNJRGtSu/Mw
LB8blBUj0lCIzobSQlA8nDbOrnE5prQmG6S9smRiVOPjGGskW/7TyMdFgNUTBqUUP+v8aEMj/+va
QoLw8qAG2jvN+wCjY3E9jZwW1D3xGXjNJJFJBKtgve0cQFSmHuxqR76vnLsUkKTzvUfZRSGxS+Tt
Uci/bLA0TE6xyFs4PuhfXDffdSytJGCbSOMQciIMAB4u+zA84vZRrNcJ+y4IL5APM70G7F5ahfrG
DIFJeMvaO6qLjSESXyhJ/QDqFW1Uj8XZCEIXP7p+9XlrHlxgtvjoEEDdf2Mb8dILUA21RGzvFpUY
iSu18ZufFd+PK+/G59eSPL507wrH27Y/EaZP12EGV6kEoj14coYcl5huRhvFObhIplexJRXxMLhn
+AEMNcFgjsr56n5rtROUAtNmXgHvIMAUerZcP92IiNfiLmuJN5dHbInHZwJ/mMPgNwgWsDD4V5Gw
GqzaWc9wcy508//wdkCZlrk4MIUKvmqZ6hYkpO1lA9VCZsId+Su1pnrpUbbW5SFyNpFuZa17Lj8w
Ua039m5dPC4sL7KPUFXUIhv7+oGXLFRZWmkBfJ+PP6X3KXa0BZ6rv4w+dKIFIts+1XG6ljSEnB5A
OITb675mT8xoIMu30EVjHKyKRkIFhLYm6Cno4+mSnfXaRI7mooztG7kSMEIeb5zuwl2xtWytzXoG
7HbVRJVoSl4jOyCDwaR7n8vDQa04M04wv7+RxfJpK0DvssJOnvtIUF3p/NyoGcvkZRs0+KyiZ0Ma
aC8LypSeFwiz3D4uXuO+IJfX223o49L4aKyso1b4Og8MDtw9ga/7MFcrY88RrYPsGBT5JKI6zkAa
XSYr/sY7MlA1CYI20ECb9LtNJsxHCm2e+ZF87WDa6SKbULZSbE6JGgOaMIID3TSCbgkL5m9w/ycI
EyGsZsX3XZjB70UqvXcvVXt9hOEwBHodBFJJSEUHXbnF7JlQ15pN7WeZH8Fm67kN9HQImvPTKVyl
h4IjWUCvLZuxswIByFRmcPvp9DOIpyi0hdhFI/4niUSUhmJOoZoO7SH+EotqPgJpWWTgN4w9//NN
MQNPyMGPDuBFTx/82LyW3aRIEkeZadHnnN9fwPFzck6wmDgOK+zvNMURt66bRekLMIGHI3mbuV8H
nC5Rrrdss3/GlgMhiTL7o0hXBmVUBTl+F17mEi6lompCLcpHc+qIyQN9MCVm+3u7LloV5Le2Gkjj
x6aJ32AS14UIY503KfBoqkxi8GeQtP1s+szXhniKFP+ZNI4c6CI2s2KkKH8bWKHNZChPiE/7Fgfs
Y6jTsSQOVpHmanjtPMCEJcNv4rJLOwztebPsnSE9XpM/i7Fn6arB9H0rm/YGwSsizN+BPyhwbweD
SvSYZtYSg+efDWXaFkTdZkTNUCEziDFNUTD13KFAvqCY3fqZDqlDYSIIzr/oYp69LZ8EcLqhomRQ
0Hen+aCmofpPkCIf8qXyFSa4g7xLc42IUdwkvbdLgo2Pw4AY9bQxRtpQnyfCi7JHYtgZABwaNG80
u3GMMy5fDIoAp5qAu+rrOQAHZKVjBLliSMD0aLwqLM66coWRnb17ki9VSZ7gqWo+aIcGn95pfXED
eQHP8G9taxPebrzWsR6NaEqtzFOuTgm18Y7+bP0ymdmzZ08v8B9gx0+L/KAkhyDNJCLqtIRn28u9
gJrwIUs0IOtWelMbYQ08rh2ElPXueCf4j7hmgZ5q0YoXHIx3rqAt69CZKflMzC0vi1Yw7EHJaFbg
drCX3yABTTpTnv6UTNbxdf8Bu8YMsiMdfoLVjzuSaNxva1SMX6MjbuCUHcwe/QJ4JHgbiok2EP4D
oCiiRN7QbyTCMPuDSYmqEKfWw+/fcUKF93m1EjObuwK7uGcYPyraGsetYP0AOD8s5T9QfCvUdqM2
90+5NRJ60e0i2+jrqPpWamWXsbo+hemazlKUQNVGmF6yVa9is5NPB/jzDe/m0RKQvUzozbfWhvL2
Vw3F46YGp/CZPi+1qTE59pXtZllaCxJHydO34q2B17VknPKod31gLbUmy9JrowFMby6G0ZFI74mB
cHeqR0V/Wyj29+4fFhCKQy1KMk/yQtTYB37BpS7QTgfxbRCtaqPMTPTvxmr6nRkdqHlalY2mEo9A
WDDkTMYZhwVi3j8OfuBPc7SGoKBEuYR06NReZLilVpwoOw+MhNbznGWSNSsqxuWGreL4k4kWy5oL
FahzPytOCqE7jnJJ1gKSy3DBsY9sMYqhyKd4AqwLzkng1a/JW9jNP2VHV0oaF9jRYGQWR1sualkW
Xo0K4096lOzcTHoeCXM5qbtNAMtXOvRGwUUGBI8m4im5Kuv8/LcEx9lzwp1XC6Weh1z5JZ3ywTK9
HrhuWqo09uvs2WHxsiB5ls1VNqDpRWlBGIJC9/VcvaobrmLR1W3dfEOEaFQ9g2ls4DE1PANomSpi
8O/UNMMgC7Es1OcoPK5m5S6k+mv8R8TX7LCloI9WGtYNDT9pwC6sJWp7Wh7lT711uEsg1mN+VZfj
XfVM5gyS62hDxUotLUHYpoH+5s1X266ACJ+Mq+JwfgAoQ1ReCBFuiKfJboAqgxxF/qHAZS4kLpXK
VelYoFTh7nB+xhXBYrdTArerrhL6vzosc74haEDDOVS2H9gKVcQg+m5tv+DDd6lYZiGEGLiLh+0a
PhObXxqz2885MsJFhYWvILPrIGE16JbHTZ8T6n855vMvnU0bmI6rBd4D2n2Sw1sKSGq+yK6FuHRS
6TMc2uRpDPZc4ji/Ur6bT5hsH/Obgb1K6kZYfC6Qvt+TVzEYt5mliftAzsuGr83CIYvcYIoca5BE
dq+t0QjE232MBC/KuZxUUG6QONHpEYRS1MNozSs0JTiNv4a+f3yBUQn6HeglrjXfaaMGR8n1LAdc
awPghsY60vudlPKtPXWwvywlqfKQJDltlhnSL4mnhU1dTVcMgc+ATTNAf+NQ4y8/926hP7ilao6I
2b2CUOdSnQpX0tV62EL3yUuciyVNiN7S29qIc1wt/vs1vS1HqmlrimdKV/Lw1lgebwmarSi+6M5N
4ZVStVyhxKMxQYSkWN9hk91un6cMY2gOWowSJIJpdcAcfMqFgtsDbGoLCuvqS9MjhpdMA6HX0KEY
+GhhPfYWcNlxsCjLvhjHKg5iJDd4dzUpk+I7iEG8SXNU6rvlf+MjK6qH6i/whuFuAqvxcUElD7Lz
4yF1xVqXLnGsxNkcZoJc5176WHGUk90phyz2ta9ffl3x3hNeNBv2XDlDUnaU7VABh74rchUm2Eit
8Afa2osmFtbd39ARM8bnyOaElwQU+07Vp7fgqCOITMbeweI92W4gffqeyvkHE/dWMljutUA1k3F5
OX4yTbd9xsZH9kVkC+TQcf+fagbPJYyt0rSMSYhckti0Ycif/1h5DqIqoJ+UJrVhuLLCIzc5Q4nJ
pvBn61PiVcCU4ck0dEMlwkFhE0IbVS/XCt5KLrrvI32mEHko3IR3XVqloC2bRaxDvUHz2Yv+gI8d
4xeCh9NWwN50c/zcAUHO8uDUp+f2Ai/CfrF82XjD/KH+uoM0XWQZX3Spixqt1oMcsvJq5c7R7Jyy
xnVcv+wafFj+vfVi3dp3qig4zPrb2Shsw9RPiupC6b5e0o7sY1TTiupFQV/U671pFMaiudbY+5C/
CMrtkd0pxBLlK5r5Kk7ElWUhyZm5kQDAFJN/ElROwWmFqCPQkXthhMofsty9YcjjemzdchxKhSdS
UeI5hFCao6v0F1hD+yHMj9EhZAZXnKjQ2rqxOcTV5Fat0umLdq528fNhYk7lHHAWbH1hBBnaDA1A
P7rIh2lvPZl/NTRj5dUvs+YNp13exmOZh/bCFVeQ4ePxAOFeeDEgBfU7aD34DzLe0L4F5rkoKoqL
Jb81mRdLXoLq+s7EbeIjP2BT9KyfCDrPJL2njL4yEShNWIhRRlk5kOR8UB64sPT6DEruga2SAADv
0V4iPr8GxiVQs19gDeu+p1VRx4s18tHbOhaq24mTMUChCOvV917t+0J/7AUo9na1Cfi6Vzu2dMG7
K1ZgbCZi6Xgbvs/L0elNZGESoUozQeL12+eicxCAIqh09NsgUQH5Yn/fyj1fGLQIlMluPDqgIkG/
eIuC3FOdU+LdElUYLq6VmVGSv/QWMiahw4hfu071pzrkS2gT/AcWRwBXK64kErW38dWUJAMNnWrg
Yfcf610uN1LD24iI8IJOa2YOD7eXyIBGWCPIAi3xYTsA912ZvCRqiLAMyhE5h9SDibF+xTaGkqlO
hnVDAhEoUZlF1N8+uAx28Mb3d4wkO0FDG/t7hBeWBmmd2CBp9rsgVPDBKLq9SbIxbZU4pEJ0Y8Hx
GcjjdQyw2KvM2TWAcCtUSUkqEsLFlUlgh6SHa/BxGEfBFnyvQZX8T+gK1Tk83B47vS77PlmvJXNh
dcJYHpE+f0LYf8pI9FrudPHzIN6K4MpDAoFw8Le+riI3t34hPhBWdKl3iDWwry/gaoDBcJjmbiN6
QuQhBPVKOpqj6JBh5w2RuksYYClhj7wEMTMCYfkBisrXmz6acyvZyoC0mJ2Vdbp8Uy/Z9AGgKHXB
QAxnQaxXrTwa7ulzEmvXiRUg0LB0IO6R0BhEbtxoyPEFH3z/UVYxVJnwOAn+MF/+9rYX34nKcv6Q
4iSpsA4hqsFKOt40brNhwYGpHon6gm40DMulBeHsfkBqHtvZH9KC6f36BjYwi+ZIQWv3dAITm9D4
/pQP17nPY/B03iTkYH58H19bfJXvnJCPoASGyESAANbLDxYu8E6OWpvbQ8N4pLinoDykV2YUIVjF
SArUq3SsNIkvhcEbkiUtUOl3RICbZIgUb8p4ef0gN9MqOR+j8i7E7vkklSg+alilBst3SplKzelm
ms+WbzoR8P/f0cIH3IPMUOiDhRbMbeeZzcsapHdcfklQJqT/2g8KJ7FHgh0XgRT3YtCwLH5OciVm
UqtmA5IILAqbwrHzV4+uBPH7HdMRYrZkSj2tqXvdxSEJ0C6JfseH5EvoOSLEyxurmydyvg0FVbRW
FHHD3PPChfcbuK9k521rhAAYe80WhjZCOMVzA8uJLczvKWewHIpoUVleQIDfWWFx2TSOHPpUB9p6
AA/luniZvxREP8UAoX924rm4VzipIPqRbWzUTfBIo7PAFsg37YN4wvqRIIuOFs0PizU2DE3jUrBJ
T8TWvY5DjQZz5T8H9PKRaBZ0NttUn1rZlWZfmI7CNvd+qn88mlY6i3dLklfjMhGXHQ671Iz0HCTY
9Wf8cLV7iQRtVgaUIgRPlqmL75PagB+rH39FeN0WZ3uUx57xHvXW6DhepdhyaXbVAxrSBFLh2aCv
l+Xaknspvb/afl8AJ8Ejz2D+BUQshriDimqD+Fllap3bGiLT+5OBewVtxWnrWdEPSkfeXL/lmujo
0i9pZOFCS6B3Hl0AwO+TNwqNz2aku2JwbjsJFScvZu3VeGQrdK2vqLPVN0sKQOnmI6Vd8RHnZ1cE
NhFktuTbY1sRtpPxauFJkEFnnO0IAtJ7rDeyyyQpAY39BIEOFNQwCjzplCD6paNO0FHZ7zGBkr74
BcjtIPgoZWzjMuOZuxO9vM822gSB4u4vrPX20FcDUWhlYBKWCiU67LJJsQDWoN9j+Ne2tw8jRW7r
Hkhvu+OWlZtz+WOBfG6dBifoUwErLXXjnfiAXhNE+U/Z6XBzMQNR7OLZ1sWQ2EUMe3CAGYSlYxYk
HRST/Ul8BPivi3EneLIAjEHlEDlGFWP2dMR9BEAwkhd4Ew0yMareL8eO8ewWb8jQyv90oFBeFexI
YKw6fXq91AtKzETZsGtDYBT75oirje9oC+gMZy7UndU5fU1b9OJKQSj9Jm3y/f+eb50VglyCZw4o
m+XgP9+S2qQKchx7MiWYeOIcjIKWmZX843ahf8L5AZ+81oT7HvxCxSUwSv9GVcGPNol7uvRYoxzI
unEWG8t/go6cfs5DLQqDxmLOux2Ii3hjOv4Jp4G3YS5aHj+5QdMdEpQwzdUgEzBAsQ4oAGdHVG6b
jVqEHYcWhsGgZvkbs+QAXz5cE8jLpurjbXRHyJptnMKSZOsAoMbr7lHmCYcCMDCp5+ZTHK1s10wo
c5ahU2jjtqN8kkcPzdYHSEDWvn7oNv6RXgEE5SjuAZpjn7P3FAd5RvZw6CZUfHF+eu4YqGTpa8a3
DubIo9RpWDT2OzmJ5qhepRVk8Z4i3TLUrE7i46hzLHIbi64XySiUf446K5oej/y4SuGVWRRe//qs
/S4wwzdN0wsLBDRGjxWiMHkvjetWbfWXS/3gXLx/VMcwAJGXE98Pnw0yrhOS/OyzvIZUm0b9iitJ
3SWN+7cQRvlL4R0zSGbP5+P3DN55Z1vtyPSPIHPrm4vkjT1mzlXcWh/oaExPZCHyf/VCKZfBIUiI
AOQ+khFlQrDCBc28qmoSufFGNKMpH0GVDP4Q6FPI4bUa0dxGdr22O+LPSmFhyZmq1Ym5yHZn4Bdl
MW50v3OTwUj3npS5DLHORxX/eNqiBrFJnLCU0LXmkcRP0RCgwE9I544kTl21N9ujw2fHaqT31lJJ
hDJaH56O0rHTq5zVc99sut4gWnjnkPLeC2G32Q4stLI54hDm5TWhAxefCtQnIfsdOzBq/7SdVNSx
bFSHCwmfkWjx3Two8rdIzxsQAFCPtlou6k7AocnGYPs8n2Ss4hmWlwZqAp+BN9pqaor4G5lAlGa8
qApcUtOKfxzXqKKKfzCnAI/fVu49VCpwGfcj9KNmbq6nKVhE4f8HFnpuSlSfbkd2Z/+SpbRxcGsm
ERXNFnBIXO6KbWNtKtzdoVnrs9MBwC8TBOexwFYKG71JSWCquvDOioEec0cfGbTqcjMhA2ycZuVw
2aKI14//CS9iIv+uptV3ytyfXY83JJTUSaLjmGfE6B5aHtElkfGRjTYse9eV3I+mp/5U/6l5AC9l
5lchCiee3uVtlSgHW7dkadWisCFLXfUTMUDe2MBdpzG2Wlr4ezK+gq/U30U7Unb2tgiQCmOCRXv7
eNeiS5Z9QZkpJ8+0db6iOCCqZLarCuw0v/+cAPZG2Dz0AkOOgu1xq7/j5D0JuQXOH9DBDTO5VTtw
OSR9253+TunDLqDuk9W0gLjEZzppk3Rm66eddHPIng0E03keIqEFWEDuk+vEJTPD1CLQNO3oU4vy
t8amqQwfkQJi2kt85VxquQHkFvR2Llv4Uu3EgfWMrBy8VuN/8gJyczNkpr+BCbyJcsaou7MS6fpL
/ZHU8Kb4TpYFGz40TkLmfVG+OIY9578pjMznOEV1TOPVQEtVffI0dnC0C2MfxrUA1tDE9Xhcenqu
wQ6hBAOeBDwvi1gHB9QZJ6wUQAShLJjhHqpOJCo+0AjeOv11+dOxk0df8TN/FtucKxeHfjYVAPux
J+kDx4ljLmZKI4rbriuhxg8RwPTMWJjBPa7uiXAGaCBkVHvX+lSQGOWbX8+jcB+i3hN4O2RUGGfs
XukBrpUN1lK/DEpfUeUT0Sz6VkwRDvsdNoQ3Q2xaAjJpl5GJ2RnO2zRXmQyHUmwBCKn28nfs7C4N
Cg2794AiHgMjFHp+KJ7VnDFdFEat+XNR5AaqIFADPwtH9PfZA6k7b1vx5Gt+23u3Ge4qbp8zfRQv
FJZLLCFXLntlh3YD+1uJ6kz8Tf8HqQqx1svy5IJc6FMaSSf8gvuHoweC/xx+MaK3wlWYLcvvnuKV
lic4zGt+pJBCrUWtfJQ0yPcZbaPDvPnsrTPXV+r6tTYsTWranI/bkCxaYPY/QcaCi1w+1eMJb6wv
HAVyLQvooLpYRYtU/c9aJWQrQLPUkSOfcANbgkqwwW1Be0UkHhvu2IBXJn3sI+pGKutwXTwp2TqC
RpQOtgigTNHCZIcObfGjCCteXxrmQpWnISwUmE1RrzcZvNUXwc8AdP1oxNFnQkXp0KADlyLXRngA
O/zcxVoJ0Z8tA+JkbmNZmdDy+k+3xerZqNqhRRRs6P7U3HTytA8jaLAptXC9KuSUVheF+WTetitD
WDPxZYvHiPiynLJUaW+zq/IUxadh2Wrn5DHKCRTmHCBw3th47yT8eS68GDp6qBflBPwZloz7g4uC
+hn3qt76sJmpF16wNJEbr1N57Fbm87JVoui1h6yCIYrWJCHV5UI0mQvljNj6EE6joM1jk9yWBFU+
t8HVmB03Gk4gAVJuZMeaTnfCvAkrdCKGIRmUkPwgE8gNAP+D9TrbenQbIgmJZi5ofZOe2OkZj6DT
e52heMvwVs05kgSYmbO933nUl5iafLe/m8xhgW8hCjYEmVlsD0G8XtNG9siFVKsIbOqWteMefm57
6pnOGTSvxqgwofz7Juvxf3GpE6KAUc3wmRVgbUK14CyRiki6btPebst+XDyz/uiBZ1r933Y0vmuw
okNjyfab3/qM4IpxnG1QowvllRHIDciVuDlHWZk8uKHpMgtIrtiWXhERIVHYbbZCVNJD6UybmW/z
6zTjfCo2n9pTDW8iD42aWnwUpmV25hLl4jJrBr6hx4DgiEktihMi8f7fpFVHZVdlRPF2oAka8Tgw
igMNonchruQBOqT5PEDAOEztRBvxKwQVKpbi5WRgBuDFbmXZNymyOCeSW4/FjcpsmEpzeUe3jHiq
nng7uXvETCIhzQLkWMjEDTyjsMUPfjQr4E6a4CDG1sKI8e64ZkDT3CXvoMd7ncLr1bkhuBLUFkIc
ZZoBnuN1YbNgjUsXZwzGNkTbq9CvHNpOan3oVQK2KVNQqVCsemat71zgWeFxO9uniTt/+xBOGKzP
a4ufe6+RMqSsH85Bv7tdTTb5KOg7oBJoUAOKraLoYkByiaT9tMWoVPXygxImmoW2U7OQRwXGryuT
8IzLsTdre/cbnhaFWEfPPbCcBmisYFt4ZZKfCvxyPszL01rTt/6ULbLZEG/GIFRTK+En6zlXXEGC
jWeD6ylYuGjuzxyuMx2Z8Ij0ummqKKVwG/2lb0PfohaIOxzHeGomxOeyl7DQOqDnkllU5tHZXaEj
+5jmpC437hGvml9gKVoQCRs3RioEB9Pwxt5coLNALKyhgV+j4Mt3avJKYowXFXyeSerIVKq/DYs+
F+664JP/o+13mrqjJMVf0gMV1pvuXaN8O3mVUN7IAjIxud9CwlcoExfL+YifM4zkXUb+/FD6Ni1N
bbFEg7HDRegZyX1qe2WulN+ngf+HLHxlUmYMtmy3vrpT2mfV+9N3lm7tSqZsXLrktNrpTxoukBci
jDoJdDmoG83XUvODPUjXMrE/BopkZvYVZs152dz2YZ1m6+3bVpdLxAlFA8tTHNwHqycmudfsIpvB
31ydXmEt/xHs6o0UGkkEFNiXpmKQHWqoh4nlhgqceNBxLUE2zzK3vkCiQBnteWywd/XzX5AqnTYy
pZUAqQGMMqXKpCNLIudva/yoxE7b/GWc0TYbC7+6Tw5kOz/i94SV4Bjn+LhT2lxmZ/ckjvp72lFh
d/7IM/XYBT2Vj5Hjm+QVZ4jNukR0Fl5r3Bjj6Hx0CdSy8XgDogRrXruB1CF1/zewFU7qDoct+dpx
zJucE3WRrEdhB6OuFENCRAK+Z86jGsXbRxYXWOpoY8PhuU3hoi8TM7B10EVq8fuRpvoaqeUVy5+3
WLoRvPpoJAXGbDYyQqgihjZFkJ3cTG6N17XQ6N5emkX4dqHM2lGU4iltjRLpriSlwIphb25Qdlif
osmWx3QpYOW7wc4mTlEkBg6ZL8pFmzg7op/b9QHBMiql2q7IS9QfzzxCT5W2XlxBAnstIsJf8Xve
1bYnjlgATESvSBHHcW9LX95ILEUX1DBPWv8gKKVMMsz3wJnrSrSXgnFi9yJbOj/yoW7SruoAmmy5
o8FSsm9AipXuHtOpcTQfKc4z5qVeFomj0Noxa4FwKUtqq9BNTxow3P5InZpw6ZHw7DKsMA5a9PuM
fagM7BpX2E2vZQckyA6UN0yBXUExqzH1PlxjYjyOeHbcTSffDT5NMNQkNQ7aryyhLEGJniXCwL64
gHYnjCLi3ZW6mRHEuEf+/DXZ9tO2AH2vErVo6A+fNFjyejeBvvfOejBO9CLXSQM0f/z8CaDKcJz0
/Oe7pezclI/3sikwizS7ZzJOA6Jqe5qhkN+igDsuDRzQu2rjOjk20mXRfg7oaIAAlfGkzi8c8zUm
7hw6W2POsk9o1nPajIfVS9y6jYzlRZBR6dNtOX5PEa2eWqtY2VBc+2GbafkznlZlpZeakKAU8c0M
wpKfWdRRN4MTn6WNL3In6hOh2ilN2TzOwTBzY/Y7H+8ftCg1h7al/SwWrCo3FAjoQKDJUT1u+7Q4
swKNQLg2vUpwLn6JSLbw6qeeQ5aQ2cRdxoEBXOdKKYub8zW5FmxCQykoi/hjKp1NhSMW2uB7Mtz9
I+GundcGCfJLFfvHCapmAJS+EAlua3ro8K4nIEMXfCogtjIPw7ykdbdropmB976KL21OPFrDLugP
lKSKLrp+8vRjdtzE/lFPVhdhLQAhLdrX+xGDwf3efacaxiq+uXPQRgkPRiwi/p5i6+oRLEdjUR8r
IuHeIOreQ1Q8OX/pkXN8QWaVfOZDknN5J4nh2h+YCRVmZ8XwzenH9/2BQRs1gbW8R2J9esC6gWMz
8pDTpu908miXLu0XJC+r4tXu13t9aOC3gztThzym0u6FyLukvWnAKzE9AabffOty7S5Xik5zeqhA
XuutSDCxJ2+/0YCHeMq2PTwFVenMZkY3A61gXoMIZjXWKGv+yCItgekO+GFlIPANPGD8lTFkIuYi
Ke7MZcu1dCE1+SbBrtON2rabbl9T5Lc4hnEeUCVwBqeC75Ds98l38RCp8RZr33PjzM8+bi4MFtBE
aW5DjyczOYAepO8qOvsNaIjD+2yl1a9aGhdxawowXK4gXvcolqGih4I5sr2OMe+z81QUw19v7By3
erMdz1/NSNbiTnP75ieM0ohlFnL0XWDvltektCnqvQ/BUCEMArwD4DoT3cirVJx5CH4qBrl+EnkC
trbJMy3EC9K7ks4eCzXpke9hlQ3Jk0XOb+knpFzzLLAo/Is/szAUSBSg3aWS+Y5wMHYK+5HO+pDA
d4+98eVIgj/HUkdODANDzqZY7PJAnnATeTzrA1CBYFnQSTs21jZ5xkcsNzcbSZ3f3jm8rzkA4ym4
joByN4wQHL1PQmLOYzxOAfi7wnPfoWMys5/wgb7VCJzQvKPMqug6cxXc/9ac8NWaFWP2o5UQxeH0
O9BilgIVMgdqw9eG9ROSLLZKzltisk0xbh8O9x2se2WvP8FEJXpJiv2aIyFPqIGL3BTfAPS100Bu
Nq+0f+hVpOUyhTtOh8ZiPAalqtG31XFFXEJWhSX7G0hycKeX1TVOk4pRY14VLa04+BNjgtd4+OsA
HKfldxAuOfmtiJS8hrs5VpNZLOAQQJ3F9g4ne2lOT2EsIDVmcbjNL9Uto6B22jx2HOXQBTE95/p+
mRZtqNUze0iXMQEWOP+4TM2QNL3LbMbocsdbtKBolNCVd4fY5kat/5yzKXNGAnoWO/qXrZKL5McS
t9q2H+sLwo+F1KPOoisAUUq2qzSSNujgU7xnNuCVX2p212detv4nXQUGdljSk5u+8PcpBxYg1Ntp
1GhzrOgyZt9vynAEuOzxkUjN6Fn/+w4Stvi1QH+lC7KxOzV7vd/7F8ryW3oZOxOHSXo8i1zLnPaA
vijmTnlsf3D72CiLSS27VZlYrzfB0ZxR3ZgYJCsjRz2mtzXDiRGecixA8PgISjztri5OVnDcpuC0
szQMCWfx3ua+rxQTT9wbGayXF8rYgeMVIgT5Rl62vlcC78e8XYs/ofLTHpyvW5l9wfitscTXOq6h
gCIv5pY1ViH2Wrai/J3WoTL00jmLU3lNEoTZLctZh6panBip5AoSXMbsTrEFclmYtUkRFZJD1YIz
Ylq9typbrPCpwZdzPMC+ngNAiCjewA03IUmg6JwJWKb8Q3/d6tIEm286NQ6pOYh1rcYe0whNhdRf
JEkljumWXgiwsms30fYwrt18+QpkBAhrsDloXI+dEU43QUaPhSBmqH5gTzpjD0+O6Di30immyedp
MyY9c8BoRluFNfDKduI+0x+orB2sCHvjCvl2jkpKv9tQxTxqU/UIUbHbnIAusN2xm8rgkCQELNtN
RKvITR8Oqu7qFfHcl2lunf0IqHAOV+3j+MGtBt9jzgXMs3SE69e2At3YLZbz44qXsl6NbmV7I7KA
RkP1xci9HtBZolwpTM1szqiTUXriZ9BIIhw/z/KpKmskj1VgxbGJ2GN58R8TyXtRa2jaP2KCRits
j4qQYLEK3KsiCo/xiLhNltBv7xSNkxIHiixcAvGfEqewvTI1G4eFzJeTUaie2y5f5WHJHAms/Ivr
L5GkbBWHGkjbyu/ZdbZVJBlRfUEOmxzeVJRbV2ERWmey9GdhY6NXzT1M2SKfdj2H2o7ad+1K0hfg
Y5qjL53Od6naMM4qKHmRJ8hpJb8B1v/zcBAhWuYnYsRVeVX6ZrwAhEIDV8Z2Fwg6Ty2klQR/2jdy
g8rVMGKWvoz0YUUJ3EzHRVxHt254VqqrzCPpnKoRS6qi5PcFxyJi7Hx/B6EQ4mmhNcyf+Gf69xiJ
shzTsiO7asFelODG/w50Thw/n9DjCkc3XbGmamXWeepyS0t8JDZL/SWTkKprcUob9VHuWngHgm+v
SPBdiLsEiaWHaM/oHvwlQfEH0PQH/SWzwD+ev4blacf/EjtKlM8Al4hzOzZMCsfPKyqqgyslLNj8
K6T8h5sEUnrhYRIKKHPzTt8a2rTGhH7B98A2j9RJb9jJNgoQ6UiEMBtXQsgV4Td2y1yyn2Pqt79u
hbDODsEVJWrV1Gixx4L0jhfsYmDOj3cgbUVsWsc7k6oEsKft8//K8GtK/CrNkjcgcU61yYqZq1NX
FbcYAMlfn3MCQ86NM57jQAIslElny4wq/1IaUw7l+XiaWM2BGLNi3P2ZjLSxlaaFKEqDCvdIT1kp
wY2V0Y0CBr7WIf9qyH7ysKOtMsPKqkJxE7vtyAUPAxvA21sWUwOIpu0qsl1nmI4zEUGrKl7yh24R
PGpQnuiataeN3aPRessSA50byYvm1XtqEWhmRlWaLWhTootaJOanNflGutB3oAgxMtk5OLQl69mf
VbotAm9jsoOTw9dD7+lqPvWukoGL/K0FSHmHoe57kma9gVLxQGVBfppCkCKK1exprZw3kBibFAzP
kQgOGVcxr7KmWgCIamdw2w6jUL/GuZcugdHmeBpiK0evrgsv0SxkvEN4tb3eE5seEQ4wqJwmrtty
IT03WkvKY8tgkYk2kL0jGR8GzPoiVNySC6/e0CaZ6xpPGHTzOgbPhEZVkQvq2S2byVz4VD/xT142
W5cWPfHgYAvqS10BNmnjnxUMVCxwy8/Faf6JXqOR9YlrAj1w+SmNbe8AwY+1Yag++zkSmxbmCm7s
hB7EwjzVLLGzXf2YA3AOoEIPDIwLyhQHHyUhv+PuiUvScG5ZFWWArTbokIl5Q6YumAP5jWHF8MxX
sxOBdsi52kI5GlhMK4knlV2UhumIWdYNkfcyUKcb50QI3faHWE9BpSFhzf9cHfLf9DlfuQzze3CL
4bp8DG3o5oYXSTLNmjwUlJhOt5CnmYVehlBV7HtUa+G1/E1ddQmU3Pv2Gav2TmUALwnli+RDhuiw
Jy2smDFxWeNFb4m1r/gdUt5VXOsPKoKE9skqrpwZ7uFGdMIrHFNtlx6aWngaBFcg9MWYvhksD5hm
rZd8rKH+SATm589ETbsnF2Yk54MV1uuC8O+u3ptraeJx+TFW1DjxVCUYJwhQjQ6WLn2nIOisVKYk
v9e4pYM6jBSLKwKAS84tiqTpIkUiUM6EejRnd9iN89sAIDhxE3+M9T8FRsXHa7M1J4gXSIifIPjZ
N/tcOt2bqtxNM73l71nXc1BerNCtiaHIx1z3x4krjO3NjYlakIMpzrYVm2s/XH0L2DzKH03e9fwb
KlHD/iPAPrEWUnchxo1nyk7Rucjd4XVPqF7EB9MdaSFLZJxpHW5JLTFgEPTUwV4onrtlSUIeGfLE
Jc2g2B+nsCe2YTULgeCr5iBIGdPdbK7Lkv5zVrnQ+WypESb8zCnBj48jYSn4OfRi/JkBtOHHLqOH
rkTcB5HJPkUgTpo8Kfow9u4+P1+4fjUGnWZZnLbtNCc01rtzVXBPlp0CFezAkrwI+cnyR/pGYPBV
XUZoj4NP6ykVBCtA9VPZjPYiFCmBq2GcSQyW9LmdJTPpdgnrHbx6UMZa7C24UMmQq3Ced018Vx4N
CUb4COL0cL0Y+uoAC9H0TD2WT2yMvXCsC8YmLXIiXmV6qXmBsj8mU8+IzdhThlz1sGHu25d4hiv0
6f+W2EHLFAtkgQGLihywCs4QWhZhRGKVMFyfP5jIf0VX55tekwlr/iQiW1il6PrjwClCeGo7Ihxq
+bwK6Cpib/SSrx3YwSICKwjK5657pOyGIYuHP+/xnkforAi7/bSvI3d8x90SN8y0MCatpnuau7uf
q+A4clxf/DlhEe8mH5ALgFxay9MvtvpZgNioNlOOpDG4M8IP2nDaIQgEHxFILV7tMT/hLNJUkx9B
eK9za7QxqTJPEFJETRdWUbIchUnphPc0T6QzAyGIljRP3fExvLoCmLv8D795LOUktM5WqOlpUVd0
9XP6pIgAln7rKRfExxHVhUp0ThiTiG5E15qvYRj6vRw75wVpEtF6pNomULrOY+YVrZzFe5eqUf8g
ma/JFJWpHoQZslDm42OxngUaXNv3Ny4+zB26XEOvUKAM3bkGEiCVP9cPcieiTV9VLQUSrt/Vk3LE
jfd5ck5QYgMNu64ifo3pvOx1BLUu5cNCMb1Ar3seNM7SXWncHYAPvU8q1oaRJ9S0Z45MVVWyrmLU
8RIbMRYjvlDxkEebwV03yUXKDKOT4Oynq4lT2o0S/MrLFUScjBiSvoLqcfOORQQVU14vzj2VkEy4
6Q1avBwjGhKKBM2Hg+kWCdQ+s3YmfMdmOAJQg4djHaknb8Zf9PLvdY8EtwV83It9jFRGtiWEc+FB
Jzxttso8HrLp/N0RtB3dls7HBlnnzrbTUd2njdhW8CD8p0F8CA6kKtzfJMPHXxZ8O5CAfvn23d7e
7T0M133p7MPBAD+NCLaKWLrWhdc4GfS5HjyFaqEaiB0xRIfKHmFL8WjXJCpJ3KBJUKZ+HuPyDLaI
DFFyZf1ByhFPkOJNq0IwP4n/vsdWDtmPTQLUe+fvlbOYBlynhK41KPKYFWYHotzjIAnMgQ0k875/
sk/RLcr6sAqk5kqixyoGuBDxWh+1EHbbHXOPdYbE11pxIwIHx3B6n1zRa8ik3l2k+5DQJOnX7ohM
7xvjwbqAWsmBNn8IKxIzo3UEx/X0MFT7hkb6mMcfrw2XhaRY+caIQXGE2+IqCshDin+o0fWMI/T2
bzHUZh2u8SUpTmuDPwJTh/gAxuzTYIYlhMYkdGnaHYMsSYR7X+2r/36W9n48il0O18HvXQE8O+d1
MHqiUFPLj1qyT4mqwRw8nubtt7KTpRTIZs4iujmQCS6ZTDkwLdFuyJU2H7Xjn/ZrOgpgmkCkkcoM
p5dtZv2Rgty0OnoA61I6YHFuxtipiWgJVrJLduR3f8klb2Em4ThaAGnXh4tS2/k8dNQcNZw1udvh
xUhZOo62nIqFRTfb7yzGfnCAw52UsT6Q7rI6ge+wZYTphgqGI26cAmkAhylaDQ7OHx3MzFaX/pic
eYjudPem04tvRBOhwMUmZl+TcypSOJnlltdyBnWp/umGBeojrGRp8PXNEsPvltqqPpaEIF7UcWlX
83cB55cnZYVLlLo0PY9BhmQCy3mxCGu+FKULmtF+m9kRrDH0sS4xkDcyp6Ei98nR8hDtWtGPzI1E
m1FA80f21OX20QolSadDN2dSX0daV2F3zlqU3cvRX7hJD9aMlAj6ObZh0LSX+CTNH6P2B+unUIRv
pm0qhDenerv0fTgDcnsJ1ixsWCAs5eg+GWCuXkWK2/AqUJ4CWdXrDLWwe5Ia3nBzQJUlQnOO6SmC
OnnHMM3l9S8XTZ7zFo9TLgH0TgskTl6+9s4nkIfqHsFJ3Bm+P4qUeap1wCyXsfZcXtCtpUtuFIIc
xLep+f6sNIxvcwJ5UIrQcP1rvJO9jFgc7b+V73k9lKpZxrA7J5nK8AaPRPDj/R6q5eH7vmAGLjn0
v6t6nlG32NpA485gfEd6+JyQjalUrq2g8nuFAc7PgbSH55ArcCemKh4s7/K7KGdYAPcwAfB3svvx
ANUl9x3njqXGGP37K2gZhsg2pKLFxe+2f50L1xFJoC4MbScSTumr/Q/TS18WPZ9GdgZGnxdHMUay
+DLdx0kgSi87N2Aq+oraWQ6q3iytb//qHMf85fpEXtGsa56lXM1PKCFU6cSCYeGICgE368hcqLMU
vwAC32cHKXv8gjWztJyrg3EVJpRNPE8pN6H6i4R5o5Ce1edcH9f5VUDqzzr2OxKQD2fyVJeJdo+q
NtndwxfxSV4JIQNMLR235iNEZvX2A/QgQ8QTQ2sHlLh8JTtq6bkznhJ1eL9PtPIrp8TaM26pn37u
r5Pk2DI9dN38iv+91xRv3r5kP1J5IRMHt3OKrnby5qF7M2Eh093ak256pdeXaTvNUdktKLVl2IAZ
31JXV3aGIRLJ5WD3XG/onEL6t5MJcUYyRb/zarhaaUVE+24k7zqLH6NRJqzK1Yub549/ZSlZK9+G
PE3IvXA3hA/wWRo6sORdhGbQ5zmck5YEy0o8iSwW59KoTVdsCMjyLJ7/+qstXyVgC8FqDa5COaC1
03qTOaSo90zi6MESeJlLO7aReQalQBklSwZWWPzYA3WwTnhgo5B6eBsQ6uuOnYWpG6WeSHSVlQWS
G4VfNp4ZXiuzPIi0ybebIAGenH895YFRw4TKB2f1fRLCJoB9M9gdo2krhQ8nnboPiso9has0d87R
vaYA/otRZGbqkjWn0zywR12DU+jNHogNeiG/rbUWTPdmxW/r+Co24tzX8NAouKVHnk6mE4F98Lwg
TDZ6aZDKLGl6ZYlS7+oYkCE9syB+8AK3kw4ZcBy4ujK4qIKoiHJc2WwaJLvtqEoK/TbSZIAsKB9b
XcoSFCqjIMIw7oRJzvuuKRUDFNjw1tpqeqTdI2kW8V1y3pZe7K1pCJM3nh69fqkuzDw5Psw4ntLn
85emTz+gCGwhyt0aKfmAccLPdHTe4Ki/xo9MWVm/3LOcpcTz/JaSK51ZHGKcBiVm19qWRS/WECX8
yowtJMPO8zCY4ydbTJUhPwwwUZWTDS28PREiA7VGsLPiePwHxVrhenuVH75VKCp4S9Ow+05ugDFh
vr2/RWcMjtPw6Zq5n7uS/Oka9Wcoa1lWKAVJZgKEVEBzthxeXzmr/LR+L5IP6AcwmgORDNkt+V/r
IxrF6AO5gnsPoS9iQhIv4uP1PAlrrXJIEtu5blJ2nUfCl8rLf4zpCPto8GbBXvssh/cSY0PJqU23
33ANMkXIRY76eeyyUuLTmMQmTsdXqXjOc2O0JfG2ZZO+R+h2bh5+HKvFoIxY7vkimy47H2+omQdo
ObIo8/nuPxzbTLC8D15/Zp0elJz5r9kPVC1gLCK01cP+IZzhI99QxyP5AGesuC0PUjDx6e/QQvl1
jnQjuOp4q4NkmmMfoF0Q+JeH9HoR26+2stNWvpO0EHr33enTBGR1/Obcc43QaCNH/ekuDcIIP7vG
WMJY06CvlDerapz3wi6YLTHsvIlSkc4XVB5PLmNau6Ohp4+KNIVLV17SaWUWiMMlOCqnLaNpMXrE
K+agvELQXp1kk/mqTJR3Kq+sYoMaTLRbNHQLb0E/LFfdgQNqXPnfOHO1LP3MNgPPNr3cCnw99GXU
bse3TQv+1u6++QodAt6Vf55sE2U3bu1S4BOEd/2g4B+M2UU7VPawAUDRSOuMlVJMfk17mT1mD/2p
VNs1vvK9EpWz1zURfVqgAEwQpKmLDg4aQ3xAeQduTqS0i00cPruevtT3VZgY4J6bZhnVE0FHk/Q2
rYlNG2J6h4y18qzKuWjSLRUrWw5kZDlcJWPmmjnCHacicbzbAR89Um75DhK31ej6oIrmi6MFqdf5
RCc43zxqTNG5I9xk6wmiK7pr+HLJMgvi0Tlan8n7QSNdMKS+B4FSE2shdFbXH2eW5HlzQ3fFlWGk
lRjO8/OEIBF2ZU1IRJd+Wym2NHIICony7vRMEi6zsFqMKCkPjVTDMtu2IKBA6IM/f81qC1XiyPgl
UrlvavUbjMOiwy6xwhAdQN0Z2bDbwN8jNJ7Pr/1uqiXxLOCYjTn1TwJTHU6g9XL35/BZstThZmI0
FhJsJPUYnusJV2mJDZuSQrz5o8Q8hD9kHdrRmdsBfzzYsqsouFmQQVlFddXG8Y48UCFzWEh8gi+d
4hsYU6W1TTH0GVN74cUwe/r7xUdltyq62o+asv8gHSTMJ85FCFfGUP06UTkT7cEoy8etkLJXSr/m
AocdbE2wGF+yvow6RYnf4tOMehlJfuVw2QBUsDJW5QooyoPqpRTZiseBYa+CMaWXMIzFELYlHP71
zLrg9v2UwPWXfbinjFjPLWslXEpYZCQZryyUuwQ6QyzlcfktKhp2yRZfHRf4Vs+EgWdSwvvR5qrO
d0Le/qMXZkN9p4J916b0ZyREHqbzAXre5fqFZYHuys1Ee6+iVm0MhYOyhybFudCW1aNOoievbxox
0G44976iUwIwkc4fIIIW9+KQ4ThyNhzHjb03Gk/S4CMIMsGsPeD7uJA34yTSapB0Sp6crF9N3EeJ
M/g34pX/4eU+zsl95wyVwb65krsr3wDFigR56iX06au6X//Xx2/zENB1AGCPznwXpIunEqPO+ljV
cEMSHcHXs3n5yC6i+67cBW6p4THtCkOr/0khp0M5ArLyx36Qzn4Nukiitvig5WRLJ2Zsf6rNB3XX
sbi3hwCwaMantQRbh66Yuwmf+f+TBC31ykJIUcbayJo71+UkZbylAti31X+VN6yZyPzrRyE4u223
KgfnQ/hAD+Nz8NhiZ3ocGXnq3uF5rLNEdi6AEwhINerFNQPLbgdXYRnbIA0D8hWMFfjcsxUw5ali
VarCLyxduSD6idy7Q9IPXo7e650/K1VQDPJBnlTA8DT0Ua860qT1UIsf1vIYOMTfNb3JKNMSuMx5
Ik0ZAJTfkKJ0oLUzNvco4MpO8HzsTxpBpYMnrw2mYDUeSO2JBF2qG3/43ERHWljwL8QxOdjd33il
C6EnFv02nMnnt0n1i+42FM2v2aRirvpguMZucsBf3qG2QPaK87K2Wpnt/mdLIo/FGoj15ndELgWZ
i2xvEl8cjcnUwiC/jWdU5BxneBftXEbdF2OzcQs++5P/c2agus3f/O0yR5BOBBDHoPJ3ytZFK5km
iFp4I25fWWsSZfmU8xqScBpErJ13GWOxx1aKqNhkgwKa0egQHBXEFjFuCjq0c+hTMee+N6trhYID
Hk383r6inBPr03KPYo+Uirto01PFlwfyyXsS5KOho5r/NEMIpFyAGlkJIYsY+DlPopQ3AzhGLAt0
2emLomis8tCT1G+jTZ5veMwTeQ1cAxX3StwDsj/cZUi3yAkHeLrfOg/OvEDEsZ6R2r0hBhENz8lG
K9ltYjOYnpxtHkGdsCLQGxhfX1Dfr+QjKvma5kTZohnldFmQwyqfthj+PTZYsU7WcIZb7NB9hkMP
P+PgNeyuPJUH2d6KnrlGHskvXXEQ6+0ADHWujLqo3w0PDRr8hUUBGM29xr5kAzZIEF89PYBvD0Dp
JiT9Uf2mi6MFk+9l7m2iy22ECwtHFV7ZmwDDe1Jkvv7WYn5q3c7o1MBcOlOUmvJr+16uPTwD+Eah
v/WPCp6BSMSPJiFOuiILk03LG9CkBbWpMolpS85THw5wKM9KzO4Y/kkJOaTc1qgmQAxWiNfGfdL2
xGR6h7iyhKsTbnljF+Vavcl3S0GCLn3+pz01P0jcHnyFmNOcFCxdSJ/Qkn0CqZ4D4mN1k1y2n6eI
bDjq20XoROefBbdIQXhMAky5doY7LuvIPlbOc4ahhdB9jOg6iRy5sBfexB9mKib8q5iECJtRaBXr
GTLIzmZuKvazFx+uMdlUrlY6TzwlhOdC0QmlgPJizeO6zZvKukk7oIyboEbLGUgW6PoftM2WpxsR
m+niEOjDXvFVPlMYsvIh7zSp7AltcatUZClSMvDJPgNQW6HbS2YfyeeNdRzVnqzSLiuTMlf8I2vp
Rm1bOdN4n5pDew74GvkS3W+vogZWX1M5aIXIPFD9FE4v6Bc4+wfHh1k4siQUJZ8kGRjzl89fXcW0
RC+HTbl7RLO613Hwig07U6ZIAhmaS4WhWTfNNkYsRgC8JOlFKZzwp2iuVG0qsWuhkC5C7iZ6Mhfr
BM3oZzOxuFi9+JgaC9Ei/3Gwfb7BtOIGlP7dvEJOFJFPnKlKhsI01SBhvQKpYKkchtGTf3r86xlS
x5dB/MFDOCkmajzt69RqmzCJXgeqtF5M1ZbUAX7gwbXZnu4/tdiIIvTfAHdYFlXCSHkN7l7rX7bB
xwWwIBxeSjz7sAtP3/0yWNHBuLd9NI/TRTtyO1u+X//vIr1PbetUj/UFNhEiBCD1CWcGKMASdn9x
n0r6Kb6t7t9tqZfm+O6t3eObAw897qR6toLkJFqz8eZPu6wtx2KCtg5dj2K1TtS7WLgtoqhMXsoE
uiG+uoDo0UtlhXrPpfHvM9nD3nAbhMPeUhd8uauBvOlrMvLB0iaxIAI0qsLy/aHA13uJ2Nz9IPYp
8X6wCNLJn2bZZcDhN8Gy1ZWj6Hsl9ibM6O1sAIpl5rm/cYgzp6xyqpYpK4FeR+2QgAhC7Q+BrGy3
zx4bfncd/v6RJSGih9cOcWapNGZ74e8mo6kAwQjqckL4r/oISRwxKxLc3f0GUq5hVvQP3BaghjvM
4+VxdbekVUqEuE5y2/mTLuIJky7RXk8eGJXRAhGybNUHsaDY4Gv+lGdYz9+aqZ3CVmcXYZtEfAtE
6icRJM1v2f4rM9ml3yj1ruzYMeTh9st2rD4qs8UUVXNRpvQ0+HiZbRn8uDR+Jp6s79wOGRVtgHdR
EqGQSHjxPiilrBIELkrtemWVn5SrmB6s+8vhJV4f5GCrTbfooiS5+MvOe+OjI6GEuEJ3VFcoo+EF
GZ8RnC2mJ94bNTtrUufpuQP1De0RUsDx98poDp9fEaVt8ZTdhbRnoWvrpYIazdFrm0vV1RoKFCx8
XgwrcIpCs4NKzJ3C0FNr0KmL7vZKQ301sYmqdRkjCtX4TiHMlqkprnWtoP0cLj6wv2MiDQTqBReu
ZVM18lWuJ9mlyvpP9iRTmi1IPUlatRTB4EP1n6Q+2eanr4YlO2JL+DwYXuC2dVAM76jMtr3x7bhe
wFSbgEqJU9lVEiNR2PEpiXCCEyoZMUWw0x4QWPqMgTotDYLezFdttGT3Ta3wb2B2mXCOaw3BG3xl
mNGVyUToQQVBtfwrePWZMdFblKkQ3TDi9lp0FZsbsnbOhFdCavZOPdaGPW3AdQg213e0P86fKRdO
iMxZF+UK3WfALCXMZ2PMEDYBGvHObSE+RvIfv7yDMEJyB1p/lt3zMaFQCoK0jUpeduteCN9V843S
5+L7mv10tBxW4Eo96y0MZJOlNI6tuSS1IJVrmaUoFWY2CfMVdt2dOEuxkXLKufplZTlGOFsCzMpK
FZQgbj0jpBxHjw54f+9Ol5fKjpKpbvJz98EA4rdLzCVxYx34IAKzGQedWkGC+FSd2fAiKWveBtbO
xcESCwYxLlM6q+m9fkNF3orLhVhewxY8WYIOaCgkgNhZKvx9nlx2RckxHHCD34fjsiC/kHN2v4jg
6hD9XMEKeXb4egKtU1VfrK5l37D/hNCan7quQwfo6Zzqg1W9EaddQ4SE2X/eYo5l1DRtTG4L/y0j
sk57kbfbbPXt5RefM5W1U4LOtkyzKZ/RoVE1VoIZKFoxJQIucSnIkD6UDfLyQE1//tD+S9h8bZAQ
R6mN25Ki/kGXoIiCPIw+4C506OUgXndmyW9zQKyClT23yhuvmZ0alR71SEj+562FK0V5tH0+Oq2a
gIURpGuG6vkOsWhRxM7RqmhWz9fwsWADUTx5xXmuf9IaggknwEkJa4puMVy4DJHjH8vZL9iP99rb
YtOb5ZbsHq9Sd4Gs+HpwWpzLBaP6zgIE87fkyaNWbdLqrktq5VboCmeiyOQ/kH9PtnLxqttgJFK4
9I5FMHrWl6rWdqBeWQIHHIDFluTTVXL0JxdsMXVjsBC2sPrSQgMPcJVNTcWnkZGXWpYiaYrh1jSj
sf8duIuebTxrAbzTCmICUZPPjdbvcugI26z2Fi7rjiznFh4kpxLYCIYxadXmmZm3GNEjTdM64F/e
KdpTzXR8LRm/Pt2hFWTpLLOES9aZA3/DUb5piZLkKkrkTrb/wIAurPm5m31//u0ACFnwr/LMhOkE
ThBcyYg09p0HznPlZCEDgqzw+juMZTDFTpVHX7cm4MHhi5muxnU5bIY5BLiVjWhhHCI+Jd+QhyLD
ywSpfobHiA5mQ9k6MS+gmJW8JaUVC2thboi6GGPPNB0SIVKAsWM4Sa5AleRfTC8zr0CfQSrJjyQU
NhsubW1kY7RORcD7v2dN8b/FmEbd7HXlfQsy8ddkVm/tCmsUvcdNU8Wx7Xc4ZYYi9VbSk6nRxxYb
jtfpGERJPK3gT4kd9whcx3dhQYrwlbtq4hxCL5Y59G+Sx+tDFRnxxlJ7P3ZSUfD5B1DQQucdbpkt
UVw5AcxIm8Q9ZTMOHbvCrDVfBgWqD0QpGhHG9Eed3FQ0h1TM7ppFRiYtZN2fmfCZ0MoJ4a+7wBfu
0FIPLd8fB7yCG3jUW6tSTjgGceS5itb4IvhF0TD4/nDI/Bv9RJnHrcFVyL44Achg0fsBXaCJW4XU
EfYIEj0fzQToUSMah+EtHE9O1h/0UYkTlGR1HtVz324TQDBmk7tsWTmrCIe8EKr8yYLOM4Dkj10w
lgZnjhOqXQVZwT0CzpS/DaCyfKgFTQBgOgiQAILvRVaf/BGPk1/NFxdqsAMDnD6JET4N9Va4w/PE
LZfnJcSw1WiuXNcLinHV0FfNJi4W5jLWyH3IyId8m6OkDXy/I3Ktw475BheoU420iVVBd8lB8stZ
jh8NMSxXc2pQL20S2fVLoJ9tpBYYfQoXOpeQALNcV02XCD81UIGhvEJ4KK+lhcHgvgb0XHSqtkrs
rVMHDBqqPtglq2EIiiFDB4EYJ93WDyRYfBTnBMZt11s2s1vdel44zMdULJghGXBpqJzDb8XqQLCl
7QI72LZ30vJ5pWK43HXQiXiI8nunSyifCMmozgtkYn8Dm9+mUv7TkjabAJlmSAq1fH+4nbnGmBgP
NIIB2CmJvbR9EUrZRc7QhGugqshLNfadMcHlhNdqlbdzqpL7YxZ1bb81VvezmyjBQ8MHIC49nR5y
Lxpb/FQsZiMGqmX/tjDP6D01V8uoj0335c+Wif80t2znkxPG5TTFZhScTQqYasKbvO8SsvzYiO33
H1oRNPZ/3BI2tu592UXRplGmdMTCawZ+iKDgVSZeilxrTxyC7d7LiuVhbeDlb24mbq271+ICTIO4
dEe5xkUlQ7/uEp3VlwwYpegbBQ7/ghnLPay6bF8pOPEyrN+AngojKRfYJsL73MM+R85cnbkDUXna
3WTiZD5m2NwVIO+0u6Ewgh+kYqzfVURwx4hf7m+M1BJYh+PIHt0dXypSAPKv+rnW+r706C9bEqCq
ghVzRKtoPrN7Trssc8ePCAY2S9NLi8xpH+jGLKeGddOhYYMlwacHVlx5yf+RS28EycPaxVoXSWUz
GJsXe7qXamw4v74lX7ayksng5yR6ggM+EmDeo58iotJzYyXcUGQONIMDmdclc8gkUQDNwY0pQJ/f
7sC1+33HRuWmAxCTPopLC6MX9JYldjRFC8K/IJiu0APQDxKSkHiTwaCZlnWuWdL+i0kP9NvENw3f
pi45wfv7P2l4+GhvUbErs/1OLBl6xMDSd5DAgNRRDDPWRlAllmiMeqj71+o8sLI/0HkuU/hP5ev0
eE4qgtI9ytZWMicTS3n7Dn7RvEU7kIhkSPwPB/MM4yl7ebXpUs62b1eLTSZhCAvJTb6VFuXNs/qf
2e2drMQa2RH3SBBVKO7X/4OK7ETzruWmplmvpCDWNj0wMf6TXJh4fiPFVe9uVspGxOUC6mc1RRjH
+v8svrIbovyZie3LuHSd5vSQw+bju56w6EfAnVbP3nePtRjy/l+4NUVjhMHbRTKGMQeHAYS7siA5
iNpgci2EggtztNAGM58t2oGcpQcIEHvLSbq8SmtgWyfhD3z711jRZUUBWMkdUzWKq3jvj95Vah4U
V+UXsj3m0WL/m3UjMTBU4wbVEliza29LpvXXxGplWJeI4L5nIviYqmP7KhX3GVc7/HEMNJTIT9XZ
OTeokMGo4hNYX8ApRLOr6vE0oYT5x47l9cl42GGXiPAcuiG/oEdR76vz94GcZZSZWLXYIun7Tcid
O+6+i7iB2fWXhyW5pvBj7rT7KJvySkU+xkOo5d7vMtGo+YGYwrjfzy1RALDxHvQ9rFBtHft1PTLh
rlXSTkJAocDXd9+N+yWc2TO7mO63L6k7C43yxxwoq8wK7JzV9SAsvMDZkrJLB5UZ5w5YnNWbL+hC
Mdd+plMFhILUuPgwEqf09PqaDWyYfB5HqPYnWQV9qfpq8AOm3VmeGnRpU2RB6aiwMrOLrUvp+2cX
ECvOFawqQEm0aMbksxRg/Q3T8/cqB1XU5fhsMaf4ko9Kr7AMAqz5HnDjcSN5ninwSiwxndJcS6bP
sWiEXWksrnFaUCRJH7+ZbYgqo6gk35e6W3ec0jqDbASA9dmYkX3aWoAc4c+azS3FKOdy7/ffGvnB
RzOQVAGeyA58XkzcUmQUcDscvWk+B3lg9Y6weoy0zcMg9VOL62IoXaD+EPQb8Crc+GP7KxXdEm4w
60tlAFDNIgzJ+yUsA9x569Qn1xqQaJa5GfQY5vO0g6WGKjbanNGsWRz/gRku9uIwiYHR/iQ+RUyr
pLj/LAsbodoFGQ9zRLbc/p+Aj1YxkcLllCo92BHz6gzHfIrIUXvefdKYnKeLJu7yMEtGYEFBI/mX
t3kGLKcfkilYnYBpaj6V/xrNL+2BwuCU99CenwgzxvqvvVJmWswQALcuEuItcW5HbFEJclbHcuta
YRPo5VPAumFChFshn/g3NHjbSTXPDkdf9+IsMcQ2ZB0r6++W4jHMA28XF0tpgNuls30u0KlSDfPG
W76aYC4Gj1ywBD5sL0+SXvpd5H3GmosmZLa7x6ZDlUpRnEm7abIp4k9CVoGVPmEuLouaE4YNSYxQ
SbwnovjSTFYXBi/n3WoIXQM8YTYDSQN8PqLc6SDDL3MbdgHZzkAUUU1RHc/aHhCOoD4aD4p3qcY2
QG7yzpkVPK0nuVqHVXtttWaZfXCgdZJdvhM0BHjj5SbneTVsfHF2sSNx+L0tNp4wqAUilhTVrdtu
bOkm2DC4zloi7aZz2qR6nWptov4NdQkpYyH21aneM1HVJsUWXHrvAAF0eClp++aW4XZ3CeyJ46g9
A8P9B0c4EErmdmYfzYOlQ/mFF3qbgoPZ+biP/CPrMk53GBue9cOmoYOR2ZCaHjh9Osdc5HGgcmKz
mZ+uyMOuDW+Nb18JUQQCgyP5nIVBsauzcbwcBGDWEZo9bxFHKJfTYBSsY2e9YfnppEwaZUK1+lq/
Rsy/P1xTZ4230S42moFqyku9LURU0zWpgSkHEOXdNpx8jtieFDF1dqijK1BEdX4wqJhXeSc9kPi4
tynk1rSpjn/z6nQvkkQfVKotnvLe1NIs7Ib4ZEJCQHlbH7ZdHttuapWD2xM3cB/5+MDTXWq8k/e7
g5K9X2+NPCp++jt4PF3wZCNRNrAbl024VVbykxK0rJNqCLTm0DZUmYT11uK9RNgOV9cp6luAwX4z
GnGpD0DDsx60q7+NFrMxYKHcP2Hv3DvZ2ULrSeLYU40+Zj3ZVpi1X3COkxrsdWYJDV6Hs/9ahTQc
5s/Av9TmNk27zmJrOBa7RWKIdNVL4ahVq2Ac2/HQvKHnn+gfIN+HXPLVpy1AiSu8JYFZULZFM4iu
Yzg7fjph8wc1kyk6V1ctzo8LYknLHEM/cm30m2C+DKLtPD65zDFn3SyS7BJ3T+Lz2WKAIwrp05bJ
cMgQo28SKBbxNv9oXXavTeNy6XDdqXbNg1W7DMljETsXN98IPzv5L/aE93EOkwKaq5knnMro4TNc
C7V1iqp8hjLA+7Ekmz6J2HvnAlLKiEM2/6W8VarF+mHw8/cLjsGP6NO5NrEtdU4YwWsy6EpNEj6R
b56xYJ5dNwFieAg1Kvj7/b/vZnCbV8IjDIIGX1UHlEuPrq6sjgkP+dquPyYRtRJ2kTFNiHDO3INO
6hxu8WibXTOc2yj8R7HJvgh8MvgMw5FUA4maK8h3IGWqNEQyrIA7UDgq9DfhDHRBJh1y8czwVtlf
BogSyQTw/SVtHbiBmibQxv1kyn76EYig2bCb38pf1pKBAnPnw9GBcWmC96tZE8RdbIEjPWJ77N8t
c7JwIEQsWvMegnTO4ccXEJ7lUe4EW8E8MFCHZS+3QMic3iPbTKBHOLh2eieMkIl6kGddXguguFwM
JZ4/kbNNFFzCYqMs2hoYfYVoXxVCplufz/CPf0fWQz8MUIlteob6wNNL8+TvS7kGgm9sKzkZqqZ3
blpRmPlngEepOyjyExzeZZSbtv5QuAxA0F4kECAIqoV6KCLh774pkAoCvpLmD0xZElAs9kM+71Uu
H+V83FWIMskEhS1s6eLDngB2Cr/pcydvju4Q/ILPHsa7l5BEVKfGKtwIKt3rTEZBfESC7EitvKys
u+qLoplCxWi7Ooy0Z8t5EjaPFou8QCFbcTFaU2eU1BtdiIU+krIQQvPWSwepf5RhAjq6Bqy1kpBy
prdULC9Dlgw4eDqcIwZcX0Olo8t6sRTD7d6QlJRnFfWckeaajac5BtLBtAcHCvpTuYNevXN859dT
vpHnKYuXm0t3e8qwpayABkHIKWZntiqMWpl66YgyuhRpNoiOaS2cLvsT1WS42uNElm3P5F6NON4B
mB7myL1g/hhClMf7GyrtHCVCUPQCu97j2fRVnpvrln8Vb6hpDaruic39J6xmIVYVMJaNB7bdeToL
Wa9skKSnGZR74YsZc44mmHLCJbLQqtNdUBxEPKvK5g+UKLBdETBLk+JFA9W4JGIgzoFxT3PQkhWd
CmHObVLviAzv6JiXSGf2Ttr0xt9SB/XXtmh6xOousLL+aWdVaSOuoBJexSZpUyb4f8cm2iqgue0M
pEP+Y5TWdwle7jSwz/gQkMh5zgf+DGnO46Bsni71PobVadWRSZySO8oic9r+hKITj+UM0vlnTZxL
82+0JmUAa7rgSqJQ6Q6y5BtKzlmmsJqcuY3xrPVQY8D58Rmh3FK9EXklFuIuWD7/sSbi/fIffY7Q
QJFBPKhjP3kdMrOraBHwJe4yiZ01SZlrbVNSpLw8Mycjyqe+Gu1yttwetZLjX+mrrq5tEFGZlMed
pMxQFkbEZNFS49mM4Cn0/qYvjbfmakBXKd9+OXQtmuqkvBMMdsyX9sj3HPzqpszJkCbKQzsGnnGV
UvlmqV0v20GGB4HJRlRSeY7gWKD5qrW+GY0T6g1G7mWS5KZXTsIYRivtETRAx9DUysW/Gg49xyWu
/aVGRyLyvmDoGBgWCzrT1wq8XN5YfAXZZogQBAzKMuus5ReSdKw2AMcMrkPvc2lOxgzMZJrlKW9p
IQ9dR5Gdaj3xnbhW06AqpuYuK3xnlXDU+QIBltBytdg78N2KaDZIk8O3AErEmBPXv8rRpi5+k3bR
8pvwDVpRmAMC++08UgXEARcVd6tin2LmihWP0crZqmaG8X44iZDUZvtFwB2IIMaUQQ+sN3L4SvRY
fFG5DqZK9o0KFHd753GLKQULrqwtPlqZcCrz9edEAiF8e8hNOhpPLUa+lWBEB29liDu1S9kjippX
78gCEz3BTfh9Mi6hUPnQ3HhUqcMMzOkP037H6ipz1IhSw38ns8Iaowo57sGozZlz+NiUUUitgKzp
GdMvRscF4OEy3qD4D+NP4p+CihNLxsqJX5ViovYORZcDCPUlxHxMVLsLa5rusO23B9N1Lwud48HZ
SwO5LluK5S7zte4rqrJRNQZpRqRB/uplCFm9tswga8lNndDwoLimkvE6pAbfryWpBsNhOyU92LXc
7hrasYGF4oafFLyzHcRYDVbE6bu2DrdBc4BDCu+Olgb/Jl0gnXP8D2VTAe6K3myKcRPXXO/+UVMx
F7wsbZ3w8E1W9qy9g4laf5aQ6tdheYk7QPPzxc58U+/8PB+cDVBuV+1PXTZnxae+oVEmQ8DzHWNu
O0Kk1j4DzhBrZgd2nf7aeany8bYHO1SXi9umtOev0dcClF/nTN49HXih9Ex59lGbYJt+szN4yZg6
YCGYYYNGHshGxfQo7t+6JRxLDVfWz3OzOf0Cbu2sgtFsRTbYwKH++Kc3hVNr0yVi4DC2/mHFr63r
Mn9HV8RpSzQPHb/xOIEAch7vKjAEo9r9hpWr3F4hDICYF8tl+qTy8XrnQZzbBkjJkAiPATWqqGYa
kMBBjWQSNyKNVZRzMsFWJMvLo9gVDAvoOvW5jqOTR3oBEwLgspXkRd8lNdQkCewv/pXB6i6qr4jm
srHgFvK08//LuubPw+09I9MJ6G/1/D86uy+zNkW2C6xCcism/E6QtDKCufyrE2LyC/MYe8LyeN7X
bsqUfKOrOOa/l8ysd04vtzYjhfRp2MKVrhOdgm1d22UTmXs/CZ+MWfhb4rXVYB1foPTbTLPFBDj4
nzFD4hNwPuvZqgu0EVPjONnl3lOuM64odZTREWbZ7yNMQdAtJ/yiHQOXZuZ383psLljqShOsm4fY
DQZx8X1KMPBfgM4KcYlz0IDo2C/mCf2ekHqZGr1unL3pKhFEuidku1eybMGDXJJ5kko5EWHVzu++
MkP0wvLxfNGC5fSOsqYNJWDmVTAMo13LluWZN3PxrE7sH5IrWR4RpvBkYRCzhaUsLyjIMpBASK9o
VrbpR0iLx9o4RabGg20cZBgmkYEKuDeAPGmLzgWQ9xHmJHPJoGWsjKB4V2Ig7MliqEYuJNGb1BkR
mQm/eYcXXpqb/7kqSe54JkPVbrt8MEuSaWak6RUul3zUYBugPCvYtx/fMtvSBzDUw9KYDWblxfcU
lE+fJr+XuErURWREp1UnRoRfLFMYs0BPg+fXfg6v7Cj6k6GpyLO0HA2yoIZu9vSMGalCdP4QTRn+
E+4D/BKUZBawKLpFy8AMT8XMg84VwD9J31C+M3iwAuBJyQvIA9QxMrz7FpFmo2/WbKaRXw8swM5H
STtQcCxhYdVIzNtZ2VrMnoE322mQNWsRTFgSU9l/jzrHR2H5xkABWsEqUTVAUtszLMUdzDjJ1uXc
cnaybcPLan3E/M58Ma0oeApA+nanNLjI4SKS25iQUWu9MjJhfE5VJLkuAFhS5s/P+LZVIWG1/USj
98kgTD3OLW7RY2XXhTNpYSn0MwWKkvxIm4CmpObxetM4BfF0xYPfGai7JYOFvSmWG3OgSd1o73fU
rOahrJqNg//zFRFRh8SXuXPvWYIknZ+E0ahaccOwPPf+lFiFD3YLVQ4H5gFL+8n2/rX7Z9NJXnqP
N47j8O+V3ECNOgbzLMB5PDJ2mK1A1BjmtHmyAEKoL9s7b8pJX1fTRyBHfziuQ3w14kRW7Zk5owJy
MR0m2Js0zPui1VI0dMp3gCKW10SwXNeJIQBiHVyBFHXodxD2xAxj9/Vo7prjd/voztSVY3WSJEQY
VXDsZzNOxlfd/Af79YqYVvLt6UbhaqQR445DpbmZoK6onZjHPI124pbupdmdVmlNMQPA+eBpJJ0f
oQuYDxLCRgiHcQ8bzl9SdqT8JXYxmM0xcdnbTpGfya1ENqWWAhb3SonT3V8mc98nrH0LypE5HeIX
iALahr4z/K1m1FsZKKWjhZBQCqZXPcqeEo1aTCV15mmnNUx4Xa+Vx9KegMFHKWyS0BmDE7b/rUQR
LYd7qwvlzD0K4x6ITVqVNPsASum6PN3UTwK5T9JpKmrz1Dt1hmswdIZlXKPa5PKzM0lIVzTG4v81
qDb2R3MAhsrXLrNU7Zh5aBX6ZcsQWb+CT6AY7I7aO/w9OobcjLe34ni4urIbP34NmrabdyzRwC+J
YVPyQby9rxburpgeaQuIloqmc59YrDL//X3m+gxmtBmV4PEpJCaW9/hzdQ0Cj0iMznDj1M1hzwEA
FR+8XQfK4Wk/i0OYLOc352eYQD52XUW1uvDLvMHWHknMUzYgAEvizIsyPU5e5elN1fQhYOb5TLSd
gYmfKnjOL8vJ4FEpcc0ds0ruh9YT/yQBf8X4b5A1mpT/9cUDRt6q6DRgFksN/uQkeSi09eusNcY0
AddAoBmGl7LRNR3moWyVXzS8c5wmNs5bnQgXbOpdKmcs2PuhMppj6bX4e98Y3RPOTkSUMcXFwKOR
dMO3yJq2HKxKBJdFSUU6Q1X0ONntp7SVKaujBinF5dJg2MjkO4PuimnmbtdyTRsVPRXYnKRNZivC
n/hIf8vmKxAh48pNgWyKEA6MAUwdixMsOq3vmVzhfEGWjUMjh2sWBNO+xfmDIFagsebs7lYAvUMo
VTkOUmNRW6/oD3n6JfzjCIgXybl89a8/8HUr2MwGBJbFAapti/1i/JsF6nKa0h55QhFay/o/xw8i
aQF7WKnLMxddnA6Sx+YaDfeqRDBAMWyTmPpFyEQ/tNIglPFkAccKYXVzvOIBVrE7VW0EsObjeuP9
ZMSbAfGGKAaMKevDlRXyE8jN6XBG38eQ4aCH5arXNl0jdn9pDhu/HUdL9lGbflIt228MC6X9ZrPs
dADvU+LMV0xDAliS8Rt9jYEoy360bIZVGXnsdknifhIJlF3U6vs11Z/DRsXIJTgFyrRiZQ/z9tcm
kqm2LXFkKiBRryi8KmgOiMMNJpMw4phasuQzsWM/CbU4yFMUZymauBqDG9y7/yjbLIpq3RQdDL4M
mYDT3abA/Ri+lylAkleWYB33NHlfCO05jh76DMwwvb6TJAj/dKu59P+wBC3zFPB9DfGQgm2x4y/I
JgVPqbW9g0zNEq0fUuNuAAlNSgdUi7zZN41fgUw1IU5A6WrOKiCD/+pNk6BS7x85FkHnFUZst2QA
x0qhoYUtxPiBhWX+gqtN/Yn9QH/fQKCm/54mw7Uw/mz3ydaTd5CLfOc+qQXkQHbJT0JLJgZa0qec
czVdEa7n4/0DvGUQYX3Ym6y4NUdKyVGvRJxBYEFHtbEmX00X9u0P7cc8jD3QIzhwiqU8Ek5f4LCI
jL70WLre3Drq53MgOqRuxEX8JF02Wx5OlVGPFmErETqdfZ/6giX4AI9dp9qJHN6i3tpCg8FR99b+
kMSBH13X7ecZwPAsVZY6i4Io2qms9hfSqDSzEJo2OG/nk3O01sZEeKlJOpX9CCTZtmpyqITEGQuH
jJi2P3LmAwvyW+TgSpzMQR6gcaLoNtQPBGAoeb3P5sYmOPz/b1+T9BhU6ECL7tO6rJs5WmfQn41Q
tcYoQl79cVTSaVQd8ZYQEQ1caqlw06WYQ8TOBgVIWdsmejmngyxDeUZOXq9qEjyOabNIB+S5dbbD
siFPcjmIxYVYvaNQcqQ8Rrgm6shLQ2vmpEuy9+hnwppCTsZvG4m8WNaHjtxrjJFya08InR/ipnhd
y3XM0Cg8YFOXmwmhIgWybHDnSu2tA1syWsnTyFi6hQ+cuY0HtLGZb9Fgoq9x8fMOPrObcDUnFGpB
Jm/iXEhURD2roOmNixr66RJlUw7rypb/tvBdoJXldYtWTIYloWAZoV6EjJ9esCeoMxaflUgVnN8d
Xl4zDSfQrOaeICsA8ZrlrwvFT34eT6rbKlLTTdMr7ISZHVn+U1SMQC3++w0wKMAZxOqQnxqxdsoL
w5H6qAIdC1bsK2fHBaIF1PVeHHzW9xNu8eHeYRj02fpIySkIAceAFNnVtUmD57y00XmQQGkWs9jj
mos99zs9n+4nAmgZp8U8NNZY/dN3MzwPy2CAE+I+KJYbzSHuAoTLfqb/ITqCUno+rSUUO+rFltVS
C+VFMyolqMBiW5U5X2dtIPADZG1YYLewHUGt8yWBruMTfiOYQ9kuHB64knBFjVqaqWxj22TLWZmJ
DYFPEaGBsMLt5tKwRVU5HzxUsk0n1AFp8+mOmALEOEkyDB8zNhs2lKUWr5BL7ohgPTg52A7bvKJ5
J2y1RgFx07mzc28/bZICgX3/AOvaiBYoqNclpdx65z/jpDYLO9nB5nKE2TwHfAAIUk15OxRD2ugT
OveWYZGsxtzxFziI8XGU3zblisKtfOveh9a5u9xYYcF7j+qzcBFtlas3tFZxjHIlOr4eq3+FgeZ1
q2Y8Wl7Y5sumzKAmvWu3VLTuabK8vqISlEOEf1efK5lH+tf+wDauu5n1RTJC5oLSdPjuhVbG7QuL
xuOK/ye9mOBVFAXFDJVPhxjGcm2yGC8OjlFQtk1WqxY94yEsxZfM+1zx/4JkRnpkzf3/HLuh9Xtu
2cl452HuJZkCIBBHdCPQy4zbPt9+sHzl+3Gbfu12ovv8ozTLeIs6X5YrkLegPgLAvi0njND6Jd9F
57ozYh9R8J2xc4Mm03SWKtha+KxkQ7FN4bFBfniiS6f97txvpk4PXpaOUEE9eBzICNmTwpDTGlpH
S89mIPVlrTYgIUkdbO+GjRqDLHIOC+XCrl7tPBkQHvjKpsVbUVyAzQZ+XwPrHOrP+U/tULPhVEVn
bWmE0d/1xHJ/8hCdHMWGitIxrtkVHU9aDNdjDrA83/3hOUTvnKjaB9bd8/ZM3x1FipCtAFIrFrOV
3Uz3txIGOE+UjhpoKHRfmSmPapY89hJ3vfMCAcQPyqRYFLBpDNV78eqglo6AUJtWCFUgCsk2KQV7
C9CFHOXSdWu3bDG2wLoqbgqOlW0Wg4V+dlfaxh8Hx4WkDOx/OA8UI/2+q+vXRTOfpsQJBqfUg6oH
Cju8s39AxDEDd9J18+MsGmZvjIN5T1/hWSIv4Kg5J5e6Q9gX91HSYq2lNnC/fBxDoOyKY6a6le+4
lRjt2veFTlVzMP8ZBabdmq6WOWb6JEhWne78docsRGiew9hIbpaG9glBQiFpz5GhaGGitwZKWBjd
iyl19Sn5jIEXJvAcpxucIG9fBZFVxCU82fmuLer/7cXp7SUK1wtR2rTLU2wx0eE7Buj0cgLjyll7
jw5dSgZgt2RiyNGF7SEsvTm21Gvx8gkH8tsXE67PClxXNWHe4IS8TgZ1Hi9xrvoTfvlZy4lAHicc
AKOkMSoaDOsI87V9Afu4eHTKhVPB15JalhHUNS4lKnTeXaYcKe106v78R9UJq1SpufIyIjg2Mct0
eS673IGgHMkXlCh4CVVe9nFTfp9ZPSQ7vTU/H7G+xf5xibSuSzA3KvfVoRGx9IDAEjKzgTWHN347
oczbPYbgBReqoQBuzxpcs3JWfm8hozaW+hTvYXRAufMQZO9zRA4Qqs2R8w4IOEwAvtpRYtOPqqQy
wI3Tq7QuH4SMC0rqvSUzdh9PH63rTqoAN5FscUX4uzqLfya/+C1HqVIR7ezeG3bMT68XhtLOZ6Jd
6k/uJHRe6TOj9ctmmiAt9zHHayuQElHMac0Za3lZmvMAHYmSp9QVmiz9gy9DUWi3Wy+FngtIMhb/
BD+Rtp2Od5jmfvtrZFyPtxZXY9NCZIvIY9YOKMzPp966pNpawm9EyVDAI77Dw+C65hpWaXMQKxtw
IZQZkkD7n5N1zwzMJRcpvF5sHSLmCDPKEXc7WHRDUb/oe5mESQOkH8k36E3G5sSdEE4VFDV/7yrx
axeyUlU6vFniQRETKfZWTg3uGBAarai24FAzxiAmWDuL0dhv+b7lZMWpBU7VY4OYaRXvHmTTbkD9
nbZLtAtz8ricnlxjofllcNaxKv5wS4+sXTTtuJXbl+2cBOOVq29D+/OzOEvu6d0KlCloXwPAv9lY
E844b2eujioS8ZL/WZ7JbIJu+b59f1uDQ6VrvYj6Lpne0wbxIDVAmsYgWJayzh+YW62Km6T2KuUq
tjzWbAT88NBxffEfXL2FSLkuHPHouX5/55m9sWBTeyT5sL0+QV5c0kCaFwxdoZCbZRAHHXT2yGLd
5RP73CIj+jnlTz1TI1vgP4UoQTwrIFSU3j6iuMnGJwowSvT1EVx+b0W0ZiaDyO+bcWo/mAer2tUK
jwYgoKUcozq+fxoeg4b6QY/qDApAV6Wi5lSj+c1txRFu04WoImdmdMQJHuaKiI7sd2zftXBMbC9i
VmMhYSLmxOSl0G0LYYaOKFL+49HcoeFRXcrTaKhICvYHO+xEpJddA5+URS106HNTS0UQ52S+peHo
S9OgBVIJzYhtNWFL5I8CnzdCIcOeUueJr00lJyj+oV9CSdxFiv0V9coSjQll8J3ri77cSstaR+S/
WOVXjpnJR1pKaHgiVyOFrJ7DT9bpgcocsOXNnyTlNuylcK8smyWwVLP640PqerEbRYfRajSQMsfp
CfEQZNkuBj2LPuemwtnm99tPvTmUHkQM3aoYaRUj7qokxmrtBOywgKvmhvuLsxLKk/5w7DP243HB
/giAG0uT0NtfcUh2S02JkDfj4CZ7TzUnujkHBeN3dlPHrYLgYspYd7Gt3wVua082G3itFRGnrj+7
QW1W3qcNA3kc2m2Zk4N7Sbkov0FrPpOhFhUa1ExtFMh8ZTA5ZgWeWiHj6V5YZ3dJ4urG5eMUOYd2
0kbzC2w3If/FKwO9ZTXICg7K5pVOq91HyeWR5ZSV+jHXBWZHy7Uy39CzFMScTYz6yFbigbSPTYPX
3ufIwM8eXO9rySrIFuZst5stbZPBEbSK/jiBQRRhZxr37oGCZqOH8zammtcQDXc64XHq5iXICUj9
SdpD0jC2jb0/xzVoTDWW7d/sDp5a/TxOWZiQFSByZu4a8gXKzJsng2nxqSp4Iyb7QPe7gC0PBqOE
XoTsGp4n7ccaxOexLA/+u+Zl+mXdTM2BKhB3ql6nHboKiNAYz66p0/XnEjTAYMG8j1LGvvojGN5u
KlDdZMtATAeZKLeP6WkGgZFxB9De60mKabtSBi556w+wxOWDIMdsk2J1IQiZyRCEtTGWCyZkS7It
CRQlPJHpCsUIquYeIRolzvw0CNZ7tVAkvFSDDvkF94YQCsLNRutxKlCsfmQ5jnNQa7VtPm3eFqRe
JF9SvnUPmm2UCyKF/7W4k7DIDRAF6IGIVUKJLX3VbYsC4Boq+6xlCpBX6FqtS8BvSaxsW6sWe+gp
BuLFwXxqMAF2MCsRW0XFVt4kjckraAQk7B124Vxbj4Z5GbZ7W8YrfETl7NNEdtkDg3/U2D8aj89r
om4zterpdJiIxDWXf2RAj/e6PDE6OlUWlZA4gI0bwSkSBzLMSJtiOb1STJlSfgcd7alpKYYEuqKU
XmshCGC0eil1HD8nGUxK9EaWbbD8J3ny8RQDkURDey49rFnBV0kkeA5NwwWIpS8TnxDiOc5st2jG
YN5PznWDpFDPcQxHmvIw2NXKUSGRJoAB0C3R4WQ2CDqoVX25FHK3Cvh7kIZ0ta580V/ow1eVgrA+
kO51KLUoj9njSWqFtSE6U5NvO3AMmWA/jc6YToiZpxFWBZg4gZH4BeBF2Xd2VQFO7MhDBzfr1iU2
LNJofCY6BCkMkYvUEj1gW/eMPQ+AAdXABRrxm9j+KADvMY3wceKvBNXDd25NLs+50ctw1gExDXVp
YByRRCZvT9sYCMxHGwhVvTQ9pX2EOot1ukX7jfHYRJcFUxiOlZLkGg7F2Y/rXmYm0ivmcGAJbFqo
7PkgYaQE3kfs+GlxzhvEe26ORvsFSCvz/HxgOjfNzLMzW3wUivAWCiRF6lsv7kdD4+yUnF2p9mSX
fWA+SmrvMsXKae/yXYIyWbz8znXTgu3x6OII/JniHZPbdDtkq6H82JR4IZmGzxjDTTzAoCkl6Yzm
3jG2s2SvpLnR/vFmy6ENX89rmB6xbf1zEJ0cSyXTIQ977rkwY/mVUOIHy/BPzAP5Q1bzU6gyd0gF
Oxky/VHAgMAxlfhfrUj3VsW4FaCh2rnT31OH673NioZTHW95/Z7lrst2ksnDLyZaIstXpj6EHJy+
p8CNgDaSloDSQRx1tXVtOONKaCq2eUfXnma0Xvz249SKVX5C3sEkLQPDr0XSapbp499VZhT94aHF
FOmDsa56BOdzgeYaRW1lVtPbKRPjF9h7CRDfl4Ns5kNoOv6xyrNR1xzF0B/6jKJpqUeaBK9oHTNP
kmWmrHfh+FlRWZUwsWpnqEkYvsiG4gMAYCYqbXEpRWTBJ4MGmN297czVUwfCR5/Sil8z/edyTGLa
pnOB0HPZUbJyvXBGdQFh0EBSOQryZqNCa3HLlm2LhCk6lV1KjL2dHRdUbzFlELpqhoWCuSwtpdSV
T8T9/1wJrD4krkUtzXn7ENPnYLptU4+so9+8B6aeBy3tcaMyMe5ymEyESrOX36hDNN6K9feuqaGj
1jCl7tGazAxh0S+psCwYU3dGAcIuEzjmDfZ/YguMAsK8HPixGCYns8uOWx4OK+qf99t/Gw3HX4un
f4EFnPp5Fow0XkOvZzvbXe03KOxCeHi3D87/ec7YsHmXC5VWRvaEULRHufLRuWISKyxgSrQFp4kK
dbKClJgAk/F+OBeuOo/0LFouoVaXPmiGflt6xsTX7/POToqLE7VRhnYWbqmbqd2YLfcWdQ196//D
8eOr51pzjQyNj+Wa6v6O3Gd8YOBgpXopSC3ii9cF0sJ5Fb9wHKUe9bgw2xluMWWo2zw30cMYh1jE
gr1EWlyOnh1l4k5QuWTe37e7nUTHM4rGxaU6rHjpPmAl6yfnyqGMDHOD//icxZYqql88z19k0pkD
syfjU5syMeFeq1l6PPe8e1tRWxAoQScC2wY3N3bSf/S6OzLCFMxW8nFo9VXyAsPHDk51UgLR3tdn
Dx2GU9QJT1UMXFe8shb8UWPtI/gxqN2kAGqnDy7MRVyfj3pTRssq9GB3xKDzsO+g5vlTzeA0UeeL
eZanGVPGhR+BFx2vWcVX2zNirt/SvvF/451aR1l+pwJsZueyk4CrY1uG9+FR/yVUtrqzRorx9y3l
kfpMJ3oVheuUK1apdPOKTHu8vP/XPNRg2XUHz6pcsUJauE2uK2OKVtnMMhsmvBoKkeUz9BBED4dH
Is8IYOb5Y+rNxrPGOYE5vYhn0ww6MzpNCvuBugD6XwAolWUa36IDplpS3WBMGm5XKQtr05t0anI+
cERILwf5zLpVT6YkzWinzSGRJQVgAhQh2ZcjJ7/tCjEEKbAFOmzu1EgoMjfCgeiw0HF/TWCzGvw+
2B+VXdAc2cDQGiJFfRBEf7SuXP+aCgjx3IlACrIoux4YB7JWMCYKJ5CyyPwTcr6bS9GGhCZ2y0qe
6Qdy+2+yxH1fjtz+JE2wCpHGHHeu9EI9EG9vg1AxYVcps9Y1JfVyD7Adj7Lvtm6NR5ljMDwOqOzB
nSJFAtCqVwz1QZoeTIt4QjlV7xccChEXtf0I7pPaHrLlyJdBVYvtwObLf/s49z+LTYyG95+j1rGa
yXSiMLM8mAycJ8YnWWtT/rwxeIWCBwG0j1rn0IMzxYhS1PBtgLvGFZvP6Hxk1lfQX1H0/YTf2XMI
hFHKJ+RRIh+GYutgkRGT2kawkR/+Rx6SnXp7Azul2zGM3MiDvWdTdeLieU8kNRFW7g7HRoQ3t37T
G4zSOr77NwHz0+gB6nooM2/xIh5HYBMx4XB6/9K3DUq4mmlkvs5yQVDpJKDcTiM0+cp5i9wdig5N
ckXfqYVlKxgDpby9LW3I6WU7lF+b7/iS1RpU60MXys0fYRIeXGqJbMArzu3O2YKmj7BN6Vs8Sr4n
QscrM2W5AeU/SyzgATwd6+lKsKxBjRvqWeDZMjIHQdNft12w/3gk+liIegerGLAs49y6rvC609iF
F/XSmFXySSjWlUuXEoqA5UOEsFCun3z2upQO1pe/E7B0UvaMFFsd2YjQlkh88bKQfhMZm/cf3kG4
7BamrZal83EZSj89GVnagcQMkQ5gwhSn1FNrfcO7yg7mBVMYu/ECi0v9BQip+WpQSwknQ88VBWe2
FhA67taXfbT8WBepxKqHjs6++gwI280GKB6xTk0gwI/44FdXwMTVK70aUommhKXO2eSN3RAV9C9s
S9pzcNP3MTEkvpr8q97BbncmlFSZDdwp2BnMZaBdv0PdOnr2P3q+8BmJccf8hEr69GVq7EWkW6Kv
v2njzsUKRhn/VHiDgmv+AXQQMEPtiNkJHOo5507mGVz2lryFnlzCVJXltxAi9wEKe3uBCmvr4u8U
Um/dznSonNS4G13jBtp0vVHKoO5e9/zyqbay3Hq7p/WKGlMywX8LGuQ96bac7SUncscgeGu+HBaL
XcRHRhyXmiKMnPzUEvZ+Zy4lXlUGWJekAMH4AtYPZw8c4hVvt7+5eud90qXYh92GpjkFwo2PsrOq
ZH+HA6uHR09lO8CM6hpB7bidng8SQnRd86tdxbOadKNCpqvkbSsuGRhXDbZdBTPsderXUw1pWEXF
53v0JGaL4rqZRT5uGPSVMkShGQMs6Nq1tWxG0ODGIl+A1FS3vseYZbe6WkWopkkD43TSQbvv8uvs
3oqfbhxdPzWxbXRjPM0bYNL1k0SrFCQBJ04Zre9e9t9bQZsGe/RYCtQlI75HSh6WxzHQGm7488hE
gKtokpNj6VCbWQ43/JMm713EQxJA47o/1gIBpknZlIhvcQoZBs9XWEthXh+kkNBN4tBOFUZWUcU3
ByRWqGMTJDph9VhonO2JctswIGu/u/p7q7ft3TgZWYm+nLcS8RUrk7atsIvs/D2Hv9bPeeEsp2g8
Sf4+RANnFN2TE0HCqq31Na7qM8Nc5ONShBp0/IiqAi33zhFP7OhK53IGmTDvGJJ73DEOEq/8ve49
6q6DO9m6hMPYaaooI3pEsHVtecg7ezOQRNY/kSnaAIN7+8UceyUHxhnuPpjaP+Yr9CbPrIEiBAiw
8kjgaRwjXb8MZq4WDXEZb4GuOUsSdv1ce4rvXPyuOf9fEABDMVhgzOnFNHQznpVa2H6IZsyZQGT+
f+/UQyfQXSN01FY2lXp42uiVTUXpdXVRjo/Qj9HB/BIZLsbt6rO6fhuS0YOfRzjq2ar/hLctKhuN
c2l09IAYdZq2HbTaAoY6otrqslQUpMzoi/1+Wb14NctYXvoZiq+P1nWUdz6P/9e2s5BjMK5cv5yI
NCvaLefOhIpDirUx7qWGJdQLFf1SaGblmWj8CoKXwWgJNyKFZj/lnh0C5o603HLO73FvwZS3z4fi
TcLw1rcBMFboLBN/VSUD4zyiuKN6mrS+EqZju+12imCxBdqs/UtEpZRk0eE7u694fv9BMUzAGYQc
xS6loGl8kUpSPhdHYmo86ylOGAq8cVLha8YPeXTLEQfqaXxJB92ldoII+CgIo27CXO2P4LKyMx3t
h/exFUIJgs6xEUZjhPWYy7xK46HXehTO22p67jUNKTqulZbQj1CWUQSJExIovoMGgOhRqsoZ2yFv
/9Ujzjr8BXemAIjI09Q24ZT5rS8Ur3dp6Q3KFjix8YHmPGwPElKN+SPT+qT6hSAKtbZuDAxyIv1S
qG6lLGLT90O3aJMJO3uvztcKuuPrY56dqxkbE0WNGyVqwloPwuSU0pwXztyI6CFZLbr4yxhBMYta
Z2FexUlN2BfIROmGYuBSfYnkelekBH/m2Ys2vh670TmKpf5/hVFq0zGKsTK/td0jl0SnSmUvoV7D
XNDoyp+0dAEhfn7BOWR/VSqQrBpv7I2FAenIMs8FErwjttvc33BzCfK7FmJhM9YweNQ3ltHAzsJ+
AG1J2j+UJ5aqMNlQAnZ59LYnWCu1biQVJHQbG01jb0sHw2zUb6rVqiTAgKr9HZ125dq0ULoqHKfM
yrdHt1Xe2UKavYFgGORtYwwkKjYkaL1xnZbrg5sEWW8SJvFi+4wLaj3AYRboHLRBFhfIHQCE+Ker
g7q2Sk2ksr1nE6dzTOLiz4KMSUeFn+70q6tvLCHuXpSKP9Y6wbcZHHqJ7glRjxOO0U8Vr+FepEy0
KHfagtXIfLWssvnA4EC5MQU9H90dyVNuIsae0aqZVWxs+TS05cCJiPY/SLbWsKFqPj5/Qkmnrc3H
nFjCzn6UqwbMQ2+hrH1r8Wr1XrO0GLSyE0tNHkSLKqQyleej2epueqEVchwVKh9k6slnxDAweFvF
8cqQMFeehqW2K5ixEwyaR/Y9zoeMK3vqVzLxy504QdNwImgYP5/YqT+9L6xm//UQ46ENXH5dqsc/
cTXsZSe+Wl/DBViuCoMeBfeB5SYqwHsw8c+nWL922Jv8SWROfhtNjtts8fKD2aAZIwN99N8eORK0
DUVoBIhH37ydJcc4ghuod7+OPc1TDiwmK8u42+H5UUIBIT4eAWQwyzULj1jPIXGRNTXK4rIxg8U6
9tEOITfQsbAt+QjWID52zv0vLdLFrQB7fsev3I0Z6b/QlinsVo/Y8OLIfGI8pBuDTW4PpadnKtxk
1juQHAyB8sijrpzNl6CLxBghVD8YqFiWxTikRp3OWFKBSr1ZakijMX5cjW1G7hbQmNZOBG/qXD+9
+mSFzooTdzbWSWfIlDZ+3rnbNAGZOHNUYoqsR0g1llhtA4nbKJdh5ck70bNFW7WsKXydJZnolDOB
DITUHgD44gufojKGtfnl2GYI9mXexuznl0jXNnN+/Mu6EO1nILI8TIaBOLIbbyz2nYN8KeJBoM3j
zBtCOWqHaxH8QU8/aH9umkHb8TRoew3B4RPwX+KCrsKlVd9xwEyMZJvF5mwueYbdzNVR3mZ6g2d7
HXT4zmC2goJ2MvkNUnC8zvnYM/uJGZ/RnVXBBOiPBibHaXkJh2LlDd17rMVmG3nUvlCbRQGxBt3K
eNrdncCaOdkYM+DyYgJTqc6lqbBvxTyV6nQ6SSb7oQ0laJDUGsLZvm/wNoWoyRyeFHlC9FXsifRR
OI/Io1MP2AliQIDjOeS78hYdmx9ynX4aYQZqwAwL6RZTM5AJlcsJDVti5/BKzGd8AL08zspJNYpd
LPWru9XkLY0qYI17H4tvlMLWNW23mVLe0atJXgc7W1sj+KgxUIpiqB6Gt3Vu96u+LBKoAUeS/zhT
Cx6cudxMPtSIh6t1LJ+sCpmj/MOZaN6YRNILd7j1IPZvodcIHwzCoqnLOheAXG7oZAe2uwRmK5pX
CrKXNV9vd7gvEr3aWvijT2tIM3SKbnPlHAiRYotk6XPh0v2Ui1yrfbSK0yEGDQcYTiTCpmrIW1aJ
tr/SoFZttOLbjj7XLU+5F5TIMMydbfL/D/9CLfneX7n1cKsglqhI01HTd1qyPbCIMX5req+Nf7EC
/zS6eg55Otqk6RClpuMROCPPF51sIPZoBZmvt61v0EarRcPEKDgYfvVzrShErXZ/47IHG735szQ5
k6F3NWVfKvXYvtucsfQ5pOVB3XPMDCbO7T4nyP4ex28R0t+D2cooCm09rXwOkMosza9o2YM4EY6Q
tJxZ8tYJUtYuv1aZpMZKfFEL//62+TpXESocsIyguzGKojxgTnZi3goxFpUBkCIOMnvTeyvvRB5D
PbW+8UTgy8YLkjYS+68wgUSwjBv5KM+Pq8eBLh4Ww1NEKXMhaUeA9KBWVcekhZK9y3eT24rFwOgX
R+Jo3+ObFMpjw5SFUGf7d8Oaa2sbKXn+XfxqQG1IjzGg47KNkxR/icJijStKlOkV8Lt2bO70z+Ht
wgAJugtxSBLKo0nlD0uR+2B3bc0oYLJXYdk3J508n/1goJwU74FoG2oU0w8BbAQVAaPGZEFk+DYN
CcTV45Gun3G/A0zdtcqqYGpLKXOfbpaUGjxR2ML0qt2QZ4pYrIyQmpOODYjNd8ujXyhDxnUV7wWb
wsEF8J2czfxnCv7AUnDxYfpbZtuuIM5nEvq/ol6GU2mt3kmXmZ5GsyrfPhe/CLUDA1P4o9Cn7t6n
8GgH6aZZfwHQWztOprWKmRBjfzHKgwEvGhcAyYjgb2H0QLalyH+v7MLQMRw5Y6My33SWhi6GypeZ
dvcZHcIn1xEeO6V9m/xOIDNKf2V/jPem22GY5MtB2XMds5G+Etimzq4icwJ+MKaiX1EN2DNZDZ5Q
bMFplM12meQBvBgOs/wk81Qo8OmZUZhnP1STUp7Ybgq31nTQzwwpi28KcLjtmFdMmVmGN3D2NRfL
KDGNUtQcA1xNysndo7uf+KKPOYbxqjFFBVTLT75EsnCgWynPgKYBdfQnYQiHNPxyHiYf/XlWGZIm
00eaNyuMX/mVIDAZIlA2fpYoPYGJR/U3LYAunprqlpiNtoVr3HbDZD1BbRHElsIiU3LJLK0qs2AR
DMQxOAacqTuAapBxUOxqNs3fJ7bzwwqE4MeyZwiKKqr0NNbUs3xKD7bsYlJxPJahQsVOAZWmiiYM
OnBcp8A5nJvZk60USbrvBXR7WpX2REzZ1ekuAbMnrW3I+22mQgtGgoqTZdb3YD8F6ZZkhLB1ddW2
/JLS0E/sKqBOAiGz76soxWQIKUWGwCIipv8qCJsdJrsuACmU2X4o89zzeHdoYKDCshZbYmSY/En8
HhYKtDM+4ENbKi4Z8jZzXo+U1DnmGDLYoeVv2oxRojAsJxg9ZRONO7oOxOWfWOudr6fuIX+RLB6E
/8YP1d86HEyCbDWaM473m/tX4Dw8D5VPeC/HH/A8fFPe+yT0hb6Ld207VBOY/x8KfhZGosrpCdmT
RHea2sl4/fhfa2UROiDxo/7mWwBItcFUIpulrlLqPuqY6N+j0d8RkDG5O3TtNMN+dp90gyX8LBk/
E291EEHrEWpJ91SRfobFi+jllb8HWM6Cypu0QdnvIGPOPgp3ApqMjSb+Vb0MVrwKT+gICfcVhPv3
PF4vMS+ZoXw6ORiM4nVl4RBw0tEf1nGy5KSGuYU3l76vrNmA1DQh01VQXhBufSOE+KLUrzZK0FiO
Uh1kNm1P0qXqortg89tlpEBSYnvuHi61UXCrSj701A+05P424xdvKXFKJ5cfOoedM00RzJYX2HxS
KssGeLEBeWYI23MPIKghF/0LB8Fe09o+/LI6q0AM8IjNZLcBPYG+OEqYK9je7XjDij31wPu9SMOh
womeqSvd1fD3yC+gFWpmek8a69UMdLrf48i+RpuD5b9QBoOZt6+w9LKbRKKKRECef5GhAnl22YiH
BbtC+7jg5u/OH1hxvVpr6gs/4kzUPWHY323xhc9MTQ69n7P1SVhI6Z5IDmc9X02zKyS+R71KEFpr
EUQTsCqijl3o7z5TOTzdqNx6VmlfKRt3L2tYcfMQkSDB1KQ/BdgX1sir/yA981HKX0u82lYiZfmS
BVRY8YSpLo3fROHRyq9K9SFgyHj4s1ttoPZNxF8rygsZM0Y1ZKfmRne5hJGxrxk9PMlujjfi2TIb
xlxuaMdr7hASzCQbi/K5w6NHh+KIyifpzDxvWEgwjHrvhVpB3CVt6+cNAvSjsO6iYDvf0AvDiWQ9
8NMx6/D8sDWbveFCyR78tpwVg9ZqIJR8lrLnj3vyNmu+qUGQs89yfYPmXMeW+Hs6sQbGAsnla2fs
HZMyaySNGWs70tVLw1d8h8yBhJH+UuKWJy5hyX8h5W+bZ4DqRbg2fWcX0k2y3+YitexQ3eSkS5G3
hDrhG3RhIBoM/TfFPz9Pp+51yRmdvmHGE3oP91BTMzH3B3snrjBQYNV3oxMGKCfrJZUAiv1jCXfy
5Oknr/VdP/TwlHrFh0NMqyBBGXWtDV7TD+PFDmx9Pn5ejLRKJOv8UW2NWGi3AoU28MLXc1reVNJ9
8w1TCysv51UKmejPI6HDE6Vaa2HDHM6OohOhEmSLIkHa9M6mVBiP4Vqqis5jkm7K72pgeul/bfJX
jlpx2RGtYboECUaYXC6l4Ux03XYkmR9fvQmv2aZByArNZJ3BzekUN4SrOWFXVq1q+0DpL+PRTymW
VZIhkunb3FRbSKdlTkvj7o+QcYiAg4W4nLfWd75buc/N6/jSUn4/5xyJA04P5gpTCL5qt3rGSQW/
M5f9MW++q+KbiT8foLy+1r756zl9QVJYp2anox5NQjYoN3KdGfQA5JB2Tz+vMa36YT6v6MJqIHyg
ouAgOr8l8KDvnKEhjxvwAIlpmBtXbNdzF1mT567U3huwQSpIoQa5G0kCdpb3fjETmmmezW0anP6k
1mWRDGW1y74MifqbNGbhHevaJ9BITmBo75n8nUM3acxoycVmqlYvILzGrioxGU8YcJVnPJlIVuCB
hpel2+gDkiSsmHUY6H33iQh7JUGeI4oV8W0rvQEKtWRcXF2PLAH+qVLql0Lr0aFx9EFj2ApaKxAR
AM+Iujvodn999Y181IhIFrb47SevcX7tQwR9FSUACmYdED1DQO+m5GXtnNNUhcjAiU5d9Vz0KTPV
R9u8QwOxfKzibCK1LZMm+cCu0FPg3yZC5ZyFho2AnIMAikn52M0TdDyJl2kT3Lgtw88Bbfkmy8Iz
odme/K552rkDb1mZ8QieW2U7Sn1ogG/EUqBivJ83r6PiztCxVo4lyT/BTUABC5mFUkznrNY6sQot
l0UvJUfpGD+29ds+//PDtHUhksEOge5lzkp/xKa/SiLXv9ho3kVf2C2zw0Sb7Isg3NyTmWlRVgSX
9x3zhKVBiSlIphFEIJRzgKOAo0LUXZbkpLCeZFkS81SvffBZ+vj6im8XhprDrVslBcpSso1Trcm0
weN73h/YzWu3pchZaDHjL/eHghBg4CIZ8ppSTvMurQIlL8jrT/qpIS+TdYPBNQLvSVxhcftZ9PMP
OCcA4MLk5vo7fKVjwperVSDLPh/+kvE/juhP8w2XuJBsidmWNT1HcVdyXWjf3tnBtqvQXhiTVAw/
l5L3GTx+r+AZ+7H9Hv8uaQitppsfTj8UOPkYjAA1Il8DL37CdNlEP0EJQoly95n79FvgNE5PQeqZ
ezU4a1GoYp5l/hm7K+pmfPM99iljiJ8I8Ps2eCOA/jkkC7EkAh0SlL1/OnZyxcH1ae3y1rKahNc0
j5XWc2w6eCKAZLNeIqmSzh/KT2yXc1FcU1q8XYpshbFLbWwsu7rkgDV0jRHTA7Zq99uj5Ts0zy7/
cy4wsasxmIDhBzKMs0WNHJlsU6QioywG5iOl6cBNziIr8Lb2T3bnnR7nd7CXSf/pibbdYMsQdJNo
fhv9MJ0EWYH8sBx1hDCp97ifwNYIdghEtN4nqVO241gECZmCjeZmD+o/RfpArTTNs5dT1fvA8TuB
Vsl2A/YiNic3esb0X4w/BXT+FHxd7g+p2PTGVcY8bBT4eVgSAvnLsmuZuvKyq7L+9hxT9g7PqVsa
ichi1DI5tTWALyGe7dVMdHaBegcAkN7ZvQHNRhp8KULC0UwF6Gg71/npzAaoDGYiH6K5kIwwdR7Y
Uwrs7C3fefGDmritcutuwLiF3RNzadoh1secHHEwlqvPgq2Ko1Mp4iyVHl/f+dVZSu8L44KAUWpz
oT7+itM/0kRu2DOCf/T9tiEJsLNOrXo3ed0Ohat77Vko1ZE1oUvlQCUO/U/TN1z5rGQz/CUJSMkL
chzf1p6EurhHl/xmtUngrw5AqvkZmQ2NkOKjKOh5G0gcgQV/UYLmZgHZvOR+gLcQN4lpvitz91V8
99f1xnMF91pijCw211ObEB0DjC++b/IP0d9RkE2zyYIbtFlQLV+OAqFvVNEUQGwn0VPdlrpUhw36
WUr179OFWrLKokg0VSARdENAh47un2qa1RVIrDtzhfA7ggDkNMpZGBk29+1mw/29WKMQonUj6Bgv
BwgqXsWqUkFqNBCthAX5fXEVA1KGwmsmjw5bGt+rdO5CDiGJ4yCsaXzZl8UmbbqsRALpuZCQbS0x
5NgFPWUt+Wwu/LZ6SIqG0ZDbaGCu6bhEpHoJuN8Ngtg84y4S70kbq1ai3FJXkKfGIGn5vUc8hmDu
8kaBzx5JR+3A19ZJgk21KBd2rX0mh1n0nK/s1tVo2up+ZbSqCsElKe8KZpi2jYIyUfdmS0JWRMLh
QLEI8aUxrSbXHMZh+B9BXd+CiIfRFDlaNBgJF9fEGjdikMMN3RJMcd7Cbb4WBLxowci4LyRfViZr
mgQUD6fHIJplKzB/dpjWXWmsBuMUENRT1Gtn9BNmPsO66mcpQ9J3YPncagXxeWuI2gIFJN/OArSD
i0dVrJrTlWqDV42X4jnhEQAuf0NswQ9lePF5h7/zd7RqKwkweCL+zN//kEf6Mpwm7dCzEYEATC7P
YqidoqBoqKJ3n2F3LNcoxiNx1+n0BDZ+Rcxf3O4wP1uk/UIeg8SVLjvh9G5wJRTMdCaFjq/pM4Es
xdWWOs+EgmaSrrzI04SYz8Gfj6TkQg0FjoBGdxRvm4Kl3QKwwEk2CjHOe0nntgL8uZIlHMnZVOGY
Um5XIwFS0p60tNadHqZU8dDtlTz3ueMSw2aLRnPERiD83izBO5+fpXu3QFd3iLAQqgsZU6sycpVV
XZF2rT791aoBCpXiProazWxE7KUQ2BwNtaC9jUu7pg8od0h9zeluKgHoW3RyRZQeuefB/vNFVadh
fg8Jg86LDFZm9c6ZFk+C7nn2ohDl9tUTl3vFANa/6UoYCR6fIC/jPfKBCVH6rFN5cdNBNIJTuHwe
u7N33vu4j1VUf2dRcF4LamHfrzcbciflbWjSjGDUGhxy1JfaS+JWqWAuBapctYPINetxCllSj8my
ZUaYdvRt/KjK8j30okylcZJDlzH7gKepqQApPEJjjFCbha9jYm+dRL2WQ5PU+EYrbrgI0VLg030R
oLmdu3R7IwnV93T3Ujd9f5+sPmFQkWYNjxIRqqmHfFeDElG60Z6aRAiN4YmY46O4OYyqGe0Tmayp
0C347yWWLMcmes6ChGf4AaCFmYW1dv1pm2nVcDWtEYHeWPwsMNQeaIlN8Z3DxXYVLnx0KhzMF1Bq
Ochy9hQZgVuGHi6jXloq0smYAX0Y5fhG34QI9/HPxFd4Se9NDK2ldMGCTex3wzYugt2juB/MHedP
15ygYVkHcZYbQIgmhk4Oo3Slk9nHZx2XNCCVm3a5CIBkUugre/UCtC0QFiXnLEfW0qCSeqhjccE1
6sCRt1rfCPC4Bj6JnX6NJFA1QCgyVeM6uW+iK8amCDc4mIDYLgCCGo8LbWc/aRNn0eCUbuLTGMO5
lFPaonPzxUozJkYLyf+AMWK7CIzPIOveihlPEwgxPmLHt8tjPW3CREm7wKBM4fStR5JYkmMvbvZf
Ed5Gk5KtGz3O0jqIoPBpO7xVw6jOxl2thGAzepPUR8hzPtn8T+Qd89f5K30lxl593Ch5vuHnu2nl
Z8IWSvA4uM5d2AAxTanJXOjN0I0F2wH4lDAy2rJXDspRV8pgIJY4ZkR1c6etDA/FcKp+ue7YHT2K
0/tD66jY/IFU+mOQaFpIiLXORnGOZKfWrQa60O5eM9Rjwgd7c8tei1c7JCcz691AORr29nesE+Pl
378oEqUIOwLGXJUSxZm5D2O7ydCNjBQbkTkvyx/wJCCccpc0RBpBcDrGvjkSl4fMx9rus5judGOo
d7Cde66q1J1smg2LZu6UICopyZCSQykwOLBOx7bbAW35xMPXshiY8k6mn8BGJ75ofjrA9OVVA//R
SdyLMP+wSYB2vBQto7kDl1ljcX9p0bb70lZqXPqBrNLwby3uvIv4P+DzvgMHC8B+vR/8ZONCnjUj
MVx1SCZOj4DeRy3ap4Ermck2bZGFkotxTHOTWqjaUPA7Xsu4UWc6ZuNwzs9WgEuoDlH/UY1sVAmF
fzZ8rAtyB8rhtjKL7FoVFverUlhRwU/XR0AgFgCsHKApRxWgP+nTs1fQcYI+wRA6hlu/dEn05FAk
b++XVglsjiYNuKMdGzfxvNiqAe0Be4QUQxgkX24KE8Glymt/tI0Ulqxyiwh8XlCctfjOMAdW3ZtB
UXmCSKandIlu6nonQzCQw2mGErdNuZ7k/in+qeKOjHL05MLyjtE7+LDwamTidAKNMKTNOl1RwYuc
u93xyA6SDJunI55l8gMsBRHZFSBWe+TRWI+Bdw4+mSafE3tR/dpLocDjPnXKxLKJeY5ms0N2lRZb
HEiJs1qpgugaidxUDJhoosQ8ZpdIP5ue57/1OZc9VQi8qQgkqQYTbJNswMEI9Y5HbY78Rv2PITRE
EFJIWUUAKDSuXaf4RRYESrdotMQLTO6CIF4W/uVi1ga2HgDIOTO42wlcTQy+63WL1YpIwgMxK/Ew
dTMtQnXjemuoUZzt5smlpuH/Q/cyX9/0cQPmdLjbOW9g1LD15Un/lJ+Tk2LrCnFigXMitaQvw/s9
7+bb5VAX58cs+rHH+WpbX94lr+3m0BGykdS3bVHk8Ml52P30vngzxyvy3gJx5FAgHfDJ1p/LWwD3
CwDiYuwjINKx+mX0GtTySGxcjnqYbdrnzAygq905xyvKgs+ImfUP9YwbIGY3Jj+IWtIS3HxERQfi
/l8A4sF1Qv6lmbOTm+uM72BjaMG3PnuL//JVgGsFOrQrvrbMJfdfsRqG/Cgqj40S/KKBabrQSfMb
do4YP6YJ0Pj1PcoKLNUBcYGkTqAPN0e2hQxHYXs4AHxpBbGqmOTqwUjjqYiM3UVN9abTzBLXjrrc
8cl3wtQiHbBt9VwqiyygN9aBlEk14ph2fkDLCJqS2pMX7cHh+bHAXRw3q7GSvI7bwzhd8eQXQqJ/
eFuDE/t1xyva3PHQzPJ2WByD1RSgnnsNjrd80WCV3SFlMxWoQoraTQXDqW5XqnWHAup2TSwHmx/O
Z2MVKVXzsT2gt6xgiK7HCVzc75dCvmfyDC73mbPPMfDKD9DyljUWJuxLAdlAthYYy2a0VGjf0oJ6
zz6P2y87OQDfnPx1A7fFiXn442YFdBOqhbTTFTYM3CkUpLxImdvkvKi/RyGg90MfErow3nzq2buY
nJjELQ2gnP+i/Z82pkin8jLLaGJ71pKEuKVboKv6eY8cBX+6HiQEKseQBnnfFibVZOuNTVeLX9VN
fwKEIOiUZ1AFb1FvBfFwxbgH7GGIRWNJrJ2192m6ZW+kbF/khaR7RvDrPDLDRmwJTFM53tVPcmwE
6lJP3WqsC6NefGfOrp3WWrrtfZW0/kcvmpLQbO1RvbJ8/TuVoUyQ1WSg+kTCfMFS3CRtHeDRv1ka
JMVcIvSyfeI8ZZXo/gd1SGqD3RKRgC3D7TTU/8tJb5XDr/CEzExKQ6I6hOMTwIEZH7wROGVusNYy
srxfqwRtIU01lsWjNx5/8JliB8HesBJsMdmgXfPY49PvBWlO7Nss+7djpMSLj7moK9utMIHligww
5yjX7JQAzcjvtLzVSoj04LN7KEgcsNS0tJb9cJqnxFSEtvK3Z3KOYVpG9sFoKPKVB5SXHpV710Ak
GG7qSfyEjDrj5gsgzWFbLfqm42fwL8xkjTm2sv5A9Ha4SsOyqmk8yfbORrxUQhjMe8iUfGTISeGQ
nID4IAM95V5UxhxlbyqU0m3Vbi9DcwfoGdfuTNLh0cnf8ECApx4heeAEPaXq3SUmORE7yH4osK+a
HgEaHyc4wpOXl9ZD0BrHT6vbGVXxDeirXNl8vr2ITg2hIi+gm5nHvNeQMTgXdD/jhDVgJe16yAvw
NrYo9ATBBydM89R5t8Shyvu9+KaPRixUNIzYlQFqhYJu31AanhxY8+r8RXF/EjHaJT+FcQKxjly6
9YV1frVZ5cr5mHbShdINwAafzIhyotGk84yH9Q/CtDJc9WOxc/jG+i0lRrh1X6T1zfEmGPIQ6crT
bB7K4hai4OSJnwHqNPeXH51pcfiVXx4WmzNetv1AaAZxRKd9XTDESFak5JYzEgS2iYqCSr3oAk/K
RwcpyDaFg2AHK2HSJO03+At5hmqqClAf4QE20qw8B0BKhbzi9LAEHUCtXq3C4Vf7jz21GMRZ1rDa
V8iffImrw/Pacm839OVpxrYHrAYhaUUeJgzPWuwdI0QzVHO9AdUKWNqnpNmlhXRVZ8q7exbhS6Qq
DsGe8JYkZ+ZqgHYzEJHfvC5g5QmT8jR+gLN8+MvneNdFkamNC3FDl90MXm1iZq4dDVwFm7YIkR25
yhMKbP4oQ+MtHGQNvbnCiUtfAsfazGauaLYbDOHmFvGYfqIqx3EvcBDWGpn1L6SKODpkNCjY/KRY
/eDdmqhparW+E+97Els11TKfvleNIJwIogDO/wpTjEMJHj6i84x6beYV0qSEsVT8Q2sMD36aXaf3
Rs6Oefl6Dj4DVXifgdBJQ3i8KZdDeQ/TsyFn6ll8KydzNH4dJdsXHmEq2QnjYKqz2usD7H7dpu92
RrjqEYhvD+BoQ8EQYkoFJ62cI0uWAZOHQnTUSA07fwbGpAO9PdGjFiFcFxPZirtOidrqpImnPA7M
l567y5P1ri3xQhCi508LRGQefn3U4TtGfXoU6WXCqLJsaq/TaAj9YafK2LPRVp/Bn5CTAg1wsJ/7
GvrTwkPmL4Em3xHajpv2oAOoBmQNHVvIKzqCJ665wiEzzGhCQVjQEdm8fuQ3IC5A+ooCxd8H6qaE
IpA+gWY08DFOTvhGrqWNx1xMaqCcAzWoZ0bEOkoQFYyY4H8tMnJiTA+VFuoe4pylJXkiFHjpjOBw
taLH+/ZBJahQxPy1ksmC+erC3ZIG3+zWqVg+dNhsOI/0V33Xan0cKXByeq74Rn1lprpCxigT/UxH
JEen3bjr6Yw7y6A80tLmSMBf9s0EsXALu8vfqLytMVxKLm/9DOpvwi+0E51aNAWWACjkQHXSAioK
G9revO1aWPyP1CC14vz018Rgmwpd00rV4JTyndRAkJtlIBkwU2LgVhill8Lx10ZuEY7zybfcy5MT
IqsO4IgPxQqZKktq2kDCUQ+YD25uXqqul9CU2Bbg7kA7U4IcWSdZ2YDP39gDCHMDg9UbFE9olY5U
uhC2DJI5LmxPOdn/1RYrqdB2SJbQSJwNNZ03UCJjtNyHmmQfvY212eOTDBikGZD5vpCLzKrgcSRK
bPvgMJGms+Gaa2M8gaFHni4e9xSMGapZM1PXLXvw3WLdQa16gMFO262mUbXIHQnbA1eGkCz8+j5J
dov86lzn+Iz4bZoDXAF9PuLqQZG9NnS7vADxvAbH5NMLtz+nli/OerVp8H5mt+fgACk6DyYSm9Vz
dNmGEb/kzRI4v5oqrSU6FnzHo9cSGoyN1mtNQgh32Dz29hQB6uP5APEBep1hmUiIrEM5KRMORoOM
r2rBdS4UmaxIkbbtlW1XNMw6tPpaMMD5lqx/csm+V04yjEaLx7DA9EjBhFUbZgWAgvtFfd3C14Z8
R3M1kNzd+DZfvk3bMvtRjoPN1AVvX1CwGZdPQJa6FGfaLTANFGimLN/CiZ5U/KXPL/hcZHc7uXq6
vcyHG4yOXvBaYEIYONvGvyU0rBvnuMMLpF+5Mf7sXCrMqHdiQ1OnhpM51zMjGW1yqTre1pwEi63S
Rt9N1f7eM7coDnuRDU7IxZfap/8jxLmdsZprCMX5wS0grzUE8mc3BwP6AQMI7+sXkSjehlqvn7T0
HH6mNj/fL8hktxc9hxFcqKpOHfMd3f8Bd7keXt0ogsADS9L4wciJwAx6FDrmx9TU94uPO68oyIrM
cXjPoiQbduM/YOVM2s+ZFLcv84SMezmM4KN7w9HH4QYXsu2WTCIqijgXjHFbnTCgLMURyeGKpUkr
zptYO+ujksiJ7xDBs4l6lIdSRmFMlJmK41/HOa8Cdg0dyBGzo2Wrvo6MPQlzEbCr3wx0U1CXgW95
lPBm/G8iSU/EPFcrlLgEQc3/WBeL1enmj6BF7R+20do7+CnZuGZDy0gpkGekHse9EAOyB/PWij6h
YU7rTn0lSEtz7wvnDJ8N6s/2v9vC1u4+HjKJ7ly9fBmwwnPTX9TT9dtwmRH4b17FGXqoOsZDCGKF
s4W/DZNXiNmaeupAOPOs9j4vwD11EuITU0JmXrmhrff8LxDc12nuoNsUkNXmh3xP22dJHcHd45eX
OueVbXqLyQnsyiPPCvN/W/NTf39g9v2YwYgE8MOKaIhK/Ycwy0PxBEe0H8Ko1AzXytZKIfhjlCwi
ZZU+ODT49SauaIKr+tlxLuKextdtQ0qwclgI+hhYjKMvF66gq3fOEnShqd3Dz+4apGgQEToPcN8r
kvO4agkUkjejSWf+IWavRguNMXhDXpDU2wMeohKyRitfnO68HOXI36e/t7MC79zIvOfRVvAsuiVN
CnJ9loBgXxoWgfKpCcCD3gWJ2n9PLIRK7BmAELFLBaS8jLb+pWn1SoFKKyG9MztH51fyYmPZKxnL
qhR3gEwqctGmcQC5e/XdE6CrMH9bUpnEu9UrTptOQwIJkVBQyXwYWsWrtbC/26RFhBxhaVX23bFX
+dghYY81wdgq/+MK4XQa7IsPmA8DVzNOMk8IySVb7rMd9NtlOpfaSx/7kk8qX5rPSNH7KrRRRgrd
nun+BX6rInpmeWQCS+uNJnRLPWApEScetL/RoYXftj4VCbNBDN+Otio7Eak/Qmsse4M+9OvqGH26
fHHTSY3ma3zChb1IgRsHsxGFzSCrtHnbMVL9B9A+vBhawIErlQ0pUZao2ADzrV3hyzp0yZ9zT7vE
ZY/vBJU7fmNGg7eSrxUyYUvpjWz0Acq9uCp6Zi3KTeIQOooQIvXg29gN6f/whV3M9AbrVz2Z3F5T
yVrRzaK3rAC6xupnBD0s3obSeq4DjRCKQV/O2vcLvqczz52VDvq4rTxxm0nwssWoevXMobmLhv01
SmITKI/NGeTzmwbdgKT28dZM9S49SkcKfMrII0h5vg/VWXICYPZf9TLc8xcTOATi72xAG9VTc58C
mEk6KvR54M2uf6duBZ+227wWcSKvZA+CVgpnpgsu7XNby6Ljm56k/9O/x9WvwVXjrII+Ir9PQiKx
XlN6GwchihrH1KcXstbxvHqzL33YWOYTT4VIj6kw3yvbrX9CCLrQoXtU7v0YV/r9L98K88bWERQq
/3Zu7Vab2IerQAiJsV7X+8/AR4LFGVamE9wNkJ/pAM2qDac/kQeGG45K6Na9nk65YNpNjaoCQyz6
VplGYT6qIsvTH46o+ncaqFmVxBu3f3HmS3munw3ZnjSTO6EOvnfji+Nl6+lcofa5MVZEbEJo1QXL
nYhN+kDc1gipxapWUJ1F0bid2PKteOL5tKUafnWQw/l2oCu1YSuWO1dPxo7TKm7atuOXdWYHIyO8
chiLL+FsryBJ65/10LMAqneMAUmQ8P/euXhLo5ZVAO4+168YU6t1EKUVBbYKnMyX79KfFMj8eYaG
lbeyVWUy54ozdR+ZTLwNeX4St1husclvYnInFO171tmrXNjd4/IyQUjIgDF5fYVeTmukB0otNPgL
inID8EnhiC3GHGFUIXzP6y25gEyCjxx3bAEK63xTs4Zsost9VSsTyrUI1YzzKFBhPNrfH1sd+r3W
LwnaxJIx3Ak85rGyfyazDMjlOxwWW4rRKVCI5SKauEJ3vDevdH+wHfOZKJdl8BWbiulhg4EzHkzr
WRh6o7a9HP1YDV1FRKqtmdLOBmrIp6D7vJaeOYNWoB44GRDUPaWy5IcT6/NidGGRrkkrH4ur/ZMd
XGBd/ei1RO5U8MWhHkOZ0q/y7ETB5495xk6Bw8qyR4McCaUEWlL1+Vyhh7Xr5G4wHMRT9RiYtXB4
IoKwCHQ24WT9p9VI2Kz7rZE2593N9HVJrr20Ai2za7ULSoOqZZidp9BlDzU5cTndru6j/IPiMFuZ
8JeDttO2YPnxRVq/eLOtw9IPuP1JYkwdlpgz/lYn5dXyJvmmbLqUc1a2itEez57A7WISV/8HVzJv
2oCKeoFgUqXfoBtJZ/SNsPlUgkIMOdhn8vKJP71taQ6L4aYuosbstdaCeX0sSHCkQu0LQrtNy88z
w02q3cR1qO9SahNlVs17IR7/TE57sTyzJqVJ5mnLIlOt5WYqWA9dGTc8BJ8uk5pmr/aLbHENDJf+
lPsuWmqaTx6MDZ5nrftgqt94hsS3EV3s8zhvM3mSSCLYm9IQYWZxiQ5L0S81W+17u5M4G9lEydJ2
JV+nAaz6UQXHuzupaz3UyxevnOQEPjR6fKhY+li+0uTDkEtclp/bOHrxtVgdcHw7mmFTY/TLyZPT
jX4FJG6d74BJWBtIz4LIVDUm4XG2TYZignhGprMQlINzBSyxMDbg7ewcarOsAkKH6KKVqmi6WKiX
012TvEN5Eo5bEhe5JwZN3c/qFMiuIZBbkbZ94EdF/FG4NGhEi9xV3ENEybxK+8In9ICVbtKRJ1Ky
6OqJJKFkTLfBh79AnUJkCeTXsaZFacdj80Ncb484WNXwgGuhEXO172lmKaR3/ypAquj+NaknT5qi
GcCbMEkeJAiciYWCROiX5mFVZK5qPGpEYRBII1Xk7f7S1IO4SmxdHEbjrw/HV7/5f7TV0jLO9YsF
SzDi4XxNzHOp1/MG18eV1seDhK8/TdW36sfo6+7rEJdhCBGfXbNKTmX06Gs8e8u/jawgs9K6HbEh
u5unonHZzR8D5W7ODj5d+p0EG5kZFRl/u31WS1j3TrFJxY0gMLp8gLHyrfdpi/JbiQ8G6HQbxKXk
GwYEu50GFZT0hI7bbLCJRL5uIEdPaFe7VG2dzLvsxhHP/Ekx8Yzw+FtkEoghhgsLPcde42MU/Pfz
2DDPRi6vlkyKA14WwrgzKZFTCD7/umFG/56O781OEe8MWr4QVRg7Jumy03Mea82pceDfRLA3u3Fu
v4QR8M8XFPT7vk+pG6nK3ZcYJ6XtWDJOzNzlhl3Tk5K+HcdQDnJL7apeGk3qdi9/ZYvyZGUaSbCf
neWQ9cqATCSSYlkifvQqY31WrN60hRGZ9WAOZQo1hapD5fMpbWbFfYRDgrKyfffeLIwjFo5UhYP7
wqnO4FKddDYo/5O/bWGL5xgjOlCh5+cx7Xgl8BkqloehZZ3mv1zrq7/+oqrmi4cpDjbRYGwlKx+4
iwmUMrD9PPqtQN5PYeH+aw5lmadmIOBf8koUMVbXWWAilIJ5W6Ovlsj+HJXpLlJNcZOqquG7ozpU
YWUmtrJ75GAXdB2arS99mw40gwelRBcHXJ6l8H8HhpaGr/amgL0fXio1p6nWNyCz2XVSR+lKOHFV
8PoB6EJ9YHodpz1I6HCRogdL7N8/5X6livF5kGzYhor7VLskekC4jrF1NgUj15tIisvdCDHh2JfA
uQYvvAlR6XWy3IORjNnXFmBguXgWwvs9qcBFi8/9mCSHg4FRzg9SgWURhijP1DDRGe03M9F2SXKr
JFPEnGnzQ69ViNDATcFF9UoxXAOP8AH3LQ4YXyvsIQmL2XErt1+SDg2hDJHSmrTBGJ1pLlKVPWc/
LJtNhQZMr8j9TehvaneFS2JTb0xIlMKNhO2bdjtJ4vM89KYwb3vGOm6/E0DRODt3RmYNzbQLzKDd
0/u4poLl5IcuR6fc5UL0tsiwsfdDtgA9xg1rzHY44OdUtRd1FMo0GlGOTyZSuFf3qVmjtF7buD8l
0qwGV2DNcnr6FO1YW0pBL1UFtqQBdiVRWvDh5EIAM5qOiUY9Fp+0iCgAr7QJQcvQwOSDVa/Zs3/j
RCnn9xrWlfs2Z8b7a/WsvmI7Y8FAUzBWOf3kFrclRUNwZYjmfKPqlOtz2XGiMcdoxTw9rO6ypSre
LLOL49F1K83F/NkQHabOPVbLJuA7/lItpn0za2i/s6VfUaVkfZqmzny2kNOtMFt3+iIa3CCuPVvi
0YaIp99sPBSbRFQPEHIdwrCV4mJxkXg9xyRAZDayueUn9C8V8MBAbz0W6VvUYZWY4RpSjVC46mLi
WwecUcKSv3Nf0WWqhlZv8j8zGOvgNMri71EpWjaxjC+h15GusNaWXN5A2Xru1OqG1nlZ+5zcHPke
ULPxTjON+nCiMoCz7lUpglTEjMkxG9N4C3y/88YkF8Q/xD8yR/moVr1A/9HFXl4yCTyfsH8q1NrL
5Nz1Z5deV7lN8Sey2hugeUgOGKNMK8G8g17eP07f0ldY3G+5+kufwVG8LheS2QatppOlihNQazNq
IZgSqKWRPX1UUeZhUhOwwdt4KTyh2B4w5dd3QFWtCP5Hz37UUyJPxloHIByYW+5PyksO94ZhD42U
YFXKYd7C+ZQqGLoxBB0WniJSReK5C2dF3Up5kIqbYf7OF4qQLV1pf61pVwFGhKKjGP0C11X0N8Ja
pLlwl5MvBCoYgwhBUCc9Po4SWIXcHyXnAAW4tPPZ4N3huM1zYshO4OgzaCM1H0fptDoUjnrA+JFO
KkPDLpHNjeyKFMdwbG6G3mmHhRk0btI+r9EkihnKdVYrzuKZCc4nqZm47hU9T0JvefD5rJtvTKmC
tcp2/pSjAmsCt7tmCxE+cjHPrkWfJfpHdp9ny8CCKtgn6oM4gvV9cz7xZse9SJ5+imzCxS2IzrWF
DLahOav+V6R13MUzTdy+UTsFbYGdw8t3MOgSzGHpQqj4gcSkVcovP9xIzgPgrQE4lc/olfWrs9LW
1x2i/BlLVzu1OQy1p8Ra/Q6kGgqaGI+4S5eLo0tafSTIf3N34peZNd00CNjiOAtG7ROfqIZJcUaa
2ks5d1O+oGimkkgnvWI9Zj9RIqUyp6BAcmgDpw7O6+UtMLNzenP/HCl62hxLkGTls+hFDr2YNLrU
tCu61iPDrfExamcnCmksFTjUd548yFX15LCzclbuDM42azpPKRMW0LhNGIHF6OnJH396EcDhdrSH
axH1o1s9ckBA+MraO66gwGmEmJMb2xzM8ayteu8T19EKw+B7HTEaGhpcuKMcB1JWy+glpcncHljr
qHfX7dF6opVtW3ZSshAQGLGTVFVNAL/bKyFU1oM0GnONFPhPzE6vF+8kBHjaGYEgeL1mt3Yjrbyg
H6Pw6JRTvbvb9ldvFqNRZ4L+T/D1zBUoXz06tzGlJ8S7Au59l9EBn9vyMysgOO0Ke9OrIp30MjVV
5GSs6YtLLFyaShJravCdy2DAanDd0bMdehwb7O7z4wAYYIc88ENm3T+t0VIXKo+6s9SDaaO0Q5BN
FOCmUTcBWYSKgzFJrliWyf53U8rBhWKralvGFgQ1tEstOljhZrw27E9ko9TQuKmGdH37AaSBbAq5
HII5buqp6iwD+LzNppWnDBPXFVXyKFm9GNQ3b8pkaMY+TRGTxnr0WCwl+EbU7jaWLv24horHoG6W
nDcLHX5Tkvw6KBk5AyT1TCDxRDSLnb6dq7/Lyg0bFYazEaUDgVcGy2GvyLKBRl+7tSQPbgt83qWC
SDyaagi0ETNknY1kqVBzo6TRQUK4w8Dpgvjcw0dfuxMSE2Zad79euDr1UlgRU63cMnl/eSzkh7XW
O/pk1CmA5+u3jwP8uHd16Mpjsn6+bkPM5CqozNbLUcOb/l9xj9MD5/ySeVpQrWrg9gbSEAf7hJqX
RRFYuuC1SXM46b7+UhCoAO5u+i8/kHqXwdU7wQedE3V9TDc+jUinp04ppN0AGeGjF1i8MTKY+kdz
GGJCYscNKrK9ApXVNURoPlXLUApkVlqm7KBZce8utk0yPnScJmKRFQhvy0O2a1VHVKinGQ1d+st0
k7sYaSIS7O8LXZAoEiOP41teqlgg1MISCVxG/8/cknJWLfeHZdqLC8v9c70EwQAC4uz8ABEthW7f
U2CqS/5oJovWwupvSEfYIfxjuhWDwr+YQlVOqd957P7Juh/+fBoksmCz28Rvl/yt0B8SDkIDxsHi
YJwAsXy7tLMkhjIYdrFOKJX6ULSB4jIN9WmspUPVwKdiywBXDtB9FUDXCbwkH5SArmvTgwJAjyX3
F9OX0/9svSKaDGy0HnV5gtdzUoXOU+ToNkeTijESsXovvjDc2G38LZK6XAcmZnxF7+ssC6SwCFiu
qVvslP4GxFvZT3TbJQzrTl3/+TYVxv/x/Xu6oMdU3jW9rnT2VfptgQtQBZVAmj7LfA8C8OgQaThn
+efH5WWjEjIEdiKt7DtCSt0/QwYmG5JSwX7BWRjghe095DQG0XhU0+lvE1qbta8KZIBAs6M1cC8L
BxpOwZcAEykHOxQsRgq1/TRvxxvjHx5X+puM5LgtDEKVemiQv0LOeJu8XUcoXmbMoxey6WZmvJDu
+dwEVHWk/wGZkhm2hDYxYlX0VT12jc2oYUXuPCwEmzWYUkP1XZqEOBDlMEjgzJ0e1krfe9XGFRp0
AMFUJrXlMhCAUqASN/SvgLcxKv+x7/leIHd35CXZBQiUVer2T8TKz/XYyNvlrrd7LvswbfvedCFV
GssGKc64/BHZd5IN8avY4EmAgNUeeo6iQwlB4CnN7ZDCCIzMFyU1mep/m9FaOgcz8to1tHXreqd7
dh3l3UwnxmP718M8HLFhOsmxwY3rKkyKHvva9wobOzGuAEbIPR5BciEUxEDFWOQFn6p+nxwFZ2wg
MvnlSrGh6vpIvtXMaYoYctCvnMPPWORRYntuXXnDxbuVoJFiuAmYlKmSrctv46I7brFnxiImLjzP
rQESFOFjtNtTBITdTzNJl7laTZybgklJ1SvO947Gs954jXj7vOlhoXS7ggNiSEOuH+Cb2GY4glPs
Dz+iChnsbr9wES2wPrGvewzDqC9LWcfWZzzxvByZZgogeaWBQRmgWAqbD4D5l+77oV152nTJDG9h
871MC5eMkV7cl79eKAhzvPjdlUpbx+i3fvexA8gO8KPPOfwVjM8kshMACS6LhRT2bhMMY3DClR2f
4Gi85LwtHkJ9QWBHl38Ccsc+G07Edl27yUJqn68tTmCU9Y4Vwzus1S7lqf7rUgXaKOqsaIdXBzp1
U+dqhi02J4eKb6p6PAl566+avqu3DRPs3cjHI8vf3bqUnqKugomXkX41HLoNanzxYEyU2gEiIppV
SIsJTzvwj65rYXEYjvis2RKJ2cqGPvslTUPwAYV9eWjvwca68X41K40vKc12nyzPBp5Cu7huPmPY
qsZwG4vNRsqF37UKokhiCYbmU/Nb94GoCDia9qkEPnJYjfVQ6/gZvxbyaYx9NU5ifrO3ANMHp4Cs
P3MieWvEkmHJkg4VxsdbtR8ae02A9B0+wfVbFGLqZTo/iU77vzFmfx6j8z3Rr8KnYOpdvh07xRAo
2VwiS2lMPt2dKkHeG18R+w3Spve0V/LCyKFqGiZbLoQyP23vtivjOxRmO2YzOgOcv1rjstSegOug
MvnIkSjYXt6jMCkFo8bft4qwNkXKUufruZACldkPrapwQY/+I27oxJUXdXJDZARDNTNpMRoN+ZxX
lYomkJoyrT9qWtO0itYQQVg6CSIfD5uIa63+59ge/O3OsYeeUOBjmUmnpcKpM5j8oDwVS+3vrZcs
fE2ntp7umHJf/95xc9UJ7/DrvQjIS2u8gZinpOZVSN7pdrPnWZuQHJV1aLnEDqy+WmKamBoXqh8Q
CgCJOnhvZ1NOuLP344y7XNlzVYpNpwxDRyf9DAzfLHYXZ3neGt5AqxCW2uwlZZ1zz1PDMHuB+s0I
VlvNkx2k+A58WVEVdS7ZMOMgLRLhCi8StnCADGfHGTcCllu8kJiJJaOemP7QHY8r090UkRZn8iqo
7ikVBBGrBfjTOSCF2I1XknI82CNdcAC3eyyAACRkdDO1EnYvj6Bo7M2tMu4QNViEecvlY8TzY8Rn
ckJo3b0PXIaTx90ATFnVh3JmK9hKONMpZccpi5lNkVkj5dAGwnw8Md9dt7OiEk+gqFd+UeQ3iXGl
vbGXjBgN3XJiFREh3zI/7paGV40+/z5li33OZDkwU1YXENs5ULGH9uu91aCsVPtXnaz4lSqH0bRB
3gD0Y2y89LiEKjkwljjTJh+derQipJt9+R7hjPU3FPGFVJc39IyfqeuHwz1KMu5bPAYo6l/X3Yog
CpTUQG+IbM3fItz98a0gvBzi4UCFJA+JSu1KQnjrlY72oT/sLltZYiW/ckxUKqKhHzhTSjxrm5Tk
Z9uKujDtOSC2YN7K16hYLxqe7UP9VxjsOoitEPqaLktURzUZYOB0qQHrICkHe7Rzk2fX4+BLeV1U
0b6SZvBejOCYbCM3q20aQ1QnmuVzsPqGsBu/Xv3ZEUpL2thS76lsFo5HfAuIsB84c00QzsT6axAi
NItSJn6/Ns6Uu51ltAipZPc0bYqPP7Tw7MVS659gaYX5z8RzsAyXxuVmew/GoqKfZP4B35W3uUgS
cGYP9fAQqj9zStmnVCOChdiHeTHFb3LLyOyM/Ba4DVcWn5GTagfwaCicg9iJjKu2NCAgWrz39huu
0lbwFczFJG2FFx3HO8L3ilAJq+isgy0bTF+nqb+4vBXOqAtlMcKL+gfmwoXh+uTevLBfUUL71ngj
kgirFHxilJRrDEewRB6dd6kg8Cc6yU7/Hd07+E2R06DIjzcZh4QI8YR/Zm3NzE8/SLEDS62hErc2
fDsxvk99nQuotDhO1bEN0HNsR4ZU/aBX2sNnpOs19sAEFbV2ehjHuMA9Mx29CURxCGmiwuy3bZxp
vJSvkbjjZtK7bu4n6LSaG+Qz6oBufR50yFMFCc2GVPR3bM23a6LIib43cGMGECYzLZjRT6mbdebu
vtuqVu8UNI09+iIPoxrJtAgyG+J/0eKPplXUiX+Ea8SarpFq5RdQGYbKGEFIh6RUMUkNsDqokb8P
PMMXLFVSehtoFEGX4AoiLYFeqm47hhk25S3hSLjebFrYcmRrKiVaHXzspvlCybQEQ1QNkFLY/x0e
yHA9uq7yxmUG0kWp0ixJLBoZTvs/R0LitdkgopNu2dQtzWVg0+g8919CiRpFkiRIj2jzX4inOu5i
mPblCnJT988w3vHvQpYUx8KhPOlp+hzK42egj61ulRnv7QeP/ODiGSlHIHYj492fgNdJN/FB2oko
AGA5B2YfWnqqOkrLx9b3Svo5c55ex0CkVP14/IN1BNNVS8n9ehWC1sdgUU94T6bWZA00s5nG4OCB
GcmbhvU6HcA0Butv91oe1f3o9oZAUw+isy3kI11N/inq7YJ2WH5NYZai93eaTDTb032nCCBwqbtx
Lw1x3HclJbGQphLIWzXv42Dh6Uc1CgtE5OGTCwE0Th5dU1WMYLBkfhf7LL/j/B4BgGuVlYr/dMVk
1A9rT8D8JJpKTX3KWY/UtV1EJXWAk0DRglJUY5EYAYrcYlXoMXWLYGYEGwrSzltZMjMcG71ZtNLS
yUfpAmVhCjE4Y+7c/z0fFa9/Ym4/fsbqj20bjDVhCB0HqSX4mxFIO2gJc2gXDoFJLGNhqqQHVqvZ
SQaRHTfFn9Gtr2PArJkbsQwu5GZga4dDzvpAn+ek8b3ufmrfY+or9tOtRbUB2puFyfcMZA9vwAAc
cBQBnW6ggj/N/RzN8igZl0AecrSBW4wdcrt/0+oF58tSj/tGcUPrmtYiY1kVs6pP8DS7FrCTMov8
uX/1DA4N+0cJH/DSrTn7qnw3fMfo0CARKVWtc2M5csgO+0w/uO+jAoLUbtnHsLmFvAMRDIfcUGot
of90Hvj0Aq1qlj2czptanvn5p5DaML1fDFgndw7nAj7IV4jX7phBmoBVwx4/gE0GhxHUAnIYdFE/
aCceFtS309Wvz/LspakYenx7bMaiAr092Yxfbly3zXmTZ2FVvAFQUCjiRyyPMeoaNzNQahH67BQQ
j2iSeWSQduFZkjNJD08Ogfi7AZt7Sk6XmTXpe6IKc5D6EIuMZM6wrS1g4LHARmdlgpMJLA19Aw7f
dXyNhSItrPbMlqTqo4P0GGVp9Gy5OMCzmbmBEZrliOveV+HZIJux6Evewzjtyev5MSSTschtTsB2
40od/BVoaSWjBlVbhuUrQJCrzisEb431HRKKL1zGn1iRkqkvm16Yqu9VBRJnuWW2DGXZKuNTrySz
HPYJyuRo3UJOBsFepJ5o4KCE9zhrzS7i4DHDxPN/DGTX6e0keaeCyQe5uKPQckLrS7lEjlXgI4EZ
/5GAjhTU5VFGlWKjv0hZg08RLE1ynwOl8KM3bDXDhCDlhdCd3cef1GZEd7PhyDigpaIIXnVmoWsR
2wkJojHSE7BTIFSqwG55oltOsTU5Tp8mGHTKZ+v66kRABPsNGs62w1zri+golKS/HZx7JNhBlKSR
w6Q8lgRVK5DHbhqE0Ml7fCikZLRoWkXOKKa1w5I1v0tFNOy/mgfcdxaY05EhBgPgHykGN6xBU8pf
I14iNSlKbmSYUpbsc9WMFr8gEzWlRtHKQZniawyyz4+BpcAOI0UAs+2vRz7aSvpPf1K4E0Jp2qG6
IJS+WMfoqNoC1r3afTuW7CLVhecXODfYZlIQFmvQ5psQPmyc6yYyeohRt57uQX6g5uspj9lOTsvp
d2/XDNNo7wqp4rUGPM/qlTeE4S6E4V2CSWxSoDQMRNFmm2rx0e5+TymUtrh02VBtjLYJzEOKpMx4
MIwsx9TXhzz6nC/AUchi9WHK2Np5hgSNyVkp0Zo4HQuqYt2hPnoXFVCLCkhmm2jlv8/ag0pXlx32
EBwCbOkdEDj8N/nWmnfh+iDl5KNJEmqaIrpH7sLqWSPteW6ssVGY7RFllyo8ry+R9HAVwFkTdoil
dAej01HMY9sC4MwtsmND/+yQ26wWNMNoE0/JrlBuA+xrpkoQOfGhajlgZkNjtmycUMFqONhAxs3Y
YoXsC22BUJrCwDtDYUkfci1NDf5oWNeVMkOOgPvAmNblhnp1C+Am48ciKOd30p1vCUvaFiw5DpfG
jtCVnEH9GeEXFgUR6iJX6hjKH9fCBloz9V8ggeSqsxvGxRczQJzO0hzaG7fE9icQ83Rguq8xVKGN
m4NtYB0PPqnIst3F20GQveWGkZp58ay7hvffD68/hnW10HnT1ZnppHz4M1zLl43PSLXdPuyS+x1C
0HCR6ENOuUKEjm5BgvaVmNvOaJ+Fryb7d5QkLRJY0IurjI/BAI12Fx++NKRAkl08IO9ZkvEqMS6P
RJMp9DpKelv4t2H01wfbSKLCwbpXYremv7m3NQeHmEwT0xbeb/4n2YoJpmSejNihy6hKtkaRNQbv
GD5ViV0/g8YPBBvT/9cH4rLRZC9F8Kt0pqrcrMm7RC3wyeQJIZVMgGHVcXqbF0L2jHyVqUJ+LLXt
QVYIKBApvjIOs7NucZzQOH6sXSc3sszm/PLQn4nCDIA1ADcxm8Ad1Ltj47DCdhUwjhyu5xGBcQSG
IAQ+IEZALvJMiIgkpxcj7jNncAOZ9EJFng/4IMA+cxEGo5PVGYvAGFqzDOvW3AuqqjN7R0lRFO4D
bcyhvXV7N29XIVl1yNnVVC6l0YbQXZ1FriwqVlSLxXuCstIgeg4XpeS/63FfcvgObKWY1BJO71NO
K92Ni5CFZ719rIL5rSdaXJO97Ns3lPVnEpCcz3hllZKbownY31GN+9qpf9EqOcvrA5k9o2E5SODc
dXAoLAZuRS9Sa2BQpmF65N4HzQT+UCGJkzJ/wI3+aU/YKzGHdG3bEpyvbsq6G0z2D2YSqyr77nXT
FlhYcz/X0lb8On7IiUObzdu4sVyjXDU4QRnZXv5xLrhqJcDh0mkyIOH3Zm7OOVX8RJ+E32q2G8J6
Wzyl7tk1mW0xF10yth/7wX4R5OIzf4s2ZeN5Bjf7Hj+J8yp2TapKCZs7561EQ8BbcEVVIj5XuYrj
89tvU6B2c6O/woCzxy3RC3gbo5WzBl8IzAm14473rSfbov2Hrs95REybG/bR+1Qxihn4XWY5K9HC
QrZeOlClmn0XyhHUU2/T1xDQeGO9OAbCZKG9HjlxSq6QoeKTRYqhs3QIE4nqmx5Ewf/RxKEb0W33
nEDj6p9ASWMHMf1NrJRcivIDkpyqMaisk2jTK9MnirD9vXBkkzYdIct4URs5+TRkR9qfE5Tim+ZT
8CDCYaxWc+AVVPHNOv/jo1x8+DJcaIS2Yh9jO0gdJre3D0oCd/nsUZLgOz2V8d64Zd2nrBqX79yU
sSOho4m1wLLcbyIsyhWQF9XWOSTu4lKxtFbDD9Y/U4tD0ww3rqiYwvP3TXrYQQ8w0n9W7ajsZ8Nd
xiXxwyWOdK0vU+FBpQMFuIcbkLfI8W/HKt5ezdDY46c09YL/RIFaQmWF49NRpVP4NwIrG+quZOn7
1F5BgfooVGXkE/AM7AC5UL7vcO5g5Wg9fkqjO81vyWkXUEt6n0CtxWklML9z07N9d+OWvAre34mA
MZ+xgycEc8JhTa8ui4iu+wV3Qj42BEdu7LTyp3TzSKNXUQ6YbG3AzsiieKRiN4os/LMo8pD+1dcd
Awi6o5lhIoEm4v5HkNoptN83SZYwnlDib6UERdvL20gUOtCMmLQbzuG4NIWSuUj5pw8fpvqseOOp
Vx8fy1vA24JSmHTE5O7abyhk8nypL8K4F4d+a+sn5yzMwyqSVT3CO+kHsM1xQiO54pmGQQkYD55w
q/Ndwg5PPKw4zyL3qZnm9xiLB/Qx52UXK52JX5+CU4F8HBE33aESsAU+J9tF7YIZHyDMUHTUli03
qLdB4KnWNjU/yNi+h9dqEdBjmjlMK9AtorcrUYL5XrI+Ban9mfAP+SPsBXgT4SVbTPZIpIy/aYw8
6uZQGF5R6ZKSOOHgA/U5lncQlQJ/Z1MjSM+hv+pQNAndYTOu0hKDU3gb/UB8e5BiLLNDA6F2n7Fx
simExozUMQV44VVSc7ShwjaSBIfUWOU4LN4KPqpWZXfDt+H/Y11EB3OaVr8C0KZnV2dmDjWiOA7J
8no4KtMjH3ZGDou9Dt8m6rG6TVOPNniXcysH5u7/LD4EhunviC3u9mIrEUNkCEnXDDwr0RSrzrOV
yxSUTCN+UIC/S2BWIESOBrJVBCVlnwcO3nm7d21XOLvvB/wvTPQbTtwYmJwTJCNmuYT/xKnlO7ij
04tPdk0+L9KXjbc8ZQZ6WVPlG3twQQyQOfqDdLfEN6OzSR2yyMxwV1saXI3vYjgsLhq0JvxqqOCU
FA+PQO0sZ/v9lNt3InpJ9Dky+0AM2XHobOCh/8Mll/lETgsd9cBNaRI3wh2LFilZrXqK7HrW6Uem
AQ4xbliCNmLOhavliqQFj/VkYrg1iIOjDixvrNb6Jp0d1izDvaxpIUsF5+PTCAzo/htutms5ejmw
zguNR8rCH0pjF3rJAjEg6dqjlhx4DJPSNAmtwZQAOL551brnoSz/D9cmMZrSYWzTPAvyQPqq7I5P
QMY129ZeBDiYSxVjvXLIMXRA6Q53Nz6JMu6pNmSP4pyDuERXkdHzutmFAsjyHYWk5R47hn1sOxgT
KbVhh7u9heJs0ItSsWTeKIIyW4rirgnc3BKuGgxiR819rxXbbfQqqojNwP3P+4sFPABygiXeB91x
858Hxsd5yUc05QpA6cuBYZy077yclCU6sOfiVN838B0flN09pjXBDcDmv8MsKfXIyMNKHN/iA4oS
9cd0eSolMfl9UlsdMi8CbhEjIOmyZaE4T3s7au7woxsDuNLENo9LygYGiw4RWT2t8/DKB/guyqDK
jt4m0/nKYkwUk6MCRru8xAl82bw6Q7aV89dvepOf6iGP9Be3Jr7UY9BZeSo/MxQQK5akg1i6gnJE
HuOvd6HMr8u+80JjSATB/rvtA0RXms50BF+ce+LPH6IqFG1+8B4WcV8FRniVgx61yuXmNoKrOA1+
VlqLcRqhSKoyWNwywjkO2K7s654Rsu3eppEkvUtCJBpm3A3IWiZ3lFq8+mqn79dPEkK72Q00Knzj
Uuc1K13txi3KKuPk1VIPgwNfnjLdSn4rMr97OOUbo5oTG1lCdk6I/46jLOF9j06BvSoXLvN9WnUH
tEN8XuaPFGY2u2xmBch50Oc6BXRJUApsieCx2aqgn0FvVcO7bAa2u8qkqF51Yw0FY2WWgxGblWez
7GLE/ArQlYMDV6Nph/au3/4orD2u9MI+j5+BABVlX9fj3cIK7pfhZsLLVCiWNjUKpEalRVUZsAjQ
ddTr8wa3K3kx+6cJAunhdXlXN/N0Euw52/zgrRdMtb8oaPtA7jL5zaNWYfbe3L2gxiRRHqLLPuo/
lqNEbUJNPtPcNKQau1rPd77Sp+r9QjO+c8RwP8VFHGxOf/lHWLn3NdcxjXOubPOHF5G6TqGT8LnT
E9Nf/jPDI+lJOBmVWnPW5phIl8AtWYm2W8mjGSpPprVL+RCeJJXMmUAwl3ZR3IJy85S9U9vGFwWp
mJduN4h88qDfetPTszdVKdPVfplLN93iBWKK70HoFDykdOtBXTCvk2DtBv+hAV2zwVNc8gqQlmgO
Tx8PN2YIM9fyvlsnPTti2Oqgy8Sdx2dYtnP57j5mYkoaFVVeAwirS3MQoxEEe6gPoBEpbYoBK1uK
/oz+egn2Pi1QkmhhF2UfYi2iJM7wu2doHfu9Knt0giJbJsA0gkTFJ1dO6icP+ALhx9cWc4zmDYOY
KnY/yh/pwbro4spd2fs5nKPOcuB6mRTkXgZghT8gwqmIvWqSjFKcxdtfkSDamKPBvXBnJloCoewr
GqU53X3cE/lSFEDXmyGYO/81y/L6FaDqiYMLizXllS5mcfTTUUaYuTTQbhUitUBlI+NSIcTVqG3M
nfL5S2JJz9oXdOF+ctDgHQj8a3WnPjaN2itdMYZ1HgoQFEeZ9tfqGLNNUKtCoqv2e8hLow70fSHz
9GATzHgAbNzgigK6x6jVljdOWls6oNYouY//ixWFAVattMIHZRLblnnaAguFLd6B2GCBUhXSPEOh
E9xMZRyXGUEUltJ44aj2LhSKy0rVrb8Nc6oB5INTpl/uPA++8l2B3FIu9aUJ4FSj3WJBb396rUuy
LypNMpm9GV4C8vISAPDlLfjeDqeEHQwAPwmh/yE70hZP4dgF4tNN0b2je9inPzdhyoRlpz2tI4Ry
WvC1xVoSVPBQEYGwnSj1TK2IcOmh98R/+eSyAsGKgwS8TUu9EUP7d8KnPzBA1x4tDOSLfDN3BK7x
JY2teAPNspec8K2HT7wh6IJrtwoTsMF2Od5fC01/1OEtXgfnDyACN1FNLJp8lMdhuc/KKNYbGyTr
J+/KAoJ/VxIWTDNBEzy/kw7P1l43sbpViC7hCQ6tayp+9nisSReS/BeKNdOYMn8ObGpHfvPbx/eK
2lD9xzYwUHkW+WZAjsTq/glwFuovJx9VCIiXT7Z8tk3swmd7nG/n5VpTbO5UmYcG3IdI+fahOcb4
wjzI7CnSO0yQb9Wgy/xAQSUUajC7f4FnXEzlfGRQpTGqaKnQagafMbcyGNEodTseROMV4AjmN/bv
M2aDnzUVS1fSrumXdIUVh+jf89ozjeDZ/dQvNs10xgBPKq7v7Qx8xRNy6DgJvC4mZFBMNtoU0ko+
Ti+MRUvEFaxVdrkiSuQO+reLDMzRCx9DqGks/55+CiYJXGRC9NuWOnPSUC09QRia8di6eSgG4esz
6iNJPQKBHTrtnSVRdqX54Tv+ZZFeBUTEBTWhtGtN2RoZYng7ZP+IlyAuKJYJ292p4tlkL82X+5XW
9PkEPFCobt5qDj37mdIflwo5hNz3Ng9Srqhf3iHK+1J1gDr35dDKvZWrbJ26z66DxJTyTFXg9RtW
PuiWOIqBNY6JrUG/zW2fUpLoLy7sbaoFLvIkqI9vRX4hajTBCeSVMdSSZ6fmJwDSn+3bu8rP8f0w
HSKfwAqBP5iVpb6/OVT4E8Wt2tuYB2EKI3te/14JUInOgFZ8irf6sl5CkoHxyQKq2ZkfbdpfkOMk
GMLdBB3SkO1r9kFdn4t30sZuSwqs/jyxspk5YG5NQ1TPYOwtyzEWO6w+cQupZhXJr7L+QqJzk4s4
5onUY3dfU46CgOpZp6IHS6u96rG/XQRSlF0pmBqvoEzS+yjVNiEtUBU+Q93C1OPs6/erxemBiT75
r6Jm4cBOYW5VV/SkbKMKnlxBd5gM180YUV1KH/YOoSTeU8W3SZNrSjUzaOWLRxxMwtW7427niegv
5tmcTu9epT+2tWkbofNG8JArQi3pUm/vCmpXDQB0TAwP01Ot5/awkxt+RnN2b2XvZp/7AfudbgD/
Eo7NIhmZxx3rFImpfXsfQAtZkYeuNc//WuikZb7cUB/yfvOKkprys5YEjN0rI6lHJQNrInW5jjKi
Qwuz0CbZk8cTQrOcGPgMS/4rtgQv+OIjYzo+7939wU8UuruR25xBlDzg3cSHdOTz4lm30GF1wKSD
/DyUFA1kSkE5rPbYMpXtgg0aRg5dfPkJD7ejm1yf9g7Rcdjpg8AUQimSpdcvBkgyMUMyBPnrAbou
MIqwnsotCznwcL2bRqIQHlOBzYD6KXG4v5IOMFY7GSHZhq0KMV4C225ykoJ4Sj19NB7Z/Gs6d0PS
dVl6r/yf6VrCWx2RfteHzvHIerN+RCSYIKv6GmJY1Z0wW5Fdsv96uN2nnUq3aN2IRUImnFO5DV2m
xmUA+yPahda+TJfmN8ia8owrMaNP+pbyktGj7iUF9kydTv9lTAd7BFu1p8TxYxEa/Mt0vWBJ2VNq
AJKJKZk3Us5bC4whHcdJkhcreamD+o6+tZg6vpoBSTo1Cm3NQFsrsrmxHncney0F2C/0cRv6utQz
J50+RkjaCyLJ2nd0rJyiJABS8FuHo+26N7dQjO3X8wxP9Bo0n6ajhgMajQ9GNow/bPcOitefHZIt
IgG73r/fZ9jF5QLIwFaaZ2jv/aEkgpudWHYDk1TmA5x3PSyfP88TZltfB+U1DPucllrlZvWxIaNM
+JNAcgg7GPUQfgGpn4rpJaS9V1/RfItUCDph0iB+B5bySq087D16PBB8CYOdFFU3Ugba8XQn4Sc0
/Au2OG0usdDpstA3IgAJt84jaPUQ18x9XWW9aVLFu8YhmZPggWwaquWgOAG1iUs9C6wX4cbVLYFG
Oser8hTpZqHbPe2icV2PPZNI9AItqr7qfKtWs9WUAcH7RmxIqGY7bYsOqtjfyMnsz/jKRDnjMswX
wLVy+1LbGCUG7xol9339ouQZukrSXLn6Rkg6FjLP+q5DBwH6vh6U6jbzJyP0UiyjjFRALCi3XZhh
Ji+0JmwBXKPcUfHslAUa9UwOHnVM+gpZq3TkssbfKxiFucHcpum9ff/WbripEOayJ7ziu1tDO1+N
Mz+AQvfhpb69957n4F9eChpSCDcJ1L4ar8mWA3wKDPA14ZQEOq3rsrgfB2ewFOp7HxEjlTN0IWfU
g0Fnz+ohR4+yIqQVQhpsbSUEMc9RjukI8X4O4DVaUOZ0NAKNKSNRo4MnBD2rwXvq2dSwgv1TqTYM
nE/LPb3kqe6UDOb+FdlACC+wOF0cbkCeYYHnOKV8tL1DLC2eMiun4wr8I0MbwfA81GPxllZY4ql4
awFOaU5+4lMIDLuwykPKEvq6jyLd1FJd3EjGvvdZL952CSoCzq/PXw8apb/M2cLp9cvfJamnHeQK
PJli0OJMS9z0ASORiTRMldUA9PGpCSHd3b6qprq6k/kMZ79WLeRLFweIcHwsy6I5wwufpsA+UvCG
7hNfjD4mZrAGHpmWircM12N4TgkVBe33ah5tCXfsPILDlhzmtA0cgykBhnn+4+I8eHGUFeoQc6Y0
JCQY+lvvsBTOEevbRngYeorOdrU1B1XPOqjuzgx57F7XAEa/CCx1uxphJ4eeLzT0nsg6NSGS8lwB
yArFSOQKNa0vGrad2+afU5mQdS1i+wfEPtZhYurYQHVFcg+lty+kfuc7PqyqSx1SyoI291Krt7U+
WPOxjz21dUMO3ISvfahyDZloeLrf5CvlNH24+RS2/LfjI2kK3WSIX1q8eF0fIlKC1d6RVbBBQmR8
/4InhJM4/dbkFR+ixeJb+UwE7m6BN6SS/Jyk5i4cLvEWuGRasJS4Y/OTenF/epkci683RhPH9fzQ
D1e9IUQ7v12Jp8vllDKHQiKWe6NlNmZ6dB/86gI5mzkho7LHWE9B+6xEN08TD/qAnmT4E9nU2C9h
7K7QnMxD65TuWzjcb6Wob26a2bJoSBTGK1KGYrEI42nlkQapVAnz9pkrxEfvrXCNjTWDXa/NrNVj
p+ByFoxkHR04WUEB8UCQSbRdYzRsY5QD7dweAFQ7l7Ien9ULUworpkhEzN1kTYwxc8f5u87EQkhc
i482lKkSz9vKUIxymCykrQcwNoMwU4H6qgWeP/O7x9CQD9D16ILn4O0uVLHytqFOVA8Rg4Isg8yZ
Th2fgnwGp/W4x4BIjQWCQAz7EVd76CT7Ca0C9TbOv1bQ8ucYLhEGUBQT6gMActgOM5nx+K8I/jnC
pEea5MKscfWWMWUHrimqPXkJ8NqFAnpbsY3qbrj+w5vc3jblIe9M9+dG1umuU51fOj9fizT+b50v
X9Abfu/yQAkmppUwbgJebgYkzFjGmBNbLZ1AoFo72MG5wrq2P4e9g5uKF5v8OpRx45gee9ra7Sm9
43xluStoDZkrgDLpTcKjmvhKrk4yEArE0Js1r4vPI6jmmUvXubWNKfulTyCHsAwRVg7tDmixv23a
FyxXdzqy9dWBG6XlgesteZyIXJD2X34vkqKhYmC7Mo8nWzqUD4qAdvsSa75ab4JPMKUQh4jc5zRE
ZHhR3ZYbFQNeWuVyhdUU561zkWc+M4aAwY1ki0ngjVYd+FoDrDAhDix70k03DJGf7R4S5XFOgCsg
Zaw0sYph/eWwuRJ4fcgUUKMQlovtejhDMHOKk52raAa/8/Vip8889DlgCMp7QJUqtZtkZPq0i/Lu
brpduTRbwSkYR/UHahzI+N9XnEPnVY+wvOmMcyzZPWu3VxCwNBmn3xITHmWTBrYkGo03I2RhQBfr
n6vmWW1YTwVIlnapqvYWyhFxETFdn1JHrpM5SLPL76R9cAt/iKWlBz3LHvUVEwDhd9dx0KjwwtLA
zNhY48qcCWzAK9in1kces5Gg/mT2pDcaqHFCuKdlLLWchjbsTAVdtAy+Qujsyx5zs6HXWwHnhj3a
IY72hcvaGa2fMKh86jhpeQU6wipItvCdDke/X0wQOeSLCoeBfZcHVVrnIj7XilVzZODcJ1gcWEZ7
qcl2k6yZ2vnu07emmOTtzLW9Hh+bL+/QUgjvbMPaHRu9mOEWMjqfxOqkuL4RMBWSw01/Cq2l+Z75
ep0PZcQs88dcnIbiVhcDBglJLsraZqQsd8WxWnBBDi+oxo0igkVHzapf0Mh8VEUp7LSfgqlBqsfN
hM7CuuPhXGLKe5YV52dZNmd1ntDfkPD2jA2M3UT8OS+PPigHqKqxxyu3btq8KvcqkftR9GDvbJhX
KgDMjPkuYoxxEkc9o3HmFaSmKDjUVNoDy3PcnjqeMO2Wfk6BcI3DTv2l0foZF0jJMovm26/TZ6NU
4Og9a4wPS7fKhH/xKobxDGZtFTUmXbMlHGOCijvQNn/PhC8vflJnuuPk0EbRW6unWia12jTumZCg
oseRG7ObyNGkX54pNth9uvJ5G4x/s5jAGgA5ZJDzRV0OYRQaz5HezWBfemJdkY5cI14VjxqDcy7m
rVIRyLNyH9pe2m4nQXmqE6FJNZG7MR5ZBem6G6HJZXD/xdYlReFsANhjdS/rYXWHuOr2xrjn7hZI
vA5rAb+AZvcgFAULw07zUorW8ydzByFF8FnD4VyPxvJQ0VHJ7Y7pxE2d2Dnp+iRvIsMT0G2BxfPh
hnReIDdPEVPYJlSAtMr2rdnIPJ/hyJV7vs95Q04SAalpLtq4XleO2WXUt7xj/+aQIhUE35URWEdQ
DW/e+/2uGaCW9ZmvWLOdvEexi8given6kwMLjpvzZgG2QvTUZULiQYlWv9TfSuxhwVqP9dAYisnw
YMg3GuiM02ElX6YVfwcgL+k0VwVrJDqmGklbRhhH0OW1LPpmdc4NwESPgfUP1ddFH0aBVtqrHHSY
HSmgDUc0OB9BYJvHFxkbd1raib7mwf2TIof5ehq9AXPZc09BmoKg+tb8oTcUnlITfoWAaNTpyMcI
fEno7ZUXKpdfuZ0nZYGq2YeddmPePkC2za+HT7GkphBatpGcDsE/57jYvgYKjzA8rgv17JeITkPy
Fny4tUdRBmxXX8wEDBHTo1DTPy4925KP0/HXDt0Vfn1aI8zNUaZGYoXISkC9oPLaNXfGbyg/859V
assyLwP9S4OHQSn7P/Hq5HSnEVvEhDP/XydKGx+HlpNsec1zMiEq1APEnmaf8VKQz3mGojjiAKGE
bEtbRw9IPIbCP+GhZrUfyyISMIpw0i8uDmtk46BNan/m9UNgKECJEBpYgCQy7Ri6nHpP3jO3f4Dq
5B0ZN8Cg2q3XEoafHGJIVuxsRK7wM9VF2o5aTaZKFE4CayjPuye3ftWBawhtkjuLdOZ97PJJ/+T2
7PsEAk9onAifxDe12KppboreiX2Nxp7OJSxfMVDXSSn9zjWNFJKN7VXlNxZYfMv7whz3sz97u/AJ
ZU5asf5HY+zh9nUBqwzD9z/C5R4OsIXPj5tcXXmzx2SY2CPPYVamMsVuxMnV5x2ngQSHzER/sapk
qfwHCZsmw3jloO+UnSFpcb52emLcxXjwzaXNiTOiIHpI49CvxgVMGUW5LJ9EesG5obaplm2IK1dd
yxEQQEhFy/TotcgLR3EjuE2yIivX2ZMPfgJjVawztM973qWou/cVcydDiCKBnklxQI6Lu0VbRfPZ
Sdr4PoIWshfOdq+3NWakNeCfkO4ZXxoOUhABaDp9CRYIhN4nL/8FdhUGknRTchNPbHhSukLKkc/1
EqVsv4Q4PGCeji4WUNfa1kpHh9HnqpXvHMM2zsAlP5H9kiNKDDURn1ibcbRaWsuxhxGHVMsY8wYo
agS9TGmYbI3P/ABFxcjlIWpQXN0585uNLE1Vs3HKUqVeiu+/yXuyJUs95jHcjnVS89sKSMFzXS+D
mpm/150Kqaww1YW/Qup+wzKhe4bT2QnaTwm1zndosTKQPEHI4/WXl3up79Bxp2HgaVFKImhGxkRA
nb2f67bRoostaOdg8fboIHDS9PyJo1xWASoUJJNFSxz9/48brKEqvY+9fymAKhhHchPSs8wCvtnE
k90hbRGhfWQsQF/tFI9Qf1F6gx/AKQNGSfak/K0KRJZsJiJqraXMWYuG520mLZ9VPP/m0MmY3FDq
avOUXxaxMLceK00mbeorq4aXyJM4Y27DSK8Wx+hbW+D6nmHzze7O8naMQrhxXH72PM0T+1rk+ncd
EDmplR1wx7zpNkm83ydTo4wViFwmYMA5dJEJCrJN4wxaxukk2n+adLDCsMyg3PCsm28fNE/Nl6ew
fnfyykyaglqHzO08a2dL1COsrHkcDLOF7C4VUvINmYxKbw+FRex/5GIEC/X6lCMOG2pCNxuNpMjl
3JHz040lJq5mGH37B0dPRGH7bkrh5ee9rp5babsxSIiYGQTwv8MFNNkmmPomS7xyYSH7tnO8VRWM
6WbmuZ7vnnSvBgxP82X9tsZwlrrZ3F4UevhRKYd/RC5gCSvPX/AaS1fpmVC16AX8CfS+bY/dUKpz
ikhSfhlBZRU663aCibA/YR2lI5v6aeHCp159S5n5DCTX0sgYDtT37KjY4NXBzyegabDbqBEs4NDn
Qc9hGQXkOFDhkEQa6cYRMyfy99D+ex8RW8bUZsYRnu77JA/OLtRTmOXjhP4jIStDBwGBr672YZhI
Tr0M+XXAEhkJDv22O/HX/oXOiVSh09SEQro2lGGbKtzKTQbEs+QCfKFR0EL4tLlVuQSlwCC70bId
VxBKCPIX+z6qAuP6Dnu5y1S+4gjv7jvQ/AwAvLLPqQSWegCh0sKkPDCLoLVaO3q3oAF3SwN3lLVs
lKhVAJfeqz0ITahtLxnT70fZmyGt0RzVjGxEVSe+O8DNXbnVml/KhhKbBsSrKfDbhj9PSqy7YMQi
X0xdjkSEj0EkMo78qC6H3kgd/6NwiBdYr+qH/Bz9GbfEjmDbMSVL6Bl0c13TkEYYw4M2AmtL2ZF/
mVDmAjy5Y9969SIo9MXZ5uwBTJX1Y/WtIUf8KVzL8Y9qEAmyDfezeuBNCemoHUkhusjQuP7dgCam
qHz6p0w2V/gFOq9gb0rqMfj2lv/SVgt8U7qGfssj/lgtefCWp5n9e7NeCmK8pyVjn+gz3YbwfwLF
aGR5vXLWfQwI2NF2d719SZ1cWWFdYNeL6x10p8HRlfcwIo5UfIwixG6ny5zSkyFX+Xr+xZ+b7ibr
Xov1t0c0pyXeajcBHNhE2OsQHkcUU/ESTSihuPkhZbfkt7VIvSna1ZZysQD7etjloAU6LmWt/w3p
fKe3y80tsaUVTr0hE4WKw8yH0clH0pcrqCtPczvqZYnvx4jx6lqIPbbX4CzgmySvKpzThc/bLGYg
qQdwJC65DIP/axPgHBAMfMAX/13hFV26hW+yAKjK+rx1+fJtMAz0XWzevYeVoCNo0RBFWnQdWriU
NBNCu2FZADYeH1tc+j1sFQhRoTJdhvdHJxMTOcsfenkWrJELmEpD1RalNxnzj2AtpyTYGWNQJCEb
Fzj2C7cNa84KZtArJdjCYhHgDaYG6xTMiAzeUdhtVlIBT6+PqP3DiF4uvMcRzrhgyXhJm9qwVmzs
tp+N/JOz8HhQzwE92L8GvHRk1S/vJQ7mseyJ6KAVMJ/pTmJa89KsEQQ/uq8Vgu/G7/NCdZusmsxs
zRviSHqt5+hvmNN+hV90TEEBWt7QNePJebhxC0hCDv9AXN8tz5FNOvKLoYmazZua1oyJOXPsGOOA
qwfCA5P9sLxB1oK0DshF8EuUPkD/E8zEypZ1AIpBZurVwIYGc4xuSG6zBtan8trOps/r00p/OufF
aJOQeHB+5ZVjoD+AbNhsLiYq1XNQ1nLKwdZhBou5E7WVV1qDpU1ojLaCv1Kwz0Akt8kkQ5oljpX7
Q/hX+FLU2/iG23ypGAK7HJTpBT+GnDBQzhSZaZQQ4MHCfIPTZuKiEw4yFIS+EQZcr7vYflw6xYQE
d3TzuFyDedsJV7eEa2s6/VlRm7ZnnOfl0lNsPKKMH2uPv6B1e3T60LMZQA3Rl/pJCsBBbrOMB6fv
Z8jJAmrO3zJxwQlGyNHzccIYNi79Szk41XT635wZOoGXB/U8yCTqX/sC5etwtWHEEf2S2eu7qTEq
xVSXw6/TbfCJJymWHy/qe1+XvJUbr/ot42awfTzp2EflpyyQ+CfY+L9ztJdvJhr3ziXYHau3t/gg
j7VldBSm/4T4QR+1QyGaAQO4nHc/Bw7OlEFkeiC0AkS13n43yiK/oz09Cd+8FhSDoXm/OrMzFFBw
P4Ctlmb7YJtsmguQSLhNTFiRG9J/vj8a6cNjerf9jBGKOuDmEpHqmqH4OvxBWv0Q9kkHZATXqObQ
WmZ5j05zMtvqycosEQTUBXXR0Jart3e5dfurykSBPm0H8j9y5bjBoEdKVE2Ev4EC4ks7uthKYJP6
lsMms0tbIKzVFPCo+nyrE+ec8+5YjWuextNBv5Tfiq3johgMzx/P8kgRq2OESRhp7baQIWNBxNg0
e8LAYEbCHr072TmHC9Hmd/nXjmKqbT+LGfbT98Yq9QXTz0HDncdAS436WByLbK3C/CsyXyWIg0Xf
LMZ4O7xRaXj+GkVzq0391J6e8fl46XTOuZ4BeqrxMIrWMe5gNFMCAzC66zr80y4dexaKS8wNv1sW
IM1dkckcu9zE8Y5Xnd3CMsogpqRFzu7qhmqmW0f5jVSiFQM6eSISTexCYrlvqf0CMCsKsTD02mKv
wcsiw74C/nJMhK4+Um/QrE5agc76alKYDbM/x6qyxD5YXcpopdzwn3k0+52Q1mbNOOV/xJ10m+W/
e7UuPaSFE8eqylLInRTOZ1emrtt6rca+/9O+YBm3AjfvExnqspT6fc4UiJ0mgaEjrqbIdRuvKj5D
SrO3UxLGoaf+1Nu9mmY4e1JSIUq7SCwjhkovgSNT6lqWcdxkiuMlkOX/ECTFeG4FtuDxeavWzuiE
4ZLt2qwxjt3dWRKyRhfnenAXceLQZi2/E10eyNSJvxyQGUCbJIyj8WwwZemcAHqTky1PGtwfzwVd
Ye63+lgLOKmlWuuFDQQ3hE0bEHIBb/Ua3s5EfaLG38i5c+8Wd4myx8VpW/2OlMoD8kN3fmCxa4Zd
ZcSxVHUpNfHSZD8IsGbhaWtHrHloEgIvSXNkZ91XLDYgYck6qeF/DUQN3agiO6b1haGIzL9yNiY9
KgUkwJPSz1E/PeXpVHHD6Q85HxiDbSaCGwUx/NcG6eKL2IpQZUGdtlLZXz19QMdKnCwF7ze15raI
iDZvYBwqvRLB8GXwea7ZUZiX1z9RcmReBS/IWNaLjbKOWbGbOhInHcNjCiF3ss/UldlPRvmswsuK
8oY862bSc2xArTDmbxq0rirjzBi3kYBtXFtw3etbtIZ/djFoUEes738odwEyPzzHsSJG0IzLoBUp
F/k8gr6Md/6UcCAK4K1i32wS6HPW5Zq9YCEqQmhZ/dlGxHEkb4ezMpDihI+Ee9H/hYE4oh3Za93O
SSf6tfrM9sMs13UFruzsL21bsl2JVccVAc9sE+Qw3CZ/HEP5AnlVIRs3BZUMZ1QJYFsAIQoDmxJE
ND/Wh9IXKl9Q09cerw6Vsi+shlC7ERDO6rtVqDSAyT8jbK3pyFELzLTms8cVvCnTRTiKjzVr1gtZ
XMJo5eABHzM2/AJtDku7Tuv9E+yixlvWDTVGLBbwbGTtMnWApEnvcSiImk1z6URp22/oAKVPzcF4
y8aam94C+GFr6QBgzt2Yp3Pdv8DoVDOVjnjPexIrdDNQJyufEFc9wfDOGthA26/lIXROGqowp9M1
v66xHLf33m5Ni70W+12L+e07a+pa93OBB0Uf2FEnsaVcJO8nCFoGtsuFTKaa39//MkobdBbJNhsH
p1vF23VgA1QQD/Q+rodjPQ7Xrg/ckMLzgyzYiYtq2xCyF98NyTCmViVnB3oizmJQCGTmCVJERb6o
s+UHv7vX39HDdn8lp/FhsFizoR+twWc2IOAazSiF6/DolExGH4yYpM2iug34n/TutNXpcQn2unBM
TLaoE0IprTwINVt2Cc6yjlR/bCk/QwZkrsDihZkBiDFnVtjLYRQJkh5anVXDtXQFWjGb8ixLTpgK
pKv/LhwxkIWApW/9/TVvKATzN5g1KjA8VZv+TGjH0HUKE34Uescdw8K/dn8ip+eK2UvvMZT37X9W
IVVjDGKeGqnHzjp88t7dMt1vKrjFPRshG7T8AiB0i4nYA67/uOThItH13q3YQaLbaeDLlguW2Cca
jB+3E7IcjnECcm7Pb2pNUk0LGB1v4V6c1P4Ko0dZLKP+yTzQ+dMjBExyl+oHWDZ8b9J2axTxLrXd
tylLQg4Y2tqVmnKeq3Y16pM4nl+F+cLh0mHmgT9BUZUpzndR7D/J7L2sQOgYyKdHzBMyXWZ9PYD3
V/FrP5+xZF/PcJ3P3lzjBcFneKmIou0Ee9AJ0bk64xKnBPWHvIbg6YLw5UuiS8E1SbCJ6HIMAZui
DVwJTNM9zHGg7d/ASbzmoxP4QjAS28htmuKDbfHHen/ufXoKI/Kaq42hGGQgTz7B9ZQ+dABoRNvm
3ozLbdnQylsQzbMvJcA1gk4PHoAEvj0GM5RC5E+GIqL3/HyyacgArGA0+uLg0fk7zWCJjii6I6f7
UNFPfTt6me9Ua0vlPgI0vDEKSyaVqUSOQYeZtkduSGuZL7TvaJwBUudjg4R7weKhoSr7Xlk5G+up
BP6j7KM/v6Ht8muQCeZ+RxnK4LqMonP/0Ec/MRTw+1A1r6E5wkYJLD7IjLTowFvt6AUz6XXzzYOd
5Zi18twAKSSmZCnwj2C4ptV1kAoJjWi7M56kLIAOE6vgv1wtwsq2CWlXTFqq13xsaD3bWlWScCx6
cs3K3In2dQu9GQ5mzLiGI76fhXoxb3+oIGooNzFlNGZzHmtU7MerWKTIgOctQi3fQUFpKnwJuz56
0NliHGUPjpBgeQMO8oDgenE/gx9vbXYiaNSsX5z8QhZdDi4KYg6ZHtL69L0EogxAEXPneTi6krBF
DUavte8E1e0KRl/M9QLVnhozvVtr4rD+I/RoJtv8xo774a3nlh1p7pHa/aItPRADOem/1t+C6/4F
tJBzSzMoBhfeLuv3NYEqQvm878F1hqI2CfVUgTn/AHjRo2NyulOcOir7qzRMb9oMJ3p2gtJaHmYh
rcYT2glFGHl8NXEE7lx8rlORfoKSUulR0mQfCH5R3gO3dczWnXC+USc28IPfq4h7xz8bC7Vu9ciT
uxropC1FVp83GbexwBFx1MfLJ7zeQaqIsOAonTZpWzrJukGe6iPhYHeYi0TwAM3kx4eZV2YYycyg
WyFWZcsPuXwzEdnGGkL/41O35B3Cbn1NRELpHZ0Kx9W3DFUc6FQpZjTt54BcWmTD2/asoQ+wiCzY
cl3BWEMJ4x7FnuUv1g4J3g6u8lnTr1Pr1M+T8cbemInT/FMALCh6zzoP0HwsJRtR4A1F8kgLCsHr
qQeMpL5TKbowx0LJrDuJmgj17J/zpu3F4ZhcPjtysKh2XTocgx8c1bheYSspvG5hL9wsxLYbgxoM
kXCmUW6Vj34jpPdj4E1H7gy+zWMl8HirFdcY+pqXXN//SXCrc3JCFK9oVjp8N+bI4ipPnqclLtMz
4C2o2DGauAjkRbBHOjMrCIKDMU244jdyPEBogAWCnz0/mFLI77dakxYPn4sHUx1JqIVV3k/0NQJv
TuegZP9L/rmXwsPHywvRi+xkW/kbt4zEVSw0y4tTdTM3Zm6376luId8WLBXRGPSNZIkNNLVaNGT9
xUnBpeDTIeks4PFp8NyYSlleh5pg1C2XJwuSBZBuMIKP6V33qgzQqnu4pWlSqZEBpsTocc02YiNH
6zgTBvxUpTpkaFPe8WpAQlLnEEcgFVnok6nWIh3S4Vje2G14p5byyCyypKyTjxdBDT6gNU3o0Bqa
ywx5xosC5UCrZSmGWh0ey/aDkY1q1CrdMWD8ixWvsSoZHWn92aAWS+mqFsY+wIQA3qpii/7Lviad
aE4SHOl+/y/PJ23v/YnEjUHqsDB0py2sUx592pAs8V4Eu6aWbqHkFknjCAMOATZpFpoPB8T0POj0
uMda1IAKU40Sw4c30FvhVmsYattqBvb/uFS0Aa9K+JZvUWm4Oj0S6jQjYRu5GaWFhyJ8C1nL3zOR
gwU9ryCSqeRKLsbsYYBwd6V06TE2oHDD4cM/O8byvz9+iYwzxHoGzGuzKPW968vJUunrL91Yy0l3
tI9Hte0PhKSLE7P1sAEOJcDu54ocuPopMW1C/b5nOzf9IpTLWXEOz9qYaO1n+lOcyQRXbs9DDa1c
H65B3wxidwqpb3jrXRLYjFArpG6d5GWJVTsy1tb+q0b5AVod0EcurjyQCUWRoVUqsgv5tU0ULV0F
gGHIuPrZLrRz/RwAj24uOROpwWBSGSiZDKg15aYJuLRhy3kjWSORfvSXKzKXq4AxbciVHF+eu4PD
2H6J4LSC2u9ps30LcgDSLgFyInJNKqHDH6VIBcnrF3Q9osxoZ8SfEcjP3iUZIy5g19UytA0Ee/8E
RzOvvKTvmzQQYusPefUiGEmXeV5iFjjeUI/1YaGwwCLmtljQYoaGHdEpXAI9RxNTXgg62pGUPM2k
ufNAm/bgZKnrCKnxCTt1qL0YQlcilojgXgGM7Wz/bVvqCMQ9BUU9APvVDbF/NbzdjhtuLHcGlBJ9
DUIWpMLqOTmQyM5NGQPcojxyGQJ4GJT7NTP3KeNjO707epZQaC/G+Ew/M01lbldHRdI6dP8fR7MN
nV/2bzxfevKepObciUsNu1KTb4rwxHM9u8yRvctejAAb4+r50NrNDWrzndTvhjC1PONTRKH/YXdH
iFoPwMCUGLCrKzGiG/9Af7Q+gSjzD2OcXJz7sXfTdPqksWa0FE44Bvd819giW9uIL4G/XqTTy9l6
sF22m1yBu/Na7L67wu7MEhKVzPqqiVjcwiySm1NEl/5xIoWVNUG6pR3uMhksJZtJrK45AS8veJjP
5hCNoRottRYgSjJ+7w45nCoZglZAF2LdWeoD9VHCp+TRxqMzgTBqP7dqdR/xUDQzB9gvhByuIkn1
FoWBBf3KsK7cNElc+kKbRYThppdFkH8zSwgiWHqkgwK9L1DFZTBX/NWEKMtHJS8j5uxr+Bp4yAuO
jxApJX8/h2s6qleBYj30cCajwpJVNLWCv864n34watvae8gpCUirxogyXgly5ir2G0TJj1nTeix0
JgJnHRcTO9LmHvZW73fMc4ZxvfR1woXw9TZvjsKdTisAbCzQ34WjYj7aTqEIsan3JU8DY/9uvH6+
HdiD5rcC9KH6B6YGOxcZhLq22pfuCmDzJsXFRMjE154rwLl1Et4jGFLH3f1cELNV+UpgfSuicoAS
PKm3UfruK9hqVsC+RwLcG+ehl1RyXfvuGaVI94AqN4N2EMU8k3RCvE0bEGvMW7c8rm11Muqr0wkD
3rKkFtYathbXICCBquL25AB71vWsD8bLlsyubVJrayAbnSFQjqKoOXRi3J5+dqZ/Gi1iHWlirJ4p
bLkGJ8Uv9+CbBF6PwdojOabJJOuCqWu39AWFgmUeODCt3ovnslX/FPd5v/4kLRvL4nE+w72pw9jd
iqQlg8lCfQhDeEB1wbfzLWWIrNWQ7tSqETw4eNKhH4ZzhDul6tCHuwPPapwxSYJsAZQ5DQ53hXto
k8qgPx+eNvu/IJFin91ExLszSRJPZrktMQdgmDwQDL9kHwvT87dA/SrWicV35XHCDGTvWNGV7XbL
T+bmLhCwVhzzI//0u2Sat8xcd7Cn3XNynILJ2qIQY/4tMiWKgKSscLA4V2coXYDuE9MDv152CVeZ
kq3gR/mkZuMAbwewSdqaHyTmR+ANLXxQbosAVbWdlmsoFMwafpOX7MYpF/qNPwg5AlKXuhaoTiFA
MHvqTkIOg966uOOrc5kKQ2mmkcfggMSLfHZAkyQE3sP/g0JxUhvt+ipyo4tmZ31ek+YqkNOYaSae
T0SfNswMJhez5Zx80vVGI6KoEcr5/r6nzhC6AHnGb3hKYVnsDAXkW9l1rYd6FLFvp7jWeGSa88Zi
dENcl1ixMDJJ2D1HvQPdwbXUEbCCIO5iv6bcXgSAfW8SghNSio0j+uoafQvSathfyUBicTjPgzf8
RZUUZOM0xau3HuPKuzfHTtX/pvve/xdtOw4QX1Y+sR29qzfHaEYZrGzy6RskvE+6SMy1yMw4Kj00
9FTKYig0M2+/F0srx6366vlVHnRAxScumbi8knunRx4SdE9d9pIdTABrk/Rmh6HSWHwLERSSrH1z
qS5qEbzDn4VWnJwd3OOT47rFHUU3iYYON3CMkTMaejW2xWEfDbJnBQ/yw4G5yQy4RXuIza6hyHm3
rGyjByD6gyrYfSrITftXm7FiP4N8plxIySP5josD8YcJBI6J60ZPDFbWUcVFrtY1rmQ8xAa1DFgc
0/Lri0VkGQn/pkevjpx0ZQnUSAd1OBMeqPf+WonwA1z0CjDgY9b16yda2+J1gwdEwT9uy/Cq0jTr
X2c2Uf3+p1pR1bEvoSZDrGsSPIY4OI8ec89ammjZ7h/m26rOrrvPtABwGDgOrgMQxGx2fi1ucO0k
I++swtWxEkynh2xvL0gBwvaCXPjWnW5lM4AlzNl538ep2QgVyu+lA+Ewk5KTFOVFjGyc8bekBPXf
WAIO/YkWiIL/4XcVUqLTWP6alLuhFNCebKpf7l8bKz/WI4jwu7axxwmzIRgjGsEBl5gZx7oGCb/K
pWMKJkpjBq1z8nVPUJwVGzv50cA/9suwQySs3ToTv5zjxDpFGEthpg9DoBwzJLVriCzn9Btl+n5b
Mq+z1cFCBuihPHvea63cIe7pBDWpvuH0MNCCfqMIB/gv/rR2ageQSTA6feG+kxN9feBTt9gOefQm
j15HSlbFK5J3SFUAJx3PYiY3/5U+QjGKJi5EpnRx/DFCzK2i2A5LpS2h1wkMJ/B1ABrlMhsj7561
zKAsTtPX3mId4EaILKxGhBE/DvPniJ20TRLsJoDWQFFzMck11witfclmXduAooEcEa3wvovbJ/Wd
IfWfAXfXQWscbJVq4uAHAMHx/jE5tjD4PfXq56jQbvM/RIN4zcLGH+38ER2rvL/xkVMathoXIe5n
xx5TbyB7aV+Mzh/3VkRcGwI5A5+wDnlaqIUIYIvbda+4WgQx2w+F0Wx3KzWcPancgZvTXHxJKuy3
rCLLLbLyYzimbn3So2wJcftrhjqnZ9HzZrKke6RxIAy1qy9ZTTJKxJMAiJcS/oS8nxVl425f9BYQ
92gCmyh73fnJ1nQZmhrMPrOVhRC/if0a0agjSB17GkK9gG5T8IlMNpnIIvl32f6lM4hEg1HGHrrM
MhbC6rT+fz7dDdZjcrlb860jFiEKAN4ZEWIgBazT3cEaCimnhLIjadvvBahBAq8wHb56MtTO/o7l
4muVBtPTqruICKM0I2PAC7T/XysA30vxwYw8mVgrIeGKUIGjgt41y8UNeTaSqFy/PQqYd3x62Kfb
+lZmTg18kHr6pHtQTAHD9tNyswpidTHnYf0huYsnWJiwuAYKyPLAZiRwUcXcmYcOT7cg+KK9vn63
yfh/2uSFGkA5K0nr2T+Hk+u/CYwtuHLy8T1KVI4lwOyVOt1gagRH86uS8A4TJ/ofb9Xax7xiohBL
XEqN7/Tv8Meh9qpr1BOSL2m4Si5LoEV86+F5KhlHxpl4PY5SmmV+XtkV510mDRUI8WCFYKf6PJcX
XlxA1Gp6PWtS/NO8kLlhP5SQsg6q08iNcKGm+yFZ66miS5Tgm/NIXQE6wZ0xM0Ic4l9j9tHqK0Ui
ATz+ITXq1j7gaPqVUiFJljYdd6BJL4vnFBnGsaUo1/lBy1faTiZR8E5zEUWgj8oEhSF8xocAWl2A
y3Sv0ioe9PaR7Xsm635hbunmXk3F5rUYxKkro63yzxbm8t6ZUpWQixEoUR1jTFvTFJS7M8DOc7Uk
ZrC8QH2bK/ljej0cZ90Hot+DXt0oJwSWCGpX0RTTUKMZluEfdKhNqsD3O1eoetM2vSQsEirN9End
zF6iwXKlWh+tAz+4q4AmEGsZ+ULQiUbzQtGLEYUdxEAz8zTI9z5Sy05sTm8VZaLwPOaQIVLW0TrB
OuRVDzcJULcNbKO3q6W2spGd15JRNmrJiVuEHg3rgGhMVN7XeJXevtwQi4z/PIeoNl2+vp6IVpNW
CnKhEERTv2BuXDhlGMqEiSRNND4GVhgO2HXcopMF/bmcsEKBxEhl3R5C7f1pH+0+c/TebLdk2lZg
vIF/QmRQhgv/U6X1n/7U3gVBQHW6JfQQO6Rt4cEg+frBYeOtGNBIGyb4m+qPRkEQP0oBhp8idBZ1
T95BIqKCB3ACbya9LpaefbvgG9Klpw6SHTbrECoE+55kEUijVh8/8MIQETFSknyuO7daiwk4k1iH
kNEK+gny5zlYF4BzUp4jwROf6bElwkY33LFlj9Q3RlpU/cKkbhJefAFCIBIkiNU5al8i6sOgvJWT
qRoOY6JaRUsCEqGnay+YDqeHxhRn0HeLrDptrZbbAj0eo4jIZVaEbKmXh93xX1Wnx5v16mwaKaRB
0SROeJYfAqspuPBABVEJ2ZemW2xNgT8Sd2E6rOQNXvvrfLqdAOV/iQ/xk3VWsQb8iYeXb+Rb8ppr
iOtiAMj4qwbjUmGCNThSaBkOlVsjWj2do1zHfPUhBvWcepxWHgoC2iozsnYYAzpQ0FoMyxDKC82c
k3blVYQ79aGkSsDC7zui53HkH4uo4NJM3zfg3yDmj8Kg5IgnnZ1SVnz3tzF8xI6Lxi/2POoth8+8
X7TeegyzKti57eZqliZVbcDrl2lyx4PVhQGqCkBbsJrhH+XiVJaeFjKB4KiYYVZ2ufgQG1AZ673y
t3L/PZ/KQyrKm3Ughksqvb6XXSusq+FZ4Y4YeImAalRsvOgjGLF9gsQOG6KENXLVRNp1xqAnCo9f
+pgqofV0CJD6YZpov+WaN7Uqg/2BZ8eZj3il2mzerZblai6vAg3kjfaUNRzomHZo2F7pLNk+t3q7
qBh/ZTJJSYel0VULi4jNti7A5sO3uQB0DvXhdyU776RX4uB3BHR9qRQj+jwDUfQ4y/ayVhPwOcmp
3mOiZ+lZ+5sz//NtYtxqA0ywSEQE4M/bVbsBiFdTNu2N8Y00Jl68rK3XEWK2P4geOXboDqM3ktVg
X6bcvBgZ5jFc9HMEIaexLACSb/2Or2V2POzRSizfIPaWTyN3LF4oiYdHGxT2ex1iw0Kwjn/6e7w9
N0dPaBCsx/dKzf6b50B8tPPXUs5ezxI9SHc+bELQsnSFFomc1uW30IkkQF64vFDy7iRjQEWenL8j
tGQuUEcqJBLoR4HS+17DVz9wLKR+R2PuqCCT2PvVYUJpU2Qcx75nzJ4efEhGP/3xZOKTWYlMztge
Ik52YVotM98wgRyWdFfpfigOuxrL4n0GQroLV/SYceAVQcS0Pfje/V6AbN/HbhjKu+nZS8Of1cZ9
YRdNe8iyPC0NxIGAkDqOsxZHameVB5rGAqTVIVpla7m3OuBvSTVdlL0jwYUWcvtuWelTxpeedbwq
z1O+3V6pwQFxjVK2s+jAmYLBrpw6ceOkZLshu4c98QeKgWn5Pe53cSnisxxrv+C2hoBck7wiZ8bo
eTrKJLm5XeGX0Yif2t6PYm8ji/btCmtzw5UAje6UBCxDpF5gZKdmf7/psUBrviTmcAHzFN6ljBiu
ev6eIoIdOCoCYlQNxls1hLmDYunXLDkuRXIpDrWufmWdxd0jYFYlPfML4Q80MCWJ+zCSS6PvljIq
axUR/ZRV1pAYjn+eyWvCF5i6bOAK0XMx98BvHEZkbw77cPHA40ITMb5DCsFEcesLL+vCp18v4yBu
p9WIoSPEEANM313Da961TdzATXtKHiRLnWVbkT9pCR2bLlStdQmt6vrEmw0ZyvsLSl94Kxgnno9N
pGne34+brXJIKY9Rt5mQW1ImhW0Ot7/7507JnZ8iYAlXpl5wR45uDx3RgVx4IjPl2sRDqyehFHDS
ROM5dDBI0CoodsyoWrf7Cs237Ku0wUVt8NkVKRJUzG9Y7m9VvzvWy2H7HCc2/RmdVV0XaqFDMvEX
1rl7NJmDkOqTRhsbBIVKLht/5s5EsuSRSHSHaKqmjWwQa3pMN4+ZlW41N+qunI68S8biZzoeJCwl
5nUQ9qyjetQUmfYluoP/JH2rXxognitujCPM2Q4pSKfTrvfaroYesfW6+ixPaI0ekjcfP0dPZtLM
lPPicxl4Qthy2nRsOckbZsDir1XpankQEGR1SNfUVhdDoQXBbi0FL0KCyqXwkQziTkR2gI+8wpIQ
pfV/4NkOxCMdVpvc4JVlqskYNHx+Oc46YlMvbdJpN2LWAuhhSaY2LOirTD5+CjutsYHHP2at7i3t
VnNbUVU9x7GhVNClvlcXOmYQ4i5wAeyQhvUfYKvVfxu4KPdILQeddb6ZX6hL4fXu5keUW3pKj9Oq
aVVpYv2mxX9iiUyWTQZ8rGVkdTrDpVsoWKTpYnj5CZuXqMxOeKfusuPQPZRzI05jipwdO1SUtZeA
pMdVkTlzObjcrp4cI9X/vYnOqt1qq69o9q+yMCwWv8pcyLcWbLPSgh0xw6DNYqNMwdQEC3gjwWT6
eD3duwDhCkAXFBmMJ7fnWvMfZY6qT9hP/oTOfwT75tRJ10fO4paw3VIy+YwX2h0FP7cYASm5DreD
Ell3YkrN2A87w/mI1vh6Dg1IXeiyimINLCUBnJ0LwzG95O1kH3q44WcebgjNPigspX+lBz2EPMXW
maMYszOhOIHnhfDbog+CIuVOLciEpaqCMQ7Q5xjDCGn0G1wMYZQp/Yw+zwPDGnmZqiKYmT2Ab4t0
1P0EG82+aKSDc+GPy4CT2cdPMg5sMvlas8jYWYdwktTia9G1mlFC7Z+Zs2f8uTLGv1ORICLjYu5P
K6AWXIQoqIhSY/GWGOhj5Flrl2PndKXZplcMddVbyOO997HYyLeLSZ/cfMvh6RyFGiB9JwJ38Qh/
GznKBSg0MEqqJv27IhpJ3nN/hWfaEnD6V6sUoHpjZkfWc9XlcVX47ogykoHnomf6giqQiW50gbuU
IndFZDW0r2qzV10EWExVEB3pXYYYFLzuYz6EOjILQpYBzkXELzi14YmjBbFnU0aKcqGv03CxpVcY
0o+TSflXr/scIeFSC1vyGPyBqreCPSFko9kJ2B4WeXBmnqvdtpbyUeu9I24/T+YxyP/gETBDU9+j
vBpWjiNdeBgr2Cd3U90ljinaenlU5ldVz0n6hiyXr7usK27+3AhEObjAf5sVCiyWPXei5hahB4G/
SCrjSl9MD7mU8ezo+UM8/WlIinhp8MevD1XYoM18hVbnedLmb4+DfhiHq4uPQmLmwbO1XVopBReX
TffdF8ppNNfO2D3MX5oMBYO2TSCNS2U+lhVGfvdpjRCLs9sxhp+ncmgS3DUigXw4fTT77rnTni7i
PQhyhmRAMrvTvVuJC8n4jM5V0vzlOID11WShK3O3HPvPyKAN4RYB1N3yuNYL24WVoZq5rQuZe/9z
M9HTT39kfsGifGvU74+pvn2kdOeVRxFEI/WI6lvJzwb4gMrnmH/DyrvzyYkhUCSx1taX/Xf1u9qV
ljRe7OjeBQaHqwlqYdQAV+gRefQVU4ekSkruP6RLJzH4bXeCr8EsVmOsYRbtUu2+gMuwiusoC/cd
7MhKTTopPLgeJN6FDhNBdmXJMrRArqBuGg0JqnAMTAEj4GvGHHJXh9v/W13J+h2oDMQNC1TfFcTp
4n5BclJfo5ElQnU++EVWz4BqUk3KhrM/2X5cnew3d+KupbfQ83lzVYJTz8JOyO7hR0qOLxmkj3sn
LJMcCrGWO4gmf0EOJOEdJ5ELr8m3/kJgwcn8V9yIscejrwM9WZU7npTLq8XXe2nOv5HClsLfcqJy
lTKdB0pCc+bzRBQQsEHZIf0hg+mfAe8qLGTOx9LnSYq10pxbgW4/3x1jv80qsSccblEyQb/Xm2qe
tFbdler2KoHFKMZ4CI3jzx99XlisX4TaTzOe0JNNG7mcElfd/iKJpX8v0NfMZc5G/RZqfpBsW/Z/
1AwLJ8D+VnL81iQc99nZd15ZcAUmVtEH3yU0NYQVxJF9D9y1h4MU/r6WzW2sB4429hKXVTBAGk69
zXYi7+oXaF+TSouIj9b81555DXJT/EjY7sz7S4sY5okluhLXeMgDMd/dqz0djZYAS6hRikSY1aO3
l6Rm/lUdT7rVUrW5HuVPXyllmC74nFOFxFVlMyYX3lQh+YluUlETZLYGFbnj6kdXMioUi5U8PHVw
AWeD0ka0xHUV5GmwvP3iBiEUqorUSDDxcjFssAOrM3rPNfrxjQi4UpqGbizdYps412jlJjLjE/E3
cf0kyxQks6d/wwXz4oniOmL5kyRlb0krXof1rjjxSpEi3drv5Qe0YEN9PA19ruC9hhCdsSn0kpWQ
MMjB0FOugJi3fzcAr2jzuqdBXycmWf7SqCw7LnJjDDMoYE4+RKDS/BNO37GFSXgu/UY0EZRoMXeY
ywzCHGTFgAbjSFC3TsXRkMiSAN1gtuwCZ6n0DBNm/lYuADTBKejKuys/5NMLu6KDXr2S9YCf5zhz
UT/5vseB4W1n3A5kxuY4FraotiKBGBvjbgRtK5x8rf9dzmN8p0RbvmHyOAAT0rtU48oqGSDhd/ih
3ZhoJzt01KkJ/ZL7HBk7egizXYfaxKtS7hQ/5eIxVSGYZMmzYwvDLV+IuDCZijSjnonitLARpMK8
+VW2dNODyuTMnqGqdMAjYBrL4jsT7+roVOMXeD6gmuw/IqDtj4s9Mch3XDr03q6qdgmPVFxBzusG
hrQxYd6so53Rh60WvEbeZRXeBPv0xef9NtXBcuCz5xxauEFgCzWLTccutz5WHfWDDlYfaHoppn+l
ugPJwaecLrZ8Spu9BS1Zpnq3Gfp9Lwe/rpeMdAY0QAnNndJBYYoD2zHfgqnwbv93qrMrXOjopjre
SKwoL6XeTL5elMFS2QzbqHWbS6MjNOJ9qf8+DnP2VLoNadveO/NFv8EtSY9idfiViSXs+rTvGljr
aD1Ju5eDYE7UKOgEm6Lhq5M9yX3g5X0c9gbwwIUx7y2Z7Rn2FI4mYJRLYZow1WsI59PBhmXaCWa/
0dsnBRw/+Lv6p1FZFfb8E7tnH7s5HgdySyv/iGUxZQ0gisT2pprXGNCyJJefFMklC67kI2Y28s5X
9E7tY0WfDRCC7jJltMDCu3yRgd2V9a2maPfgLaSLdQTs7jwY8+a6xoeVwX8ZphvmoDrE2lGm05d9
t76KWfaj54FwlcItTEn91Sfz4594cbq/FancNZg+GQ2cvDH7twZV6RnnrqzQZjCzqxo89mz0xiR8
URPmvEl4pTmBvmm5BQ6MtJhCggzHboRsPJvZMwvilFuWAISoQh330ghcAdxDs2DVtbOYXau7Puhr
3nsvnR7jiTSKRhRo1YwakwxgIptF1s8x2r9PYBxeAQqdyZLCHx4ewxl8/Xthyi2+ZT7+mc2j8hvH
XRcCx89qpSSZYcHrj+jxFucN2WeMMPNzDDaD+XuVDPMA1BmOA9IL207RmmkUv8D9Y2mXp96Y/CEm
ynOESEs64CKKJHNyz/amwHKOf74jdNeVcsyqkH7tXDFsWTntX3j1NE04OytjWhJEXYN35usvNEf4
5YlJ7Yy+2OcG8a+Ss6PItLJYQPnXZLimfh70wTJ9/tIr9XA6imBtsazG0zB7JBQciNSFF9QMiyth
Plis4DPVHdf0shNXmxxqcj+flyX2amUw75JrLJHVwCOmQyzXE/YnBjYBErP2nwkhpPtGqHZ4eaY2
WaLzo5129lIPA+sI+6l73x4cVwP24ZcgvPqpbxEM/KCWTc3fw8KVjhKfbCbpMVZ/JL5lqkux6U6t
z5tgWpvdutb41h9oQf+w7zcFHjAbRH9TnledsA/jRba18ttkFhjHhI1oOZPf3uXcI7CmFIUL9JNu
KTsfeZ9pUyPMGsvLKHu88EvbfpjSxbYLtwmapm6wvnHc0QGET3RaGaiA6NHGqukHtPIqCe4OF7Ba
PVDq6RGWw+IOE+5e9yndZx5vW3QoV1iBshjlDRFHwRxQcmAxUit34WY9Y33gQ5dj62WjgrxruYPx
YyyWMWwkhC216AduQd9tZOoPfkWO9pT5FOipP889i1z/NiBRv5ZW1wRYLdnCzzErz01/vrNz92XW
ZxVjsfZstB3FkW3omd+YCYyieIKLPY8+Mv3ritqrd/M6x5i5mECJqGGllNiNEDFje1JaMnxlPtKo
qjr5bYXEX0bzmcPc0HUCTE3KmBMFgVWk89N6Y5FzKb1GXB7sV6jNb/tsWrbBAHBrMPm37FM8g8bC
sjmPfk45BIvtMkM6v17NjHgbI+VlQ6pkltho3NcEQ+aDptIsigcnrBQtInj6YMH5YQ73x5O0/DZA
5HsSIchyDc/2Wiq1ON0PZlFtbzSTg7VJWH/1BqRKN/hEqWnkztulAs5mvpUDpFdI/A6qmcShkoqy
oy2aozvEx+CGkCo5EwpTnUHj8gr8LByKu4orn/uUR8xSVdLzbtFqqzrwhcYr4bNoPp2taJ06Aza4
o9p9UBvWkTvvzoqiGzYC/nDsYGO9HU60j+f9RruJ3AtMhhCdVriH9M5PNEpXOtNqBGvD4uUqvdoO
69t2OB9EEOdOMPuMTKbGIwsIR0pAB8DrLcldEZ+F0gbNBMvUjP7/DHnukVTnQz1bOaq7ddjb5PCr
DNTOH4zs7ieAL/ymeoGqUR2kVDTcD28Zdo85ejTBsqps47NQeGXeJVTVnL9Hd6uYW3iSHD70CUUf
gyZlMYqvon5KQWUkgzyX5Ak3WDj3WLOdh4crF8/9tscRiT3mHGxCG8HoaIeqgZ9dFfPMeaG8HSxo
mVe7PHhAzqx0rfaVivqrI9fiRYDmMEplFWK+kl9D87/yEcWvGJ0iCJ3sJdt26um26ieL6ENKygyO
+HkcM/2xs142HyqkUd8rwrvHtVYBg2AKMP1J0hhbxVKTchWETUBuvpuN1jAFn39Ir0wwqEf+0O37
60/l7EdvX+saaHdyY9e3v5zlVbLD43b6oFTg8RxPZnrW7b7Pu2AMaDyyjQ0KVrwcwm7uRPwkDLuc
9o67o9d+Uietn2gn/wiLEVtiQtAjRb4kYLpxXHzXSnSfEvzudafFsyYa/CMlNMJFQ57iwJxdoHZs
MjNV90sa/ta5mvNKG9vLV39HLlgy56fK7GqVNjzz36q/yPtcOhgzhDO9HLQHyCn/IOIdlSJ10EbB
MwzeAGTGfSDYCIiZlFdsaTTQSW3H74xvLZ8iqYOUoAB0EY4LfC4DJU02x2TvSQMvCA+iuFtf2U/g
SOGnZ7cUx//OcIDgzg2y1HxSWJWLnkrTj4oN0wRVSTCW6bxqQFq8RkSVeRc9FRaeFrWMFCcVgxB6
0lNbXPRzL6nAXI/nl13r3hHMEo8nYRhFELiZmFjjW14lrIWZZAPd1JOLxvv/w2+/dzXIYqe1ko1J
odenr7fTvbzFYprfZDp6aEKJnSIEswZ7gJLzjflLtL8vDGofdLWeqSqsrmPQ6mMWXvx0DpI6jjZa
L5VG1L0WYTgOww3v7xBUph4c0JNwJhESuXMxByxFzwtl5JNTyZcmgSg6lNX+KbmniSHFzijXFFVu
86VsiyI3FI7WiJEhlLISrEctg6FZld8RZuSAVE4eX8nllPnZdU1AAWkX3eF2sAspTWhwntZj4yb1
3r0i/Te9rPZcp1FmR6JpO3Y06PIO+tLCl661TUik0qwT3UaU4GY4xhptldkRQhRaKCyHuyZXxoYc
zYLk99BlKIDaMY7R873mbCrP8EhG1Mpj7u0pZEMsttzke7m6wQ438Z8Iss+MogjRCDpf9GXzvNhu
gcbfj+V84Le4dR28ARmUs3/4RkvQCwuGJo86//QzujdqjmKMPaOBOiqCNdl5aEpym3EbH0yqmksI
hb8ZRstq+wPYrTK3q8CYxaNbojjELUYsI/jWpyNQWkkWIHwRf7DQpueITNEQLhaMqjThOOLD451f
UG9VyeU6M1uZDww5Hwe1lo1WuZ2KuRoxKKcXMnZ+MxDu0eGilwycHECz47SbmoPc+8m5WtZlqAtM
ch1UqekkqO8idNK6jQBJLvcRmiBLg1J+D/Tc5ZMEA1IFHAaaGG8HOYZS1HoqnvnRqhpZ4IHlSP2r
tP9x9ic4cjBwhQcg31xOLqSv8OKHposo1ON18zGmyLKnL5mFhMi6aRaMuCvpbEX9vYraYpaUIWxq
DKCneP8ojFB1CEufETRM4omvJm00JD8vbjkMo5g8OvQ7leesY7JIPI3tehp7AwPQJD4xqO1XrMdb
Sg9aEJ4qfmcd/IC85yINnvDRtFESHlYZ2pO2aZODB4Uio3+9s1boTfTpwTj/xNfHpFNd9b8WBaWq
xHVYCLxuHE/tGO7DZQjvzKudinHonw96fGn2JVWARCwP2R5MdF4akybrRneOdOL+I/kAmFA+xa2E
u55LxM9cxwys9OSeoKGX7RVbqzvFnIU9JlE8+ihaLs/QAGJuOAmun1Bcr0Cpr6xB5EJAstJLCXvv
j6se9QU/JgpwXGni/onnCmG+EvWj1bRI0J/9YjM7npCKDs/ktlVMxCcD7G0Ib5cXedkRJ9koBJcg
GhS2vcAKxcMb9nwFA8V4aHsr88c+8iyl3E9FW3ghZPkKJUOQ0lOo4ppYysj79Hv0jTAZzgxxEkLn
2RuA9eWZu2ph5iqO7dKsjZpLCqqlIog0dl3eM/EYCImSCuUR/gdH4EXThEYajNbWfFYUEEJXJIpn
9R0MYMeDVXuT5O8OzP9Y7X/uClUDREEzTG6k4ZSyxYrWy+9JpalgWZoljSbmosfcMucjrgWRwGLb
s684RRHgPQpgOrnbqGXrdFQOcCKfSHlVDqvMoJGy+N1uHG2sMmEFjjHTwrxA65Oo2UdwvOwszLbf
elUclUJrEgrwU9CsOXp0bdJHmKiP0DvYT6DZCGyaWxd7vwcOaRGk5X7LdtSSyfNywDASS9gzhp2l
DmTwmyO+6kG5zJr+f52njV1HSbTgZrp+qwGo4k9V2SwuALl3IUQ2xhJzPV7s2Qm1gHFoDKVGm/AP
grz76zlt7jPLEgEzlk61aA0dFUr5MF8anqAwtAxdoAYVCNc9jSv2KyrUjJ4+/vAxrQlIYTU5Ti2I
ySNXauhPiODICXSDH+1SshOX1ahbL2TiCylJbIogvKcoVOE4GZxI25SSQPkb9znfqOZcB5mOMihl
QV5VUzmYb5lcOhjDGv7qTdos4CaSn8/0ekPMaHmudXJXxQSuZgzwGq7J8k2nOvH0VkUHyPnAf5/m
j0yst4npfjuz2KaDPyZnm85T8Stcl2Eo9vw2CAVkuAsloryaciaSysxpYAzp7EAwSQ5Nqxlf7W+g
kx/obkxXYVTPJNutabJ6QuEE/SQKh5/Uqp7Tjerx0yyOqITeLnl39COKzVlUwxhyNISxlYvvS9mQ
SDMgufL+Kv5kie53JA1SNCUbXcZ7M+QSwo6fSmVXOnnpOGv+eL68u2B2KnauNSp+Lp1dskkthgaL
SiffkpVR0sf2iC32tZZaKEueNZmvUxLr6kSVJNxxxtd7GB+pUsOC9qIHJu8mGeQSl+jdiLtZP5ka
vXdF/LFS8zlfcDmxUhyAvIrSobMAriuboCz75bFnnV1vXIGr8Szn39GDqjP/4793sWSdVn027Eax
9cWuNhSoPqw5YiQmTt0eet4UbRKuqUYsRNFcCE+egkOxHyA3igjNr2kGXT1QJMtBnJpNPu6miBtV
/3NGK80R7YSuQBWRR9CN/HUlg3mwtWrl+YCMQjuCzdcI/Evur1e0J30jLPSu5g49IhPIlvEsePnG
PD0QS2wKKzC92tflsiXLHvEW3BE5vblFlIZbMFW0jWYnAuX+48DUOxy/GZjuDB/oZVk/23wALGZ6
mSQ3Z/lK1tbUkSuOdVie9Wm90JliUrKpGiZXAONx3nH0aDCfkHnDSh6UAkF92OusxfMtF8HBMDmH
P27SCeb4T1JpDl6Xic0/F4KMCtc0q4wWcX6a9eXHjDFJ/t6jDxCXJGJcr/Y5A/uQWnCu/325JK67
CO0uzOZsFUbb4D4Vz9CeuCmHYBzwR1/Q8vU+FpweSTFU4xkAYdW4/iV1B8D4YUvMDe6gseTzyUi2
CADw98tMkUKHwJPuwZrlellC9GifwE7NG0Effa3EL+3+Dmb5DiBOHoLb/mJ74o/s0jj3d/vK453r
nj1luVpGBTcK8+reKWJrBZ4hVKBs9hebdPN61jGB8RuxFPjEBwkrSKtUWDW5pNPSDTtBuz5oMj0S
k25d4UmRqsPdH8z208bQBMiRv2Q/GhdKtpwYffbSSIsyBMX9OWrSAQ1b/BTSLF2xH3DxPBg05bZ2
0nShaFHCh+fB6YeHVrbJKK8pVyATXaHzMflBs5oklVBLawKP79U7Wv7baCtK2lsswDKu+FcLKah1
4cLf0K08JyNdfyCq2hd1QooEppdo61Ua3w7af0hG6h4oespeycXnkLl8f4qp3kOrobeHccawnf57
3aF3C8gk4fIWR3hw4M1CntGI5TK5rBiGfyB48JGQdzamb77aPhYbGUZRXgYIgLRMH/xy4tpMEfDN
h2Au8JL4pg8vYXupmeFoFSTjl7la7tkt1AqcV43dcyQXTb5n0lOFbszBXYVfEGAF5FlLM9JYy2kU
w1Tu0TGkVAr2kAFKKI9iu93w5lIy1vwIzUyhwzeQKN9xb9If4Qepn8vXKtruN7RI/qCI6HN1zC9Q
EquWt5HPe7D2F4BdZ+PYXsxb6b0Q2733XDyqdLy0ec4a4t2yA+Z6l5rZnjhEd0tPaAemd54BENWp
l77Kt9E8u4Ot2TGMSK7azScVs0jCwZ+M1vCmzJyyrPBb0EjlX+QxreDR93SQmKSdxYAR2PVKOIem
Wavedk/dMCuV2bEcBmlC67JbRzppmbYeQK0j2PXrL9eQpsLAYe2Ixv4fxAX68ByfULZjP0QkRSl4
gaR/5z1ZhaJ1wD0Axqzwh8W0GrtQTG4wKqhSF8Q+lUGd6/p4WVUmLMYe22XSj1Pa16bkQVaDXki3
wydGxeCvTpVlgw5kr1QkgUtIKp1ZkIkxiuqoHio7+9k71xfUpp4PJPc5FcGhB2Kb2mXYopYDkAp5
6orZsVh6+O40QoT95sT8IB3aOvOr4Xz7S4qj3I5TDu7Zg1KofI3alr5FrNUd19Ypzcx34bomW72z
BjToj9ilNwcxjkswdaJckwCRMuUv+iR7JQFGnM5/5V9zGYYxes7dC5gRsbbmGN6oPhBtG2bKoZcR
roLMvxSk5moHJ3wLpPouG4bD19iyj0jmXwOG438LTGD3vfjCJTuvyjUMOrutY62DvUNz0v4WcwA+
LSXRsxx+MmKs5e+YpNLmEMWbagFVWLuGf+elU3n9KecmN9siEjxhKk6256XskNtE6+uaxG06lbuP
8T7hpnuq03CBTHQzj7PBHTXtdi+hps01asIeTKeZyk4jZRtenJrF2ENmG0qaRPCvmc5x5i27Wfbx
uCGbYb9PxDp+19cV4Lh7PQEoUp7FFt6gy0KEM9tj7RnRhvHSSzbzWqXocykXI5pYYwjljsQju4Vf
cRD0e2c9/IHKVB8BpFbLUR99P8bTMrrYeOnsOrjxvaK9N7rfK8znHPXkGFEnM4vXF5Ad9Tzc0yEG
TCGNEmAJ6YpHaeZKJiuyAiS/ujP2xKKhB/qiJrDq+ylxFhju+eD4AJYKkREhjZD0cVmWBP5BZF1l
RoEovIP5nRTeaobc3rhw+LKB3uD0DbTQiutVVqRUXY/M67lBqjcqDjYWfZN6hvSu5weX6OuUHoqG
9yW8lZ9cKg7wjcEG0PQlDta5NTiGFXygxyT3b2d5c1Qglntl18K/lB5nVJxCXAghWbqcOFhLR9Ar
f6royVyqjcv7NTcDM3GqTfgWv4Zxcng+kdhqPG8cHURalxqXcVshD7VpFAV2J5itUzynA9Hf3/6U
ci5WVgDO3dScUWyoiXDTubm4bDX9xbEiBuJOfIxzQXKSeYfYbM21yD0Lzw0/AJFcHhkC0zfuXBnP
DqhPZZMDDk1PnZMZ42wyDgeWdoFyiAbLbcZfR1aV2PF3+wMTTbPoTIFExy8l/Lg9HYNclxUGhvHM
uQrP4+igIjPuDGkhLleN/7ZMAQlioNgEJH0v2ILRWM9T4e2ivKc8Jn++a5Xfrynk6u91pEx6djPD
KHE3JyY06zE+XDOqUCqDHJuENds8jQFOHZBYU8ln/tI2Ygl0mSi2TZDACji7pvI783EWSWrLa+a4
8Lf4uur/FMe0ek/Z2QHKMyj/XIcbqy2wv+SU8IaKqq13fNV9Wi07sBSHIxyTx3nSfGFRY1MiafXQ
1gI8SC01G2fV0NcZBa0uO9yLRb8D7k7ZuoMXJLVgdtZf8jyr+LzeD86IArdzxGFmKir0ksS+rFb0
cCf3VWVlH19oRpVh5NC+e78XOyNyBHCO3DK7y6eS3nkCzV7FC8OM3vsRi5DcIpun+OGPGi0sAIYb
18kD7el2+4mu98Cpppfl8EwitBBmOaQC2Xfm03spVz4+N6MslY6FfCnZZkbn3RW1c6WCZ+sNfv3X
/RRns4PnRuBBjm+2X+NRICX8ogJBdr2cdy/VSB481JETMU3B/xvrvTMH4PN8KeH9iJegRV4yfwim
syKv70PIBG5jYj/9e6XzdK27aU+Zg7E/TxH4yhAQ+jbiWUMoABKpyIQ7bJLv9VAX29RkcSEm3DLZ
UY+hjRHD3N04m6iDteCfRDGNMm64fLLOs/jb26axPFeyzNC3tQjwNExoYfPgI4N4/5lOZH91sxKy
UZ2LmTjC7MsMWQIlQ+l2ZJvmTsGszzTthkWQ759su/qWdVN5o8IR7DWZxYV2m8VAsha1mRsMC09M
scV398s6pfn4h/tZltxhgWhvLbYDptcb4+fLNS8MmNgwpfXqGxmXI56ZqDVRN5egQMANkT3jUkh1
UteS9VS1t+RPIF5uxPKU4/vIYKtLXmyNLkjS00gWlL9ta8svdFEGRf4BgfeMUNs8gtHquCQJ/i4z
MOFWeapZCRBoU1yDjG1Pgki3lOu04t60DOaSyRclf53SElLldhUBw84oUG9BNHbVrGMewpdpRw89
ADSLA3rO+W4PtbsBRKTrUihYAl+R3Cra+GZ+z+W8TORk3elA6MH1yplYXAxVnNCWB1O534Y6nG2w
/llVbYEx842OmZAAbaFViUEveZSq3spsZqyxsvvd9ee69L/glV20B0qlOoWxtfDogb9gKcOYN5/d
m91VnE7cWa6kh4fpSYM7UONX11ne3lM1piWgT2TEmF/nlS9x4ze5w69wzWQ2i+UUaEmlhzTSHU9M
A3WlyERIZNVWsdl12839APvXdLrsTwEX4VhTIjF8g5NC/3K6U59oWX7PLvH5++eJUIUFmbZYkEBx
5h94e1IprGL9Ylr79ytGCJo2ctKaX/irgHiSb/0RdhxGvYGmbZdK2wCrBcU6dUctvlTKfXkZfSV2
gjG5dKITgccRWDxM8E9fmBhToTs7oxsXvLhCM3jAK6qZ5mc7Z1fRJP0/Zwu7fkyOSHVQCO6hhowq
sFLsRk7rk/QjNaHYlCy/BYTgBxjoYSS9odTGcP55bl2/I9Vk+0g0blTFyCvxtTCxqobsjeVX24JL
K+cqIvattaOk5Z35nnwpkLDuSNDnzXtp0GWVAJ/jSAvJm3rfHUOP/MwveC+eVCm1lCMAuL7yvSOo
lI9h8JaoIk44pEMJxz5Drl3iEh7l0I4yImiUK6jHABkW+ICS/qr0lI/dRrFbwgsAvzhyqvW1Yw1H
Y/kze8ZJIyo20cr37IKWknMZ+/jPShhJcEKLXBaVvOUPuDzWkEREsD8xRfIlF5V2ar1ykLbiwid+
MFOwUHjZ/BtQLgheTcNHwMidix35QjxjLsP5cgd/qUIBYT3UnREbos3hgKZuI+Kh3JD54dvhMwKI
VU58jYnP+RHVVMq9VetsVEhBy9SL2HKEaAcJgTO5/Uhjn16F4HJhldFlpiPcnVzkei/KYPmrunsH
oRu140ydrGYd6yqrfrhPXetd9i6CVn5LIWfqgid6EMre32b/pA9vd9kZdrSqbevmIBoGu1p67oq3
qQ1x6LRY5Jxnc76KTCdDEVWKwJorXlKyFZImRLrWD+mVPTa84IlJCwonSNyA+QNI5tuyANZpgIcW
gC42Xrzu7j5rukYFMuf+sqo7PR+OrSbROUBLgBpgbjDdjl20tw6CSRB81H2muC8OERlzmheeKw6g
8c+SKlOm8iD3qjirHt5G6+aF9/4eJfH6d5UyKhz3B1LVoW0ZyUCTbIO8CARpKwu2xRiYl5v1a86I
BMqql5tlfiZde3rnOiyKs1pV/85AtqXhBAQeUsW2vQhQ6llEW3+ff3PO3m4g18MeibqboCYS3hIG
UqFS784LLdUEplYsoPvvO0V6CEENQAoeQ54HXeueTwURgpMCR1y5B6fMiWck6Cqrck6hZlj5xLoH
alFzH0YanYY8eM0/OKtNqh5cRsOWXnWJBeqzYFDpvdPDwasH0B8xCqJ2ODgw3YVuymrg04a6TkqG
eT55efcRsi1lLKRRvxqkHAtgiPnA/IoGZk+WzkIrHg1tgKg1qHjGaBnrveHa7Qhc4ayIAKYfS8A2
0hU5o5+FEJ+aQjvrJ67+q3BU7wCDyBLxPS4DAhw1uv8gna6Y4hQzg0LGOQGAN7+LDlD9CU7c/Nle
Ren+WCgxNlH+put4BrKtNmTnn1BsKjwtvg8YRqIHbFs+M7Ta8C4E3BB4PZjDtrYn9wlvV5KVZTDy
0b9C7KJRCOleleVAXjhBGDX6Oflzog1JQJXq82SvaFW+YpGIwk1JZmhVmKEyzBt7zBm2HRSK+TeT
qQigYKd9+wOVqIOa4XmmFsHqagry6Pxv1aMDc46AR/Aix4C6k4Qse6QlNw0C7wg3rVcCX3gteWYk
8HLnFJ9fwqamZvpv08f2clAr2ijtQ4L8gzBRQWaWnYpFrdoqpB47Tl83sA5Uu1ssTCqYFgpcnGW2
oXZI6WlsBCka/aOEFdzG6vv5hmuWxUO8S64bjFEcWAvoKsO7Ymii1ysnx7/6ohw8xgL6qkpCLKxx
uQ5pquII5/NVmtYVHndx4EuTyRnvVqMyKQQqenCjImb+kXU6n/rMgyVO+lmZ/B6V0UuDAai1DCKs
Tx8PXzKOMOJsHsBP+k3UhoG40WA7Xq1sIMnSrNvXMuSzPZ1NvIzLS2/odxmaH+oEtLtiF4yjfUu6
6vlr9lM6DIZq8Es3v98vcs6cNTRpSh82jqFE0L9GDEEecai3IAiJSuiYtXLsaFLqrUr3T9LI2rw7
EwlTv3g8zxnB00NVgAqrN5rDr/xpchMrlMdbZQWoQz9aNs1NBQDEtkY7S6CY58sNheTvchKjDhdq
M+e9aCjXRb0Qm/idJ6pcMSzgw6PTN7yPo9xM4zCkQIGwd7KxWUs+9f/d8kcD/LB8XGAGPohnWch6
qpqe4wepoAyDbHg8qbmerLLlQ+/GNIR/shL6Hp+pn8i+zbCxIcDvfrNkIx+24vaes80fQKuU1vXr
F0IkrfR4H8Vr2U60TIa71WGSdivFUnS3UdLomHMP1gq0ye3oPMiHEqGcuc+5YbUw4fmGRMKBn0v7
kkhTtaWFJMiWxG6NG2QmjGb9P4rDGVXsqtu76+jAYhKYjoCVKTpMrKLnsqlNQg4vxZU0EBqaM7Hv
zmPeyTBt/pE6QhnGAANRweO2fVGndmNOj5ztloQivu9G8NBcCVksp/kjhpNwGYarnacfoPR/0h9D
c9F84FPC291hEe/61k+tThSpHFuEQOlEpi97hLV2NsxbqmLqGUU00m59RsGGsi/+JnleGD6uOjI+
0s/fpDBE9Mqif8gGqXA1tv92Bxmi8yP81UqBT3CBUn8oknlJn8MPPq+pgYMhB8uxLzXAbdqFkUST
yaTCintrwGqKWk2HIuf6EGFTvbE8gtUlLVjZROP+9GeQmxDr0QGwCilcJ7/OubuHZqRlmQ8T/xL/
HGc3QIycGL6LS0+P9SLuGXhs3tpOiauwVD4K+LX2REAh9bJtu1JCdacB6TQgFANnWMdOVf3c4D9c
xeR5423+ASkW9E3wDfr0fnjct09/oTGOnm6GudVx8NPlFpBlie+UtRlxrx7AFIDaxYykfSZ9Tr9I
DN56X9xmtMScwCGo4FSBfZLtG5HNjNe4tFdPg8mryhpnpCdrUTEuCz8rZEaVhPm8zDYrSsNyCoUk
vL6kOAVNfQQNoIy5Msyg0MxErbq4XYJ/WZM/YdJgl2huoMOd5e7dktjiKKvgZdEk2txztcpCFbeK
ej7HM+2QCgDM1j7lQxnzMX9A0ftzQMzudHNR4AOiWK3crBF66GBg0BSZzrEioqQe/drWLslJlDGH
uyWAlFxMBwNeKPH2qHys8UxDWndYkRwWuTiBJgU/2joNZbRGPnNoT7D1HlNu9fO+WmikKToOQSRM
E5ZM+wHI+qTD+7JRMkP4jZrRJxx+jcGtqDghqvc6tyXi1PrCBQkDHvdF76dOv7MNMxDn5/zELeyA
g8Uck/I3jnAfOwOw40x3AOoNx34AvMdzrtHQgD2JKq30LwuHaFRmz5BMxSkMzO9sy8miwcW3T/P/
TQyt4Cxuwt9dmN2d5yLwovPvG01nL/z8IIBIM1J7qr6ChE4BlnhsMZxknIZGNItAo0RNUlQFqD5K
ufblwv23dhQdFjkePOc5Vmbti2d9DLNaFW1gPiN/0RNT/9HEXfyqhEAEho7Sv32zNRK2JdBuhGkq
AqgwoHD8HXx8lstpyQQ/xtYeoebcroQWHC3A8fLGaPuP2frKH+W9Jzy39DLFZslNA6tSeX+6b398
v4i2QTXfZj8lksaO/sC75Lfuo373oNxSGdImd9W78wpwP+yobEcRp9u8pwVuqAbRmmWzzGhL+TCA
d/z7hXz4gnBxnOvm45EKnPE01HN56ZxmNHVZO1dyydrxgNTmKEkFXjR+7eYiVY/UInm+fb1s+6tg
CDvBybj8zL1hS7MtaUUhgwVIDM0ZXJrSjEkliz5O5Fe0xIN6NjwQmbz3GWVKSshCrTLOF9uGBh7/
6MJTNyC66Z2CLPik7AnV0JWNfUJLMij9lusqzZKCAqLAbc271SJmcbhpRhxRBMVKbLmC10HMvR9s
7ksB4IWKdSVOsSvHNGpuyR+H1ZD+7QlrNWtQJGaXb0D7cqKuYPKV5J4yZJT/v+E1vgHJiPQRxlhJ
KWghdVBkgQKME4fP8c6W7LfUfnh7aHOZW5flzNMg/I0zQDnj+wZr4Ho5SRgKe65rLt+TdbxIGpB5
jtOI4NGzdcvHqiABq4/M31vGe3lkFCA16ExMupIJbR8UhTKa413OI79LaMpn2stt8aqNULRQ9qeO
o0PAEQNupfGjBHgfHbLpoRiRIVfNXo5A3eB5oDbmrrO6ouPv95HNqOtDvi0Nrj8qvTbcsup6+ZiK
GMrFCj7TILXBgEdPjBSBJKXwG+tUFmc/ss2/+knP7w4Lt6+Cu1KqMSZRp+QkHwjcZcVrBPqCWoAC
IzKRWhc11rrPp/EyuHjJx52Hqizl9Sb3WfIolG5uJgtETKXqdXbQKUu6Cg+sdVnfDajbwh405IsE
72jnFI8O5vMjXSKm7ErnurLF7o7iSqYMjgwYx3GBLWvklEpki8ddNPln1XzxiF69naDTYq/mhkFl
H4Jo8SW8rL7f10zz50Hmofm/dMu4hLF2wJs8kDtA4d6nwXsWONGDqkgr4g6FGwkLgNu81u/0GIRG
JlFkXHEIIFfl+3SKbfrjHQKLHSGTBsqP99pySq9EwghUkhpTD7j7M8Z5iKLPYQtGYAeHnhQJVaEU
jeHUcHZVWUGBbGXm1AUStf7mCivw/s1s2qlYF23zlrtNHvBkXrh3LaM6s/ob8M+93216pw6VwvhY
y3gnRZqy4dXPVy15s6J8NXTXsZ+llDuorgtDk4yb/CtuBQfSBOjphvpwxJlgY5x0dYuXkpSvNzAf
BXYrQUGjtZi4lqzUjoSJ+r1zIeOGe8L86918DmumtBiXGwSo7aKpjHdPUo0OweGH3KLkAgqxzDDT
N6JmLKDs0cGpriWALf+zZBmi9lUBss5O7wUioRfwNWkhsBtS/sOEyTsd1s6g62nOuFQR9WfB4yvG
bC3aAFTe1p6EoTtJsQrAVQ+6N+QuPNojBj+sjqnfJ4Diz6XoDb+jo6p5A/p+dH7YzYlu5npYbtet
CWbTp17CescrqG2WtV17Qk2UDsr+Ji/mbeAYFoBVnysxn0OJ3MsaEVFVSW1XzyzNZuuVrcMqaaRf
9QmTN1Npv1qSi/ejQCIbV1vOoesae7M2vC4hpaIBr98zGO4GhOdt2swLMjCJlh4OV/wap8FBIZTa
JsF3XCatqoIpt9yd98yZK0srVkeHy0xBpuZiInZ4R0P4xefFB+ctmO+P8rUc6L5xpfLbQBoF2Qh4
7L8ffeP6GhTpolV6l9ta54xF0ptlcEX0pbXAjrX1guP/NtY8JaXBE9fln67BFkMW6Y7T2ll91Bf9
Uik8d4b6BRYoiEINbgvV/OymXWTRV+1IEBTRzLnnPF8drx965iowNG9Nlwl/xEBq6yG7QRdJEp0l
mO+nLqFGO2Y1TWQyn0HhQY+ypNUCs40Cnec9tQZr29xhgOj+Nm1ALy99/nIyYK7YqL5fXJfKxFb8
KS78I+j8zO4zdH/aDNV99OxpwvVLlsqEo5f9w7SirnBfgvQQkF7Ma62xGpqfRTgd9+tDNIZKV7Si
CDwLgxzAkUBelU3TWsiGd0w7O8AWfe3n7N+XFcZD9tMuo7O0UsKDzxqZv8jkpJXDAQUBB3m6u4Fz
vKdxit+OPmI3hEFvZRjUHi/nooJScuCc1I42TcrOPXzZSdaXC5udNUKIHCnWJ5n5kCk5IFoCJV73
wjwywM6I7CAzOtxFLf3+WyJoXeOVaJSsC0Q+vtR64GQBNMNvxPSZwX9Tj4T/Wot4Omtf+RSCPqUd
0DJ/L146CoxYz8ipAUeC6Swrl+Rkr5MffF5RRMFHSqv2QorypqH8z/Ax9ZsWnPLoAloUoNtuBAy+
PT62927/MTexdnE5IPQyH4tmmAeslaCmZ6lxwq/WhWtUwT8ysGXuGgkEbYM8fqccsqRpS18a6O1S
kezOPkokQ280/8Et3EscWjglR9TwpZY9vowJUkHvpL8+XBnQI+c4EwW5qENHM+xiDGv9QBBhdrI4
jK1y7FsLybZ8egGU1IX9KCGvcxUPh9sAat3AWJoV1We2V2v36sF+/U9eB56jekvnbMPgUfGbisOv
zJmY9iVxNKxanDv0PxokdaSzxopMxOl23cKlV7Ru+nausefmws7wPhD25hngnlVnhUgSsCznkvGA
lHprxPEjWqiDfsWS8DIu2j9CvhLQv/UX/gr+nLudEPQxsY6t4pkprN/EkzLFgjuQSpqG5fcTOMgx
FTF4JHA1mtZJTNOKnQELFMfmyGNpqv5uwKZvQX3e/CrILo5JTjWJN6eP5p3/d3d15g73e07vtkBc
oJgGDGEYbSr6IWwaQsLkMvfchwV+NP3Pz4fWvSwvrDpZByh1j2vKvhbO+9o+LxHBJ5QW4vZ1DYlu
4Zf4dEEk4bIN3f1nchVpFrHbY4jNT5r2hgGmQY7Q2T37V09gJNx+JI53vzD1RMgT9b5DtR56qg9h
71+x/tmahUYc47ymgz8O/xhX1CFVS/POO2s1DLtcrvxY9vt/8F4rGaKXIXgwQ7+6K4e/q5srSy94
eQKAeqXecuWzOjCRgxeZn7GR7iYqklmzMzTe9FEyaqrUKRq6+fyv0AeZb6SzRs2k9iqlB/umPjWt
Pu7P0yeAQrIRz9U+5uqpAhevl4QZQx6Fp7wpedLysCzBFHqsU8UifcgPFbkQ7sEIQfyYRt0zOT3g
fi78yZ6hhae8GsGjLse2hW2XGq+xtCZom/j6e4V1Iqk8fKCz/02ZtfmoXFxasRnABT2GjBHZ845y
EXd6MCHIGbA/WaS++qD4nm+gd44c3sqaDIMp4++D4UZXdyR053+ZvReDOlGIRhODnGc9okbVSTMM
Dh2cPlDgsDj+MivzBno50WwyaZ9Kwhki/gPYdFZkYbXqxey1ae+w7T5CoZMCEpjfpTCK4i8rk0hc
VjvwMiRwnc4S/9hVGIaFebc+hWkK9BTWMjHNiY7NxwvymQtvSapaeRJN0xp35IIW51/tqCJD51zM
pmr6K9ZWWFt1LAcpbkMYg9vxnxan4mXjVbuAwOmGZJ3Oud1nPG9GYffNyVoL68NChh0upE5kjg/f
kD1ex2S4rXfEOp+wS3LlSP6YDXLALCCgllx2zoy205Mp4zuZvlO5g/zCPbu69+6ADsFdLg90UhqU
yu8Rw8jH0of2Gzsm71lHUSFLct+NLCpwq1MEXKholHE3Q4OVn4E8N9/wqjS/cWRH7a7Qq4GXjOTI
OYZDJyTm87vj+LOStyX/F31EuvP5ditTfL/AFkUSf+vaPaZr+FavP9sYfZpwtXtZBmVznf5m9rA/
vTz7oI1mK8NZKmwHO+S5gXMY7uYTINfRLlEAPEAjvCNm7RIP4VtlXga9WShzVNcf+U+Riw3a0YYl
LkG0vLBYmeTSFtnF9C9TRaYpmEGrOLpLwgaM5UNdJOtp4wM79RbZCHsDzV+o/MNfZivHiZ1emxOH
mIfHEdTIEaw7TuI2SG/A1ndRuySDfL/TTH8lvFQg8CV+AANSusSdWfQ0yIcJiMcmgOtVFubGccGf
Mr75bfNtHfdK0kk9MwvoHoAsd3DYo1o+ZWWFoxtR3DMpLsSKS2j30OlZTbQBcd9aX2LpyDQ5aB3n
E7ZPGapiH4u9dxocBwe8kbJbf4Szglm9FszQOjg2K1bU6iS6XgFydV7Tmo1ZYk6CRJl/Qu/DOJr0
hcBrwR3XcaMvENH9ySvQlqOQDX3rz6QG1SK+eM1oPTCHGDja/+RabJCzmmGNjZZ1rnNbW7kVOxtJ
IdS6ScLQvLJCe7v3Gsiegle5XqFs8GSJQH1BrcVLuMyfc/v+4Scvy4vu4Ag2bl+ME24xBgETWdSY
Mh/D1wk7lxLPVY3GtK5B2IV+COnLb0gJsHawQzB2ohAGrkZkM8OKxZAGW/wZK+ms7qo5KhXM7Ivi
8Dy0nvB2Trp6dlNVyJfgip+RwfywkGAundBG8I6l8j7N3Ly4BvHsODb+tW7Pb7XlFBSVRqxt/bjO
PIO+XHAyryzhDK0XXXA8HKodZDe+wP1ZrLyliydHu98SWrI0kp9WrdxJswuP99eXcBH7Oj727O2o
8m6VGo3DorjGEE9358D/xjAjRR/EKWqEHmkdpGeOn0dgc3IuTUBpcvks+a/R63rJPcuh8To8s/yP
j+l7gcQPbeOrbt71krCjwiUIAYBsrVY+WvuE8f2siRY6U1hohYOT1Sgd85sncMsF/RDO4qJ8LP+3
BRS5hrHFdtR6gQ4BbY9wO33vJXTTTHtUwLmxaSaHTZnEF99Xo+9F/Gd4L7uPC9nbrysV/aImgjZ7
lDbgimUFfEe9TC2PghkxGi2RLz66LeF4/aCalNk+H+EYV63UB6DYFRwIMeQsEtO8eDr0yPvQ2LwI
HI6kuGVKhXJPFlcdN5NIqBZHySsKbfC4Y+QVYdzoUie3q1ykF78bpjHXqmwpYWdoZ4O8Yhd39QED
bghlhd6RnY6uBOVcPR9xaeq3HDfFiNAmYG9e6yLTDdjH16Wz4rC8Ifs/WzldfeOlFmk9Ldhez4Dx
wPvjOTm00S9rwNy+XthN4l2lvew40X8KitV1RU6IFs09PvzJrSZNu0+Gs5bDhgaRiksEfEG1ZUo9
kxhdKNUM/0QxFtDion9AkGGAqyWVCF6Z1mk9FNUQnx+9CEOfC83T10/hZQB9ZC9dONYyRaKYGqQI
DPef/t7q1ux4miLIX1EtIqEmDsfdiZmcuS60EnzSYu03GraivzICawqq7bY27SaMKmBrR8mFuDoV
Vj0NYoqO+/56tvUDyzXnywkDlvT1eaNSY1nxHCyWKeymXq5SKM3glvAEQdgjsy2O/DSn3MMbk014
/Q23F9V47ZkgsQMYb2Ka0CrJ9IEZCNpOzw+a20jdAeIiezdgJ7zgwyFie2PG0KeVPMdvhUtFLNRn
QniIvNRR6jlLmf7b7kRqObA3Wqs+16T3mdGUkAzSzfbeW9U5v0i7KLlW0A24wPtkmHYweuXXrXRF
LsY7tAh7QCqVK2XcJATU+w2HFi/7rd9lOk/fxjTSdB8192zstv219I1wL4GGrSuYowuRTR199kJH
E/y9z0kWX/AH1uXFB78SoxkPfgkuKugEztYIw9+KRqEWoEUtegj+L1+jWniAXxJ+IDjtVVxP9it8
eL8dbNfMEhH29nm5UDe+ulUS8iB0NKH5NZJg1d+v522MYlV10cCqWBHuH7s1ojLgYF5IoZqNlJmR
xqKRZP6TueKcOHK7exx8GjGngEF7mGBLTs5H9h6PtCb7lSt+vFyCkJejrO7lbs/jfEN3CwRmByxa
1NQCTDCuVfWCZVwGAqIERQ0Sd5bfj6vO6LO/J+cT0K7hhXMHNrPJX5jSvP8T9e3/meF0X+hcus4Q
eZ/QWDXqxvi5dzY+gstaTSIBxx90gFgMLysGcWAviC2vRcpuR805qG4rO2YOaytyiSigfbU9cSK/
l6zJSZ0H9bcCcwmI1P0kYxRsGfFhld644gQJax7q6g08D7BJ6sxXM/Ur89NGhg2MOH1K8AHtAIY5
wpNFzLhWqvkoNyBSQ6dRlZ5N2GkIcjGAdlx2h/XCEu1a5wdlk+Zm4VH+JdnKe9G7lEDvMHvPheoG
y3UmxZWk5VQnlAq5n9Dhey0AFB6jWoKVIkqQnOz3LUJ/hZoaWzO3i3L52a7MhYSKPMr12CZpLBF3
uAWsB5lw+aGrtH94KeE7ygAq9MctYp2UJwUfFDW7nh9UaD2pV8728BMmbB3N6Awx0JOxFEgcvcce
2+1wiRyPinSLJYT12KfNwklt8wIi0xvYTr9gmzjBmvcCa7fj5VHP5qN4yW9BYGb0L0jjrSyT3uyb
c+P/PSKkoFpYQiEaWemiZwJ0rcG9Rp2zL1nWudQ3LwTuGfv0pbNvoXonjvhVjmwVOcynB1fcRzKh
r+FPvlxOrsycMgA7Z4vsFpJFNg8hL9xobOR068ZefKAUhI/AnqJGmhc2CQmALZAVnQ1sp6Rxy+TB
ATwv1fuVf95xtOpxX10behVZvqkB2AWo02VLNTrZqQiEMoa9FAq3uGAR3KDqosb59JG9W/go+rGu
FtPrtseth0mX4GVp/DYfcA62r1K3NrSJ1unHmN3yUMR0ekGkuB83w7pqa/66kItGMiE+q3Y1HWGA
EQR1MlPdyG/Y1iga31yFWpGjTMkT2URxNf3vE8/9eIt/F4Q3HBwbF0EknIvcWiyWWu2zUKkIhFgO
44i9S0c5Y4bKRMwWWlY0Tug7oHulCpY1AZFfp/Mooeb9S4WzmpkYXfx9kdc3QNeHYi0JfPhSPvLR
TrNItcNY4yyndfOyPXQaaewgtLLPuOOBzhySqtIKV4PXNazzm3yAbtpt7eoAn0S3W/kSQjeGdbz2
jC5N2BYFRE7HBalBPmls/UuWrAnO2PS2rofsc5m9IYkp3RSGfeyiwKlHAB+SlSfJrO8A/I4j5rmb
Z8ti9xEeUzXL+3d6hhETDrK7hu2jmGwslH4UbNWJXfTWxlYh/Wq9YveHbl8bBiXGMiiiqmqrzAOd
I+SFy4LjzrM2J17F//OOHtO9xRW7O2KOPtvnx4mm1a6JbxY5lvjHfmtYcr48JI1qR8Jl5CUP+qVC
Njo+623eBpCaudrlaTzqAt7+2ElSEATmktacbYmFZ5Y9P58gH2qNABztyUMeRMhMI8qaRAbnBGM4
Yvl8MAu07TvroTo+sdfQLhZ5nCOkWQsWJ/K4W13eO1kYfVDbvyTv9O4vQAGOKZ7xPp1Kj1u3HMiC
Fa8yPmD0QOiXVPwiXsTwqLYGdi6bG7ENY3eNykgMg9JHg+GaI7zYKS/MWMPVFJRDgwMWFkuCrcCT
3wS/abIY/RyuZZvOTtfLYTgLZoaCEZ8oOoG5IHOVkEI+U4AO8xyorYdzbxIb9Yr0uXYEy+0UDyVB
6xtotFXRhrcjlHgwsvPJ22mw+zYFMtpBwfH30eDnXfD0fwKvj5qE8O5g8BNFQdIHkuQRUxnjUDGI
UwcAzsx/y/V3c4kkFkcS71LWrCoHFFWPPP78grDPCpZpW58xLSpMjCWme39Isa0IHduiczBsduWL
m83sVyYsPlTbEroJMxOQuJwBR2iUs7LovkCfowVgVbEsJKn0enXQPde2S7gCdz8At1TuTjxFBrId
VXGk8Q2QONm1QWUO1AkBQnysm6h+0GxmAVnXl8WiLkVCrFJEx/9RsPnBfTZzaXEtY8mho+qPu99p
ktoUm2cc6/W6R9BMcm6Dja6SSkBv6wKyMlV5O7jhbBPZ7v74i/v0KKMdyXw+U3Hs78mZfUQNnBBq
ceIjwsCII/TPRIFZTUdK4OOs/ZWdQPLSeJc2HiqGCugXmsT4XPGxhn5yDEurd8+y1zErgis79PMJ
aw9KKacMXIb3lvTEeI3Kt91xKvmKN6Vhbm0EwzQR0+3mei1LKsYXMor8PECJhAn6puyRGmHiOVrB
tlfMzwgcE2cE2t3HilymQNuJ6hKg1eCXtG7cnspkzy9d1o+TAHlFLYN/obLydUQEsCimX0IlYbS/
j5RZ9skIYGx7+FmAvzFG4wA2FFxVhXNrI0JdIyePmfxa9BpmxctnSXdAH8a5iK0/t0CEt/gMda4I
oRehtjn/KOGSIiE5YO/d1gPYJxmurzJGinyc/FdupIerwAMfqIDdvq1JVWmJnAO+BbiEcetFDgtV
xAwLOkP/N4myX0zZEAH13yP1mHxi1eH3/lk9CQwUXkBcS8L4+kiZWFabeujqvzGg1MYZ0iXVFwPu
EJQvhX42QZpH590RbSgNJW+uaDtUqIHRpkLiswH5hUL75u5l+OHbiNtm6r7rd4iTJuypm+O8y1J0
ZR+B4fwMlDFIGA3t0xF1fppGuMqMyAuNP6oNyF1PRFQFRmUpr4NJP8erOI5JnBwggts+gVZFLHKs
AE6qqENZj8BJEfRCcERqjtqd/Roy26nZbRjSNELDlPEKohezCa5IdB5+wR0bW1hby8e5nbH15PQg
oe74U/oSfpBj4LZbeVCs+IXhMziMdB8Ab+CU49XCSho+ETPfY3RtrghTgut9hafsoGa4CWioIjd5
MkusJ2YAUZyiQMz9/0gNtd2/nrCDQwDrN9LmLHMQZ+ZDLBiRr9h1HcCZ7YoDktpNbqepxIkMO7qI
0nFqhJhEsT1GdPku5p/mTYuCB5/9HmYDN7RR9nRv0LWO2alDxbKcU/ZzN7DdzYctettssP0DHB3J
bKcv9FCsDLfceXCZzsHNlYYcFYn5BEqhZaBA3VKBslXrhucjSa/MrEnerl+blTQipBwONjvbZhhe
LJCoBGJAKyUitlwGNwnj9UhZBQVHjO4FlkrIn+dyrdPetI5EBj8yZw+PmJGswJmrdt4Gj04/p7is
/tJRDwW8HAXmWjsV44H35d2Vqc28ZQM+Moar5ZQWZF6cJ3Nyw3Pa1ks+/u23RzzgenEyCI1BSqFl
1w7FXjvE/UQYiNUYO/8CmPvrkA+BJqgWzrcfi14RJ8Iq4rQpmDL6GB+V+5Dt3745b+vMx3KN+jWq
TWAObxN0vKOTpIBC2TVW7uu2F7AErlLLlucXUSRRhkuzJF+mWBhqS/udDa1DKpValSk0QOc2pEmg
HKsS+UZP2nzriB0G548+GOVD+So1LAW06C868vcGFpP0VlYFVMvguHe3u3iFC7DCi+VbLVTTk2d9
OzV5OZUbJLddmG4r5Xcpsnn3Ft6knVZkvpw6EJfbh+kRhqwLAEtax+ho8z+9lY1GzLF1Btf803+u
QTMyYZDB0DF0lFj4W7UxzWZq3GmtmfMwzn2rbq2j7rtkpm067PqdvF6WJu6T9WoGa8u2HN9n/u2H
ICPwOPiXn0gQNFTcUfAEaQ2r7P5J3S7C8gWkt6VMwzx2TrUdRCDPIkcOdx6YhOkL/vPgdCS5b1gw
wl/u9S8JSmuM85jzL/jh7iAj/vPk6hpxHMStsrHTyllySZNWNNbC0OCk6vh8ebGfUeIJ7cBpUO+P
PJ/hcWPZxfwRCmx/MfGdvRuGsJCbW2CcXoGCIqvpW08Frcqjzw4JF3L+iK3XMuqGS9dy39N2nX8B
ncqN3L8TcMFndXRr2tYL9/VG6rn4PM40H/9goS+WYB59GcyDOxmWQVumR+RTIoHG7tSiI9+sRgjL
KJdaF21gP6MP+eetA2Q5MSXsqrT78PXEB9S5jtpvymoDCqvOJsJGP76w7VufMr11X8rIEdS8UerV
lpfW4j0kbwdRDYW4OWGwEJp6M7JD2/odoj1Bx0sY4eI0UXvXVTCeDGIbP4d5Vsi2NceD1Bz7pRnt
RmSwcXRN9RWnH9it2WPzQRQxiL6zk2rfTH/pvBpL1sw9D5as5hzupMZdG/T+cEuM2nLfpmJwjXzx
qrhC6bXV/P9KKUtZzNtiH2TXv2MRFcHaiTMOfib0bAcUN4pUl/7j0CZYoAPQ80Nyop7WQZ3uP54o
6vSn7ex6Q10bpcfoAUixEu1aDZ95MrKkB9N/feuwWaS6KpK4FTVU6ptqI76btIvndxZ5xIKxtW2Y
7lmaPpfVDljPFZRgR6X/aK6tmr/4uY7c/6+WoA6T9cKw4JT5YAMUUurM/lrkN6j3vjPnxuQaCnaa
v/wMwLHmGTSlxK3fUfFvPC4yylYTzyzteoYJ0BYY12d8m5OkLVbR+NY3oTe9E2hCV1bza2WGe8hX
L+/nNWuDsejkh9jnOQXFFbIDfMSeLKfQLI8bGpeRpRNBKDVdV7n/Sk8ai0K5i+C8qbRY2FQ8orM1
6hPchUJFdfs/VvnDII57Pxiryp9hnYvcoZFfT4/7bCJC/PyIwWS1TS/KWzARsh/z3J3O1MXjD7+I
kq+/3jRrIQcY4MEJybqiWnWMJSAnB1DyjcXf3GEajpsPh2WOCys2X6Y/jL+CU2bX2jbqhsCR2o91
HIBB4MUo9GrOaaQECCD8EGaGev13wytBn8seUI3kT8Mz4A03elepUiT8axvd4V/iI5QntrREZKUn
EEOlElxQpAqKcFdLC5a9o8q591PimANU5tw/Sf4o/NicmR19Qy2LrFptQel7cUXWCLPL1otQ6i9J
M67HBYbJN4Pup4zkBbjvCNf/US3HflqokgHnc1DfPLWqwrL+dcigD6bnIaU6Xojm/YapmjkHQXB0
yfAuRDiprcq0JajV4Jn3Euotk6tu1IIwzFNJcGIJ9Y42CxasrBlvyUv8L/io66gc7k5qmo2hhx0S
FbP0PnecycQjUpywX1Jmkt3SIVcL1ZlX9q6Czjff5yVV0Af0kmdbUjuQ6j+N0HAtm+NH8SWfQGAG
B7z2EHzKe6PaIq+Z2vLYe9dErsvMUys2d1Y0Ju3Ju3wGsw/Dg2KnEXuEHlXqsjfTKqXnMIFoHScH
Pd8fgaY9hONGthnmMlB0pstEZbiGc2LvpuQLrjdxvkfz8RsHtbGyO77dwyc6WXSV0Qpu7wI4uwfJ
FNDHAtU6SSwcWCMen/CsWJ9JfpeQH8UF0VjFiwXaDX555e8h32AfaknWsZ4yaearYMTEASc2aynD
71HCUYTZmo2QXSsjEuHMc2kX6J2MbWsG8w5Ql2Iiv9OjjEZPkNka3cY5HRz10kbUxeT9MmIX51OG
09YpobCZzHewtuxEhZ1dJb2QzQAzO/CpNnIcjxIIBW1nkq7XyAba+NFfypnK/ajXad6ENipDxrub
9zws5OKvt2hIZ+P4kcIoHKpF3jow+jQ8ZNjBnGITnbxJtBRAJ15TPVBi63GDvVBwkD9qT+qW2yuo
tQtVbbpf8axiAtVqB6txhl+AtUva0vwsUlL/IFgkEHmgPOV8RruVFnZoZEhTv0Rm5cSWpscuKV4O
q9ustg9xwpnSE9vLjY6Lo+MbwarJ0K+eFQdPBm18JOIMp5JwNwO+Lly2hLd+OypRcpsZcOzyv4RT
VQrkbBMQIGsXh8hYf1IV49XOAtlKr4PVzIDsqGOHc2D5Z+3HPgo0Txy1wSHrbGqdugaZP88ldkX/
p3NuJlmFD6O5n1oyvQ/pDo80ruisrUnNNVS4GHLr4GjHzMNZjGm2kTljrmVn63i38PTId951Vnp2
A6V8sRx/wfrynzBQgBlqok2lAQDjgoCU/thPRmnHbB/uAt0IbyIT+tQvcuOuySTJNqjFBwrI9jZD
8vKQNVQ3abpppMBznfXS+f2Glo9ShmKnJzEQMLtIHCQ7YDieLGCLNaMQ0gtl7f7ypF+4lFR3QlYO
tAbe9APG1Fa4ZnZ07y/jVUR9Gm3P8AUZWe3t6+k3S7epIbHtggzfc2yPfsorNCYPR0QaGsC/1DLL
Q8UHj3f/TChT8Ve5Xlj/a+hAniQeR7NH0Abldi3B/a7cZkwP/05iHL8B0f0y49cFoRAUX/om4ftH
gy8YR2FiPc4da0tZNQJU6fGSrnoUcIY0Mv/xxwE2n7jKajdLt/BayH26D8+/bu7kgHNUJzqeLfjy
uhKTVgnXHt6+HEojd0HHfP0g5E4w8okJI/SqQ+tjGccB7pm3FMt5/rdzu6tZhmCLQyTiknw/YiOU
s26Tc5sASc9fbIlkRZk6cTwDhDHcHAmQ2C99zPKl8y8P6hL0MJEZUQbFTltx3R8ZStM6bKzPe9Ft
1HhafXgWnBkRDhC8wH0+bArDFUpVtAPK3nKcvN6gKv0Ej8LDTmd+I9w7cXUlCwFG4VrqmusoTCh6
sBenIQDiTtq93zj+03ft9EQXEXsr9ruKwKV0cx14zSVF/MvPRjE9eEDsRDopljNscnoYq2ZIZliJ
7MmLyIOlzZvZL6plAy8fnVsdgxpuuFs1QPAeg1lroBK/iFgnjTSakkwaRseRA0xwinKW9wyIedAw
ihRkZ+WgBQ3HqjZ2oBiLgX7QtwXYWIY6C2dso8wH6rCAuK56/KuqnwxYzaCrAXq2M0aTfqwhWeg6
TfBcdQDsNBoxXRlUd7L0oE1+isBRxTvsID+bLCvJ97T3BUwNE6Tyj/ExGGo2is4p7mEjGT1LaC2J
Uf7AOd5676FT802ULTarKyPOC/cq9t4myUfkOAFCk19An+JtZfaUhrUbW3Xs1U57wSnM1qVSF4Zb
+JbWGuV7tqONVZreLHeJ8/eJpqZ/p9UzPQIWGvz9eQ5oc2vJZosC9HM8KKauwf0R3nyXwW2CMfqw
JJKyei7yHTXClap7cKD9UKXJG5TZlLj7aHF8GPVSHxIUdmDX2/FXtFZtCQv1pDyP8bLobGdKNYTq
Llw/FkgLPKKBMbt2beiHzFkHjvN/fJCCiETp+65RwxZHhuz57g6lpZioKUKDMpSrusNcFAnH3ZfG
2fjjOCKLf9OAKswao5wciD8IhPH4In5RI1EGv5Zrv7a3+IXpe4JdOiyWvoz/7jhJgdXIvRTm3Wbf
KIqqv2pb5AYW5Afoa7r2HASXqk7hPhMG9s2sJ2sIMB/+NSh8NhcO4RrM/QvQsC3AL0qxCgPUmAGJ
/xML1IWj4iyIlWF9WZkRljUWAdA1kkQrUbXB82EfYCecTBTEgQw+FjdVPkeRuyjZdfzHUFnytFBF
3wU2xLLfy/t+D7L+d0TWRtI0abxabKCZ1Ku+1jDoStNaVNbiYDUqzgr03qy7QD2CWs5T596O67KK
fh90qK3YdOhCueu3Jf6LLLeVa+XoR44WAocGju8OXZzE7ehWvBeGjWezGXUoHEa0HQM+JWfc5O7Y
NIZ3PvmGqBztQvEewNVRM+djbfF9r8zIxG0flS7HgLUSjfmUpbohi2BsZxkr5jstcsqM3Hp7xzEs
f75yDHygw2yUHOKAnw4f+Xblhx/gHfrpFwrGnIAfo2gimAsww2OBB+a96kTr1ddhgGTCqEUv2uUa
AL3Mmogfygm0a5Jclm6Q+SZfLaUccoq7k8bg3yNXJN5vBRRk6d4qc/RZrHQ6Zoqwph8zQ14yU8Fv
nZBSnGu4e05TpcuekRlh/h7swJXEJN6rL22V6UETl52MYhkDAK+uKd/p0tGgE7hgM0fEyzrCqu8L
yqVBIjB/YE3s+ierfSQGY2ovbrAWWMROH9m3N9k3cJ3XutI6Eayqm30k5CSKaoUNvGdFYFle8Btx
wuHKS1nHNk2ndyxZrIrrD/4S9BBkN88UQ4UaE/Y2rq8RXQ5D8k3aE3j7FzL0cMc6mTRNvo9yJ0Hw
V4N6pPYF7VT0YldEtzYkWlZ/KkriNdBRSEFQVUxemHxwNKwYyQ27RehXHA5nOHABMlYtwYVrqkjd
jX/FkYOn5PXFF969C1EWdoXFOnVyfQElho7lw/aWn+09i4+iEav5yimvJDvg8Vw65zi2Km6/H3cH
hhBnWlQZnvfyYZZhKN9ZkC7wGuMpH9CsYcQYNEaWtzo32eBoSkIfqGdtVnADSB/lEMBQo5LjMbu8
7warYd5raPRrPtnApjTLToFj87KH7JkUlFJ8YyYyQE6bYCgnhbl2Iv0v8LHENGMR2ruMnS5Az5GB
eNjADpyThEU+b2ub+/W/wmEMjbcSHhDQElBD/EDdNEl64dSVijTLSIvXAOyhZnSXMohX2QIGyE80
itQqAt8P5LKRG8nT3YfilgbY9XtoE+Uh5ZlDrD36BBh5KLlLBZPZyAO9GFwn+Ubv1km/GJevGzs9
ddjyFM7BK7l/gnIUspkOPvJYUCnkYtMupykrQpuuD1dgxLLlJAW2QIP7FYTOAsw6zkTTg4nbqOzy
FGaDLO9u3lWuSP/YEPAziOCJA0OqtI1uQzzP2cOvmikaOysbd84Eo3M2OQLr4UZIsf+qxdkfn+81
To+/Uy5PflMoObCnBoO5prZiU/Iok/Uri6DoR2Yu6VGgcc0aZFHvEr6y92EJqSzchYx67QvTEjrl
GwuArpUnkY3QeXmZNZMjOB3Trys98AwxVjHApDR0y1+gHT2yrZ/boi5fB2Q4VSqk01py2bs4tRXt
fYT91FUiLmagPfUTTjVHXFISDcsZMJYTgeedBhh7B13fBrePotcq0kOt/+YVIVZDB7cmHJtdXVIR
rdb97tuUDnZ7j608c5W4kLDWXWAxJLYfJ+Y3H52pqxDmOB/1JAEOAX/rK/DkwwJtW3OU3+4+ekHM
VOpZlePrcTEui3Z97Rhw/Ys3pwcv9HJFMbzJxlT+KGhJfxNNGKFvbqPQi2Js2M9JkdbfD7v4llQu
j8+SIbE+jfsVjYnF6NY6UEZHXl4tUKWa/q/b7zPrtE544UHQ6ututlnIWJ5PvYtzCbt9zu7lzOKr
5jfePkUIzBgQokV0JCMruwE5zULA9Bz6d0hbqEDaLDtBrXMhigdVCxb1+KECnH8meeiF5VN0VfbX
JLmzc3whpPPUE8UJ/cyThBrMckaeA7XWjwSEMMT7Tz5pcCdqZ9M1PsrRRgRthIoES8/SSeV6ukC7
FFTNCWEtBzajrsURdy5GYCD6H1z6f2TQXYs+OkUILjTY1aIPgLTvQtf3L19bdVk4De2wqjJey55b
Cuh5XTWZkeAtS67KomuNnRMiqP+bYtQoXx0uYAH5fNqX58ehvYt6vS/QPrcTms0JLCs9in4PLOX3
usCty36c6Arn8zCl9Y5o9A34ihb5FOsoxZHAOSBFO1Y9j31va2BZMzANjvSrj1JwnCmJiopjnYyz
f3qTFTRoBHUlLNi6E4AA5t92sDq0Tz6Yq8XjBVOY2ebFnoJPNNG1kC8pPi+vqSa/fuQzZ8nOzFFz
orY+qvbqRvTChEYxIrPgg01jb7QkIm6F8zlOGPtpskY1fhDudfKuuW6xcPQxa1u8rwACdM6MuKNC
8fxmSLrlocXe7YUn+6fJO/TLXeqkO526OExcxe9wf6vAn60wLdzV18VGOmg5MS431+CeESK1LDBe
W8m0aR6nzA0kGoUh+kn9f0QLRuI437b/7A24jIPr/poeOQTfwt/yVQNo8fH0IcxPP8asYbng0RM1
GUc2+Zs+k1tYHQ6ydpoNoyejW2Sd4Y/u7jNQ2rL+GCmINx2it8mFHq8fVst845bphUfiWDG8e1Q/
w2eV78z41UbBeOIi7feLtVw4h+/GNJaxRbXZRUPwt/hlDkn9QWhaclns70eY5uFGK02ssRTLWbYU
vuizBde+5bqq2No+itXNkif9+YxQpZbZXM2Otb6k+OR+j+PgtmmoY3MehXqp6qPqKnJUOR/KPNcz
zqk9xTLG0ZQzkuxtkCqPJ5uHeyzSpF1aeIJmYNh67atNFX0+BLPWTzRSFcgTHLzXGq57waLcYmom
wMqsXf7skSe9T1QyrWhuGyQN2z7EgfLqAzfLduHh7LI1lr8iCC9laUxm2fFegmVWwVkfVSitSR6W
zfqRkPAnBsib78HqEUBLuBIq7EPLxzaLgOf8EFHCogdvJB2gbSWpaDHRAWf4FnmjBeH3dq7PmiIn
ZwYDlbMDceuF7La79D5ryZz3qp5MV39j+QV+wmYBQar+pk5JQUXSa9+qLlnZJ6Tn+YikV8TZTe0b
AqawBPzgWNgosa5S1MBnzGB/cTl5rhcaufPARAVLxHEZ8aFQPW8pHvkchP4e/Ki4zwr57dQiIiZP
Ru4/YF35WwG3v29BOTuUCO8XMiGYOj8wzAWmto5LYBMqjYZC5QYcnmhKoTgw923G7koWhjVlnfrY
7H62tPjv90UnykIp+eOfdE8ZadQ7p5zG2Yz+fkBGkhEK7M4s54f0JZ6Tcya+rXAWZYOIUZZb2o2j
68fHs01yO9qd+hfFcshGNFnnIfTJmNcJ/M22SWT1mdksAinM71D0fKSMoCw0SVaz+p3x6QDXcTjr
dMpgsvpypImbjnq8O1rmCpt6gXLB+iwnH6dlBDpT9wAtof+a76vOkD27jrKabex0pIxiybxucvjB
EqTOkU258DctxfI+zt7z4+tXcFQTiEKMJnKTVUZvNNETXjen/D+MbqW8GDXXsd3PVI7F0WsEChQv
4uKXHMSD6folJgXeHAVkyMk0MPyFQX7lRLshihzwQsL8kNtousIWFE0NsC6Ko+tsrd77JMX7ejcf
NRgwJpao8+XbuWXuDQ4vxoWA1TgcMOMgcZnpuB6wZiSXhmx30IJJRiYtz7nd9pe25GNVho0hGl3l
5qUPufyw9Af8zUOLef4Krl21Kf1IDrHTDKYn9lT/D13c8c16+U4YkUVyo7NfeLhxvOL3qqn2NFVT
+HhIvMr154fc22imH6AqX4Aa1NxexdGE/LbcBjHrh+VO3S6zN0Kre0jp/jFl0qR0GoADWaMC8QDa
9Qu+ID9yZG+qMxREDerjEdA1R2TyAXHqX8UJ+ZYbmm4khpEsA8hbUb9z8ob0PXpV+cBaxc4kN8cD
0JYglcGI3IzYwDh5a0Kry6oZovjsqePh3QRrod43ruUorrziOU12DdfK/iKZzmpOo6wtTrkTox3M
d0vP5abPceL5X9itppmSF9wzkdzCb+JUKSvVfxSUBIBiwVXKEqWBg7D0TznZZmdCKlXETF8VlwOQ
JgGRzPnThyBRse0e7w+niRwhNxn6UnPdZk94SwOLlRiP6Fp8jlgVjd+Y9u8u21ozsE90blDQiNKl
unrhkEGpxyIhLrSQAGowsLvUo2ccB20ZwCHZDqifxKxsagqCGya3hu1yXxypk7XPLRU4cnEvmDqQ
zk2SD6dqKYxX25wcuUeo2puQdGIqKOrGMlfm7TKOy+LQNDGNGL4LKSHT91199U6fv0q9JsDlp6fK
BVk3HuJBM5X3II/lIoeAMJ6vy7dPgpI4fRq254VWMqwGzxqqhec2iFFuBzGUCDPUULJuAt/BNruG
a9mGw7qAG7ZRd6excVhWYQJdyRic9URZkddiB/fyofVZ/aHVB/IZI5ucSvnzkgbTCLMbhNen0zA5
xhxzo+KqudHuTdWg0bC51EoZd+0GBaqHrgZ91Smr9DS1HQUS3yFWyyPOF40Kw8hdJcNGB1D1h/th
HlBUHlsyOqP845DJqTUyY13zVQlwQFkXe4ak1gdOMqsf6+5Ut/7YqnIlCb7uAnUXhVHnekStYN4e
nPvMJoE1R1DtU16jRZ+pbhgIYenC+0sKB2A/SVGwHl0IYI743AAR7pldpSA5fXcexNDFCITK1DWt
65XDYyjmYM2NfUgxlIcMxz1YBi8vHmfU77L2RaWGN6TerhqJtxtkec0kj0/NE1IrFEILKTx+7cjs
bchT8J2rU6FREOsjgRH/0FnNk4MUgLaQCbWRZFCG4fXYcDzcJnVEwHoxt86VS99FEBvmgQKs7IbA
ljm/0STJdDIzgyhA3TFfxl90FIHRs2Uky5L+rwDA37k5y5IkO2no572waVsY+vLcPsqtYju8RmoH
jrS8zL8ZgevgodBZUwer4dYFHu7BbNYYnUKoNhW7u6eq3+u65sSlgg6QpLlwqMkDqRjLjlWQX3Sg
fVBvSyL6uvLf1/sDSKS/s00ZX6nUTuOk8MH5h7PNsVRS0Mj263qwMxV2TJ/n/wWGnk5zrv0Xx2Vb
4g47IzbeK7XcBJCTlyWY/m7GgxeX2OvQ9Yl1/AYC2aW2oI+e3SeWaRG7b/E6/XLgOiCNySmcohHo
YnuUAnckFN3LsGaJr+A5c6gPG4ii45bN+YaHsriYWbkd1cPM4aElmcdSyAP4FEL6nWE1XpcHo7SR
mEpw6hnAQDnak9SnPqDrdd8MQo8tPrYBHFaRv6D8wUTe4tUToCokfI1xFHMW0EJvWPv5D9fu36g6
yRDOqzVFcaCDgg4/3QGA6uPZZ6ACR5+aa5rQVwL2A0y2se3aSOYGBLvZT5rSu9AsZaPQr6QfTG+K
ZhpvaM1ug60tvP/nZd8NTAzksyoxIavgMQMbrkGpWgJwJVQq6X8rAjumek7ZwKkbnbs2enk2PoK6
dUSkYq9/P8a3CcIzGAkLUzxPduUYc9YMd4WAO4v7fllHZuDzzinguFsmvXv99zld8vPP9pyQlyAv
JZSma8NmV7AOFp8j7DQ3N9MO/eCskrUBdsdx9IzQwjYp9/A7q8ByTNuosNqBDH5QdG672fbcZEm/
TzJlybdD2eYJTHdVjnIEbdMnl/Z9vwo/vsa/Go37sx3OS8hEcEsCzltv2JmYa0mINvDs1jql9fHL
atQyJFTiN1MRNp2iFwQT9ltu/kGlN24zE2xdeS0CNVvaCIVLuocpTLHI9SSKL3NiNYZ53F547o2o
Ie0prEN6evbTzp0QIdoN/nCxrC6gxMTxvL4PreMBqElyRRKICzTA+UzCg9rGVqpSKHfW9o20Muj/
sx3eNkX5SeOc8I3hAUQYeVo+l+QFi06x4KflUtGRgPr4m+OQ3K4O5+rdMKkh8vBgM/xVRNlvpInq
MKEdlA1rTKP+Bw/CmLmndzAC95A7noP1thILqShSSQbOpfNAAurLk8Kv3RuX0zKc2lMyJdukViUr
O3FrrasY8Q7UbLsXykpVl8VIOIIfYb/QBID7wmOFVzHSflhgSFvs5W6phyRxYL+laoQVjrtG2uo4
C94v5PWoUk8fHOXcvEWc+rmlOys7vcUSR7fV1xVeSvrC6i284uvvgIo4pjfdJMlWc+i6zA8XULhR
hxR1u+sTuW4R6Yvb9+z1+cB3KXo5FduB18GUzg4QkE/lkhAo8UtYwQ+0BdoETeKTuRZAV2QSY+Q0
QaTpdF1XRx0DPL9IshKHXUnOcXnqa2UoJsdfICR1LCCa2biP4b9dIlu5iJOJPPsqdHlH36uUyO0T
eeBU9ZaGvPtwvJqrZ4AjxE1xSX0OGuVk6tCb7n86fzbOSvSMDMbAHEwOz0c/536zoTqaehTSX09o
Jel5jFH4HNDAEsiGxjoGZb1dxLgHCBTAlG972Xzqe+iA6ZJtqoPyQscWuybc3jvG59P5XZeCVFq3
H3aeyEtVGKlmmSizsot0VWH5n0EB+O0fk0XypGuy9aoYO66CCxy6vyEG1ABbbMDDzm9U37QefNM9
n6SYAjJYMI1TBZNF87fSlf41+GhY3OnFy+mWi60BDFzIHxnwYd2bx9Zii1hh51XXeguSTy6SQKz3
SQU937Y1qSFbILmOJYeDh8le3EYQvTBcLujcr+s5VxKYgvUORZags0gVYKtXNg3LCVOzJfayA8Me
FF++ewKnW3BoJAIHpYW31BaAs4/+RLSdHW/maWefDSXsw4YPV+74HuOVBdOD9jv6ONvijFsGZyb/
kyrLKe9X8ACkeqmHemWiZUVmJ0yYe3yo7Ug4oXlHFrVp77wOYNsUDK68ubZjEWSSsbChCt3vhBUc
jx/QzgUtUgN2cBgScxFEY2tx6g/lZtYefzf/54MzmI+UbBB1iirSiVVwzUMJ3e7pA7jef8+v3DVs
MaO2PZT2Hf6uORrPtNgPVn4CiRMb3CF/RHS4Llc7DSbacSpG0l/REtx+R+73bcdbBQg0b+WrmF94
074mB7ejctj+VJsBXCG8VgxAqvvTHkdTrW/+KosWE5sGkzHx/NuM/2HCRngcwAudJyQxNffhmLSw
POx/gOe3ZGQmpp6qFOcU2v/8Pq22tsL/UGTrvcyW809uqkrCxnKBJx8I4W63wmBZAq+tO2SjfgxG
X2dmGlv3a61O5ZeXJfb+mcPi80qQ1Fmn+WjRM72kaIRkxDonarQo8tLPROw0c9OzCSmA+XghInjt
IzlkDt9fA8wdoQN6eyZUKUtYAG8Izus/sisxqwG2P5NBAl7O3MRq6hBmUb2cjaR6jEU/hrFriAr5
0bjNw/+29pflruSu+AD4qsLox1fTDCcLqA1D0d3v1ENCGjsQfXoWVryBr+hr/Bur38UK9MqnXzCa
WKerlu1iIH+9SwAgJBgo6nsqvJjmV/2SZNk4lRhzEf7Uurr+tcy2MNI8EoxlaTwDIPwN/9gHJ0EG
/IEQsH0FFOJt9szQXh/xFBJ3uW5Vd/DDUmCIuaPB5fVIrAsr5B0SzLG/MN/7h/D/0CrC4uV3Wl8v
yYLQl4iC3B3bI3ANqek0S0H/D/LgTGaJI73EuAha3mEypX+u1UWbNG96+r5uUuRCBohwTPbDNY4e
6tSfV1fFtyd5cdAxgtKm9sx57LLwaSTWdhR6ErEnMcskjsWdGT442zF/FjCKCaoclfXQyzHVheIV
8PFMLG4PsGz3H7047HM3Git73XIyzhsJq2n+xejT+qd70UUgG/N6p8qf9G4lInB+HsZQuL1KWumk
IxqDPJwHBsiI+MGfMNvFXH4ZAK2T0F7ua0dB8pl0pNANbe0nIiSNpb1zKPimjxXkIUQ47cL4GX2E
gguCy1dhcBRS+VUTNi3Y0a8CqK3W3XfCS4MJ7uwGpMrT3855q/ocm/hDItVk8BGIH2s+nr3YBBG6
dUC/XtZTJCChBUnglIRH+2pqD0+IOfnb0ncqyry9gqej7CC9nsf0sJsv8j+pIqi+wHuDv+oZckK5
N30dYUZgNzaEK0SxFxmzuvrvgzDgvKLcmY1QUEgC6uGnsQRV9RQ/Wcv3CDDM++oBb+lYuqzW/01G
f2YJP5enCBK6f22cvcdipt7cHpslX9l/uufLzmDhQFh/lD448ZS4fyp70pawSxO928BVRGL6xr9g
uzfAXQ6PnTc6FJLR4QmFC0OfjSg5L97t0xvFKKywkIImdB6mD6g1KQIgqjN+lFbYVWrH+wP9Rc/c
wsTBZkJRywOImw2Q8cH0Zb+BjzkCs9BRJUS/98XHS7NoLbTB5u0oTcCpk/GztYnRDQoPLyUXDeYN
+kFE3xYmmhPi/WlqO6dxS4Tgy3Gg7h5uN5z0l3N+zkgWBAhOdHOVrpdtL4/v9sQkkJdz3PYzUhxS
KKPGUD1+6XpKczjufGJWwNR4vDIvdzR1LNlvUljm2lQvb/e5/nzMOHBpi+dZz1UAYTPEKgAbTn9V
qG5u+anmjGu+A1Lc1cu3tQtX9j2t1MlsGkwAGnsEdJApQbx4Sp2nKx76hrTvB2lPGd6/yxx0JQxz
ryDFyhExX1EC3/Ea2A7/wAcUQuWkQWcGSoQPIbmc3wKPKBDkd2AI9OtNI3E/9qdmzYh5Td4uDOHz
acvrL7IWFsdqQlBp56YaZj5m8eJNs3DiyOuTlaf/MrSHLXJqE9lnBtn1H2tGGd6BFTb4Mh4pcCe9
xQcU0Hivp9SpNkFuGpsHw6vQZmFBq8JWLX9VKamasH2+N/MFKsQ1jHoQuzxgEr7f2Y3xla9B0jvV
8hiSvDpe9sHFpMzVEVYjEdgXvnTauUATL9C+B521BVv4T1o0fZ4ZY47WDoPLghiZPl9bhm+ZwzOf
shXFhX+nz66QYlwyTPB3GtQZQTzoqgMkW+X8zEW0++FD7h1N1Um7aQ6na66qVtS4IH7PE0//8MVf
OTfCP6UCr+UhRpTuq481GyhBrbmHNQe1yhel840jbS6SmZqNc7zjUB/yUVRd8JcNlChary+Di8K4
q/MvjxVKW7k4fvGiGsmurZpmdxL1kleKSR8m59OJ6ZuTqc7Bz1MnsanhqUrnO3EdqKlA/uY0QjXE
lTR2aI9PTQ1Q+4/YrtHOdehdMmPMEiALfAjDckftJELa0s853R+90QNdg4qECEq03PQ1sRMm36C3
cxBZ6vLFMVkUAitzg33bZ2a8PAQX3ja9AnXK/yZcMi6uogCvuLCIjoD7lwPtvMQRrUUlC64ITe5p
4svBjVwQW5Y4uPr35s7Ntk/SEdkBbYfNSOGRDVCFBQ4fyMc5csWEaBpErPuLzK6Q9Vc/gsWlMXQK
vOxtjZ1jUJh1Na/0g9YzjCAdW77n72M7+KNuluYYh0Qp5R+c4Dd2AXIxqi4DMuFMu5KXRv5c31EZ
M6p83IiIjg2juaB+GpvS1X90O4exEIjGTxy5Jl7hBFifXx0TnSCbFl9qGkSi/3wDRUI20/0Px9W8
uOMaoAqMTJcGglBCsC4J1CKMY2hw4zBVCRjgm4nwBuRLhuHjgdFkehWcRx0eX5ba4OVMQKLywtA2
PJD6SwT7DGRwK1reGQpKLKZ5aJ6faQbcsO/4WKLtbzCmi68NRYYrel1m+d8XlXWY7De+2jk0Jfgd
8kO5yW7wAVNXpPkO4CgF354dWb3sce+QEbxGE6B+DMLBeESjYrxfIic3Qpwe2EKtGe3w9sL9TRgJ
IqBsdHiCGaj+XsaA6ivlA7xM7v8TMeCcQiatabGAArMFsTt+JeMRyauC/Bq1yeCav/2PfHSZgK7e
Jyo0j7q0UWzyyFGhkdjT5uvAZpbCYjyRsJHREoH1rwssJiiLhgFts9jmYwWj3Rxv41lGc/TXGsrZ
LGUFs1ygd+LU45/9W6r/2bBNZqyKfJLuPcRsyiyV6wKX59pGZeJVpK1Bkvkmg9jxUR8W7VForzEm
+O28cVOD5IuIYBZA5zFEzphiHl8lgzuf/tnARguqZoh083mV81lKnijeqhbIJL9eDdMtP9lpr1i4
poF4frBQBMGv5PrLV1YogHw+rNTJQL5romKar45D0mvbxSvH1I42CNNoTXm4fOE38bVpmjtBGoBp
BGbmE8oQnZMBXBtHQs94tUIlnCG79gcaw+mprjMzc/rVundAJsfPo9G4vBkEtyMc3VX8N7MCKy7a
1l+w9Z4JJP5H/rc16ymJGjLxDDf6SGKhcumqsqD1//OvxElQNfpFRlr5GL2A6Bdq7v1pwHNhspUc
Yeryf4qZICYWjNTRZSsZAQ5hRZIzE8kug2GlYPU92Bl1LigUudnXuYKwiIuV1VAB+msp54ec80v+
nNr19q66IZFyF4nQOeATHDzeni3OA4b34DAtc2tYjZMIpokbbKALtxb1vQEj3sQ2h+rknAduD0T6
gs1BfBNvU4+buq9PWEQ7V4GzgelmliZcqz1/O7mgkltPRjdWSxxCNoZVcTdrmlZt/fEalWtrMlav
LKmcnpi7SfFVT6j+lmdnd7lemmhxkfRSy7H4gbp+WiLZ20P/RTeyKAtqy3FJtq4H3sAXTOrUZCjs
OXz+FfPs4J/Mi5FElygH1D3N1ml3+a+0J8WESynyV8uWeWlQAGjkY1fasQg32anX8up6UStFKQE8
p2k7e/dBGYDkYYaGqfj/NMqIsbIBZgRabLk5T9O/+t7+yHV8dUzn33GezFlzeeKnSPPTfBu6FqnT
/mHfRRjgfjO+Hvyy7s+M3C42aYVdM+bAEpBRH4tinkoLB/yFQ4Z9FIEnkJodbdXtIC3YPX6InMrm
zANGlyd/MSmy/ZegWs6CFq1ll4mrRMmnLwW8NLQgumK2iegpcr4kz18mpSdb4uz3gvk3T9KQ14Uh
KVpI+ddtZ1zwmROlAmQTJG89niToKw5InEVuzMUZztmIaKd1TbjUQXqOoha16f5hcx4yBwgrRPNV
oEZmt24ZqRaMobmttEsP42EeJHL62UXTXNj5794BrRlc/cFGONcg93YSs4irt4WuuOV1BfyirQ+P
UZTaVlTOdU/uikSCgv3MgGsyd6YJVwlZipOOkTOBvzTHHAUwNlCPGkI7bc7T3lxVzKdVFVXRifw/
Qt1tg/KU4LviSOAhFo2b6B7DlregQG+9o+umQxyiBo03LjAAW0ij12kr/IWSydaFoPQyO98QcGpK
teG3G5+XHrFDR9GX5orYTIU9p/wGdmhUw9xQAypzfFnEFydI169FndiireyaIb7rAWdDZiET1sJe
5VmwDPBsVgfWSbCt6zF4NHd/Pe4PzGrLlJy+VhBn32WON/+H27Fe4Q3uGePsiPmAdq/X6SqZtE3A
y6t97mJB4LsTorFjHBSiBIWLtWi7ciPqQlcPckJqilFOa24PbtZRNGUEV2l5bhe384gkIeh74BtQ
68gMJtt8PjYJZ0dbZvtgNb6Qjd8r1uw0arzRHk73oxWMkLYVfaNV5s6jy5KFn2qpwqjZBjJYjuZW
Z8fRlIKXWT/C3MpjiXo5ngyxcJiRgJaNoxbcwit1IcJJp4xnFIF8T0GQ4z+NGNtyYdp3PKWYO04I
cZ6djDul4xftU1ZGFoBircPyV/NOoxCDchj4us2dRAH5dLmnNrd07jAsQr8XVHjR+tA4bem/oVp9
rym+wuh1ljOofWsH4VecHWaJ12TduYcP6MX1Jfw/qs0ihn1wSQQzZWNkWOkPiwCebFcj0YVgKyYM
ZT7DclfSYbVFK8nmjwGqHv5YueMParHbDhOWkhT5iOq+vZvHsl8zoE5QQ98W+mOUBA1uXo3Y5BaK
zXu9NymVzlnCXynq/kRXVnaqBgz4bCAeQcuDSIwVMNDgEZjyWkuilmpPwary1ZljpLrmTazLLpBn
yhJ29s0xGSTVYtuxdrJzW9Kq2a6lA+YxDiRMOrg7KYuiknH4gxKTgcWBT9U4q/PCfbay9SUMiXH4
i9pwQlUN1fCfWTR/3/wXrXLZzLzbNY/7LC/8Dw91KqEMLrn5elW+WjDIaSzxi1M/lgjA3ckUgwn/
FRo7z9hpqsog7cQUv0ATamDRsZCrYbJRrnQ/5J9CksWkA4fICAxq+EAY0NCpp9IYcbiDX48TwVfm
0mso6PT3XqODQnIvtiED5njot51RQAeVlVwUBND3ts7KXWmkaFCXFbztajO/tDss+KjDAkdS6eef
mCSgeRpi0tAlWRcU4LjWR3hGZLiiibgNbSBxjj0LvOfJjNlDtmvqqUMLA++4fqvx3BqeFflw6xkR
pdUYXc4TapcY3BfEWju5Ka2WDOiuPKIcldkwQS6eGmnWlZBUYQF6NzSFiXTbJn5AVw38H21J2Blr
PqNemzGp5gHBwgCZMO4gI9K20klc0/8TFBm/mVPNsoTl6ahpz32gXmWXOChY2BJwm7a7zDPigxW1
Md0axJWB4vf3/jRmyVPupEM4FJgO+XubWOMfdMd4wyNlpMBT+Yp5KeJt+GGlrEnapyuT9M8QKla+
UN8eDTLrCzCrb4TW2fCMb6BXOAkyoIx6mEqTSQAMjDn/wIxB9unqovuuyhHGGNTKQZI4dM2FGkBM
wgY5zRDTkRqHEBOeQuVVuetUvBGSKuTtLdTTKHzXJ1anu0zaVJhE9PBbzXHGMTb6hZNCPaadApbY
eyzKGXH8vXjMiShoKdtnHAcqFLEYQKRZmTtqWfdatPgOLxFmgyRIJ8KfxYXpnwrRE1LIOwxakzXP
ItK1FQZI5BmAtRmMJFOVjUGHJ/PJzhnFCN681aQQILLmkRsXo1BYUbOBHi/9sp+Wr6Y663W2oris
6hd5KTjG/cDf1izpfY/NydNdTyJZYhO1tOELqbBivFZZfc8VEcaOTNHw+kYwwqTl+ceoIZ9EToxZ
PL1FqKgqAMW4i2cjbX4uC0NaHfwxpDYUp9dEyR90jArPUkZY4EZyQq/zFj04pzjhUYmiyfzFeUWy
3eMHZpkAgSnhrM0O7vAS2Hgji/1ZIvVppKSwPCRqFw63uf6t2WbTNIyVQh42UC7ATHjOMLGIvp/1
OQNWFf2a21qcTkIciOG474FFGR5CTvNNtfaQ4X55HOhR1pEZO3Xj1NfNsOdish1Jvz37xyk0SDgR
uSRg1a7pH6F+X/qWlavlIPsX4TIvr3Z6LishlEFr+P1ID2GIzCWUaZWYN1T28AngOS3jilHvpMCS
YSqZtLkOCYjlsofXPlmpcag5nW5XHxHnTNBneWe4WJLVADM0cjh22QuiMZxknS5w6zbY0XtCZ73B
9KLabKtWurqGKhng/h8O+WSk96mZX0P99unopGXXYC01YOjO435HTNzemFWvETHyue/4b8ikJFN6
UWmfYR5actQmeKNbjtdblN76HuLZdLk3wmATuCz8xGqCgXgVmwvHskaFJzIW18L0Ji6f4qAQbYMd
uDLaHiVCuk0npAC3dzAfw+NOvDArDVBvrGmXWpgNFuKjXo0Xiodb7PnGeHzl9UeQg7e09iHrLa58
l42+f81wJUyrvVL/zgrIHl6Djpq0VuGQZTxaqVJRXoSxhaMMFv/DTk0oi61hbiOvS/T0QdZFsVK7
B7v5g1fnhmKG1hbx82ARxy/kyJWV/uYI/PSqf+c0KjdDUByeDRE4oU8sh/OL3m12VJALKq3zu/2d
OzhsyrcppeCy+m8IvApST+YKFDAJyys6HpA9ZYyec44NrtDUkdyIpVJ/AX2ufx2rDTonjgzvJrJe
ZBxt+y0ZTl3gD1xuWhCyxHqA4YmkJa5f1RartcIip5DNYZYpGP05q8JCK3TGcbtZj0J19ggstRJs
cjId6dOBlvOsbEMDmsqI9uU7yRsSCkF6SypMtdxUqHK/NPw6+ltbPZ7HoLXxDV09YMJWUJP40fjf
idKKZwjd9r9FIYQ4hW9cBZyN95YgnEVWGYbJ3Q9xx3HLPWGG1/jQYjKW0OMHnj19EJzD0SzrWZ4Y
5dP858di7MC3R4AKCxqouNr/p2/k3Kyy2dQwGvEo1XHQV37GqHDZD2n/RS5p/S1i7ymQ6ZKBc7gh
82UlZ2jdH7UhGhto7rICFDQ7PbcrJujmCNJnwtcpsqvxrKX6uqriRSJ3He6scevVxPWeRkYCNtt5
/RqqPf2tKDL3lZLPgje7l2zoiKayp57bPi3deZHUleAQTn7DhhlI92TXm05RQQr6c5zT2otMsK0R
v5COt2Mte5FrBOoOggqqWyVi2MOo8zx3V5WVYkmVMWJAQ+zZaYZzURED6lp2Fji9IEkwMW9eGaoE
E4ncJLPGnqnXH1zhSoTJiXdYT5NBdN9UY1EENozix1EJI4L4Fz6/lZ5JT1B23VsZTZ8yv8TV8Aq3
Web3hgN5UbB35rXtSlX95YJQ+tEeoXQDyW4j19z6SHkpnCe5I7aX1pPrCPBQHSTrhUI7b1+RO+1X
tcMsiDxCgRCTXNDIofYm6NQF4abpJSH3VinjS9j75j175Q07xPieWbZvOFm6Y35cgV7ajRuqzODD
Zerd0YSDikXz12HjPJJkAUnoXSgWV6bH6QuxY5R/Mb1udBQtgApdVq/GwMZpDskrwRdYqOKHKWja
87LcE1jN9eonuTf/5ULuvs8Of5y50iuZPdFnBL8CgSNCJorvlk+OcHkDnrHMB9QPE1n2KQhmdE1T
nVkpyyMj642+BL3Xh42e2/TsVtrx/fdMoJwDIega+9SW3gGQpHNorBuXnMV6mVt6ofgZfLRgHzbr
9abvwImRRvkqq4WGlUaV+0fsxo6EY0Y8hAUhS4zdmUPPbXWozo3rhHFe/lAiK5Hl3NPocEbwOAzF
AGkNVmq8CybK0b5I7yYN9hBdzcnF1SYq9o3IF1dDXf2mzRFUfEuK13z7h3/d30+2ibe1roGhjnIf
Y1P7N0G1bynpW3491Sr/dYiI/rXuxqZI2QYio6XWaZGlDECqwQIl3z9KcDh3bDoXdKwsTf0yghp7
j1OCxUpfyihSq/QBnVyd8OQ/XGOK2cMKxEuLhZqp++JF/ptV6/6PIX259QQ+C9l84VO0CMVIw1AZ
F5AC0b4YAYbyoQTXxU/xYIwb9PLHBw7WT+6QobCbGZmnZ5wFmlQtwKtx+n98bvO597nFrOi+EYAX
ttZgAgiz+aeEcPkKqwCMnlSMyjodvu6ZtxUBf9TJ1vD57QmbrBrTTt9bjpOfn+Mpm6he2WKvWZES
oVcWgpUG7O8sFlpBmM5RQNL048sCwFQFg1xRYnl8wO3mso3P5662O7D+NVulBhpCh0IWe3rcobM3
MIwSxToNEVKDq1gDOULB2+wNUaDz0If6aeM7bgF4eXtsL3heemXUOXfYmtVL4bQKhOlHn4IEXLLZ
P6fkl3+fmHDYa1DX1n2UQAAjCvIiFrqkbovCa6J9tT3RhJyxk1Q42cDAecsn2u0M51hQcjYysehV
QnQP2U9Ti0NihNxf+Vzgu01nIRZfgajiVQwBa/QCb7poDX2WvRBRbZz4jCF9Z/pRfmiRjEQP4sOx
frH0ktK9dTzQoWdJ4VB6hM+/kVjmqfCxt1hTn0UfOHnSVENLu4ZAt5jhQjNBIL0oDLQvJr26cg3D
MeRv0WcyvBH0kdJwg7JBZiou96VVnlavpiIOnDDQY5KRjTZ/al70AdAFkEhsOPZgR+3SVXYQ0wzw
/vZ75aqnWu02QrjbV1TkcEztN4HTLIPWCuJuGiP/yiFtKFoJBC0BMyEP2Y6hOL1iCNo7v/0QNBXO
OJyUQADkEW+7pjSMN6eWPKxhw7mGMaW7WKHQIs8WM5hWkv2zgCOS/4doC+CzasnllQUMjm1ixQSP
+WEGm4bhUc/hA7ohv9MRxVB8jTXQ8NfY5t/XGsbbBeeJcXpsrUB/Sar/1AYGp3EOkuDoP8a8MnXB
Jr4zA//KVTqC3TneNhX9h+kT6+QYfdd18k8OZE+qnr4hj7pcpeEOwBEOlJdLtOGuPZGwEZl2Dd+v
/riT7n5Pu+ZHw9ZwdbXGZKrOOJZbYxaowKE40BuNEWOZoJpzPWb+NxYFEMrFNotVRQFoUEsNbX9E
WaLJzlrnge9I7yXAhVA6mA69fAY99yJ9QWwc6qfUpLQrS+u55tROdEDfDZViKw1Gr3jvMGnijiGg
uLs43HFSfcApn576HvfZ8NGLQamlbil8YnV/j5YmNmqPqGBzEayqzkOKMz4/f8u10QzLAHJlf8++
H/srSgQ48zLMeO4YgdppRdkFtExdqF4zlKfjiXkst2vJvQJ5kCQ29NETz6O7QBXzgG1le5uwP5oJ
jLZOYk2ckgod7WqagIxPLIQoHyTLbtGzo3eArbm/4sYMe9oagiJHoOncNoH2sk/WVbkX7kXN2BNk
ie3KSr1TtWeZpQKbWBeJTQgv4bGCxzbAWT0GB97yw/qjRBUDlr3iqv1+13+bHEYIzb+1s7+D4CV+
CJ26ZM6OoWWkjmWr2AzrfNu1eSSdAS2tZ80jYwJDDxZWAFJRIk07VdyBc6yMz32U6Z6fL4TM0qtB
s3zLpwf9aDIx6vloGsWk5vv4upIIrjyH+vyaq51Lf1/KpWBAMjX50HPWmWTbWoNRjrLtmeQ05+AM
djxtirt4cUzc98wmP9vhiP81g972lr5EIC5B9jiYKipQkcGhWP+x8V4pDoH5CLj+l4/4ZK04+y06
8DMjfbD8xzFlwIh+WdjffBdYGiFhKD146/ApPGL9cPFDZQMoffhw3SGyZvuJ6LRFQzYRhPLymf0T
anw/GGsxjOShcebqKiAb9Fi7KTmnXo57nOG+5NEvH9GCZ9FPoo3p/ybnDGXdsF3/SWi/9IGriWX8
4c2bNXFZSDyfO2DUwtLNCFWNO5mQ3TZs2DlBrmImkh2u0fAonSYG2LkaGs6vCSadteLxiTk7TlYR
8UuiyxnmKj2omjk6N1KfWN9Xbv8Dr8AjvOnPTo+xS5NHBamvvfgovpPy/lU2pienDTYrcCFAPl8T
snssNaJN/ENxvvZKd2vnCr3gb+6sxtcg8mNBZGhhXp12R90gt+za70GjeJFwOJsxZCdzEz5n4uf4
8+rnIdhPYIyqKHYPQXorwNlKBeiMd1NkDzBFMNS8NopRU8r6LCPmIDOidUV40wefd/TmoBWeyIDi
o0GREkcQwSzF3sBKBRgGNs4OS42uxPIvdEke2X1s0cPr2CKujGGK8UCx/XNcFidRMPucY1S4tJZh
dm1ZMMTc/laRxZg0+fovXr+geNE/yHDgdcejoWro4QIk0UjUO2oGg+2gEqkDzMsIvrxxvyD8QvZX
nCW6LH+wgPxxVS5PTKsTEcMErv5oGs5lVqLJlXE2V14InVP/vN5P60P3V+FBS2Q+fBN3Yn3t/ISE
2MLpvyiHxeM9TnFdkAQvz+ukRlisTrZN7HkzcN5YKowNjFu2h1zB6lJGLQ9mr4Q4U8S3bgCaOooD
vuPY1Q4IQMP/zZ+BT3BMD0Dw9rNaeKT8qP7oV9AYfzGTR+XEmsXUdsQhLg90hyirGdKSy8bOiPFD
5sf53StrQPOKyKS+kOZyKC3+nYJe6J/jbo75kbnkeWIS6hXYLFnl/C6/3MpvXno2zYYkcXa6sWoq
Z2G2wfUi+uTJaSdWKJHVguLbwUmGrKMEplHp/3RWTmfrQ51HG8WzO38pVTJGmsiZWtxc00jMP1oa
Grazx0FfV2ZCUIbi5hoYgWNkUf7iZrFkvaNcqOahBK8H0XkvORr4bDd/G8dz3ElQhE7yoqqsDLZ7
Bt1pY7q6AhQfQJTohHLXsr8E98zypiza7hsD/W6kHqA4tsV3HryZRQCstiMpGXdx8BSOfZKzYlQx
Ktp0lVdofRyvYZCxChOtI2AnQu91ZAnlFpfT0rF8ncndAlqdXnGl2jCDRJ6Vvf8rp5BhyiV2ZdpL
39oVbgPhTWHiuKaRn2yqJcyIhyNpcFuPRxcqa6WJcXVQYr5qOoZqeF+YGb6Sx5we207/6RP2JJxx
fcphS3gx3mYiUbzPj5BaDZJhW9FFM25HKIMVjrYVBwoMgMenAMiY83ngwBKYO/JAL+M7fDzUBJl8
2pGD+h1uIGRPhMm6daiJB7Gnj8ARsNle4xcLPlwFttewBuHX54dN7EDELSaEFufWBvo2x5N+0auq
7JMhsWjosRLtf7mqDTWE3gD89eAlN4KZE+2vhWWqlnd5mSKIF33RszJd/MwNoc5OwuZpj060AbNN
+gt4eeYMFTPjUnFQgqXq+z3o1jr2xM0r0jJN3Geuam08JPSZzNtgWMgp3rz/TXpkUxR7UylpcQ7E
y1FY5beY6gABA3p7TY+L0724aJuCpA4Z6fRK1PuFu6iI2rxPweQLegkj+1rrbaeLbSN1WRWgWNPc
/eNKDH+Oki46dTSBd5b7ismkJE818WwfOHsEYPykTwKzlQPcWc1gi3QJwQzIQyTzDmWfH2J8hjpL
cQVwE/JRrl0nDb+Obzb80KRjH4tgaAWVUTGKN/ho20p4uqLrJQa/Ojq6ycbTuOo9tUomfSvLIi7n
T9eg1w8Tlxpue9TI/AXxzIAmiRoynMsTnPAPr53YetHJXPlKTNz3yzH384MkCpJJQoptzcenAv3C
My8BkhGmupWCQ5PNgzJ5EpiEeHsexDPwnJUYtUQI39VxqFQjE7ZFKuNIhsNGi4SylarFIwf2FPPS
9iJS2seX1yD5fnbt5al1k64NrQ5Drbgm7MstlLoUxtrbZaJ4QNUGvL6zG4wKCqTE1pbAP4caszzx
vi8vfT9af+saJtDBkpkSKBzbWKqbe8qZEbT8CpDzQ0hOn5HimfsiJhCN2krqPlHhjuC0I3QPpAws
bYYuvUk0NOCi/fYJlg35570fZVsElwpFkVTc6M6x0dhLJO6FAO8tfVy3r42CxhzmZfnB7U2ReKnN
X5Me9jlP9ZP93Qe3jNsgOUtkS54optms+cA1kdLSnlLuW/Wh8TAuDDtGkmlzMws0fB3QZIk7/8zu
VMrfDjvae5UMOg14ZMnSKhjgl0RAIliDii2HVxOiRKf2psksSu6GR6diMRMsmApU6KYc1lNrNxhK
j/PlS8633dtaBSi7lYt2kT+GMMIMgRiU/dLeGQ7Jwu5LUH6758beaXI4EIKqi4OdiUWNBsVWJj3m
cK0zFQNWm63/aH2ATYiTfUx3K9gwjjEsnZNhe0d5X6S45skGvhPtrV0RDazqcrHtRYFpTC4h7par
WIxbIiqk2a1+b+pZzqe+mPfnbAiG0TxA4ohWXyX7bzLwcyHHX+paDa9yUqPB6p0KyN4Q2zvZRgOl
tQiIB6GM3GC0wqQiIqY+Ixi6XU9CJI4E6bo2hoiIGjGkJnLiY5DBznCqQiRzjGb5Az2IirkKMrWn
hwj0V3SoVEcHSRXgQOcepV5+kezx/Zlxz8lIPYvsJwTZLTbIIak1MjEJiFQtqUPi2j19Zv8dTSAv
ldz363yeCYD3pHQp0mnLBdvc5cHwnP7Zch2m4BC4EaJOQwt6k7SZHrGGKnNboo1d2rRzKEZm3Csj
8MC1qYB0YeDhtFRLwfT+Y6zHGsbxYHF75gjKGcgwSECeSpPwKmP+nkZyP92ltZefIm1WUqfVWX1b
ek3ewwDI3j161WmgYB28ytZx8rm/TTCErg7gKrLnve/0QlTGztPsHz7ZbQnqmqSYJ434aYpewz/5
PO5WA6DbDBT6/FPBgqduLFIe6HjPXRta+JA65ZbaI/ny3xdlBm4mHG6wB6l2PmxgJGPovw5S8p4I
ZlyvcjkTqTNeE0mXyluun/DvvJ0Xk6iZ1VA9njcNBUmfn7a/axuSK7j5nxaCiqBAsjEEz44+gQH2
8MQKtzM1IbboWJhwcW6fTnoajuEDiq2mzAn93NRUIDpt6gnT2t0qcxAFikdbHbD6S/kC7mLX3tuM
YigfIS3aACDb6RaTN1IQ1Si6HMxkJelT4wqaaYr8m2B47oBOY85aZ8pSqUNZ/wgXOR28Wq+YmtKh
4KSMRXeyRdZH/Gg79jpnog0dijuRdethLv7BtZLPfTHUZ207kAO2xmlRmIXSXzVJQ6yIWTv6uNns
s7QawcQgZXIvMDzjIEHo4vE7+9ZpT2veMJDD6ubPxMZlEt+RovYFfpQUkOQa9IbBC3Lg9OZIXDjr
/24qxDssZ/ByqZsWIrxNSsMvx0NJ68nLB100qSOEkGUSzuusiKIXyQSEswla7njmQGPbL1ksx1rB
DyxovGq2x2eGMH6PoEdVMhUnHCCDOKG8TiMdXUrStF4UasLVc0IdDiMeoLeHKeJYVW9TZy6yDsa0
d5NrraVORXk6sP995DMfB8JizmydncA5eyWHUqJvcpK+F8/1biSfEU8LvhgP5TE7Bt+iu8HrvaGj
sIEPDAmeImkIOx4sXFKrHFY4n7CNZiCBeZq3S/avxAj4Q6UZF+1RUvlKQnBGYqvoNW9mUwa3KyFu
M1PzaRqps5ShKQp7KnBsTTaNxv9Jtoip7c032x9y2UMcRjEQFK35cNgvjn2AkhzGSBgkXCPswoC5
gUqLY7/ANqxAbnTrFLJZAytv4IJlbXOzrZeoqDx5Sn/m4yT7LR1kkt3Kevr94VcAG/DBVvElTDI/
worqKQADs8oSd2AjJyhJJGNsFCXMvqMkDrRTKcKAlvv9Vk/vgSBr09/tZMimZr5aqP+wdDRBclBu
scNJ7X1DmOWXEyPJyg4Q6w7PFV763ClnDU2iH/x7/lrOsB/k6IHEVrMhZFwrdsHufVDW4mg/XgJt
lNih8u10HZGcX19rQlbO8Zw9t9SuwRg5xAmGaGOjm8AEe9K9heE2Wt0HnK3ecZC5sif/75hKifgl
kierb6BZFvWy0UOZ+beW/qEHADjFwC7YTJy5mQ17HEJRo9ToKRm2BCwTJKPL4dPkfmVM2ODJoO8v
kvg/+3ENBvp4tlOTUYbex49/cHZz6z/0ZsX10ngNh4cc4JmcIvyFxSuA0oGzZArPw+e6etZtbAos
4k9+2FhpLT+LQaE1xvMvfvXLwIKP7DA7g//huJP8v3OlgslFts6+aw7fDsgO1z3VGsHUR4pl+Jys
Es5zjofI0b8g9mKNIB+i4E//ToQ2JBr8allaTirs8jjGuGh8/l7flcCv9ftliZBBilTd5aXoyoIp
hum3zb8gFtES2H9Q23GhgU7pNz47brY0O4wIgHaoyJvECCAY75pp8uKnH2OHP/9TjxNHzUvUDhML
TVPk6R7TPBv0cIhFlg2z/JbhqQ2OFBDZ+xivic+xwRH9NPJRUSS0WauTNVzz2Uti3bqsLCKie5xK
k8Hj0VltLUKYT0T3Tv8XY1d9LwZKuQadoxBFrYFVdsPza6rC5Tpbx9k9+BLHXq1tlSp9EvtgfF0l
fNduQvqKvESAhmB66g8pYKtVB6XNZaA5xfB3YzlITng4Ssl/om++4pPjMvwcbOxU1H2+yLLHPkms
9PA3YnajJLIfW6DSzlHO1F418KTh+mrgl5zUU5/86uwkpjSxQFrXuavlJWUjN6mANu+U0VwgW4U+
n8HGUrWWZameLGNogjBRAys8jF4mGuu1MuSgJf+SV1NTphyum2KnqsQ7E/pLHkMiuP+ZkNGffU2d
EENLGojRYqge7ikg+uNkNDBoBiVLBxGKzLrqiaFjm8px+tW/7l5Y46eZXtl2dUgBItOxAiujH23l
T2uF47JsjVv/eBuQhGwubfOD443Zlr6JYdDjOME7vyRWqaKL4npaOxIakkR7YZEKz7w1r/R2MsA9
DG3J3lizpmF1n/u645loTFSKYSOVs+hglfuOd9i5qjvQ2rmih+QCQkZK+U4NlfPnnl9q9aTltfU0
gYWRl/xmwcPZTNtbWNSXdG4I3HNkp1xES29fcdJEnjcLBDU/aogdB7xYxD3kzqjZPQkqyRhvUjwz
sJxXj815BabKQKDtp5VG1s58whrwFIFBnn5hnKRPky6Hc1ziDNPCjgz2I2LxO313ihFpzbpyNIQj
wO7xzaoIXbwbUJd/jr0mJsKowkpd4c+ooZPQdPBWCcB/I/jNLsBEjOQmoLCzodhMfOSvClnfdIDd
bECzNwrL0Mk8ZUD1aMaI5uK08fw3fA5gkY5YKOdoXVKZDqubNNEeCMVrSnExAx8vAp84VJ+L1MR+
JrT82dRTaF/J1yDXcpL4CRyH5hjuVmo/8Bnx8nsEzxI/CRVjL0dg/Y7DSZ1ejL7i0oSnkQbmVi5T
3P5DxnRQUM6lxKpI7gfPVYjFQ1decPa3KrssffWDExFubWhS9oMWOYoelYnb8KzmKx6sYqO47Dd4
Awna3sxX1vp7CL3ekt7p2GU99c3x+/3YW+SgMhtx+9x3eJSvCFM/DVS7AUrXBgeUUhoAW8QePYB4
AYT9dNqCHHA5m9dCz9fNlP5aYj/jaw9U9atc/tKmVFErgcye9bLeu8qAd2RRL3UcgdMKETHqHvDc
CL7aGDhqwGH1UmAPCOPG8/Eb925FKyl12yq7mRfJTJW3jtdFHWsa9rRnxuGI0P4YlgYYQmXlwnJV
qU8TnQvpWeIXMC/ZAhWxXPK1POihb2D7ThESP25b0KGhCiIWEWE7NoJQXQIH+8a4An83ojdosSyF
TU1mAntRQIyNIOBZa3IOZtI+A6+R6YyM8s5DY36tgG1/fPdijeovR93v1+TKQ+N/W161WujBbhau
bZCTXU36aBwPQXkWOiXExpKtxQIE5vBQ09xdTWgg2jyuOYjHbJIPkosgW2QZ8W5Qa3r8XOUgMcCG
inpXAwqOvg5djtjC+Ux0y5eeP275JnKHRFjtDM9/Z2jAyROisbG65sH+wBerwwhdNQt0MIFDFauJ
gHPTyYvlF1HfshZ2j9A+AMx3mgP35ATeYRwL9bmQkBM3qR11xufCTzvMGiiq1z1I/K4NS5uUWn1p
z6YRzdBbRJWaI32nORYVKozD8VZ5DceG9w6mfKYvJdzWSIShI9tMGt+Vj70fsuWNAySyAqDLz1Qm
kKS6vEZi3tw0PYqNCk+iFdjdWdkc79TEvRfhWC1BenBeDpo+5L0FShSE6vIpVlGdGqg+BBuZYavJ
6R11GFB9UnztIFGa1jn8pEKBicF4UlAOtJ2v1qx4hwjJZSaaxVVtzgadKFXMvWGbc87rGRBX44xs
+9pK2B5WXlY7uddVK23nsjKruhjduVTvXivfuVrL5dwNkTwOxlOWJp0+YqK/rUM6B4tk9NM64yE+
JBEh02M20YwundGFsZhISdjYP+K8Mj0VUox9ckbIXwFqcq1y1I6zIGZ6eD7XfHqAVzQ0uY7lyP9O
p0At3jB1qXGcRsuykrGFyDO+huP1UlZMX8RfyIOBMN+7nMYnkEh9DiB/odUTU+CjHTaPUhaXEFut
nnLTzZFq7Ofs+TZLHh5hEB2TdQZ2FvtIxUkdfTjBgxg63PWMej3aPaNLysEJBsXfIqreOPJ2KuD8
53PGb524UGHN+kYxmyv8nf0KXynlJDnnIAWKKOi4UzfnkcOoPBk1TWtfXyZxJHnoJYg3Q5PmKe7d
/OMcolb78sf7TqpyR22UscFccnBRqYd0GUiKu5b2Z8IDZCjvuISt2Kmh6brHPpo88KJfrCqF9chB
5lWpQ5ApKOf0ruSffPc1Zd2TCvWsymlpVV4mDFM7N47KC8i5VmIc9kl5FzsvqpAUWALMXzpib07g
AV+Yf3wQ0EQvaUi+bcCC0iSoNVj8KVawDj8m4bY/qW34kec32s0Tv9m4fUmEmH+KvISdtVYvJWny
FfaYD+KOoBi3JIsTNPkg6wBQEr7H/dzbEp8Qc+seqoGieOioCLpUxPSRyVUmiOHQQ+j3yp9EoKYr
A3iqmYBTf7BmZGkzjKUCgb/fseQDG8Oh+Hj/Fs9udPkXbZ1dtkJ4hfyxOZWXSUT5suJhMeFeznWg
ztjthWtBUHgMpwg4FHV7vBMHcGt36IN/rKAZ6iPqSkVudr+j1fQG7aMaeOrB5WexT4K+xde08DCL
wtKX0Dr8ZZmShlAuwPShMz4LM6IC+u8klxE+2tF9plnWove7vyzmc9ABFJFgGt5DIXeO65djLHZU
Y3vJH8fpviy/BmY/pHKDFu3U0jC7yIaNyYYZFvsbTAt4UhRG/sC1NwutwtsMkwvQJuD+0RYhAZ12
sw5k0oa9sFSmHD2bE+mJJzC4LtjoCymFjfkETJo5tjH8mI9ZET8VFz+C8MwQaggpLTN1MFhEERIA
zDdWRYucpJqQbd8BwCC56M1faaJZU2S5axmhM3V7OAHtOZaf3JnzoysZyVM/LQYXGBTfHSNIZHNr
a/fgWB8x+wI16/yYepIHfBk8SC8sKhQUNX9yIqBhgblQsTcg0hhbQeQzp8EILjW069Vhhh89fsPn
N4HEpVvz0osUmSHzzkmgU8z2oD9NvWPbvxrIKSxrM0WhAn7ehKLKWKjUhRzO5xfd46Huu4Ugq4y6
nq6j4KmBCG9YjCE2lxLREx2sIwxby9O+yBtPMZ3dRYQfPfrE7X5gmNURUiMeikkKRrpyUkx2Gwf+
oq2r4rPMvSKT/K1LcRH0U2Fgl6rheMg+fpfsLsjmWPU/To/MFlUZKd9ixkZi0p2wyabw2mJPAhhI
nuoNA6Li5LMmgAvZ0TqBaYx7KzylIJS+flpOH5pag27I3x55T4yEZe/DJaoE+mZPlE3+AZqAWsaB
tOWYNYH/Fg/gbeXTukJPga+CYARVjZcjjGNBwL5Z1Y/wmF5kDJXnG+NLv0dX0WM49P8keE9c/rAE
XJ5I9BOAhXMqUfa1LhiGdk9+vePehE41EBrKrymHOQiGTlYeNuh/iAh8N2u425JbhzArXulqRrJD
xgvcapKjZ0E68WvjcHDh5cjp/o3P3hPaEe+x3/beN+hmSFNyd4tDd2kNuxAg52hLoK2+QWuGO99N
nAFFlK8sG6BUkO/bQKelH8Cdh3qBYNdRPoAiocrB5iP5jTQJpqe5P3MfH2tXyiHRzQ/BeV6UMQe+
p5BcP7Jw4ceCkoNG4ONNxJgA0TqKwVm4cyBOnJCtl3EiWozluK4H264i4x75sysMe26dl7cVlO0j
xamPvB1WXujQbW56qiOdkuKOHW/h4wpvvJnyrPxZZcjvYtkK1L5tdloSBECwsz68E1dueN1Zx1mm
oHOOglvLI8VMcZmDihLE5pPu5pmE5J28TjDnM4iMIC1on9484uScl8vZihc2WWKUWYTPWKKmthYI
iQ0ibNhdkc2RJ1N8TXvGHroDqH3nP28+I5Sq1BNe8wwTpYlduVRx+IsRYV2iMr9bRzom5f4kX7Dz
WhnkXLvASo9e5WdVU6I8j4CSVISvN1A/J356HM7OynEY/wf6g58Ajfpm7w+awYjhrc9IlhDELFBA
TEBoNWXJAEQB4xIow8FB8NaS+1GLZ+ytZnXRN/SbbUoYB8h0xj1d9UuTN6AC4EF1OmhdZiCVUpSV
Iv990Fy5DhA9UPQp1i4FevQafcZ8VZ7JdLhUDRc/LODHuTxcj/ZUcAjU11O9fogbZgKH9Eat/9vQ
ESxQpdpb9hRQLEGx+u692WygPMuuTnYqjvv0W1/wCv8iD1XOALitC/jCb+0LkBiYZBHoJuyoESwL
LIbhU7eh1zqHCWwo2phdRAFkx1USNQIoW4CsIRDvJohuD6qVZXxJ/ly9g1WhNUN53X51IujWDEjD
wqvdwd4ZGTRet4gf29tOuOrlI+wQ9djgp3wsd/gS4MlQEBG7jQajhQbLgg5c8hMV3HoSz0VCRs+R
SxamFrNjaT+PNPknTvDtdo/vni67+tbQayBp95dNNVNWnBmeMAbZ6d2/m3ySg9XpeR/GrjdKc+nb
lGVKjyycNdtH/TDqogkP6CpiVyLLJMNu0EYQY5kJU5zA/6gPE0gQf66zBHhJzhv64fKLhrhg1bjx
BX02zcVuVv5rMyrQuE4Ji5V4/9Nk5RlwH7iM5unafVO8myvO7ON5qBfTX3D1QgyozKoj5TV44SwP
fuOqsw9z5qHlbeKNMtjk94SP7dKXPtkqgEwbUuc5wySGBYHOKSz5rDrARrGtNzMBeRr0k9wxHKsX
Ctjv28aIFDyF0stXGjqT/Xh0MeboHIjj0wwqobRtq7TUbX/yIsyF/IoSTG8W9woTNkoMJ6f2Qt7l
eZYnlQDDe7IcYNaTeg/Yb6Wg/eORj1NzTYhegCKJbQDRIH6bQdF/wM7z7mX1pF3H5hzV1wkUGnFB
bA1rIgb06AQES8M1aK+yRJfuL60VFThVQVr02fcn8cNZJeE2x+YEZyG/rMk/MvbHFGXexROxsRMl
tA1NOeQ7iAKp0Ip5JLP4H7WQxZk8/K+MaE6uKiCIpE5jfbwUAqtX/v6o0pGvSpUgbmC0XVnew4H8
7kKTQNnpUutn936K00qtLDpefRpKoXTCdFz0TpGYEdWCJaX2Aw8PQ9h5b82jPvWdFvvx/RVYXaNj
2OhjiocjEL8K+zJXEB7YozOE3mvzYlTAvhg7VlmERov7ncjwEDXKB6Om5FzoAESkwC7DJkuKpBP5
KcZVIPEHrtoCx8t0xXH2cGQQPhIoQZlYMpII1L4fZNZZ9T1tM14+BaVsBJqvBu7rBK81DDk5GTaJ
UqZUH6nG8/i+9gra0SXQhsa4PBLfnstn1tuqqgyrvpb0zsjm4Vpt4uG8ejwEUO6pR2cMbK0Hur6g
3sg2OafIkk/B7pVT/Z5IHEbxrCESaGViOJ0T7/HHQpi54kTIlxdD+J1te+Ix+5f1HQXMoy0CKQZW
ouYi7Pt/AefKvWAkSzQu6ihHRJPzLgmHBJFooqPljTWNfxjtVbQibZw1cNodkciBo116F8jx91zh
8hoOPrkiGdDXRvR17eb53x9TV0A2TSAsLZcAWBsOG9cP0Lc2mqgINfD1rBK84fI0bMPBPz93GSGY
7sVkl1ODkX7ZDTuj79wkBzRNMB31Gt/PmlOkPkRJ90tb1+XCzn4aJNIMSR209tFHb6SSwUFfjsfo
yyS1oi5EBEZAkZe2Pm7bZjpP7fCY+1QEREPpe+7oD8aswfs/S1lXFUm3FM//qU8RmecbB3OI8Hrz
4bAglKDuo3rfqS71dNhKCcADNnzJ9L6L0IqO7McFGy/5/cin0kYkF9q5TZTGYuby8D7QE/ky5GzE
pp/SW22vJkuXs5Wy6Vndaf4E9HtQgfsugHoo7ACJcFYVyA7zIuZt+UdVnvm1LH0O0CGHMkdrRAnM
lYX4ZRjELAPL4fd/2Z9nW1Eai4ogIaIanFd5gU9P2pHX+gMJw7jIr1XlotDKerfBI+9p9Upy+S+V
p9jWcm2JRcSs2QbJ3E92lGfBKlMT2Ihg+mRX1e6Au+PCCW6EPqww1sBSlvPBLPC5kT/utMBlKcPo
y5frKzHMOrJ+f3RpUmZQ9bm8NxSdxONqGgSJAo4pCLAMJGTwM3xxWgUfD5QHKNvVTj6RiugWcYiE
skopmh3aSC0++1q2DuXz4a7L7hiN3RMzll1skVm4ttaQ+GVm4snAmmMFqhYwC1OIks+4zgg4B7ob
Z6FLnf7AkX3E1Ficp9RU19g5qRPsUYZUCY20NAsHcpQwHfp/501DBVIHyltg52fFQBer7heY1qT/
QXxYn01KVXcE6KgUNRATT/gKQ8uHC/l8w2VS+ZLGKE6Sc7q5YAXOrUe1Uw3PoBqqCmZD2i+S5xyx
etkUX9eJMUZeSzyICGqojH/yGuM2Ap1+8U5SL7+8lTr0Q1spSriIbEyQTd3J8YQeB7QsUeZBBpls
5F+Mwyo0S6EqwrLDpjzRqduyAcO+WzaDuKCuYNMsvtGg/26sbwQNtqR0JsFelm3zdgsm4ptzAwTL
ujOCvVQpOjOFUFDHrO5isp5uv5ls/5nUpvIcHUK/DQHjnEDjV2uQthDF7PeXt9fRQsmbD/G14fCc
TUWaMON4mk9E4KDJ1VlAHtWuN7WUvocVnX1AIS+owMd7XmwLQh1SLVz44wc7ZFZwiyPA1gCXunQe
81FiFkgnYmRvzGuKNS0tEgQ2KkxHOZo1IHvCVNJE/cTPtYHwCOq8fG8/hu0PXruOvURXZ723KOrm
WaEl+TEibul19GVdlMLpywrwKFT2KJ0zEHinc5JRI6OV6Y3J0l5cDdohWyggcOZvRR0te7Ee0M/e
rQAaweNB5JIuoat2f0FZmIB1fPWs+N5uKNkzI7mUNL50jtk0ePBp1oCtQN6ocKSJ1nfvKOH9iqUh
wgWrNzdM2oHu090D5MUpWRuEY5SH56QAVSEsuewH0W1sn1lqmg9YOmiExdcGgFkhwdiauS48btT5
abZlQCvnt7RVs2b44+vYEFSHqF/gXupVWf+K/Zp7tZXPouLJ5HOPY+t1kF1tvTmbswADIPN4qbm7
JlGzkLBa8QCNgZSd/IPFHECZF7AHsrA0UUvB8e4SeN5j2YtU5L2f5wuZLbMPQmJqYiqmiVkXrzmr
nxmmPBr4U2D17CqEeSHCEFw7kHmxW0xCK1G+jl4hgmHf6wFC0HhYaIqG4NQeRgJ5JcQgNBAffwQd
zaWZoCwAbDHpptEObD0DPL5V30/birDD+3u0UTxU0mtma8K4sa4xImuSjs7LOrTLSGTRDzn8SkJa
qMpw4jvPHLMS7Lb8AsaNj0RmtDGYtB7zu6GhF4MREIUO3Cx28enkMOSNrE5dAR3s95z09T2ucBLV
GeA6VWVjvoGeP1Rfc/f2jv0Nr4EfEaxxSrA2yHH4CNN9D0JNsE1Amuel7q31pliPluuX296fSVYl
RzefhDdBaa6UeAUaOZn7PCTSLIU6OHsXnsh/X1GQSBB6SvzjcgQkrvxwPXGqOZ82Z3DIQtaGZTkO
su5TimUaeqxPD+sxpo7/HnD2NetpNrfgNrPtGs/fwZYy4paiaufSXPI4lbJCXHvjt6LaPmGKLE3I
SF+Oac7OtExJyBtj0cOLyX7aI/rrhbmZPhRwPM6FiIPXZQ5hZZu+eaDP1Tx8x5Jgxsiv/Y/YypJz
wWMN4oniSov06eDckx701vUXNx5inhZX/sMLTJfGdtni2nm4R6+KAcWb25WcYurRYPy3jSzhO9IZ
qqWrr+kQoOC8xcb7T8rKDUAmibnZRVDc6kX70JnHJRVdrObj6DM5OxBIL2AMA5kU01CNdOEDXNoI
VgPJKk0CApT1Pqct6N56QyUCBj4k6mRaPYvBdeXQRsBF0cD3n7Qi9SWtZ2TM09239KUALzEtiVNy
Sh+8i2dyk806fc2ONMl4lmiTXImZTNR5V1y2E3DzsHWiEmsASqy9+lZgRE9bG4fXUd+1RZb7XexN
bfhLfuhqSRh3PMBBFdHXS0fIU/lVdDBXAR+pk8ICRnUkc1MzHI0sBUHfkMQydeC9PDRy+wM/hRpt
4QLlxa6U9vhZC+YCd4CBQFrTtxrrtxTKhy1vWFEJczdlfOp+N9PzJmrij8OZH4l2ExWsix7c+Ysz
jiXalLFSk5BD5WwOV/ySJecMMKqRl1AGzDqkNnAGtx8N/MsqRk5RG8P3Yr4kVSyCqVgMRQmaMUbm
+dB3BKKGJYCt6Q+aWxlZZUKysB9r9h4nqy7Mukji6K4RtL4uK4HTvB1DKsRDk6MQrCJ0DSf1wnWm
GmlYkfhDVn1Vh0jwlyiYKuN25JgN7UnSPAnzgXWw2atZb/Zo1NoRkvP69iA82EQiEFJx6bWCehog
LZV2UoU8RdpT9/DymbRPChDr0slbTrXfY8K3K/4Aok9qPTwQJ7Otan2AV230aY7FKdUmMpNuY2Oj
iB6AOV1mGqi809XMKXImJnufzbqzs1eBCQr2RKoOw4jCCzBSa0+OjMmT4ugtLtAQJoUOIrbh3s93
aPFmI6cwivSlnEA/By8GgwrFaafjFmHsLJZa+7e6chvP1m86dguhEuDNJq53+LRHyXUyWMM7mPU9
jZ0dq8TUxuZnwcuLC8y46F2B1+4bRV+b7DdlnQP5OTe/OAVvAu0+8NoLzyuLe4fCAAw8bktBOMb/
5QJRAvfS4facoXR7/IKoEx7MyxGjsEy5HJFufD9BUz1QNPsXZLZdzZqHA+h8crzgSioXeOmpLzkR
hlvDzlN9Esr6WOXINWM07ddEsAcNRc64S+YnAeH2mDHEFX8a1rtnAWb9xbLEqeN3p1nDirfWSFnq
lUW8Xnp+C7Gqodjwp07RgP7dd55ZGM0ULYmogeb4zRqqP5uLBWbWIqaKeoxxV1g+CM+l10v+73e5
6u+42GRFpwcD4aipxyT0y0jxAxCLWSW5oWj3ol+8dWuyHruTF1O2XiOuu/LXmBLfaXEVFKUzcsUP
GFskvBC96F5Tty/FP5hrn4G4rYoZLmydar8T/TFkKKWthWzCQ5Yu2iLndoopchNp9QLFznqtnCSw
Fw+YDksvX5CGEwmhyQiaTAO7rEHYiCBxTb+5tqHI5YSOsAh2RAwE7k2FrSpHBmtrvr/4/06feQUJ
zb3szGV3Ye6vQKeqeTGwaz0weRavXuoKx5M3zq+BOxAWYx8GpnvQEdd2yBVmdWgCVdZS9aJIJfPw
BTFRXwn4TkUkoXqNE4YVQ51oxkF5pNvxcYLz2PINqPxo/uScec2Xvs5PEnLj11chx8YgDAbBc3wU
lb0XSWSTsnLAPDTL1yWib4BTKw3DCjJBMmMspxOyVJZ8SOw/GdLWPPRR2ODLAzlz2nu+Rg2BTvK2
o/k3RgvkKP1vqrRSYNyNVk4LNwzOn5uhb/QDpJB1ewyqJLTnHikHjAjaVsjHywpdyUTsG9JrKgBW
+49+fp/AWr+qMmEVFKIVw3kv4lEFJvv91+CdNzPXl2DFJYtIhv3RDxTWFrKTUttfxCtWqJ1VQ2FW
JU/sgEelA/wwymF+K3Qzk5a6YEgs+uctIBkFv5tt6CsQeAPIN3Tqj9YHvo27G55C1z+4Ix978Lba
u3ip5+e+CwnHwe8S66qeyFV5vJB5xpPLIqNLvxaxAyMWFzr78UvrQLs1sNypHVwfbbH5eESfdaTQ
g5pN7JGIjB8658NRmVXKinYkJ557hd0zgfQLAmPnVx3+H4+fUNuzS/XUXDi/2iXWnlSFF7mqh0T4
thEy5c4CO0Z7uJWOXPjs7JEZuKYtcetXB3U/42hjgLs73z1Q+SskvPv82Is/0HL3fRaGeMLse4/V
peY7p9YEbDx1qRvU3b8Z/appqMMZX22fV2RD98ogE2JlkekKdtOzqkzXTeEHR2xiDUtD5L5kEtPh
lbHXAn4XUJT0f08G/bYperml2PDHCUMspXibrudGYBIP9bL6VRyd2OWvo6/Hh7yjFWck1HI24Bzz
gSlI0TEEjqfn09GoWTU3Ox8HuN9CDhsgu/4KOIjoUySdnFVIYsbXeVm8Hc1qwoq+z151j5PKLO4T
X8HValqPE3NZq4yP5/CSjzWS9+9rO+3zB4kp2uPmlwNGzvTqwjQfvK+d1hbKHlqdDbl4vUKfxXBr
9IgkQGydXn7pGClTnpC56HjOeNEBmYCB6Vl4v8M5rogTc8Q249HSeIHzz0v84WKZ22JsGiAyjsqn
WHjEwgF8sNuFkke3hgBXs/hfBEjChN+1kB2kOD3wCeJ5m25vvwjRIFQO0Q1uLIrpQUf3rcb3SQ0q
Q+NjQssKffyh3dBiKw9z4AzerxPkQfAU/AuAd/mfCIyeykixPllyvyogAvxN59A5KSChdNi0CXna
A7KUpZvUrSxanGd9+1qpjFSZmwX68iICk0umQ95kttMOYhriyamAscmBMd5+VjvdpNuEHWCsTnob
p9UdRbngZMPTXBiKzVZg718JvALy6i/qmUykXJoVeoLFaGMyEQKJbYL782rP6IXOPKGpKW+eJvyi
cXySzWfXWtcLax9h7Pirom1ZEyy8t7dEjVn/PNmtMmyZ2gjT+TZm3hp78bRpZaQ6KOztsrm5fEjq
P+IIOiFFzd24bd9HE+XL2bhkynvuCNI0nnmfxvsXiFbR42XyaE0x/WTycfL/1ASNuESU4/R5dDME
Fh1NNEAWMvcEIBIQzZXfGII3A0C6unJy0tzgXwLIhV5bOzgoROQpyC5lP0Wbq4KqGmHXrxePWvMz
TgwpT7gF6j5d7PJe+y0e/GK9/AhzB1dvUqB2YgltF+F9C+gk/CjM48HJCyTxfaIaHBeKW9zomDMV
wuR88AqINIju2srKjYCYLo4f6Mz/WclRM2bcyIsRvdWUOEdy5a7RBfbduA42cgHaEA9Rjrg1ZpRq
E8ZJvHNpeHqbI6O8inIvb9F0vo81+jfqTT93LkRx+ttuyBEmJ1U4qCdpOz5SeYwtgXq3TLQpk/ZD
tPU/rccefCVnblZfeaB/rGaqDW/SNLpA4bTf1OQIAAqQLBBttYcpHC15YDnAu1EtlckyBMAeAbgN
dLGh8Vcj2wg6tVRZgcmUs0YkDjt0kYBrAMU/m62O053CF9RuIxaQvrNRaI2rB/Gzw+bl9OLChCWb
AVvCJSqdmO1KmBG24no4qFTYQd6cURAf6lqRZV759ex6V7OrEgiTlOK70jdrMhEaPu+BPGUhisBB
vKUS3y0rhSnK1EmLzUtMIX2dxb+c4gWOpPUJN9OFqv7ps7YBhs1VTJvVpuNLD2VyYo2fWGrBug+r
tDgLruX9d5CbfbLFo+r2VqHq9V4Vl9GuB8e3IWKr6GshA50VQVJ0VkWA6xMJvmtSOLQ1yWTy7Z3K
TGtJ+2ORT7omyn4Gjc9+hTdCDu07O5Dd3gG7+azl9rPXGXoW28Bv6kuiDg3NMcHkEIU7lhnsdMqN
UfGR2nNXwG2ux7qXSa0LVqLYAgg/yC3t1sAL9f+r4prb8EGIQVbMwZOcstqq0nS3VA59r+nQ/HVN
EvY5yS84qGIheeh0xA5NeoL2aMnmRohrBXuOFGom05hMAdSBUIg70vUjzBrYQINb7vayxU/V02ij
QI9/y0XS0LTYSF7zAP3wXz7UKUlhL5qTa4IRfNN/8gMfOROc9ESwXFl/z1TN7/dz0lJKRFYFlCY6
MYCoBd5L/y2KFf/zuLGthIJrhBgNiklYRbgG6u0p670Q1RZ+iETONyXAY/Ar2DPsBoo60tA93BFQ
UEs9s+q597jxoPso4pH5KydYUr0nN6J0ZBl+w6W9dDSR4XeODhZZG1dMTgSirWR1JTjcGF76eP16
hViQwmXNtYN3LRo/yNvw2o/pj8y3VXbrbWgx3o72Isy1RB62mnKdqaqyoVEuWozGXrE8pkwrOJZU
Qjkwv75/dMjjrok+xEcgFJpckTHRUdc4HItHb5CLQuJC+SVSgVwaET3lg1105KkSoHhI2Bs3GuWr
djdLtC5dxtRaB1UdwC4rdn464XxS/nHhpi/vNVAUaCRtxPvc0qYOMtK/ZxKqSEcws7HgrIA+rBa9
8nVKdoE5lqbvixx1XfcBR7gKO3LO1sGCsilPRye+kgO4NgX8Q9/zt7lxu4Xrs7038v+//visJekn
9AkipB5pw3bX8/3PN85LAcStE56pAnGkez4D47ny3Tld2jiCZ4mdYWN7eC94Z3u67XBNiUOfN17J
pAvzw55Lkqz8bXdj8s8EOT0jFmPMNMVcJzsDwIibNdtZMklFfRY86kxqNoCWduQJoSh7hAoayffI
gQCrHUkViSGFUd3GvKEUh83VaEiga8EU6K1wdxq0f9QuLNbj0ri2Yfj4UfTqYjZ8OuhBjKTyvsub
zuC0wOVh4iFXeWoIZC13GNeCLlxq0T6MrzfffcUlWBaZBUkK655Et4o3WzKdAgnfeItekyta0lOF
0ybSLdjyew0Fx7+H0Ya+dRm1NSWgiZrkBtME0KB4u+Wr50VYCEj0OAJ4NXLNmUBNQyeLzAH/71oD
UpItnrE3o3wJWbXrlV6DiQUxoYcyRCAZv1ohcusvS2Ged5NdQPFzj88xPl+Haayy7CysiF3ixQXd
uCVu8RyLqLL6OcyuJunb6Dq72ufUTiRMeCRfb0mpdZYa/NLKaavB62CTOFaWqceFq9ceKIb1oVg9
VZ6K3nOR8tzG+o0e8u5Mzduj8TU1DPzyOluvf4VDSyX/KS7b/vio437hcL4Lrg2q4WvoIPsfNiI+
93KYvG9CJ2RJLdQ8xJphwEu0sSsxVIJaeftDJVqzKceLEfDTs4Mmh80D6dhpzsvI6j6TzEiYBW6P
Sa1ncbVKIUo/xzEH+1v6fmDmEV79KOTUQwAcruDt4kfcEE5lZ36eXPbVQ27tJ/AvhGAbqiUs6IsR
y000cGZdYqRBgybqZjEzH5QNudIgj+aaWaSrcKCtpSetEfFMX9XFEAyh8rhOV95HSQ3eicFSU0n7
R/ATe8WxcK9o8HQu5TqziNthRm/2gf7gjBDiyBkUoG1NzQyaL5jnPoQOIo70I8cP0HngpseK0h0u
dptTxFtKpUtoqMYKtil+beuNL89eGEzbFNP8ck+GgmNUc3vCaHzG6sFYB1l0YqFW88n0wOwPqta1
TU9mRN1KEoI2xA1YISsKIRbtSuY2ctAc0+xdjlHP2WEp22IXwSXdRBM1oy1pHMrGr7ur7wRwq4PY
nhD4edjJOdvl1+BwPUPaiyY8cez+94QOTBcdRz016nThg9xwzphtyl1bsUzeGGTKL62Y8zCWNAyK
HuMOzWKkYE7BFhOWjXmfbAq32ri+m5braa1uZTOY9OBQjKT3IRRmAMZKvpuwNjrfRbirIU1S1xps
z6txXslXQGqR/HfMWgwVmL0cQ0vcKItoibCBx2MXKLaSFYAObq70HfXuZXFpJ2RQcJSXx+CLNKtc
JKbNAX6XTdr7vMLpbQXxnme5ijx16I4lu6bIE5cAIbw9RUNxS7qCzaSqXaf2SM1a+WAA+EmKDYML
pb/e+j6Qi16dXq5tHUwwOAbXwjccXtW7M7tXyQ4/q/NniW25NyurynJ9aSid0EWKU8yDoVMdJ4tu
m3wB5exkk0RYSLQPwaZirjBpbayT/pWS47vITRjLi8tCNs9qXy92jbKZ3EyIJVRSqizhqRomR2K7
V5RxmCYXCvMLsuya480kT0Eqb+7Y1KT8utVWC1wT1NCWPAobpyu3vxf7HhVwoNAVeKb8yq04EiUl
f5jWHIrsg9jbHZJkonOvdrMJd/ukMRZkucSPuURdISN2DqQebxSOVi6O8HPU6umPvksa/XEOWYXq
EcxnEQmPW746nT2kLQMGE0uLwrRv6ZUzQcR/RG7KItywCOdxjCUQ7dwjlWDAKp3VOqn+L87+v93A
R4yAiqH23Mq0k7t4oHtqkYZjeUrrt4Z+yq61bEnyzuqIO+WiMPfLRVUbdXstwy6TXVMpd/EkO3Ke
PLAhuHSr6sL4qpnt1JYFDynGxgvsYy41of7xVZpO4qzS5fYAiJRofQ2FGoX+L5e26HgXf9kmwFfx
LLAypKU+9sZb3QhvH2hQnTa4f5Mmwi/f1STuutrj20BmkHXL/Os+BA9q4xpyvH6h4T6EuWw1rNto
itpXJxvx3o1Fa7yDECEY5wV8trn1CPz5pOShI3zbZtvNTQ40MJQFwTqeZSWtSaMErGdQrSXwZJJR
XlQO3vrB6SunSAwfsKvni8I/W/9VZvr4DoTtQB+p2rSN03intmNf2+IKYhO6vQlRThFEFgquZtDk
IJ+To179hgIPuwBSDWCmGE7N+3FATdoJxniU57B2GnDQrYeVFxJAfSpYZDG607tosL343OCW1GEC
kyUqv6Nqh/6PRwEbSXObOzwahu9PJDErAfBcqFyjeSwaZL0RtrelpR/hWVLkZ5nBVWR5xTsQ32Zg
O/gBLdBQemKwZe27n0wViSSkq3coJh9yx5aDFhUUnWv48jbaa2ZfOuiZRRssRi9KHw0fAaHbbUPe
jz4L1poC4wxGX0xLz5rkbJDyAYZ7MFnW7pOmaeEbPpgqNkpbUud8C3QXvJOuIGmTPKbLxKpz+PI+
G8fw+7Gocdn1JJagnIN/zQS3JeaTptnqpf2Kbgs4YptlinUpleQd9uSvxXn36R6z28VCmbdV+Pj/
Y3YUI27JvbBsHYXXBlWW4RbpTgfhEU6B2JI1ep6bT6VVwMmnUr4ppCq1gED2zx6pE4AjOSYtvlR6
X8V6z9hDcAed4+FJxLlk9QZJWz5JCKkemuRYqAuEElncFvZJ9a5TJEl7YWI5KMao9wTLLkPURoXE
fgUieCk6yeU3lysiM7/giCk0sR8Uuz9lMKhv/UL7ZBzuwB5Jn0YeyIhi0QlGebTyfApdGfkthR1e
dU+knX81JayNhvzw9KZAN12xildKg6rkUXMO+LworELo54lX/uOfh8dev57m7Di7BjdSJ8gTrAWg
RxEWyXaiDzxxMOZ/GI19j5OqU+zVVCJn1dgCTU76e51Ko/Mv5eadY3miRXy9KSRlNVsRW1dhms/L
g1574ZxPL6b4NAtbW98Y5Q6FAg+abdK/+EhyzRvDJ6Bk1nbKa5XR4xvAyW0+Ytigfavam6AyKB6H
Sj8dC5EV4bxnExAVI1bIuMSmHMcIShUguB1YUsfqZ3MdV8AigJweopBlwJxi6S0NWU17UGyY+okx
f1Lh71oyn2j91/A6Oe/bWUy03vYIoipKVlzMUmnaUe+QUwARW9QDO6nyss4ts4+2iFCuzBJMd+KX
cQlkpC2d0UE0WAqPa1KbD+prsegLvt1p1Gf7SGc/3iqxJtcijCxjr2I3Hz1SxqcgZfLidCMshw9C
nJWOmjMG+XtDS2RG2QJF1ES+dWinXSmGXaVAceH2Y0cXY1exCb9a0iCqjDPZfpqBB1qd13ojzWxD
AeSC3phUsZkp5AXFG/03rcuoSHkOP4QlXwp7zB5/JVDOf+Z6TSGfXOrOY3/O7Niw0pnQjDDu0bEU
v34ABG8eFK3p1Fqmk95d4dp0JDIdTzZRl0oD2jD09hok2X+zqQCFvvkGC5XN/uceX8Y8PZsEGKgW
4cpaupsnZ7HLwZ781zKPoT52XPZwMBx7VNM2EyJ/kMNGVwGxHEi8QJfrZXvuPSHAbSmuuG5mhI5c
fioPtEjO1V1zRaoaZ0h4FfIJMeVSID1I/mOs/xVL3rJHv5aBQu0JlC7GLf9K+nnm5sCSzzPxTaoB
ffb60rQSELS/jxJCr8Hf6ZneNhPQrYAMbx1UfctV/HaFZC6QAjYYJr8j/lD5tIQZvG/DYfJOFgB3
g2yqApYDVKd1Au+SdbGOmaua9RanPsa1S7LhstfAYyrDwaEoe3Z7afwTyYWiF0vAcZjfLmL+F2R/
ySmTdbmT2nzCQCzDvAaxStS89ALaRriGA2KnD6JxSG7dXcHsmUeSZW0d8Bd35gOafwZUpUPQm4dN
ci5Xe9d9fNIu7LmS80U9ASgMiV0lpyOSWdXq2YmRIcRZX17F58Xh5+cCmjnL2NfG3LELL2uTm0Zu
1JZracTd0Z2b449Yo5ci3b0DGvnPLl3SqL9Jh9MKLEnDe9boAx0x9+r1ls65CtEvDkF2fxRHqI0J
+uJD/VQJ/lZUeLwY4qbJ/4hV64mSUq8pmUqJc7+rXl4+z9/jcU8NUbERMcmen2wygVF4iIu7ay8f
RB82PNInSwDT2hhS0r+vfu/56rPhRMY6iewbfIhm+ba3N0O6TU8MYDr/7j030tKELoWyhsRVuDFY
2nprzv08aLEM3PCbpSt3OzXJGQBar/jZa04Uf3xVPzEmEXMkeYfiKSR8H2GvKZIAF/wyCoVTC1kJ
JaePJgp3vxAbaaghec85M7/tS58PcKxdpplDIrXV0DzY7CmN61qAP420bfep1EC4VLEg/nE9N2/Q
dgUqz1TSbA8DNyaedr4b6EPdghtoMFZxUbYxUc4Cm191E6bRcoI+xmXyKzUzyYGBHChbc0hw1GPC
pDTkbLHlknoZycqFsRE82m/Ruicr/A4RC/meJJCSH5Rf0BQ+x/cMqEVp+KQs0BUYT6SDTmC7SQoB
kgl3I9kCP8XjUVhKXaOVKgJy+pvlrQaXJwTKQVdi7L7mVCAKaG5gIovpNhFqdPTxGXeJzvqUlCx9
sl3ladrCfR4OzLhbewUW3Mp5cPyVeD5D5+jlLmgaMSfiVJy+33bUWl6Mdcu7QirB++AKWIfHG31x
hNGneaRRbY0ZkSGdgFPSARznQs4bOqr23juqjUiOp5TDInvE9bLpOEQKA7lvPf5h686PgFWRt8fP
Vpj4muqhqQUgZ4+p30ld31N7ELJbS77m6JNT2gjRDoPlgV0VZRecW719AK/fB8E5jAKoEy+0rhFl
Tl3Ccbs6iNo8CGuzfaFu7L+wr6+MQ3YohfxCnqVDfPTzCFbyFSn3mgiqsBOBHR4bZkrj3O2d5NSw
au8We9bRL/Ygd21d03cSdjkVyowL3l0va+4W4s+tGyilhTPg7TpJ7Iu312tJt9281pGzHbSFjpKC
+ZB0GvoEbJWsUSh6mPuzRg+GniBSCt39R0QetnwBoTq7BTqPedA1Mn5oDZk3cXcxAHFPQ5F/k4w1
yApaveF4Rfl3TUoamwiIieb8DcnIIGluqF0tbVBg99fCi3JJ0vipxcODoyLBXHFhiX5KFJkakjPW
dNk7BOFpmFAH4A1Xr+0reBf+Kbp+Rcx97rEgoHhP7TT0wuo5UNConjL0iPFIbCtb9OXYE6XkjUwf
5gUjC94M2Hwg5+FpuMeoBKtI9j4hwuuCh35lvHxWsYgHAj0CBBpwfWd8XrhzmbEQ5MIQcSzovg4v
zu4iZu7LLQCf0wkvmrYrv5WV63kQ2Fwv00bv5J5nY0GwBSyKHPjrbU7wi673wrtJXX7XqGKCO104
nyNt3MqON2qTIq0ddPbIBPlH7zNZRf1l77ExaRHz8gK4uPh0iCzHRp65SYAOxCzQUWX0E0Gi47TK
6Ar6GahYyCuqsEhXg3JNdB75En03t1+zaI68gj5arue7ZqL9ZYuTIakXSZvnrpZSAtJnwQdpICfE
9xF0joFPCc8B4CQBju23BdPQGV19VMen26ZDnAMnZAFXYnI48bst0f3i6/Hwc3twzlG18w+P+IgR
y2cegzM09zd2uqWf+nfmXvSXQu5+k0g74Qh0amtCdnkOlr1RPRe078k5nBfsUfBlT6OYZe2fi0go
PkIExlHUz4u5GEWfs5rY1BsMKJ0RUhsp27nllZCVOpsl1jBJ2EeHpAEVZJoYLCSzco1B2MH7umER
UecpjaGqMY9IR1JMyN831haUDSPtOyMS8xKk9MlYRKDxMlGM/3KGn0l9glat3s2k7j/uhrXSusDn
wdNKxozgTQHeCaJw3kLzwDTM1aKWH+1fP6/21FqoYvLJJGONHjPcKJRGtnfwYRxDK+dtzVHlNr63
VZhY5XIDQeLEv/Yz5wRh1g60CGDEYHZtYJ9xVObcR3o7/+7LBY2slKHqz/HfJ0m0XSdKz/TSE4dE
1rJn2YYX22pOxNmvgpb4P9QDyMooqlBm7ul+W1uhxCJavj7Il+GuQoLKOyCPLYbLTyPVId2Bo4tT
CjWgEGaXVJXRmmMxPjoJGFToKzvIiioM1uvWNbGZmrqAEeSW44ADxyGV2IkWNNsEMqgOQsMsvG6G
LH+qRGZZOA4Mp3UIolueSmNV/1DYksfi87ki5A6Xbw4G9Uu+PMMztho5mmPFsp+fWVirY7UOpWJr
A8ZXnO0F+oYEtf6q/FZpWJOG+Uk0hgU+tvJA4JKSJf2CXdVeAipomKfJGiQG/gzaOLWsGPm9k7+Z
vB6vRqMwCmLPKoq2dNbxB5m/6VIsLeKAH+PXzN0EIVrrULCxiNWlmYNhbmJ2sLRNoZ5yPnLRFyK1
/Ij2a69YqlRhZEiv7Ph/jiXbFlJS1EVym/M9d2c6raOVs7AkIM4XMFC37uvQIcdGHYjnn34PO5Sy
YRxKWWFiIkW1smnN5g/DIVD89yDngUINClqv9KxA8+TuD6zZGCCb+nzWbzOei4TgCSP/jhqYLiOM
Oow2aQZh9aaWPcajgzcsaHvsjcZNzdwQVGkqvzoEnAbN7YKdEN3fvUfVpmNq5IRKZeKeXg5gCzbg
EDri6/v4SOs1W02X+UsMReUwulg72ArKEWgt/OX3Luc0bDunco5caIlK+ZnVtHZ1y5iMqjjvNT9Q
cClE0PPaIEk3/ZZ79YKBYkfEuY3Ilc9BGKCysM5u5dUoSfVLEgeSspWwuolUyvJNS4VTYESlA+4D
d4NfuO15LCx+Ai2WfHAJ48GCQ+BuWHuf0RR652smjGgX9a2rF/LqygiOO/8VL8vV4LlV0BBNP3vv
JJkkELaDnRC6Sm3nIPprGqa/9CYfJfWofV+e6HXbOzp2/ltgWd94Fz8aA9tZSdYGeIrJ0fnmkvnq
pp9VyBcrLn2agNxusoQG0RhGBDT0J1/BO62s7HAUMJE5eEP5h8qjYI5LMQ0PoBdYZqXS19CEY5MI
UR53FMcjLVIirhbWGm2B8yldztgny9CZMQarXBcqQ5DVqJo2dTHm9uqdpS/hNGfgK7b3lqc05lqv
KgQtswVgNxllKKDl84iUxDzIVuMDFBVfU7Wm1k6Lv9/lqCMk7p7OE+HUCGUaupAyRK5UPPWpM73Y
AOvz2TzuqsbfLTIeFOLQQCg2fAeloy/m/CTNf5Fny3cRCPleW8i8ArrhdM3hdox306jlcnCUclrV
QG/V9PPeWTIn//yO1sErJznsICVWZQBzhoieXoW8HVrYdmH7pQrnDt9Jdk0fzqkwCYnla3WvneRD
/PKuzshXEYJqKrZSbMpGVOsM4c0gVbCrQ9GKcAYROrP4r+hJSO6sUxDoDIfxbTbogg/5nb4x4cGn
g2y58hN8LCVdAWi4L2ExxcLsJRxCAIe8GcuCkYIbJLIfYI3XbHRkn86zo6gO4Qo3z+rE9hwSgN9Y
R8Wp//+9AoiFYQZcHOpwefjEjnGn/822l4py+txxel2Z1YQlMpaXfWHL3as5a3YQiqBBljCT5CnF
ztY2UL+zwjPOAh0R5AoW9Qtbhz0zrWSwqjJHSC2TONMWE9bt4PGwxk7Ba945gPksQODa+5Qai0Fv
OA0xJVEKLbxxYKmu2S0Aoc2xctjBAjc9JPEFVbG2Zn/FubK3Hr2IY5FjCHrVwbu2nciRpiALGNVy
q3DhrINW24lokvUt01nE5v0t9x4frxatI5NHBiTnud4yQBqqTCngK0HQsocgH34e2GsDC7eLBobd
2tTvmSRIWuFOpdBKnNXCnsWdsldYlZQ2HgBpJGzxvCq/33oWpbvWW1Qs1PVpKAn202Q3hXumOSUw
8++ktkOvGUFoeYu3SMxC5rSvn6rsMQZVDef6apyD6p7XRBzkb0lizqHdiziAGwT0j47CIGmvc+j2
zLRUzh2PAaBtFkeif52/qKfukIHJDNfRbEacbvlFbKwRqw69UBXOB+Yzv+xoNTMBNAj/0bZ/pNSo
7lAaPvEtxJ/WZRD8BvV3q5GbnFhWlIfyxMYxw87PR9dCXQuZOH9KzNAxP8fALQgXk6Yu31JbQbFH
fRpP/606TKAvjr7f2sxbo6LYgCmnFGt1NcAKWjxDx/v9xGBUVMzKbJYTKt8jZ47UdR9/VVIn8l5N
kRPLn2hXqMq0hDED+Tv7QooNQm/vErOJcWZIEL0QheFCFGoRbDBB5f+WR+Emv/2gPTfU+UllNc7p
JzOrp5A1C7XjJJZT98Zm1+VY2CdlODG+n4Xd/IrLY1+i2lZO/d+lzfbBYFlIEdLzf+Q1nEN+6ga3
bpu3vxzJp+0FYxJgGMVVOESTd+TE4+iUEq2xCPT1aaSeLCTt3WJc/1gBFKIy92Z3aWLgKKQEZm2t
o7VBuMXfS7uISzEw4vNqLwooXr5NIg746wQTrp3fWqGkQJjOAq6jfWmjmp+HUwSnOATyCbxuAh9K
H4CkHs5B9k5EJ5DURJLMJe16/6114G8StpGK1WgWNmVD5ciOVVX0ZTabr2+bNsWN9UdnZ2u+SfU+
kNhH921Ob3DF7I62JT3cp1ufjFJ5b+03azAfOqjLkLM6IhSniccZlPh+X+Q5DxCTHqsIg/80Gnou
y9i1j58wUVgeCO6S8QRjRWzrY3jZrh6zuHpHvQF8UKXcFmBPhMvnGvHo9rwpbkUmHqTdn639RQ2k
yJQRewJGtATYI5pQOQrK0NiDLiex4C75OJ+TBbcn6IfMmNm3dQhEcde7Vx0DglrNQX3HRjc3KuuZ
gpEOq2fEXb138WM+yzDXA3NEHsmLm0s9Xu37zQaroV1KLcMDT4Xw6IodDM8qbkbV3kKCSE/eZ7xQ
K6wBYechenSkjCHJ0g1ybzHDq/567t4uey84WQUa/YrK4Tb3QLp0hGh1rUdUKLBib8anXrsvRuPP
cVDsNKqzF/40rHCZfGqzw/Vl8ed+RHGdvErIGmhjFDp02YHJbipEHTOIyGPX1wpHh1Hzhi6Z+dm+
VQYVWVXxHGi00ynMVaUU7Wzfj/+fpXqWeSUwPtWOSgJcIAcLpwRNe5HBZNbUr/88rQKQyhfRFxIv
fKs5HR1Qe8sw4JzfIWB3FXfIQKB0Y7ddNRTs6HJHl5nLJE/xaXMadl87FGmAnqBu79fwuhWte0rL
rOW5MiN/thC2AQXpUGMwY6E/7kODEDN5VcAHCBLs5bE+/hokPkMCrkb6d022m8aGYuN5DGVoiuST
oZK5AoyCPVIuCC5FJ3MHLJdmXPQoyswOJf3GlcPBXzoPC323BECDPdXPdQ9OY7IHftN/mupHQbnj
lj/peKqZQff13s1lArvL/SrBgTef+1FsLnkNJIrByPgOkuG1iTuZkROc/CKGeLq5Fyfmg3Zoq6WZ
ccKvH3wCHJMlgiMuM7MXoNGMny37BNF3MZhRvuwm5dR8lGfe5zvA55tGdHKtVvunkSlAmI4/u26n
f1IkwYqRDr8gisBQX4r3+oJQeSPTlEHXV1qwxHEFSYpR4N2Y2GEgT+q3sDDrKJTeu1y18S3t0isj
hOZe8//uQXusptVb6wrCpINIhBXAsFpu3vmEcv39BhZkH1PniuSeJgckdwZS8cM9QENcBgsCRu0+
c1iI0yI5LT8jNDyKek7KXpCOFmG/GeZTwgylFl/DcwXGO0YT7XWEV6isebUr2l2QavFfDes3IxJd
YUl5PjlP6C2rI1qQzE75a3qbtuVAE0ZULMYn/JUxUZC5i7H9JvOT5xXB6YDRSoPNykgLI/nRR5jL
ZCphmPO1s7+zGcO7S3/3NuWbB6kAa0i7BUExne2rH3Yi8UO8uqMvYjcraQ/COfZD2pGEqUVEPH/u
+VZvL8+o7xJtLvzdSsKyB7ps0gC0yW5P0rOiYgn5ttB+t///RcTMCRLfas8Pjp/RAEL+xd3WQkSO
o907+1NuA0Z2UbBzJt4sK5dSNP10wHNt0BGoFhOIqfVqYFJeVpbGpcKbjN/+fk5o8uNX8V2mLtPT
bB6XXwAjFrTzceisR5S4GDaw1HIdWjctEhFB/zzMyNZClHKHcxEB9/lqWDVqWqODqEAPS4FuSjYM
CDwJVuIYeqmdSYIuClA6qSEeSTvosC94YyzPmwaFnk25JtlvfRetmyv3Nynt3fsJI8dV6PymVFas
8/WEFPkCHdqbYcZ5pYDf3x+A5HF4L74RBvb933ZkjnWbnkRH9pdrJUGaEa7k+R4e7q9qgDbd+Kq6
5y3Sp8l+X3grvmGUpi4FwTMhFULKMhVMPFUkZkXI+rCt0L8ZCfpbIvG6X7l1iiYOSXY3iXXGcGcn
F9QxCuzfcZtlGgbF/WVN/aMnUOLBdH/7B7OwWM0+OkrMh+jJAZu6mpkszVnhbkKeDfS/b9fj1JC0
PhT2OyX6i+sbYqsiHO5Suzqk4debBT47VG32d3JYES/4HNnULYNCmDv3iu1oGNvb3nHk3cRh7SEq
76vGDcfzM/u9vd6j5+UHyq7Iw8lKPBh2bo+7pQ1WV1l7Ct7V2PEPZHK7KP4Jc1EgrNfrPp7Tw9x3
imkCbgiAu0Lx4GBDV7Z7gBFjt1pIOOT+6FNW2+Gk4ld2xnh4hr0KGvtJL7S0RjBQXsa8SRCyRwfF
x36XSi82K83gzWaveiHhrfgs46n9Kyi/YQjZKQCCiyjyaKeS42yDNoY8C35s3v7kD8X+vaivOEJ+
9gy7FVATIcHZyrgzuFDMxMfFyCLW83F5OoKHh9tcwiTLULrKvxWPKP/s1dWNDffKwHQk91zileSu
E2ZtZSg499faJAAQH75QZ/jw/YRcptUndCYbznwVGdStT729JxPo0lSdYew6p3k48/r15oaAcoMX
mvuDVolw8lHAjXUbLzUU9Buizg9HYRUfKLrJ/TiVFdyyWw8dt34WhUxfkbG1oUWBCrC1E3jfhjt0
oqHswK9yRFRt17N3jpzvYKRtTWpatIojd27+ZREZuSSHhUz4RtUdXPOxJD+HJK3j2nYNEN1icL45
w71c7AQtdZEgRYT6MZuWji5l9r6CgjRDUkmTQp7sFGhvPUDj0d+U0Vov5XL1YZqns0erAIIiUNq/
jIonDVWBACTwKymn6cRWKDGFy9hxqU2TDtB9L/pDtZBOhjoA+x0I6DLcXHZ0Qxw35Q431m7X1b4/
VGEvLIT1swnQO+Oq+lXBQFAmO60RaPjIkMHk/kd+LhB3zfhdmQiDtE89FmgFPJ54sPhTbT7A0MUu
XSddj9HWAuO7FKvxVMb78sxrPjzdqvatBRXCAp+9mCNvW88Q6PhVDyljOBQscd4pLLi6NDMadr/j
0k2OzUTQjNtwNNfY3pTfa59GwjjyIu6YO8CE6oHYGE+rrtsQt6KtdyhOMnHlgmMld/OrHlVbD53g
uxZHU/YDvPpnk5gJDc/idd5Ftrq9IVwGACSwCVuEzQgnH+VFsk1qGDcldgm+x0fWwBsKppmbmJ9Y
lKXSQqLpb3hAUesKK+AoXKQGuvL2zwqbzfueFrZvnf5dWfA61ML2vQFLT/IzUcbUN8n5q+CrmwQr
z21Ya/SVKaJc6Pu8G8LBgOBE6meo9S/r/38G8NR8JxAdRIaj9HQC0uW1d8HTD/RUE32HCj01zO++
/ih9dzDbQog05aI2mNFQO4jnH5OXRBjYxwI/CbBvYNyf9+vVViDRFWB6GHRZR8uFacS4hw3UFTwB
qh0OwgqT555HTn+MxEHCG6dWs2H7ZOVN6VUBplpx6edXMY2Qhxs2wE/mpk+w6Mzb2q02LKSEBvnu
ShcgS50Nj4uUY43Di6aiJfKjcEhWzLR/lApVSZ4Ct+wByrvq9CD47/AkOvWW5A4b8k4DbIKdxRe+
NBFQYHr1QmId9A5OzGSKQ27ww0Li8OoZvlsacR9wL+cfd2sePP8f8/VBLhQrHhOHYa1QZHrMtp31
scFGIIFIZYDTKtdzx5p1q1vbJ781zVE4vTcXL0ggqzCGOqzSPNw0sEavlOfvGr5t5k1L6MZNAk88
awnfrjmlVJTRcYhbYOsrGlei4Ye7a7QkB0IqrbREDy/0A3IibTySlhb5WEWrv/w8IXYAoavMbtoJ
2pQG7XO/GCecwAAumw6ozXfKkpNkZ51XMHOqRTy9A6WHQZNwLQDSPiSzKhhnBo+l9ACelRl6iSEp
T94D/hsDb8zw1vsUovXP9ELrTScFtdk6Z1PRAVcaMGU5+akXXbKJlZzx2RVns8h/IKc3QfqmelJD
6kxJkLRjE6qPSC4p+Pjlg/MXZvnU9Q8xCzHfsxIGjrr+btksecIo2G58BXqjva69a5o6KdVZlx4m
ppufdVw28PqLMPQ0PVW4tDt6aEgFEOnrGqdcPoVYEWQjLhxNjOulPQRnfTRalF4NA+q0MXWEVbim
8veNCAPHo07YsXuhiPKh1vtdz9il9x3vweFYuqs75LnUL7oP6OR15yRMcz9DRYVgXEthwD+sOkuw
ItPIOqopyCNc7Lwge0QpymQAQYJ42MW08w1b4g1YHnpHhVUDgmLirPT7RhSv/RbaWp2hUDwdmens
KaaVamdTJsRpRcTUX4xB/qezaevXq6lVcMnfwJAWZbax+i01gnzQrZ6ML5HFfXujWrMRK5E1YXpG
CvQZeWUySfYG/IGlATypztMhcwX1z1MEwTWdecgWHKSR6/6gbIlHB2uD0w3V3s1ILWtgnG58/2QW
9kP79s8UdD+AjYYDh+TPhfaNhjWRRdbeESRFMOq2vWDVOLq7p3MkWIU9eGmMnl3bIlqYD7q3cqJZ
sHwyBXyVwNa/+jq9pMi6LS7iTyvwBV7K5L3h00KLew7Aye18HOVxDge+oUp4LENuk9yQWYbRlxfF
s48CydfIG2dk4sSWIC28ub1OwW2cKhE9oQKdM32rVGNGhQZ2myYLq4enWyN/3qhkmYM+xxGwGeM8
iQIbrEAYGn6fqxdXZCK/SbkZ9VR5x83qkq8pFT5wEl2dtRXLbpUjPZ1z3iioY+3qFjpwpD6MiqJt
Z/Q8l9/nO3GLVC9hhiwDfTxcXT9EQmq33qXRMyliWvjjgjXKgLVOYy99KYiHdzDp7MsPfVUzrACF
UWdohLNP8ufRQW7jDqOAiBEFcMsP1qyna/ABA628e9KqlXdt5cF5KeqprThl8nRPoQamhTfW+32+
iWjAi0ls1AT2bUVU7BPOEGJg2GQstYuCiRPdSXcrsPhyRBnjGeiz7lGA00Ez0vBs3S0DL5sHkHSL
s3qR0S+qNgRkYtQMW7HqzUSy0Gv1iONJPkEEdCM2ps9YQfNuGUrtvEW3ZfFgOp6PCW3sXwFtR/sA
s7sP24GdnZSkyUqqW6MgBlovxtGWwSXiQ24NP1YxK+9FZflrJaWL3lMvmQBD8+AYRb4WwyYFj7X+
d9TxUIuBjttf0kPhM0iEi4rzMmzr7gFhDOUOW2gxgA9f4bNKlNvqhzYR/i+VCiTMV7w5UbF812+3
uWMMayhbFHJ7GuXozZPFxRjb9yvFLquQK7MJl+eV17n9xLqGMpYvlcQ5Bj4sQnxofmXVVNDtEqLZ
BSoWqJELBfvb8m/v8RnUH+n2fodFBV09l+8kvbxiN4m+6hm8I/AbSR4N1nBlI9Fw3rPrlGpufo/b
sX8os9fNUw6JWon5P/D9Lic4GaTop6UcPy7DZTS5YjnSAvc/IcTB4I/NIsA7c/8SntLDNHQODKS0
aKotsYbseb9c68DPO49AS5+NZyYLjrlInqUSsv8e2yGbCOncVO9KkQmI5kI5mwz0UkX3mSDXFKEA
yWlVRMQ/OszH6N3RKFheNfJAojjpviYt6mcmi/m+Knj6Eeq3HHhhdpSDs0Tb4A7F+aEZ4ixVeSjK
sNLCD2dWjfTUO5KDJlNdXWgw4hAneV/idpiYktG3Z8mdiOCjgTCmKUiHVXASOYyrl0a7jHVQSubm
DqXFgbBG13lXSxb3Qo62WuD5rrc2ozdhLlgATihWWPXtZHNl/99h+vuqAKEev786ce5xLG4avlDo
M5DGzT1wUrN1mIpbNVwJ3LhyL8DTW/s1UptjNim+mmCJJp5It5Zvt1wA5fJTcaUoY8zBXL5YDBNl
1sIEMei9QZ8wYh3wGpvr+h3PCHSNFqKv/2z+xaaQEKhZne8Jkf0OClUpI3bxr5cT+0Tt7eLNo4ga
sIvE/1xIv9e9oQM5G3zpYCeew5pvIDzIJKrg8e8E3koJfyoUfLAXXOFUnK8o2owimwPDYjyzOCwg
jg/oxu2Qi/f2UEMBUn4iJKQvxSBAYGP0xfwkxp+WXm+y27hzqxkWMHbMWipR6KeDokU8WhYcJEnx
G+0XeZqu0bbKZs1JIUtz9ngyl337Ql4bMgsBdXydttb6QN2obIU+wENk+G90BzPwBA8YtYZi6/qh
11F647LOoj78TiodX6VPLY5YSiWM/zrBp4hMhNM7gG+uGfZfrxN9YBaJMdfxEKBkG8n1p5lUFcwy
w1QvOdqpmgpySFOGmYz1ollvGupZv7ZUO0Vf9jg5rRxXG3yVuYrFzP2jCdvZi/WJpKcnv+eKP/3m
9Yh77OcAT4rSjDHI5wj1FY9Xciff2JK9EymjkVKz3iNl/17r11Ho8JkDJJtrAlrdk3/LTzpa5TGJ
azBbmTQ8sS7NwAr9s8Ut0tvZBhW9xE3mBG+uf2VVMt6E+4jolJPF1z10KTS71pbgDNZ76G2sZ8vh
UYyVBRhK4L4UwFSarO8hX3XElIPXCnDAmRGlTANtsfVKiyTN+cV7jSgG9rO/LZ8V15rsk3nHcvuu
kQg0fioBhpLuu3NWqHTizADLQWiyCFVFVCuKjGEmhm4XWHj79d5F+k8DBfH01S6AMxpwuBko5I6N
JSyQxuoTmf+en/v4P/DvMmmqKMiNoV5DFhkGfkuWKGiLLAFuSlbyeqcKDFW08VNdYc5UkdSKFe70
5TDBk23Jb+YUrkCuyeshRHczFZh1dSXO063uzapPyaIOMN/8w93sJyjs0oxX3UKukbLk1LO4u2ms
r32VTVu4oFYtgLEo7tYKfMuQPEGmS4OPaLNJWSElqhlNLLE4u1MEh/lTTL6IJCRQy/n9O/B/CPTc
e7p8azML6PDK3zZXppMUTQz3nUjHRiaYvIG4j5FWOpfnGlJQGUGPW3y2WisBzTf/jDlG6WV0AfEi
gqDWiqb2g+/S4aK9znSKJJ+RLs2KzOvTG0/lNNdy2XAOaXkx+Oc4xu6qdBmcDYTE1/jTG9rO8bya
pyva2SsvPiCUHn2VQDvFvlz1DV5+kwlKKIO3UcpGR8TP83ej8kUVJrL0CzQJvDDT9jEpL71+Yjv7
YV3kE08LxfNNMJLoU66NF6n6zNn7MInVrfw6YLoM+CFEeF1d7kC6PeJ0dAUSgyW6teRbsHKTovEZ
wVpXkzE874ppIeMFgY1wO5q5intunb6A25RNbRfbbGXDKUMXiadTG10cNK1c6yu302qkLV4fkqYC
+QzWvpkHfcWbLCN71oM6VW1zVdUObx3bVEErjForKttZmhe6uX8KOXb4vwmZky2X1Tl6ntpwLoUd
7yKhNn9f6N3y0TSvytm2T/ZrU6FuiVtJTkjKxJQ32pKWe1HhLjZnrNJ4XDIF/1r1pAa8dhEO1lZo
vcTKnNHZoRnkFmk+S+J1XWrOPe87s5V0Ggd79+YhoOkSWYZtwq5EmnOdlCYpwfuNDjF8ivGpP1UM
jNUvGNnLqZ/2qzeYhC3gi5SHdurMjJdP8Dg/u6bM8diBcU6I4WJgYG9cfD3O+hY+qsEsLm2n3aqi
WPRWHp0pCbu5BW5azsJaBiQMAIPXsjcgV3xfguO7/7urZdhMUK6AzPVrtQfkWPt/xkuCjx63Ubae
9IbuIIy6IFe6Ln88/YLpLQEkNRxtbsU5vMboWMdIjLeIsVTu/4bK7HOcGaCzPKK3qd7CpVDxnQxY
iLW0q933wmpx3jeYaY0yCLmovFHyvw8H0ab7Zw1iHkC0xYi/YH818T8aieUgXo+lpD5EhX48Xzma
a2ryBf4H6cUBiRdrty9zq8AQvInRKuNMFgO54YUJ4T5iThh0XyvRt+lilIP4E0tOhZTAWeRMaS3D
erI8nXTzWC3eQOLPv+LX0KrP3v7gW5Q10BGua4ti71TqCnZeRaPGXz4OtwUAVerM89oUVxpmkMhY
0EVFc+s0JGt7Sn5gf1V4JtI4Q7c0kAmaz1nIBFU20qaLKWPZTuKYBFY5whd3Ja61ag+yMmCn5KvA
Y3Bj+CfeoUoe4iYE8Jb4XMcmwz5SDWwPbF42XzfkcVijL6jImqb9kW8ewpTbQI/D0OFlVfPnXjZy
mki3JeyZFCIjF7qrwSdqHd9+4EYY3Z7e5Stuzs9apnZy9nOQIqZQMyz0pTmhCD61Fz/kpIRKAYS4
j6Kce8CADeco5tk34flj7YpOy925RB4Tu+5JWa8nJbqtF0Q6kUPRJzGlshGQk0SGQ47Ic6EI3gOl
ySm0egsv7yY81WWNK2w1TT3ioglWitXWGNNUsg2C4Hgh5QyQmRG0CqsxSLhsDJtvODgtbz8QT3Ai
KEWHHtzHPFLrdo1RjmOJYb6D4WhvKgDZi7OvGpETTujIJxMfyrC56Q6W2LUYVX+6qI1Lhpw+iu9b
TR5adAtPJLmg/ZoFbMXqyWRynOVKr8B4UKAVwk/GDfrJoZ2eenO35aIxX1ENDkv3zr3xFVyHhj3m
hgDKuIpY+FnA0YAqiGGDGiErGmRFScIxPjMBgf3i+KowsKNA/tWwBozZfbPm2+2nNYpEFmqurXz0
e47A47I5pqzTg08jebvv4cPYNoT5U5F5ewpwhCH2DwdIA/03bDTkfu73fbggNVhTy0NgKc7Wj69A
9Nic1IjytZSaGpTUXRfmo2Z3om+Laf5e1GLDSkgX6CO0zrxIpuQhWPsG8syT9mMpXXI/dN+yle32
duwf/KQ7cIkPVe+ASQph0KDryA5XtISOrF+0YJKRg3jOGsIwrro/xlvJRMI1AbfE/ZYCdAW6uu7j
iJ11fEF8c3RaTbu3jyU+X21WxpQoqUCIbNGJKuSIbt2U6lkINxGVvUumAazN/A7KEUbSxek9xCfZ
KhK7r8ykufy8dssm6fIq9dCy6jg0VcA0ok9JNS+LRr26pZeDnxWdl/nN3osl3F3cSVH2JqAphVeD
Fho3lr+zwQ612dUdAPmn3ANYijiAzfWSDx/PaGAQJvdnVTbT1iBOPSqlCRgVmOMJdSWzhPdlbkfK
O2e59ycfn0ybZJDrr8x7MCpR8yFshHqxEsBfEZC0QonTq26xJX6p/V+HOXsBh+zTdRLqVvW3zTLh
Qv02yHsZuMupSJkxEfjvx/wup6YLFJAXMJan4BMcJHHAciFXNroKRFk08sshcayKew4PZmrQxiR1
FShydprTA8N7GPL/u8vAzYJme8w2Z0OIh8jIzDKs6eogLY1n3Jhn5Y55BK5BWR01KXyF61KgG8dI
a+K27T0iNmBZ3KqLVq+vMUfhfdXGiZ7i/vNKwm/gEnSQx6s7M8x1VJ9Co3Z1KfH6CLZPbMY7/YZq
yFdOnFoR48uPX1SaZcmki5tVWri6/iwbCYNMOCENK96JNe0wxgu2Jhn71wZ661RATti03+CUZorO
YX/lIkyXGf9QIAVTPUkDCJ125vPgFOLlIXsk/XD3UNBkCrPAZgAaAi9SrlbRSZQf/jw/r7BgYjDK
PVZRnLhfWIDnmkcUjwAuORikctgTK6EYbm5O7nBQIMlcfQDPydvGC+5cYqgqGrvS6eiwhFDUdP3a
JQnHb9bMHwa3o8n+9AnGCOQEIEzP6JbBHvwNdVEPJ5iZpaOD9EXYAQSFJWIgL+cLhkd6NFoq/aCE
3Q0eueuFeEBYz0DXNKM8/8mkBGYtPGizc+Y17OcWfpAr2kUgd6X5xI/98Mx9Rzk9D92+CkwkZLAd
+GxVQ8zm+Ls5bBYecX9dHbQzNbzBxK3fpOWLem6fuuZDQozR3z07ugjhbD5I1Al+56ixzz9zuCPx
5Sn3UDwLO2X2SSLlyvoE1wTPGWs3UqV97P4P6BALXwKJq4GZmCs77wRrPk9wOypLr4Won5QF4jU2
uTmDskeEDxQXzIrkSvZpyLRMoZ/PWPN0I71HFmyMgguV3yhfSN6Yh4Q1IYad7rIVcMSWEugJ/Cuj
BuB0tzujG+rJyyl1debdcjzwjn47G1PimbaSs5GRQFdY6YR89/8OHaQPQVxzvEuCXUN+8bvDydH1
0X4t57oPrdfDcMz/VC43bB4Z7d8hyj28bBsG6Im9sMeZFsAJ8kmjJiZQJAUcvwhLCXDgTel69Aml
Aez4Ts60f/GUW7TBtbJNm0yzg1w7L7GGE/elHuHGztTMLoCEww6i5YjIYQajRqiCyq9J4jBRfuDr
L823+JRrwZY3/bxBCzUef6/X7g6wkRfppltiU8tlMNRsgXEEaTpMzuKlOg7k2s1j7oU/+Czldsa+
ZbgSQF1ceaMh185vc37jOfJ3vUZRqkJ8EtwoQeAsmWhx/lX4Y1A9gf1SdGJzzyIlv4S8WNL2j1ZR
2t/H3s3D8Y6xI3IdWmKXEdQ9sWyvR3Eee01B2L5UMH/Li8JWG23nkJyhOnBXX6hPach6TOp9bwet
JxibSC0Q9d2BXKOBAL77212S5q/EF/jfNmYbbD1SdVtYHHYV/bTKPDd08qFh1LH5N3BYiF+ArpoU
JZtGKjgyLuQkHJQkyllxRKXcmcGHvxGRWeaZqH4oy632UXEVHJXuJ9FfFVe2lUBR/q7vLGbuleyc
h7JcP9n+GmfH8xtjjz76ryJ97DWHsvhw0f0MbIS0dKylRU3Gfa1f37ByzGkjp8w1tiKAx6EaRD+H
4H51dq1qJcPLtvVIrDYe5fdpJcpElOHoMxWL8O/qpb//66ewXwLu6zpa1T7fEvcrF6rEELzAH+E+
sFkvN8zijAsGYgeYo4F7EFpTd2x0oHOIpYnV9/T+Dm/ym4abuDpr2P9bQsc/yF3OoZgdpGdxaInH
QrCoB94CIh2toD1EE9UEXGHI/pS/Kf7EmhWGLVWZvYDPP3HpG8fFBH6/MiTkS9UBoqHcAh9W60Q+
FwogrNxR+zWOjyhUslnL/nZBJ/4dRxGIx7cY56G/qofqJmt4WLRQRcDJ3voMSWwsJcXAxu8ye3az
6b1DqbM1EtAQ9s1t3nTbanZo1v+wayyyySETa4qj0ltz5qz3MH9EXsg0L1+/nWb5sZ+l9HC3WgYt
r619vsG2JX9BsVVRAVOP3eg06ntbyA1Q2FgeKsb3Pel6wGSu3HK9b6bxm51giTxszr6QW5sDMrR0
paf3B1DVN7jhgqjjUIpg6QSHsUEf5f13Ymah+HNy4KDebLhVQ14YvnLpZX9MwtTvPeZRhssbMPh6
cEQF+SRg1rBwzNGV1SyG4pjfNTa4wd5rcF7FpvmQ03YairGdNXccSaGZRGCD4yUwWDhxLtMd2DGC
Oe0/tN587lsFWRmZOxsw7n72oHNU9Gk9TCsJIEUP4Nd5RZDT8SVriYvXrfTYm4i+kr/ZLZi0QfUn
Nn24bAMfkZ11+XTB62Qbo7hKB4bTSl4rl2uPoLWdmV2X7JCtBbdze09U0nc6A6FVn78qfCtoCCCN
Rqf77P+UcydY7cZpZCFXbu6D8/zBx3vdWtyhNeLY0wCZBM167GLZHA3dnxJ3XWbxdN+KNo8k6wCZ
765YN2HNYf2e573rwEarztk0GaOAiJqLqHFYZpZSHvmIODD9cXdkd3Iwy5lR2xTxAD9K/mGaOV4g
l9yHIigMHzqNvc3nLVdvrXXMWAcPT6kdd36b6lotC0ZfUukcqEaKpdYGmcwaqCtS99e1MAWoUHcY
Uh2nr37jE0yNHw0f+BiO7Kbe82n7D261vh92ltA1WWoBePgDRSraXOtkW2pkV9xwXKhsKBVPlXUp
zsuZ2yB2WcNTraE1tnSE7bu4AEzGO97wyAm/hPo+L6nomcGJe5bca2ZvCDXYKzqeLAE/EMpShtsu
HXyv9M4rylUmqpzyRkSFmU/QOnIKFJp+u5nTKhrcXlYh9pgMn5ob2XW3bkiUiScTudC9TPIvT4v0
4XrMc67P7Kn0hwMLljkb9KLqpe2fsPAtBfiInz+6znKoCQCcer+iFFakHrDISxbOQYcRflk3sE/r
X3zhMQocpJj5wUheIbWzRBA5AFf8yqfa4xrSNfLjy9BC0BX2vNDYJB4tbbdK1tM6EbHXWy11RV/H
UzP8F4H2qFmPU5duZV84fgRLKuUk/IJvUSxF3FjONtkLZ7NXUdLDSK8R5CG6RDPwV8fxq+0NDhvc
gkXyNVAuAWdHXyhOt+fyRz+HregQ2gfRBjnb+eYfjLot0RjyOmENFv0kX6vptCDVt5qU/QflhNv+
QC/77DGytE+ZLJ+DhmuBRi/BBZDvg36kMtdtmh0cQr0aIwren1XlstfdgAr+GtrYq4tk9RyxUJQ7
534abjmli3KCML9wzcinrYfQeMkrTGg9MWegTYgEJn0JJn5dekTtw5a9v/WyCMQNkvH2rP8ORjU5
D0knRoWageLkG/PnRtorK2Nes8ppXLE6nKuErnj2/ctaJfy4cVTqsIa1moDG3gSvbpj7Ao3poQ2Y
tsLupR0nVU4eP9+v8msjc7DTdpn4H5BiFfehENK0fyS7AHeiea8o2AmrR9QDIeiKrwiAytHPBe4k
NP9ardK/2q7RzHjldle6teHEegdOAOANwm/bdYdRhbQ8G46mwoRULucJpK9dz7snsrIRR/pRo0SV
BwcaefT9+6lecBnXuLjGTlvaeFmEpELoaIK0dmcRszJg7WT1YPAf8ukUeoIqLCoOeEk+1yZo4u9X
iDTW2zsLeHrc56P7DK9UVYWS0ZK1s4ZL7zE20YhJuIIQbNJ++tOrVLh9DP/AR/yW7MUZ8RlVcqL/
DZTlELqx/S7JHcWaj/ATHJVSmoT5N1LJMVl8N/BlU04JAQJsRNq7p+XGVSsApsL0G3v+pZ0pCoFU
FWaIZ5VatLE38dYugAvi82NR9GMgZTMYU27IZRG3LGSXhaAC2Tbs5BQo/Uc4XBOygdqGb5p0pRgB
0MmcXcFcC3M7S+irTPL/PG7o5NRoUNtWMZt/hzySfMKWn1fduMBGtV6L9XDBMvHrQLwnlowfKnRM
Id4UybhiRLpsu9HG5ZKTgU8Hn/SzGLBH8BLtfR0FoR8BjqyulsaGm2y7JhBRzLe/m4mdx+XHcxnM
sJ3OBvXiUKc3iQdt71oClawDiJPyK68EHI+0SbYES9ncPxk+bBhyyzMRMVfPPT7VjCP8eS9StqPz
9O8NwznONfaDElTyE1Yq2hHdInfSffgr+p6bK+FaEOrazupYd1UJX2iw1l5njYfSEvAn/oKuD1yb
aVVzkgTFGbzdnmhFIWgj1GGjN3In4uDnec4g97pfPvGUzGgwP3QwwTlawwcOzHaFTIcAXEcPDrtZ
K4kSB2NiHHBFQl3J81XTSVGeqRE6Leh8zFeKPqIE3lhMLVTGNIays3vV7J00R0wscKzy3oRu9EiD
vFjffwCdSa0kybl4Jcv+Y0ItxA70hTAeQUfhJpeK+0XusI83GUZn+QRF/8dWnGTsVLw2Ss1j/ANY
REddWZJAdKVLr+dV5gQ+F/26tB3/mg6VY2PJNo5mA8t4Nis4XWoNrg8LeBKO32NWOBf7PP+rCO5i
kwiXxdTmf/GsRPYIXYaZR9pWHw+n06DlLmDLeJinzVBy/74dsr2HZxQ4fjLiqP/CdVbAQQRX2vbu
F6tGgD7RHu92m66Z0ZLy4RvYaTAejyP5RhNHtEdnQWukfO5UXr+em0yqNeupxUEiCKJqFpDKtLcK
z7LZ1RQDZITlOtE8fO1PcgyZhOSY/LHZUTewGqgrpP3cMjPvIS+AhfQThx2suXS+SviT6O/OyNaG
KSuyl6aCmwO6Yd6S5RWdRJt/O9ttqJPHK62xBZBQycMiao80GbOE/mWg6O/yS5V7knwLuDmBr8zA
u3qY4O5Zzae4ltr/dlDp7ncf+vz92+rNxNvP6tWPCoIAHnBk9EHDXeJUfdAdUpRdcJLD8NPLf08R
HFh7gYn8HOLhTcvOBZAI0DNpmYNXvzikT7QOUmOmCGAj8Wq0+1gIMTMVhdzXvC+pYKgWuxba2uwE
sqgp9cy7do8pXxm6fzkKAM7C+bzuexRwcf7x9YZ1XxHEG83p1o8VJTe1pzDN4ua0irYsDogiRLuy
PyIbwhAw5VNBE+4KXW65Y1kDHA3KSU8tAdzEV5iWpqI/xFicVGHjhwZYigNyBwp/TSxNE3/KUsgV
BT8l0bIXQLm1DE9Apf8nLzQm0ZcTBB04vC4E0TYkJI6orfrZ5ux9vvPLmVcwhZMTbpQWw9wc22ew
I08Mjj15Etq9LnoITLym0DSfciFI9eYnibnW2kFu6+opx3YJuOr10/87u3ZKb4umqkzFa4xfR047
XeeojJryeEGwn0rAWfQB6Hi2s9vf1Uv2CH2kgf40I5U45741mv1gjUaK4ksJQJNoB4JOkiP18Mx0
DVdhdEJpWbJxKYJnD5/eqgJU/HEF6YzQOMpn/4B9XKneJKmtPZQPb2ambW+cTYH0kq1TnT3DoWhU
rtM/6UE6CWup4oXFcUiBW5Tyuxe9U0ZZjG35S9rX3Cm/73rd2GNuRIfVKfL8xgsqrfEQwyy0+xDO
jaUESs9LY9zG9si+V9ERwq3BFMvNNr9kftOPp6VXqm3h+8VYDXfokMKsmn6DUr84yzDHUX+eaTFw
Nrhw/eUqU6ZUbCh2Lb3BWFC+VG9jtuut6YzqsrbW2Ol68x0gfzTnEvJToLx0kOHiUy5L/mYeJ2fs
CJLf78a5+0x/OGOOMRKZORqujUyYk4MOCQ2RfWZGR9gayVbgEDhWmjOtGhCsu1txMURMDgExOwxy
nDzyY7gnLY4kwX03n8RkJH3nPFDi2KerbFCJgeQfWJwj5z0hnquqm4pRYeGlPJ8pdJWiqlrH9Ty2
YIyfO1mSmszWQ7hxmpt9uwYY9FxfOZvJiEFprnKt8xjb4Hh+jSXNq+xP8uMjSGmy1Q7+EN02OWiA
beaOsPvZN/xg5Y1oFS3dy1sP+Hr6qxChpx36a3y9/QF2YcaVXiD+Vpt8suXHsQY/zEaS92p4rPMI
N6avkKBtuRw8NwsQi1BoMdNpj3HJ6USG1+HAYsk0D0g3EdhMznmyjLAvTUI7BU5j1j1pOsxKnJrA
MVynq9OLJbtgeuc5xDBHnX43YXcxOsaNdRasgNXzS/LEB5iT0sAQPFXgkSge8YVdV+ixa/ytP8+u
wth6HogzrdcNP76ZY4zZcH4rRi6y2g2Ckma95P61glXOhH83+RQrDXuqjXkr0be2STShJ8ot8OAd
Vd7ok2cqwZEI6uh32tFXEjHotQLrShFFMJQMJi1VOfzbUaOMqgBdjWjpaAHXD6/9lrBXASSrBlw/
eWQ/246vDU0Q1sWi5FmHgmTdaRmMKxFdTXsqkLQ5Cojr8CiBdw0V6WMHsakz4KEp6rvgbvvGxFvl
LpoUKVf+dmnF2zdO6AK/nvDZWLj+AFF4xvFiOcyPdoFUR7YL9Xmz2GpOWZ39GbMOBFaEhILMEv+n
V1kkcV4lDuTpgQBQRn8d3p7Yikq3jZCc9WAnTOWpRpwUpuSsOSrrohYmQM2m9ufWPSJhj8SOUhiw
Q59iI6cKoEaWzrIGKdXencRayZsvnQL0uRJBxLKf5TlnY9GyI7jfXFXfoUr4E2tUo6kUHJ4hO6Sl
JkIL9xazEejMlNFzx9kv5r9hJ8S613E44ke4tYaMsC6tR3rIT5e4tdr99dmzGv9jRAkYFvS4Ib3o
o9oPVeMmRzBs3VWbRvfYh+ABJl8eEPm73qGuHJiIlA7lZWRdi1wuMKzBHvbK4YjqO5aaENrWqTtp
T55wIHgCxYHOljvyUBrCpMi732eRVtaIjOuQLMqQQKAa1ZeX3PGIOHmzsgJ07YtDNvi9ddi3shtj
ivaoMMcE/0o4gDfXL3yW8H9tXwNXRqoS4KWsOUgcEMitH4dzfoYgzYNMxWhZzWLD5y+L6lhvpbCt
KbrePSG2Xrd0Hyr13VW2EzsXTbJ+kl5saMGmDBbRZyAio4qWdn5BDl9BWETLng6aG40azrZBXniB
5SZYeui9IwAy+otvlFjOEX0poHB0zldTUA3X+wSLYIh3eZ2O2jQkceBca8mq09IQAYBklPmXBWRb
KahLCIY9dRt6UUEWkI9x3pK7YdqFDoWqa+P3m/Oqo5lIen+zez1HDGHUF0+aausMTInLMd27WPn3
qT9v5Q2W0DDluj4B/O9YvAe4ik+5aDQ3RC8Nt9KaT9PElGTo4vWCyodG3gohqlbX0cxJwBIuF84B
BCsCJc3X6zoqEL+FotZhK77UGXpSskR2Whd3OOKZvBF6RjnBASH8362a6m0EuF4FedJsejznPIX8
iA5Zxf2cczknq1Nsjm7AoAYLbIBDVI17qA9QGKLd5l0kAt7H/AItQr6JXTCdMDWGCkUDvJsjnVHW
tpRJsxyLpa4cdOP9pUpPgWCSz33fA+d8HCu4CxmMlsjudKOcXf3tZs4CZS9WXIXrBGIoGI3vZcMh
mm9jn/wgz763+i+f1Ax+MripBqzUFs9jveAUlNw5OLBHu3aO9IeHqiWbcpYd9RzVbey51FTTPHIu
Ln2LkFqF+uKfj01NKToGAsslf5XUTTfbfEAqA8BiZhuBgEeVzrr2glNsgWqZtZZRZLslKMuQEKjf
vcp8VQkpz8mjbDMqERAUBG+k4zfb+69LThFDxBHTA66jkf9YdR9iLtf4u0x/RHvA8HzTTt6S0pG5
x+9U+E/vgntZEbSp+YKBSxw0zvSjHbQhiE/Qly9xlXROMenAGY93BqLQ5hYngATEDnOCXN7pwKKv
eKgQ0VPvscPT6qhpDGfCJZd5ykF5kza1/BCG8tFfcB3iOmqL9lj7uFVVtv4zDeZZimNck0K1x+C6
HhpFev0I9qDjQJIwQfQQqq3t4UmoSmvS8fjhvBdDT+9E587UpYEp/V/EBdltcak7DiBAnuI3hrlb
DNkzQKPzgJaTgWpWJtWaB/eYA1iJyY7z23O3YoSM7gbXQPJgzH+WLWNJrXFADupDb/9GswtBKGQ/
wb3q9YpJRBR+sD93+6v1PVB3IweKxIdtS9lRkxnrjrW/DSlP6lv+ctvEBZeGr9Z6T9p+RUF4Hl5Z
ng7tIAG56XmiV3jkNrEBQORbaysdDu+YAt+4E2GulDXi31NzMmf/VG74LUNl3wuG+Su7kVuBUkJO
jzNq6Dr/HvUqm4QbJC6cY8Q2URui/BXOG4E4Yz+VkkI5izq3XreRExKYy97uv/4STBo+CV+I4zEW
nJuaf7ToLzhi2yo7mUpaMHzo50MMHzYNSd8fyNUq/V40DnrhpYZfq1gnS+VzLmfRIsJK2KtAeHLS
sbfF8bGP7lTO4WF4vdg7vTLPnyHJA1XrJ4thug06rTxLxAIPKZ9nMoJzRd6dP3llHAY0MBIYmBrN
zvup/rSZ+I06/vRwNDqdc1Xnnb7F99BSG3B7vtDEV2h9JXwyWOlpUYN5FsEsnhheOv9FaWsybmQ1
aAKGTVh8lb50r/RJ3hbqypqWDYyymZODD750d2mBARDNZ0W4YPlFzmx+OSwukS0fYR2HqadJl4m1
d2438ZsEOF/LcKYmIBKR7ZQqfFgXLMcv+WA8JbWdeK+xGGfmqaVAqwBKXJodvtnCaekpRoXB6dA2
XpPvdqx8o4isjmIbhd8nNC9aACiXLXOlFqs7+zmwhDysKQTg77+JAc07LWOg0zfjbz4+7M1WyFTd
U6mAX4fumC4/C6MqGO744reBMHE/erMDULbmHnJv6U5jo/JBu1wARL5e0tg2mQOtaTnpwMCecN1F
BZbeMfXpHNgH9eJPLK7cpruaY2ZvRPTTh1WPXdZjCtVJcUvHPWec7fy1q/zuyy9u3WsRByBZAiSr
M2vsIDNaysrFEmNhSOWt67LxuXCUll5/pNX3RmqxCLrSBG1Jyk0YmqBWavAFAPL7VrDi+5uKA2sc
VB9xYKOuIADjJf7WvmM0Mg2sz326FEUKB29sXBBhm9tpvQmXoG12EkY4yiVdPms87yaZCWoVICq9
xSadHsfvK+74BB8MMh3MGgp9Av3OvqtEF9QRQGUrFoYy9m/txdckPcAhb5r92igmF9QbP47g8RlQ
W5NfEZa8rtFlYuRpZ+ChCK+Vw+zv1RdU5ixdVOb0tlMAU0tut60j+7NBjXjTLSbWKbzVv2Q5/5/w
ArGpttHDRfrm0buFQe1AxDPJVyUelyD84ISRm6/FDhgvMETCC4hNKAg0SGvdlJhxiHA8rupydM3G
sMpEZRrHi3GTR1SOvjMAPk1Yv9aHv/PwSvyEGNcHTYN/f3T8CU+LfnGz937OVJfs8DGH3ECmnrDs
cye9jvMjQ0EOSy8D8/z97Oox/4pAmuV3hVt5xtQJDXCr8wshfDaVy0C7iCiQcCr9CPP0Xxx525yS
4FtyJ3rusrXUxHGThgEcydyeo3nhXVM2CQ1lpmGXTNXhHMMBgTZd3JWdlZtJi3DYPIYAiyiN0pM8
MTjcdQX+BNNoDo2nt/ONqExPsbInpC0/QWGXBnF40qcTKoLE3h7fpnaXP2JqVVEL/Gxlev+tO4GB
fWV76hY/iOatr2ZGGLzrpvtlhawbNpRLe/NcbmbCsVebhOonASOJiznddSnZz/rn6RUus9GWeIGM
kOetS3wVuhw/j10X7C7s/vyv/eYD39Z1nm9FRlZWRaHtUjaLahyKO8cuLJH+TUOsZBFsDdJMASvq
2TNUYCM13fa2MsH+zNm3xfDUzjvkgyISwxBuqQAXH0XToxHNgW2zS116WsaT09bCsnZ31qDB3SUT
E9PdTHq2TQy0VuRVC1BDRmErcEEJysnCZ8uiWen/8LPbmJmhxPBHd1pRtcWCMgiZlqYBfKuaTHK2
rvLA86DBrsm7gzcffVNw1LEGR1DmvPYkkFTSLFKfEcz/BMJptqDTlpU6ykYvHDT3SEfPJO9dm3ji
bQm6gLFa/F/9RVvZioBiNrk5PmdIMmv1oUYbe8hDfGIYxEYHMrdYC5DZPiOyvLLlLnw8MRjx0gNT
J52sfkA7ZXL++/d0bWr7O2m8kSZNQpraIWyDkoLok1cO5MSh7HuoK20i98ghlAAi3mVCKJNCWdKY
oBe46t4gtfNO4B+EOqZj8ojZaeYycUapvrkQnsDf79YJ1SbxYXKG3D3m8pVu789jiFI+izERb3dw
k+RaCS5ipAtmEOKKfItCvpjL+EFYYnjbEpoIeZXKL3aP/p7OS4GJzAnGOuB3qcdnIuUZ/SwjcEMw
PMHxYn9ypb0/ODQdP05zLwGYKmqKH1TZoVO7H/IZUn3CRgRz/3sScAYymdiZSa0kB4D1ZgYvnkIb
kdDHPyrTcbsyTTMLNh3AEFQd0TkRFAMJhUc0ebe/RcpPIrcke/HK6lRV5gsjgfCkNIiv6J38E7nV
mrEVCI7vBeJQX8r1szOoOrwHy4vKsmealgfx1IasL7AxUlBqwSa2L2EO6tLiQ5OaRpIpsS0fANix
kh8Pl9TdZcvBooaKMxu7kzo4oWWLZGFimFixPuZazcgr+HOnW1bOd2ieE1pbHW8b/vzdZDn4SrQO
hDqriXhYVOhJv/zeWMXxjWOIkj/Bj+0jICvmwwNKe+toCb5WBeE+Tb/VXiqg857/xyXD4rpe6Ljg
pxERQV2+ouKbMi5dzNy5lKpQSveW8VosAnoOjAzRVtIxTaPYKbM3FfO8qBokR8EO2SqiBTVKD2XL
9NEuxKOJgZMKTdN+rUXenknPP552ObWIqh+pf4SDael2sZMZ18nN92ya48t9E8zw+RKhzwMPZfmG
q38ZS9IeLSbAwtYrNHR1RZ1m3a3312oQCdFys0RUJfK3ajlHLVGXnCcSsjFzW9Orw5DYVq5/LnbS
4HdqpHXhnuv01gXnF0i3+qG52Y6K834H+tS+rn/lPr8xPeXk2v09xn0r4Q52ntSAQLmj8Rf4muhC
XD91d6FYJQsNgxwXQ5hDghs0J+L6Ezc9ARL8gyul9o1HDqFt8ELpa9PEZJRU6ZdQr5jLbq/erphR
G8npx8B+KKKgmPu5S545E0ApXLKPe1OEmWJzuzNlddqukDHdQNWGKpAPFta4uUx3KdKOtfhldza+
lWL4hmp6HS9IB46M/jFfNq/7UvNcHrYL6puBlO2CcBhdMBtCC2E0kdTlU14RHMKEuHETh3xqsZMC
aJZT4SPP2xjhtMMoEXtiTiy4F3EDHiBopazVX/EuqvilBc+QvvPbCmYmX1P9tw/r3JFBh0S26MFX
WJsO4wiyr2pnzxHNQnUMFhb/9N6w21LfOF/A3/CXzXGtpnz0RvOlSOQOQxFPpezVvvGaZSjI7+gW
DqXG6P+A4uq6uMJp6WriFkBY6SWYfk3impFeP+5umkOLghWFxuLJ/XLxalscFR6eekggTVPKvjwB
xB0taQsFofJXB0somlcOa07qFwyXpWcZE7E1YhbttkbJc5NMx63JUEcmXXesflXl8M0OYhZx9/H1
WrELMB0kmMeGHo4Sq2LIlP3uX4T8aoMQ176n+x4AlVJtNZdyLaOBLfD05+FLVPHnr3GUVZUqz5dK
vkza1h9YqPGFtqklgMNS4UX87qRqh2pMBxeu6smDEtDJeO/MpOCQ+iXeOY/Lm++vtQEEQYbIqsLy
vQYrIXsRs1epxjIaL5ecAb+HA9ocYY+6nS103NHT/EtVcBAmH7cIcuZQwt0ST/rDwP5RVLewMI65
Ma7WOzPL9AZnVAQrrfLHTz3MV1Y0NgAkMQGhtQRbWGxtZnDaNgxZeIKS0w8694iWPJ1U4VKdKYyw
SlfLRoY4CQ6Air4GtiTMhSoFkaxGV/mgRT7zuOMuoRwejIE0CVc65DEKhACWTyQgLITj8/+7wU0j
umUpLkmMozyMMIYtuVi9EeOsdgsQWZVBlHAU83NL2t27Qotuk3QBTodtkdBMIjSViJnuh68hip69
CppQoFratLOktKlpJfwca4/Qebd1g0pqPNBAQE5WprPm9TRE3SWPoDeW526gk4DbJxF+J7sMP1dp
Nf86ek3ZcIYoHC9d3N2qLZoou4U7tDbV0azNisy1tEG5bCgkoGqm6qUtRzL/aSw/jmu6Jlgo7uBo
19Je/CoxwSHkoEeloaAD5PZn8CfP5iun8AVoI/rgbAbrZ2INA5Hrq6Zps+/mdBzyHssjdLvzT9ZO
upb2gGYtmnQsF+efAEG/p+MR/IzgC1sHWqM9+xP+HENtfapVk3/+nIMiapOon9Cgy8gdvVPSXg5T
LvzKMBZsRwPM/tWvKf5AIaFxes6Zhsdh8PvtpLS1SIsZcP5bWHXzaW7WZdgV+1IdSeQxszUAkYc5
D2DkaFnn4Xg/c8dEXlAfIF1NmaCHokUj5J8Dhch5iDV67gOQbr2wz9P7f2zILWM8h2j8MKOhLK2B
gq2wQLk2mYECJH6Whz72//z137m5Sz0APBUsY8F4PDc5tVSASm9jP7F5LuBXKu4Ds+x7Qm3ThAor
oGV+GJWuwzX0L43tnP3xicUj8lCOCkP9h2mjhHm/Z3ABFi46lW+if4hOt5weW3S5nTEAeAJdwUR+
P91eZSc8L2rWeMcly7jMXVEwdEbYVYX9+U/MCjureztfJFNkOugWUo//l7HsWmdC2zqoXs0PdMkF
PIB12VIfMiO/eE3XDUMaRk7b5xdjTQ5cQj1lL1b36+Vap8645spIITgaKrKfMZQQ178CPmRTXFS8
LGfQ+EykNYUS/lcHdrXsW6mBKaIvdSX9+gb6X87/EiH1NcEPRv4Oke6m8x6u1k9P004mTxRxOye8
jGjsJlY/7wWD17ULeRBEs3H0qZcpW4X9T7S7347IK+137B7TkQjlAcVgeRlUEFG3j6kin8xZ3dlK
1WVE78swPSe79SQQot25rZbbonWjBJsPRXJgDT+3xuRoPMoPnK7f88/c1vjb+9wppqnJykm+/gT5
NGGloc3MwgH4mbv5xu1FNjMTgbEeme4rE/aWf/JOXzP/C7L1tqqL3ifcgFb43/5EUDbt/i1IcJ1L
KyJIuaRzZSz557thjwRWGNUeaY65uyYOzrBkC8hsxilagvgwYlReuguBOexo2TOCE8+hXqioDzQG
r7f6Jd1Rr1TsLf8S3Q2d4i2MSlUr4/GCoOTq2MskFQ0eRfqeJtPch3fEemwSM3FAgpsKZGMCHBSs
OZ7ER9iEKS3cGxjIgNlnszlCF97ab5IWX+HzVzgEVZ6CA4x2WTtunIVBZ1o3k+TP6Zem+zHiSBuA
u6rGWVMvW1a00DPsB4ld3vHYWeUUKGP6u/E3iGHa97fLDLV8emjf+o/AA3OHAZg7IsPpADTdqoYt
rwwdV6vT82Kg6ob2BffJmHqDktUMJ56MG1zyaHKYxzOdLAyotjAlWfmArd5k8+MtgRP0FLYiofW7
9d3uD7Dh1m337QZGi/Al4u9V2OlS8U0aT3Fhwo+KSVvz1WBQLhe/0lpQfK89RsGdpNYBiVQMQ2rn
kMni4odLTCYysWRZ2SVlqzEujoKWGEfv6GgZ+XM5WIMGf7zAgHYYPANdkvntp+byBXrG20v/OIP/
Xi0igOGnnSywA5hutRIyVzLrywS7huFeVC1qmfKfbH/uGB9NdrF26WkC6ut8+FN2Q2areoG5GC+e
G1fU8TWm2LI04Gb895wfeWpa42EGjqlShpFZ+wVGa5yF33bKKtyejR5BoKQFM96s4+EKsJL+dEm5
lEwQc/+0yqr8Nj6UTTtJfWN8BE7NCtUlTHfpoXi7qN5weARbE8BE4SVvTvYD9c0gLmJ9fpFMLFdu
s0v1VXEM/qsEZ6/qR25wbcQhiOsZFfmb9dP0I0XO8yopE6c67+gvDIhl2sX1vVkmptGat3xzVvSS
hcl4Km5lEkERwagCvx+s0F5DU0c2o9Y2BL8tp8cb12F42IIcJGba3g8a39DPa5oEHsSmfvAzqAT4
6AKKJ6wxZWV8ximN7XRgdk+BK9llJATMpY5CiqF8+LyYvU7nh96rd7014z7zf/h45gNeIjlitz9u
NjYTkCoSQJyJkZdvgoQ927R21tuebD0lF4g+wAx6A5hlRDe9ou09HCgeHDuSf6wmuFCpbjJHf0XG
sp0oXpGSeASy6Q99UjyLuko8J/eNeGceevrp9CN6aedieZLSI+fjHONhOIIaBg0+ti+Xz9R28NfD
DrDcsyhfummxU33iEIyf69Jpz081hqngCjfwB7xYIHa+lfvkqqVNHpTazN26QMfyC9f2JOUpEYsG
lzj7V76rC+Lb8qfij14TGt1zWFzqa3lLUyZrftbsJ/dTVNduurmC9MkpE3sHt5MOHlF1ce8ebH7o
pEzrT8Sxih5xak0U+Y8OWiKzv+UtKlHceQDHmPCl4mAlG0rXpKkdFrhQ6xOsUI/WF3jzc/8J1kmg
G9g5fAm6HDAQyVj0BrSIaQsnmba1JpR83CxuVE6eeYotvL76fgo0pfLzgeB0NA68SngovQ4VYjAN
pa7WMW3FkVqB/uGGtSr8GdqZv7exreRNiPGu8Ht86jQ+hGhPsXuPZRZHUBMTHUFNHKIaysp65ZQe
7nba39qpm4EofOCEXTD6Dm6iZR4DBVGLdNbjH+II1PXH/9CyJeICTQUpEJKlVdKJMHsCMSf3fTIa
q02sx8pLEM6flI8d7T55iUteLsg0qyq8HgM6UB6aOgdvo6RE+9lHT/tj8CJPyylOb5rzu9aoxf5Q
+I0539XELBPtB9AFNeRmr3TrseLO5FWvk4l835dAxh9vVLZsDVwojGD6Ex+1YEi7PYXlQfZhltFV
SG5j877btBYbzeTCkQQl+pSTeCKTp8UGNQeMEkxLAdYJwJrSWmAOvck2wG4KSRaLgmLpxkjHhclB
2kyc4oz7zdOu7Z7wGAO3DYbYAhAiiutjeEbFTHwjo3yojaTMs3v5cuQ5p1GmOwk2o1mTrziSiKNN
NavjhGt69S7GpuU2Y0f6E+RrqqhS2OYc6Rkxl1in9XHhhZ+SloTRomYEXwRRc4Y91Oh7NKZhdXg7
L2RnVncPuMQ6ILotnackJBtwQ+5Ue06pZgidQZxberjnFmz0rdkQvQ31jrcq0vDyWzlYPuFVPwwg
HUatEEwcs7b7dNdzqjLQQpVw0iPAafXdCtiRsq5oPBswJIkIh+cq9dsqObmd6gKfiLFpk8ZVAh8a
o0yB0h9sj8Y/xFSlhCcFC2C3yqBj/KZuA+2D+a1090lsq+P2/OUHLntUsZeer101Sig8gEXBr4Gk
fPcx/27KZnKdE9/u/IEnna1qmm9cIsXALRkP7PlUreTm1DcY8NltwQ8TBzTEfvxuygrkt89juNfN
KCWG5ZCMoY4vizZmBmhsgOQGf9J6m7kFaqv9nGw4QD5iMW/ZafBEJ1fmO8oHq1C5ZlYPFNb3GzIQ
hTvSY6QCnZ6M+zaiF5mgSvshOtwtkOy5tOtnBV+8pGmurcAf7f7rlhZrOIxMWej0ykABnbwTsVTJ
H+ndFY7hO+OJAXx/Dfnli9necuHsTcy7orH+yxNy4yJk9zGc0F+OPzXgPKpffwIfQRT5I7QD+sv7
q/aBA1Uz1JTXSqo1S8NROEfgGd0h/149h7V+xKaCTVu/wGOJGuSzggSaYRWe9vocyp5MBQargVGw
aTbZ8gxWo8tpP0+fmDetwvlgGjSPtHKOfytpmvFoQkMOVpJC3lY6xKnRrS06FVEqWikSH91awhSz
mtp6dYHzccAxpVfE15tzfFu1VzfWXhESP/6Xcyjgdrla0cvr2lIG2l5IiPcmw4KvOm5ADzUD2Xwg
N2GDitTXxqDcKfNGgYuQIMCZH1Z9c/MUBdBOheHJYBB/20s26nsSe6WuaAZMmBPUXbq7kMxRB+Pj
ztjJ5xN47zwNHCtXnMvR0lTw3aiXaE7ZQNriNc3iqqBm5P16cVaoOSStiGueUksy89fxLE7Ko2jx
42eVnwFPuWn4kh09AWudHw++jkcwxjVk7e/8cBfw6EoHA4dzvk3hLAWrSVxf/PaqHijXsHii8e9s
+lVD3b1p0A+0SCrXWBnpkltu2iyUrJ8ZxOe4x02UzIbyrJY8tsFRBE/nLTcxcLG8B3MAvgSgNSzo
P/aMuSY+Nr1RfJC0rah26l9QZX78YmlLPWubIARYZXrOfByo/TiQ+7z+9LMhFdVJimWfA/IEryX7
G4ngHxJcQq9Wc2JmnmCiVxgvBvvHW3RlgEhRUvyvpdl1uKHBS9wcp4Yv2TB2E9NHYqVNNUBvgdiH
zZm36MfhHBrI2e4B5pTfrMiCbWdZCFDFN/3A++SPKrBqC1c76npzD0qvv44UwIT+qypP1SJpGVeh
rrfXAcBuyGXTDLlnyp3WLh0xKdXFHCEfR6JquKmcV3NfqOpJmr8BKVWYzvqbj6wfTCyuqk0YKynD
w5ISiF2R8ObGkiMn9U0jMZ6UmmEZvDVGrAcGEspAPmdInFtnaodPkTFMJWBtmeyKXdCrDRyWvnil
yvkErb7NwNo+Dwzu5j8FcywawqCMN2KQbsS1MyZT6Tg3v5sd1dLYkqlpnD926J1aKVdMxxIphDI6
uTrOzJjnI3DsTyb4P1XRULdRiGKhHCF1SXZfNzou4AADNEKKlPTjyH97CFB4k0JIeu8RTD7Qlchu
YwhT6tosC9inCCrEgWKSXFK+p9h0mJAl0Wx+xloHygMFYMIgQ6IuKIel3o91yfVjIJdeqQSshOac
06yrNsJlHRMsrZ+4Qx/0GeT97HLBLcRSeV+4WjwwRL+dIpOx4TWWaCPjiZty4I6fuFlOfW6wZ/cy
OKZMiTJviwAryp2JDE6NxXxMcqjdjY3JLSv178e3Wb0f5O4+jitsDasgl6GBZu2A/FljYRsdZ+Hb
35xvqqXjy7aQJLWIF5/5j67kPdk/oRgMl7/dLpjXm9rQI24M7xofEnfA4sgRKhtDIH3IrTFdxdJm
GbixdoUOJ0nNuIkhInh3kZWVQmDmvgiyTqavh95ss5Hm/N7ryqviTxQlspeNpWZoXFvBBrWjRYVF
ZtWzt5I+F7bxL0A0F9mhF71H4H5e1Gjh9oc7PYb55q9mG6kPJgau2jcbTZPjjMmn0g9DN+7f9jEX
XOUSos0Mca19QX2Enek237DJXSqZmuf+xdIaI5bgnX6fcGynEd8JAQVaf+2YfB4RYskB9WVWZNFa
mf9Fivse8PmrFDI3ZeOEU00YJqYUKZpP81qzvn+JAVPpO+gy9e7waQjf6pwL+6P6+9EQCaxqMjkJ
PPyJg0ls92jY1iHaoLbrpj4HxvO5ioWHCVHwJqSiRH9+R9EJKrLEW4KSE9FeMWtD/IM6Cb7N+kkW
vF3cCMs6/XPiLljtKaJz3ufyaV7XSS0eupgUKJ2KvWGddY/uAlvVxNSu4tQA32HuVOXLp0rltjfA
H3Tyl2aYlGCcn4LTduamyZuJopm8j9l7MZ95a1nJFzyBzvGURTHgInDz+9Rnp7r16M2k3yA07Hiz
7rkdDthkB/BFGwVWX7vBRqQHGxbAAFdvR/hRDes2fTJ/tzEEF96VhkY+eeS8qb8g0oNYPaJRe0XB
Sr+Adh44oMpx501VF+8hAyImqPhbRIshmETabiAqK3pU/toNZv8mRh+3YDS15Lq/PtJTGJDMaY5y
7/zR09sex+7qhgKMzkZy1uRDK4GWDQtwzJhqBCIdUEdxH57c4J6niy4+wIw7hyrvMJIQOcKshs3X
T/SQlpKaon0WQ0rzro4zVYlt06Y0tuI4nLPZdYfmjavcl8EMCo25KxIIkzNB9lIRKGBs9T3IlDwS
WQpQ71Xod904QdMqQT/9++/RhLUuQSMrv13tR44RYN5SfoMQtwwu1220QxA/v6u97YKNQ6rRFygZ
5Y+dfwkTzzoW+LKrWofYwoB+gswOEInNeZvRA1eQLUVeB2RjRZs4qdhd2ThPU4vVsOuo8ATQiZTH
QjK1b2Pi9nOypR5cLGqQRfflq5DucgJAMB80HPLU09lDiWKJxnDlvlHBAxyhsrcXa4cZNha5Y4XF
kSteO1ccydsUI5rmDjGNqUN8xtuG8LaWWO0i3EAKbGO/lrkUFCIXe8iyvgNJ0sQLsc8hGNap4Id8
rltzsLPGFtmUPpiljeo+F6vGaGKEIDEXRuZZUD1l8KRNlm4CUYtfjyIjfmt6HSCeCKVthFECOPiW
GKmIC8KMQmFao7CKPvJrHcgDrWnHvOgviq79DXQF9pGmep+lXv/BfQsS1whAaAvJeddjDAFLjmNM
0mcxPof9UyPEGPCZXVE7V9ZJhLD11dpfFgoqQVVKPCke39fcpO+UA7iwGl/Pk5c1opoxCb3sZxPb
szj655ZDk+8PGIy5JtpNmzXTTnfUQ5aX2fxIuNxsGXnCqg+J/Qztbv2Lo5g/GTQQvdDDxMrNa+Cy
GN03fs4NFJZlf1/SW+b6TE1MN53jznqcNkC+7IeFB7AspqCNXf5a4z/SFY3YkIY/iRbbJ6xM4l7Q
9acosmPfpA1ukvPFj6KzR+yXOu0ou3LRY50ptlRUgwA86T/bPJo0YrddoDnlvpZJGPOyFCt+ga/4
GwCXAN3bFASq+mSIJYWnQlzrzFRvLGw8qfPVY8RE21W/FfmW9jmhEVzm/1dkkuhEZbCQOMsAHmZ+
e2JnddrmWCRvjRl42NfredVWe5zp7SVTAUuzAcbxQ0EV6sENja+f6zgptUGnVQB+widRueBn1w93
BCva+WMVrI3FHy2KRIq9WRwkbN5B+u/3Sk1xHFMFTdRQls8kLzmu2MQcAZuELgSX2WRKl2y7RCud
UwFxwY/UOS2x3YqsrdRvGUF6n6hzMfraaj6YUeCeIMhO6Y8PmEXwLnpRQ2H4eBcdqoCPGh9KnweY
zR0kwIFMYH9G/ELCMrwp8L/5eBGDVca/mT/7ILS78CJPR9sTbUbPBD9aNKHMG+2qDlW7Er+EHYLT
2hk/H2dFdvaYm/R+emotZb7janELpHapSOgGK5N6INcKRi7BTep85OE7rRdCyqswfRr9ogxGHUC3
fafr0Y0pLLfGJ6T4N8sCgs1uaYKlnL2eaoh1JN/YqDJ9HqmBPPGAbojTayJLhrnAiZ0F2SkAl0Mg
sP06F5i0KXuqicQgGHd3aSij0+3aU8sfVE/xY6+q0LW8wkaZ3TpxmBHZoXHuHuEfxXVK0JWRDdZ9
yoREtB9Y7bcqo91VdCfspL4MDNo9osgpNjjZjA+nAxpvDAWaaHrnIHK5nU+nIgESKH58NL86W0+h
qe9GEEdgFHiwhsuLI/tbKvezwk8fxYBdPev7irwl6R5dRHRTeKa2jyXeHNHRlvDk+2DJgNVpy387
vQC49OF03CM7SyaX42uVTswosf4rX2di3Hrg45fyg8mTyZ2Ke2DkYtlNu/J2L6liPjOjVBsreMdj
ib40AHjNCouixn7sxhShJHqdXn9CbSahtqwfV+goA7IIgTCy/x7rRcMMUG5pmDHLItFN87D2scvO
dYDyayBN4MZvSuTvS6QZubn4sXnq6d8oGIbRj1R3ZEPeaLEXXYjWRsiKoppGtFxnbCZjwA7aM9lv
GatM5wXmI0sPSRYO3Gr3ZUUQTZvxgzb5M2S2tPbQ1OL6SPb/Iv3nGJzXSEM3tEo2cWEPC8RLHkXa
YrDFS3kxtvmHpdnC0H8TQnpdorz+HDM0d0CAip+TsHcKW89s4YCUZKSYB54uOtja8yo3FCMRQkBU
DGRYcjiX3+/gOu9EwUdWYYn2bcLBcWu3TM/DKtOYRfl5RMyXsaPf/cBy6uhOisqlEYqfwKixfLpn
sUrlJGBNuPdFR5Y2XFTLCdIQDc2xnGZ/hT1KhoEQFEkhFOBP/Gd2MIwMUOzo8E1eoF8kkTLuZCZ9
aacTWTO/3Y6Z9QZ3DNwGdcb8PcR30xUiKtwgiiHAapypIVRbT8Feq0MTGd47FjKRItbUv3IqUeUc
gvutV4qaqnbyXxRkkrItOo0YbW2hOncDgM68d/fLk1lRLgW+SRsk/1XqmKEHD1BRfqjrBZH3VNq3
1pfHhtnpi2CTF/a0MbslDSdDP0hPj7+tJZnKHdQ1AI4U19tTuC6srtcGHClo9S1enqdnhZzvOZn8
eqV/5FulSvnmcvcWlFg0uNMxuRC6kebXFg/bi+f3hwdLkWF+7NZ5+7GgdgwJl0qMPLGza4UtNYR+
rTn6CRnu8yqXtoVdVQ0b8V2HbD/pG7x2wsdFJwuaAa+UV3MLXwZ2msEAEufSgHOsRaGYcemRYky6
Q68aqHyggTINzrlS9dOW88XIkhhth3tYwBfs0Fk6oLf0wFDsg7zDWBA3zeR2guFMswNPjWXn1PcH
KIYbf+0y0HYGP8dkCdcrH7SLBQKdI+E2FA7OhCX3EWS0rbrxABt+NlJbiM44u6kPnQdnsHRq5cLH
xZX+yrjfDtmZq8ZLgr0rInOENGzXwKxmNJtEOyczZChAOm8WbQJE22w3DGx0UzXMrETBJJdpGt25
YRVuBRfzJ6BhLUkbEwPLWY3xEVBvlzh5NpzROWv8e2dRp3H+/dnDiuDa7RpdtOQjVokz++2K25yi
jZ1N7gNZSmpf2PGjEiANLNfOE2bT6/gPyaJEUzEQOjDTWwh1PttdmVUmh+kDxaNhdiY2+qZfZl8H
XxMBo219Nd3YHwD0w8QmGwy4CK5K5/QXVhNQwl0Ttc1yjV3kwsknOev0vi4FUL2mw8wb4DM/ogcl
sAUiXcY4LWUQRL0GKcbdrtgeoaN2GNvvrZ/kwidFs05cYfFErY9rjDeuuAyfHAUTQjb/fdZTLWe/
6uw7yovqxBAqV7MhoiAJL3t/CpwFmS8KUWaOq9bzZPHqukS78mFmkM93oTY9qYEvFP+4v2aZSorm
wMKSyjnJ4C18bDwqSCsdUOWAvLJXYCTEyKQeD1YYxj3a05Edxlp4c57XbJfNdLwywnHxbr0IsymF
7MCoC9GhIKA75BiNgieV0gqOyHUTxKzNGF8xIoqlBO7q2wO5ZsHGkluH4LhXF3Jo++z7GvCKWm9H
rSwHaJ0AbKAGx9rz3Y3gSejriP7rfqX58+WZ7pw/yzwiAC3DqqsCt4QyfpXjQ8Yn4o7L4G0YEnW8
sGnByzN//EC8IDYkEj9qZh8C9lDQWR8a2Xlc1iDjZs8qPAiHBaXAq/KvbgEklb2QEtbFEUjVSR+f
AhMhvWgbss0KYmu3mblUqYOPZUGz+GN56nD4ehWPFf3/mH0e7hMeUbLdzuvscG4dxFqBq04r/vSg
nzGhvLPqDxLGBMlTn4s/OJeBhbO3GJYXRWy7xoq/dKxkF1Edm07nOESDKc/H8362hlM2PByRyN7h
92io7bWvHCTcqQDYwBeS/NeFjwrplb5xTcfJpvq+Pngd5rc7+vce/c5Jm+G5xv12nloif5rFMQk5
/xhiZu37xRwHsh8OQf5P1Y1Dv3dgNvIMyNCTSmHXoKh9UpR9vulK1braMQZXOivCK5Th8Qjq4UaB
5WSkrnVu2DXz3vJsIJohlnwPafedPQjm1qR5MFloKxCo+ckABKBpasOI4lhhPLF4m3NeZjzxJ79V
c8IzAsBLoomE3oJyAkj7EEFGX63C2UZBygoAVm2ZSg6djTytR/OKYmk1qf7E6riII3cT8IG7vSJE
HiOehzR2Y3uy/i6w36i0T+TGXwRTiSuuPxVsIbuaBxFRcexCgqKqzGmtwKCryOb3x6dcM6BOHGIg
jfAjASbLa3oUPJE9/LN7KC7pD+6HZ5Qnhc1olRH51yNoWuM1/sDB3BFUhSoQ/doy4K0daY4EM6Av
NiT56z4fHe3ZJhNa4b2tBfwyPsc/0o1mrkZ0awHBYRDDdJ8XZd9qGchP3IflOGp2tDjRqb+7kuXR
SGCJJna5IkG7qX3wZYyZIQF1cFKkHB0jF4i1jBy//+W5cgtNFFmNR+pXduZ1FW+rWsbCgL0bZbNO
MfsFgtm8MCqoQaktyrK6JyC+fJlaF02uDhwEVNHdjbwzycy2CyyQMWmk4lEkuuUYFKbBvU0jlbkb
PMcVQCCeZR2O5IQu0i6Nv45sKnPxEkSIqiYcS4GTF22N8yuQMVQ+kM5b0izmsWqz7zGr5vqoAyB4
yRLZScSa2S319Et/oq9uE4QyAvQ7wBFb6S07vs/qe9YUniJ1FZR2MNpkqzItrQIpQEXrkPDhjknl
xTuit6kpTYZTTAvySBlagzvAEJcKmJC7Kc7T3Qw1ReMFfXIhp+HoBW5vxeNQ+zlZjDIY+9rlxJcL
cT5nQ3BjXaCBOdGUlesAI7z9G6Y7z3pEewwGNBaLo4N59nWOG1x6oJfxNeIvCLo7ooepqSvXax29
R3hILy0nJDdnknXkeoSKQzJ0ruFzeSYZHY5hZIErXfWMSk7P+faPgywlyMgmQBi8r3hEiJxbkYl3
FwYcqfu03XtWtie7tWyRX6fMF4u3+ft6HePWGDjkTUDyuv6i8JuFcwotm032iOirePodyC3qjsdp
whvorb2nKYVV5AOH0BmAPGesvoUvWnYkKz0Y5+jF0LAiYaW/Cd1G0FwfOty44fQQ8/aDpdM3cseC
dZ4aFx3qQsTvLYk11HY67PTurxvVT0LT3cIELdXZtm+zsNxTOSCUuEztsjMYFlqDio4tetruabab
B3muRQCz2kjk/smFXmWVj3AxoyZbjVv+lke7ewmznvIOHZw4msoKEIYkIz2k5BsUBhRzlVMDG57C
4BGxy2VavCS5Vg060bL9sdFYaXam9DK8ZyLekM8Qv81CGerhSIIN0/f38LpCeb2sphOch0gY1tti
Fi1Oezg4H5E/ISoCQiDHEYTMqkn3sb5E+uum+tnu8dmfYfw+toSPJGjMoqejEwH33ZUbMnYYf6ER
K2sYAskVpz+roGfzmdL1/JF7YrnKMZHtVdmRhAYIDltCvmtNfMQwHmEWXir2sL3zv2z/gv+N153h
BxylFJOUOBfC5ElCSJZMab8HOLWkEnsTWzUhQcRUV2rjeDr6unrKWYmTHGnFo/I0HFjyJoLwi5kh
hFdkf+koSzgN23dk4bJfmoqSEQbWc39uUHgjn2GGzDLFvbU+8TdMer36VJzIl/B5osRplTnEE2h6
oBV1nWeMhuioxZXHcKj8AKYm+4lOZqDGt7Ky0kEq2SJAhf/w3/AA90YT0Y7v/VIb/Y0sULnUMhDc
ImFgzCVbqoKt0434YUNfx3QLea34TckEXebAZeDlm0jJAQJ+HOAOUlBXJghUAICh360GawcBL9FE
ODf0WHlguw5cVDaJR9NnNRPKQKhlOioaJhsDbZ5Xm60seRcQYGTH0IXZgwFPsvIS6WBpjbMbIMky
fx+bDedqhMQfzCcP/TjLI2/TilrwSDX4OpRYCFhTadeUui+CmzQGbebT/zQYoj35OEbZuutlhUOR
D7j7POtPCaGvvbyvAqy4ZWs4Ok6oe56H9aBLF9nUKn76IMSIvhWftpWo5+5GGUim+NWTdmUCIXdC
SDZHP6AxY96RkwAUIqDjG4de21heDksl8Hrxt5WZDixxaAWjkwp53Gasmh/ilD5TEtqQ/6mEPE08
OLfBvltNLsHt/NGdPSPDl2fsPkVTKQ9XDjRNZEpxY58Hz3qJZGvhodzRa+60DATOZz5SIMczMorG
A5Sq3wl3gMkNTHQ6Mu7PQv+iIY2yJ5gz3oucqomHJGyWk5g3k8Ydax4b9LmEFJ0aRxqZxffpQFbw
GYX0ko46MAbXZpo2OxwWR/OCae+q7ApDpRNlWIjROUwMRaHKFZH56KKoruc+oKlAS5WmOoEk75Vi
RpheI8M3TZx4h8ZYJylB+EkpVaG8LJOi5Sfs667SMCUAhV3iP/dUA2853RaBspD59VH9Tv6I6Gcu
X+N81OoUlQzOiXa60btTtJ7Ig3wwkAMh7OVAmNTRUzTeYoyfltDPyq5D3PoFFLHWiXAi4XMQgimf
wQXdBkrXT9LH0UFkysirXJu6a/rZSqljELBZkm14q7D3lYsldnhiVQs+ye/WSqV+y7HxkUeZSrJD
52qgV+6hOdfb1eFXay3U19odn1kcSw6NvzR1KwXnOL2ECt1Ik8DI0emNfhpK/5Ft+JKP+o4Jvc2s
L0Wvo66WyxG4jvLAP+N73SXBhyvZB3qJ8jiqFI3q4bByxP0Hpak4PubFx9IgKgZqnn6uK+9vGQSQ
1TYjs8pStdIiM657qG1rLysdm4Dc//VU8qtAphMu/ADrC8pqdZ2gG0hV/M+RpYSIPrbC4LlkDrQa
lysj7utpdK170UbcoDijeEkVimgkp7L+ZA7AmYrf1DLq660F7wxq05DxBvmJhLOn+9MISQuWg3fb
pHf0pRYracrpeKxt5cjCzc4MX5/pxYrE00jWxMMflDGx1vJKXskOuIys/u5v/q/YoyqC9fG4RYif
eFc5Vne78fiOtQf9nZxTA3Dikk6xV3QuwIQgwGHAgE4L2WuOH8eC4MndtvmmVF0Q5eGQDFgKEqAq
30K5gqh0TeoncHTyeJx5bFnVEmGPuGRCIRfNfHEWEIhLAN2CgMRZ5Fu7qy+rYxR0z8tkQDLRZBuX
KNMLrEaNfKwJZwbOnmemmWwKlNEMdpb8AlURfu4cB8egbEEHtRyf6vWamlmknK07bOe2hU0CNLyl
3lD1r6jH6PUUl/JX/Xu41TKvM2T+h4JXSzkB158Wl5yTHN/Y/qLglLAa1LjTrk4tfY/B06nYVupp
Y9PixmrUyUYaIIavRf5QWsCsZ/PclYFcAy74LIpavOkvFypImYhVAltLJPQUfHyZ3YxK05/5HDx4
HVy35qq2CM9nc0VUsWkYNz5KuUv7KhOTJsfjBwFx7+UHhKKmBZWoRZKHXAuTs5PSZQhyxZKWO03A
rzT2LbbiGDYqRJLITwtefNNU0zJfWlWuJNGaZtIgB94Astd+GlgGldi9vz7RFd3MfxeAFt8eDGTh
t6p8ecaTwBqKMrVxQVlgVUa12KynGzXanKcaa/jySzfrcVZJcCqw/mohNKkcbtHGbgIoyzcSG/NN
K0m0/bJXb5eeyQ+bBcWeWKEUMhBhviP5GZe1xE6VEDJghJVO+RL1DJ7RgpPArW6MDrIiI2C3KvUg
x7BnifEJDUXxk+tTREtpsITxuiy8DaG1w5DZadLVK/gLbfBFrNyIZ6KQZPmjFj42eDqUPmwkdQEc
dShnsHG3aMKjIUykiCWQAt92Rddy/I08Q4EqtgRjyZRuWkcqQ+ZqionXqz6qczetbIKk9hBpI9aw
JWFVzSMHHhnRB0zfqfT8jeCLJmxJIKqcyDmdQp0Gj0THttsx6OVvbAchrRblL3x+O5C/sYkWwQea
NbbNfdYhJVd0KdHVUg0RHx56IMxup4XIQl382P+O/+bItHBM+zKmnppoa5yc78CZtysLvr5pEjx2
8akmGiblOgyGhQVUO0Is4LIOdaiE+vELZYU0467/wptUlTlH2Ll7lADZGuWUQ0I0W4XdP5KfUs6+
vvTjmRUuKark1BNqreL44FvhyoL4I4/jNrRGx13MyxdyouuEVNrLzqvDp8DhTjUV1gOVcNSMJlsK
k2026r0VLnkykVVFAv10dimpbWbyQ2TuoIwa36KD2XKYPc+LWhYERPso+w2fPlXU0V5uGCNlC/P9
urnLH25j+SZMOq6LkTvg2mTRrCg7zQxQik1W4gMBbUM9W0XCz+U8NS2n67KDdgcBwiG2CEym+4to
G9whPwo2ETvUQH33yKyCXVT5hZhtCKaC18pyAwxpUGuNz8pWKDuvAGtGL3drOstWhrO5vBtirfBJ
DjrUACmp6dQantaSXdIqN93hRloNXuLa7X/uQ2twLYWn+mXHharTqZgVXVi6N6KlY31NLD9qlyWp
oyoStRdpGeWUu0wMekMPdTVaki4SVToI8MDAVKXNkRIiUGDql4hM1PiT3nllSDEFVRL+Me6ZNPbW
1907i+G0N6dDF8l/3yinfJEuuNOljWlzb16Rq9oyj5uG7Vd0pNEzFQJFz5PhzBY3HNvJKSWlJkEV
2SYkVxFownM1r57l8ooNUlQ5G5PLyoWtNfeh0fMDIc7T0rz4xIVtFiAjbXkSlYkGxgTzNvJQTF8y
PUKbj4rbsAiJRWd0sCHUPLHpQTqS6wiVmY4a+f87IKKBcApAK+KY0GGFVHFOZmM/WOUwayvk5s7X
8HzbQNEgWVB6cfnRMiurdSozO5PwrI+gbiyLqaZhIGLQh8ysWqOv1C/tF2b2xzhjA/7ggwKUFSrN
czTGmalWzF7Bq62AnaGPVfa7rxoEjSIOU5iYXQPrCsIjye3fKEqV9mLx7BhCoL4E10mhBKopZass
39pxxWFk+CbQFmAk0s5NXtCEnc9Ll4apD4wpxN21LNpUotJX7kiF4bZ4ecIGVxH1w2fpC11q+2iy
f7PwV3d3O/QTpOOyLrUNelMa3TcR4FgboSl91uRr5v6YORkK+Io9STMNeOKikZy0lL7P1guix1OK
YXBUf6Ku0nzVVajUNjzR3pBepsyN9OfWR9W+E+t7bZRB41DI60926yxRk47ki34oR/EMN1MVG4/4
rxcG74CgO2EkNzyihRjf8vVLLYWWCBoDKCwB9LrkR8yycpUM5eUL6e2qs45JGvpN/SZ+rdpVY3fa
QpQgzoNQR2KREZ+FboRM1wl8kMasRjvusr+K9wiDMq4nna7KMcbTvidw1SHqyHCcnq9MIU+nqS62
RIinLQSPynS1ku3kaUJOCAb3kVeWKzoWBTp0JV1PmPxACFNSiaYfgmRtTAwShVCuiZL5rBx1Z4B3
sDgi1QeY2f3IRn/cUoQGqheNuE30AehfJoyZtsc2yF0trwMiHNtw+z+Jy2+OmkCnCBFUoS22HWeS
C1DQmdmAOI89DI4uR2+aYeLdMLMmgapsUPYo9yzbIy7W3qtzMTWmD3uR9nt3dzudVuxKG6Lx0V7d
gh6ccb/BLJKuhetqUfVcaGmqaS7MNuExLz5BvuN3EmdgNK6XmHn/DmKsKvluQXHBvxwA5HI3vibS
y+DQ/7DAaXOXVRyjjj0unDQcm1Zw3njFNlO4g3R/6O02as/i/TjJLa12MZDvJRcOA7X6tye0AP2/
YRlLSFJg9cOBRCu0gMSUKLZAqTm8SFEAWESbSdQyhgi90aprM9YgIrRfuEsIOItwxLFqfXmlGGIm
AhKdJ30HcjStCRZpZp5+R4Y8fcAUOGNRNErkUadZhUERnHHYs3DIERsLg7/MFPwJyu4tkKoovvZy
MJTCR5ODt8CEgZE9k7cqieLeLk9A0fbRSuA0OfxzEFhqv1Du9sxEw/e8hPEFEhAtuoC5hXjwYBey
Y4Fwr6E/98AC6c9c/tAItQjG7Bj2OTonSE8KaOpGAIRG8vdwW52AjP9w0mIFSx+NYWPWT0q1GqxU
BnJUuMnpbW57Xi29ZvlJvaMGASZpLJSCjdlyaktCDPbDjktif3kZ+wkFSRcqy8NtKqHp0SHn0l5+
Eu97t5imlK93993+OxC6m1VkjxLUyS84jrou+GnAz9erOr/bQpQH8V7g5BGWbnFQum1hwDyCFqo5
4Tcdm+c4I/e3Rk/pFRgdvawsOlL1GZzpFTrAnJAtL9rkr9F21mcGqPYgBKJy6nXvuQsbiZNQNuiK
wPcbsrj6mmt8kQXo1zGZronb485/+JU54Y3DCgN+v11OaFs1IHJPxdQMk2pmvKOfFyLVgJBwSB0P
wJPOeKUrcrlcdM6e1ggIDlJ8xpS+RVvr1kc4c08PF6RSxyEPHbvo8pGDIEwLjBM/HBPO/SerKfr3
9AZ+ozzOjw2yNQLHgx6YvYZ41Hpx4mz5wSQNSLYob+DVI5HkYk2jDrAl6QeqFwnRHdwlPeL3aEko
Rs2gIR9oGSKZIwzW1rQNVQzDq+DZSUrBcJUcvDAuTdbewIW+ODnXEDKzoHSC07lKXwwqBCCEIQwo
BS02A70X2PB652yKGDabjkOflBdYw/R8x+TrUJzv4BhKhdeswkyrQLUWXZdpKQG7jmSuJrl19k42
fHm2utF1ibvQcou5Bet1sdWM/T0BuWOGbcf4+PYt/mUE1/Fj+UoNBv7HnF4zNp2F1ggTn19O3UA6
bQctGKrajemPmFi30bHvwRzgBcPe/jczscnmqVatgEyyAWb3jN8yfDnlRSqfPP67XBLkI84FMKas
PVE9yxtalHRCHdCVuKAIwnZ0HBpFEAcVpgb/nz11s77KMt3HgDPIcSl6vwqIrGnl7u6kDFrSs32/
ExvD9ymt3jU+n5OrN14eHLJoJplveTRrRg7gcy2sGT/xUEDlYXVngrrwJ3r23h7PVMYW/qr8pfJp
u+tDutuVp/h9v2ajdiGkNXCQ1vuWBbCjdxfdF7I/KW3zN2e7dnDM9r+zQhtd9vhkaszDtP+5gUvY
uHaTaNirXVojViMSMmv/H0lf0iDUgk9qXJYLwpGrqIxrNNvJR5nWndoRjKtWn/R7AWUb+c5QDvbH
9/ae7sL68grsO8HOt7/r606nnWQXFNVpHguOXxd6pt8j7qsSR3qR/V++i2kRcDL08QKyTTYicALE
KVZ9Il9YbedaX4uC7jodFaaPNeaf8vxwjaGgjBv96lBxHPXhxA1fAAMAWLf9O17wLrA9Lj968Coy
xOaw2mIPnyqrSlfvLJEdlny5HczgpKfh9KCQWgHuoLy268ADoqjjbt1l2OoeQEvDp6T+9bJ9apwz
Aj0GlTZ+VJc8nbD0+qYF95TqXcirAfyhsbJMq+cO4o5TO836JSdfXUH8rFc6ernt+51LkIyJyY+V
rjlvL8t/2icHemvJR+VJYBPQsVvhj3qYEIdyK60fpOlCJnrG9kpO5qG6d0alkwRHHEY03aGohvTf
jnpiRfhiFRD8OpHFAdBTF1gG0pDF9ozLy/AyyScLPH3Ha5X5vGX+Ap0rIMRzV6jvNXhPNiGIiFxr
qB/uhQn4DTtKLS4ZOUZCzJVZi8uhatU0Aylx1c0eqGbMFhEI5OHDGyEMPxayY/6eelhsUofOgbmZ
tjBRgCxK2IaqaGlBHfexC8aU7Lv8r8xwgBjTyu6K/YqTSXteu3EwvJgok6YP9dG/bOzGV5Xl5fvI
3Z2yh2WyFSM5fYSpGVNGTmoqk9bdlXX10mg4hqr+gmC3Qo7RW1vYufxUXPaxo3uBmU/n5HzvpXxB
76SWj0c5BZ/svaHtJ7ILrYzgZoSG6wWIm/3OtKcJU+MMAam3Sy1PNS5roGGMOiEmKses74kR5AIu
rWFQuq7GdROZ2VTZ/YNTHFUKqsX/hCepp740o9Uez99Qv6hdB9ywIexIGRSBTUAWpE87EcmebO7D
eH+3rwjm0PgzT6Hqni4wHaoBRMaa2W6xip9RFLmIdRtVWAPCGljkZe55gAkFF1fHyUEKYK1XS16u
UvQ0obcxB07kl9TLMOHIwt2SyQhkHjzQu4LcZahmn6n5ImHyogiGWpijcjGpWbB34yk8eCKI9AUS
Hfo6aG8o/RIRQSfVBRavKWWAaiFfGTfnJA1ADpESNBcHNiI3Ixgxgnprtu16OhSpXL29QUtV9XvB
lFSMhPSI1bUnRHNRPPQlskUc5fYXpFH/po8EnNzTnmehW6MBqthP0b1zo7qeFeCQqNAmkDoykDx3
W2qJMQ5kLNRm9EIh1qwMS3kSDdlBlmOmulyTv+1foJamanDealAcGH43cAvOfgC/4Lg+irA948zZ
UMpxv7Hd13la3Okn88oq0Lff/IqwYpDojD0X9Nu3tl6XGZsyB+rb2o5O+/NH2a4ptSHgu6hz86NI
9YS1H0/tNKOtohsar7uAg3ERB/mVHhphwyjOFbrtUgH/79BcttYMZobhYaN4JfJjQBZNtpQlaX1w
6nbd8W8TWYhC8QxHMtsMChGrNGyKdqT/mRY8JynbeXXxwOPACvxYbLb9S7dOCeUNaInR98rA/8Rh
2qQZcI9k+6ijtIbOPgwmjyickzqzl5oSD7sxNOL8+5RhkNTvViKqCCczAat+4fZLor9Js7WngADX
YCPBwMQThflO9Ts2G+g/fNiop5tFsuvQ+1y8Bjc3x+QkVKKzefcjVjFMqfCo+XvdI80O7XdpJOk/
R1jiocowjS4pmjNAAAWHpZNwEqDoGAj1Cjo31jQI106fL/WqMbQfwdNFKcbR+dZMbvZlwGhVss8y
lLiZtJS89mGicNv7j1xnfOHyGZS/esmf9n/mNkfItG/xDQDaXnJYZdERdsLlq8VR1qrgqL0jICiu
LtQm0ZkdJWwHoI4adzIrpKY4K8zNOTogEnSRaJcA4IIHMkAEJ/EXl0IfxnPBLPNRCQibDYew2/Wm
/0xFP+6N2Pc/tPjK86SVbm/dKj9lKL7ZIQLFDeBJjJ62F3ablM9uUUTs7j0+aYHXQcetwg/RGXxr
ib2Dn2Ik+vHRjfZiI7ap8p7KqimddJtHDOzBHRM6HwoeyVvNukrm2Ph2wK/dtK6BOlpRjhvl6PBn
xciLCOcpSC/D82iyTs5FEfXH/8lZMsbQqmCWYXM5hnYQjEXgGnS0O3onZeCZLHYhxs8UuWoBgkWc
Q+ecDv6tOsfH8l8/mWbCnE107mED+bFU7PSD97GKIODqMhqePJcyimX3/xeXKrZ5Qi93js3ho4n3
Ftno/wkYKP9XXFvvHtXo4NnvwP5KypLSKdMY1CsvNA6ngYRwb4+bGYFlO31ewTdc9tivx+o3QB3r
RukcGo4+w5/L2oW5Qrf53VROJIppZNqs9qKV7kVWZsRF1LvdiPP8gk/ZQdzAHWw5pkUhatoMXrMN
1GsiHRlu/mOahZVTLmYlFXdi7YGn3sl3aZqOFBcBarc1hGenk8jfjaqiubbqJOCJwpdinbwL+Z6B
X4a72aKhxGI3r4KaMHstVJOSPO2Vx7/SBbBWtlo6oh8Bu6zt173QaO2hyL+9JR3q/ObDNORcPRkR
SXbXybHMwN834WTMQC+Bxs2G6EMkerezyrpkQpgAU4xheT5wKA65bkFs7DVKZWlhUVXVwxdnc6KK
LIVbXh0NR/q5gzOtCa3RbmIkeVv9figp8w+8uWtbwe1HBfQNb7pI7eGj3T/n41yaY7MjZkRDtGOd
AUatAA84kxMCiAED81zNls3iYu0ooNlj+kBC4qn3/WQD9G+HAFXGgd/pVNqpGBlwQuWZhJuiVA57
cVl1kUqPdAwbODuMA2M5uhweGAcOKdnslMW7PC9U5kdcGm9dKtrcbaiHjcNVvX95U6dOziWz5KWn
l4SxDAA9/ixGgWeEWMuN2v5eQo+EtWYAN32wSe4hH61VY5T2EREUw77gt1zpa/X5j1+MBsgF3hKk
YmizSzMPYdsDfGEkay3X86+NtyphA/lY86L0rtfCRsF6CIVC6HRBEAfaeQ+LFPlYU0NkKrfN2ZuW
ljEyrH/75yhz6GGrvwvnqBD+j3zAxvPfaFI2/3uFi/jW687My22HW/T5NIGDgajZinfrpkdFuiNq
MsrwxTO6evUt7+NaE0HP93K0eNF7IaMG6iOPfya9CWLzNIDCyQEOdx+WzsnblDTo3gmtW50t+JlA
4f6AC8oOiJtas1UinamJ2Gi58CL4RLWVYOzIoYg8ugodjxMuRTqI8LhftRIdUe8MqY2j8TRRigzC
pb3ulTDQkIm/yoQ+sH6yMmmkoykZVSC6cZMIL/zS3Gr4lnvXlWa4FNvmSbAd9W6ieKdNC4X7/jEn
g6aWDOBM7XxQ3zXFlY5OMvCFHAKn6m4UMc7aD/ShIatLRYkRRu/vQ5apXKtTbQoh8jVPcUhVwcEQ
i2ZzOyJ6asna8rGJSJoxKjJEE+mWueqI6YxB+DQBAZBwyRqw1SqgVmQ9NFds1sAVx/2L55FkBbPo
Nt+MNfRpcePkKXTIm+aBJPK6xVu7/zlADh8UR13zKKTHV+J3gJd7yC73jbmYtk4ADDhec2n/4jbb
VJ7D8bBzF+YzaDdWaXacNxLK6cPAnyKnEh/qri0yqNRGL7dB9bReYk6GRaXhw0zDutF959JvbvY9
rtEHNl3miwVABczIMDKJWZdzwTMwjxvnt4VzegtVZiLohTOeQBvHYbLKWo71GyS971gYnJ5luAOR
OfmZiyR9PWd2NlZQ0mlzGozUWLO/CX+EOYbRxa4VtC1zTzDPtIQomVjj5xFlPSafEpRWoXPdHx09
cMXDe6uwBQ4FqBhldWcGqDbzazy9qAr7U5Y+ulLd71QbwImW9l9p+h9858lw9tyNGPlVrNwK3a3j
c1EWxKc+o68/cW5nWNPQYp089aXOerToQMzWYQ+p8nXELSGz4ItJixVqkASXJ9PgUWbNsR92MDLi
xcP8TcP6mx5ECFzbRyCcO2EVCrzoHiU+UX0K3elI67KosuPu3iCUXuPaLffKbRaU2MF/1rJpogzc
+IfSo3RLK9k1aMhYVrqx5U+AZSoGk4VFZF5Ed8+WgTiY1RRaVDDuwYQ6FRHFxin1EqltJBxtRteV
Ql1npRWEJ9sOhHvgNTWhllR+8fwjo1mZRh7l5pgSjvAQg9J/cDrXOIf4bjPAEELWnWYZIe2MDyP2
fdOdXWzBjHn8krFpQ5Fc7lU4yZZmsiwsTeZO3EyVseDJLiY3LF/K9IjxiQjjo4hUGaCjmguUIBjm
Kw5Rts+OXqcfDAAMw/DT8i4PMwQ3ketr85+pOQOEB45WeoXKUJi+4C8pMBzSyeJPoY+0UmCDe9f+
oCUXKKg4UhEV+5DYPOp5/0CHs0GvTsCIlcPwDFS19L3nWxGivxgKNavikBj0wHdRDonfPLEWfQiG
AAMJWyR0XVJ1WOZFd9p2yszIVM91wsvtLOB68lg7sYnbNbadQE14ezs59qMWc3Cu39TQBFcKn2BM
U7Ju5xs6C+pIO+2MyoppTmtPS+NTOFJeadDxq94ukBmbvny60S0rFGKFcxjzIndom2WeQaDD6nCZ
59BqlkKZm6meFIfTTz4/imGjsyWN/PagvhfyeuUslZr3BGsgXHrgBqU8BoJzrYXLA4PkJFvB+UnJ
Kc/9n1oOPP+h/msr03ADtMQBswoTeJdXZ1CV/8hf9v0Z/4upTGaLFAgtQecwOVbGPPCNTQLAkqn/
/mQD792MJlJUCYqTVQIDcs/xvjxhg98ReGTcvpjeRw21R1/MHLQBSGDKl3gNeMGOFJ7tLbU62Xqg
K9xqzSjAD0ZbJMC6D1+t906EQNG+zTMoswYAEF/EInjHr3q4MVhvuSLL11HZcJ00FA6kzCjhNbv6
GVw6Tn7cyrkfLE63Pfj2lrzRWXDXm6qW3KKMzAWfzvAPULm1Fu1s4Mg3/L0WUnLrkmNzzS+fygft
wEqHfE8bkxv/vq+haQtJfYTyQsiAnF3xwjgpgRM9Dw3eXFTLhJgYuMZMmL2gEUgM+dFlFcBZEdFx
sPoINDoxjVWDuXefkfKSau/ZyGPGYvYsmmIxlVRWcCcYOQGqjt7Dj4UN0gHZGh+RlUF7PeomuPZF
Pgt5B4xV2ad9zM3Y2KjSx4CnxpJTN6yKppOjcN9Ifj8Mqd4fm3Z+BkDQA86i31ay7P5BWbLaBHyw
SWdzdleLyVSnMltl0TFt/ldNhWkmHsL6zFkVX+GTM+fw2mJQhGloOVv7fAdEJataS35FF5MJ8YU3
wOKPWR2gb22bbJGktat0Hs+RHPdOhVgaenhP1vZr3ZWaJ/xcKxbIiWBUwrX4c71fMcoXGaEWZLW6
84he8JG2eH7fRN30ct2PXnhzcHdZwK8FiO5H7H+JAUJ7yL+8qJroLvgdOEeAbFoVPR6z3EnKXOHi
FSwd0oJPyVDrIBr9DV3CbcDvmcxewSlm3bTFOxCsv/jI6mzZElyuEN2yuag1D57/o+x4v3ZVnEOe
G5PP29HH0Zy/SV/OU/LKKPlr6qwb1nzhISUv53fTtjSV8DTyH1PobaWtbAvr+vdnFqSWtOcSt7bJ
dOpraMLfnSWzP3N7tqyZYJJ04jQYFpOU990G5mIbjpmgokdTprUeabuZR5HgSL0mymIA/qZ/B2vd
+DYf+++M7FVhPBatEsJIYHiPCW5B6vGiykGtmia3eVNks+3AH28IvCeci4Dd4L8TdOE7CwrR5EzA
IsaeQBTYcfnl1ueLekHTJSaPElefPsHD7Ar4DcX4tGnUM/yjCyLR9ICnNxagSoS5fSi5tKP5WtG6
sZRU8q76NAc/sIelS95JJBRN+avUtmdMKXe7D6SxGoBXJ/1mfBoV9wuRxLva97rj0QhjgYrG2kdt
78soCh5MODGYdIw9qBO7G6GdMPXmB2LN14o0UttekbolsWiMqmDugJzZykPgjEz3Yg+1hIxj9XC4
twjgYn484MIP/8L5zEl9HPUmFFxsOSe0V4pwS9FD5e++RDM17LPa8OCAaQWnoub/neCFBRZEaUH2
wgjKOH4KQCNtDKhHMzlVvL/w6wCE+UdMXlMl/lYThSrZXerE2RHvKrFsMEiA4BwthbxSrpES0eyS
+FueD04F9JUNsFJLQz+kNwxrVc0MusMeNEmvtTY5g7Klrcvrsqzpveoq7g3UEZylBs7UDwhp0PHC
zS6/G/DIgFyOf0wGvIQM0xqOU9KG2TFzJsDq09/pVor/fMjrm0QMnLmZlt6Ct+mLxbcnJ4TIJqep
1kybD1w8JszweUhBjaVktm+kon0ZWSMrFmalTmxdZjKaoyDcFBF5A6o79IlHJZEvKxBNaK7iCaxJ
G7UEs0ZsO8m3HlktbX3bMQIGypB68eytfXYt80d/QHPHXSov9RBjWYvOPrumfztVSLsUmhk8lyrx
TtijnYIQe+rJ4u5kOL1FuZoV+yzaKUc69sFkVmJT1AI0LPCFamFkqXnp9EAM9IDHFFLV3gLRxfdA
bezLm34+Ed6LD8lp8ws0NqGe5Bdi480t0WBVOrbwCm4AOIOi3gy9QjnZsiB2eHbF/AbIBk9EmZgp
KDO72H71sse8qamf8YI0IT27qOu3Qce/8IbEL/J5ILrX+J4iQ0j1k7FR+mRx0vwcd+mwSUy8OCdN
aA15JTZGdPNbYCuFKcBD1ImxxK0tHjEHD94HlrzGqfW/3daWHEjnOAHhEeJLTJFEXDh8UxVZ2uAK
xnK7I0SBSUt2YLaX1PhPBBqz1uMCKBtKMljjIdAgvyElk2Dsn6UYWMuocM9b1gK7qolWvdJZjmrh
h8E9bnOnhkg3jWH3jnmLp7kkFo5GP2M81W435oeuxJN/HT0xTsUz/evN7e1IfuPT3hRubZe95UwS
se9HmI1q47s5n/jZzbjVpXkwb6LOtP0r0MtrCKAgAmYCa0azHFIbqwhAmdYlTH8IBR70DXLCYWpQ
aAqyhmUQ2GGK4ZjU5ovUNZOtsNLJ5kXeLXIHmVc72nJBcNL0wUEGUJlzJu7UhNhPOCOPx/hU9UAi
gDqK+KkCSYPf9Pw2am5zkhcliYwCuqk51uYDBnFxk8YiATEet1S4+VVrjKAFSDZtSHUQG8MomRrP
3kKMeWS99kCcC+SgV/aW5WB/Ek/oVrzqqWGjgupYxar/fBtVbEcrXE+V1MpOTXHfjhd0B+lQttXH
1kLggx2QjubbqJbDMalovtLoDkT2wXQCVP9NF55gHIbg2zHm+uxSd1nceUhezlJXgw2G7t8kP0AS
Lpu/yOnyX26oiyVOOrwrBoPfGKmKyruHCJ3SNDJafaUkZUroKciko9b7Obn/L95CIVRo0ssniObk
kauY2dYC58Ra8BP+ekjPAERcg6gbQh4urYFwv95uUjsrPjk3JdUDQYLtO7s0mK74CfDdQkgGuljD
umKjteuof45ZEVtipqcSJZNATg2nLDHsRT+/gMftQt4pvO+MRioPRkcB1whuHW+GLXgLazQOhUfq
ExpQnWGgKgvsd/0l0L0Rc4Gl3ymCsUV6eNT3Tnw5ywQKTfyQO8wCoZDzwObA68JF2oT2Mv/w6EVW
+2Z44fyKeaDw5O2wULugK8Mfy7zNKqRlUI+5axCWpQpampzn3cks9UD7xvODJvGK7JWwJ+mFbNAJ
2eLX+o0xBuF+jzoox+A/KGuD0uyFn7ABoUVCVK6GJcJ8alAjrYD7vrJg9EnMaOn1UY0nzkctdt9K
8uwSijZU7ht8i2YnTTqufhLqM7GVzsrrVsQZaFpmAZpzkYMHR5QEZQc2v0vyH6TbBOWfYTXVosR3
I5G+H2aIt13XbwGqLBnE8lTYTVtz01iIqIsBo2D0aPwlg+71FrTa1AMG2uVpGlG7GMYUfY5uAU2h
WF1+8YXxDK6TQgMibGGqMmN/oYOcr0gCrKe87Jc4ROxisR+G8RCGp3xby/EOCnQgpaK+8uEkKn0O
ZIdOeVzncL8bVXNqdg7Vak7iSbHV9ma7L2TgJuyj01uCbYij4aSz5R7TD662YuBwVSFxIfV+iAI9
D7fNLT2ZAfU0cJccmyNCKJuDTTta6wwkTsz0ZYsbGI0x4pn9Xv9dGxjv7QA221Z20jRObJHTlFZ9
SZQNOxqs5OeEMpDsri6dtvXpcGSenDrRSVYimFjbcZThBDmNysXYxrgLTMPejMuQbPDrHM+E7wG+
SBBFgtsop0pX3WOeIUyrztP9sMWBrrV9Rf+4JIxMpHhlIbK6j+mBd4bKLfaVNZCR0U2BBp0Wf3jW
VBGxM6rrvFInkPDBl+TkmNnod3w+fiZ0iScERF35UmyfKhXmUbDyYhxkVSD1YANOwN0a6/K8sPHp
uiK897OQ93ot9XJsq0gY8GOprD65Kw0wb9md3hSlrqaywmnKUmhaQZZRoNAgTIRsTJNNxlciB77b
QvPWxhCbAqCYj6gZoTf1SMBmGsQVWxjewxAT8GvAAF7PVdK5IqtMumk6mxn8QEcGPh06BIw4sUo1
pwy1RpVhEzLGMJZP92TnN2pkSA9r86LGZQ1aStgAfRR5yy0bnVGQCpU7lThnU0QdBoS6dvGwK3v4
N1SnNXBYq4xYsBqBSET+TOsKBgwto+EQXtwXYU4uHLC6kI8hQaKU9sNDs+59BD27ib0DrzK73Fd+
Mvg1RtOYvknhXQ6+wwlcDwx5f/66+F+rqOeVxuafg6NFBMjoWEeYHGBwGJYCyn7bXlWb2oEFGK2U
L7JXXXdY3DQ4pWtvgHis5NMaE7iVE3QyVdEG+QXU3EeYtHKAqPxe3/CuC6pFPAAgWPbpcS1Bl+kN
P3zJIB8nJZv80maFsRrKiF0wpgj+C/Z/AW+eaPzTjgyi7IADkMs0VoKy5BBJB5LIzd2yOCZK6k8+
2Zj7NjO9XR5G6TIymmC9JHxbcoNjNyHtNPz6mVUeuCFm7pS5DRW4/PzsYJ7XSW2rl6FKag/aafl1
+uXxYqLrFoX9oALfKCbvQb8/2T/Ip6/5C+OKkDeXMke3frGJepXfmajb48OwngW44Ppuk2Pae6Vs
bkUUOMQpyTVXz0y9+TO+5pqSQgghq+cl3oefrFehSrYVOCpO+gY+/OxVnpQaer8OoSsbuS92RYsw
1Rsav7G7UCHYYJuKnHgScvPow8tYJjy3UQlD0oenTcfIPDP9LcsfJtDyBZEFVQZDQANtsHv2hq/A
3a4nMrvGyXuTOoZPDHzC5E3PQbiKdT4LqqfcjX1J/yMvYP/2YtNcDciGSdCN3OTGxKQwG9pfWskL
TpNQC4XQBSbmZjRNKrweDoLR+nOb6j/pRh1zzIG2fuP6K5cWg6ZQBC3c63sNaFQd5uqMsXxO1Faw
V9QPVdcFtVq8MX9T6VVmbfwed0ROV6LYa+XPqvG0aWoAK2nnDrAkpJMbM2Hicd5jCqjpB6te+/ub
tl5nR7h+k+2uO2z297HIL/oFDBvdITxq8dgPbDFGIzCXp20wIKpqthB/+aA078q+yB7XcJDRoijd
+N8iF/YW0PV6V5Drvg+Mqf660euLChAxD33ujkFCgN5HKbrkNOeVxL26pQf55VMf8zlEdJ53u0OC
vmaBXWSMiIFElAD8NAUnjJgAxjHM2ZygaqzPgcXcDouaUoR7f+aizaJpMNW60nY5WpgSjJoFwW0s
XVUy1eFCpapjMZoxg1xWs1pCVICzto7RZSpqs7V6FSi08RyJOTrlJDlE+K6iUuMVLalS17GXEf7w
sFmzygC7TxGEO/34fMUdYU8uF/Pwm4y0VV8XY10w/AWxMVjSVFmFlIX7aglFmHk+Wk/i53VYJ9Eq
ndXK34YyIWfgeTK2r/zT5y8Xg4DLNleZXq39f3B8b4NW9CPM5FBJIojpq3hw0RTx75nW+j5KBDtr
eCMph3ghOTaHKEvDjbBuimDBc3e5pGN/GYQR449h+JAFlVnLVoXxvHE0bzFqNoTK/3UungcfBeM5
TA8XXTeEM5CGQtoTJIK/Ax1gvx6FEsCMy2+xKNZK0q+Ph6+jfAy2JPwFxJhjDpSfypwtRJes1u5X
ZR+t0+DVC0lTpj3zY8SgT51t9tlbVyZnvLCJzN556toW08ST35gU/Zo/S0Q8ndEx/6/2zadUxz/9
u2nUeZKDZCazPSqVrDwnX8vKH6rfTwdKnddAIT5izs8Ia7ezNOaItLIEUOERKkEBnFzgxDnwwLZu
9flaM0qHmlNrS1VHGZKJ1YPOxZOeOducqMcSjSSkksZxMxUfTCeQKKjcnoZc/ZtAYktl0q47Xqzb
yFQNSfEtHWt6OjYsX0CX2BkjTgjsvrib6F2GtLDH7K8+w2iGYWs7qh16YIgV9sCarOQ6TNXLvOQY
nYJTWos1D1bvjVpZeHRevHu+54kur0tSeL7tlNdidg2SaHwwHU/jGjoJW3hgACRC8a0+GvuCVbqB
d9d3OGq+5Tky596EvnzSLBFn7ng4HTMeg1GwariaPCw1vSHUD7uxlPo0BH3GzcTnLPZOzvk/D3Ku
7mGb7NagjofYkkkWeuHUpVEyPsreCdEYhFQVTy7qfhXRPdSfDC9X/cT8mRAHvktrjNWTpHranvyr
xVecFMP5GWCItNR1HrnCKbk6mDqk52TErAvumLP5xJFsGZQf/6StgT6ST20vAUBq9YC7qGdGujkY
EU0V0OPJ4TIkaWBuroS+ZrsjDuNXmN84r/Z+bFFOq6pVWv1KyiKyxxPg+RmMiTJ+veC5W279U0v8
sr80AKnIvjeDhkrjA4kdaQeSOF+pspHpNbTyoj4cMcRTZl1IutIKkjC0vOFqtsm/uuQqf6vvIdM+
CU3wPeyC2vnbknSwuj4Q+A8CUtlQ7ozXZk9Y7hzNma/h19hwaPQdH5rZqvO0844uJM45yRB+A0gK
FgCxINJa0UAyrbXtjF47/w3jg5VM/gnaHscSQdPJrJ+EvwZHefOCRydS6wsDeuOl5Ln5iu7mQG+F
7KOhpKSD0yevtjwYSJCQmRcHLHgg2ooZCDy1Cgcgy84vItYSfvm9q/DXJF2bGRWs3NocNp6GCzYX
X6Qom6zu7VBwQJuDb2PDx6GLg3hHgP7mkju5+PFV6hgi6Z+uGMER+5stlRhl8NVzf0wDM/BGCpXa
KOK5GvFEU36k0snaVWREE/PC5nE34qvy5asBY5AMKXJ43KuEkc6fo7FpUHX+B6Hw/gzZa49QBhJ0
giUlDsrSRa+YMGqSMAI6Tnz6E+M3e4EodziNq7GLpH3NHzZvSEl9sB0Xgzp3cr1j6PnHBXFT5/z7
Sa4E8rGviyYAMZKKnruAaHa+FrVBRpXw5Vr5EgKP8SDBNPspFdbMIoRNBVZ5f/XSpxO7NdwvtMFg
rv1NFneNkhYIw4/W1i4YhTOPnHPFNlOHBm2yCHjZMUevuT4l1pol6fnOId4A92L4PeCnFPngYMfS
X+8GAmWon9jXihZnaWhwb6DYHoeQ1pElj/JL0nem+2YWgLVYb8D7RLlsxQUCXN/jZbmu2c6LpAbL
A/rYJ0wkuFMhXuhovfEgaW++bKDgPrcX1XqAtot8EdrDGi6TkbmX9Rg3A6D/Cuu8IUCq5Dr4o9Vy
4nrZF7W4tDxn9TjuL6HCSHQ74flHSh4hyg1qj+KNZFMtPmOpwLhLN1RF7O6TwmEoxgah5V1L4zhB
t/BA5xjobkpo13c4876LH6LvsE2ragz73x3cTDqNypbzmKIjAKkgTJf4rzDBYJ9FFmDMG5XVY2ay
O/ayU8kyoDL/QchKq/zFEX7P6JOMbPIOpHjyZoNQNcRiUVwEHzI5VUsAWg7bq2tkuRx5rGCrCW3B
sKObLa9gCkWNsdUkWk6JwqcAR8q6+KEajnCGtXhKolMOQctSWADc8N836yeY7p1jeRLCc8nIH1YH
QDduhm7jGtNpl3Xt0BqvE8q70dNuXkXL9Bgkxb5BOrIHtoVtsYC70Yr1rijPnRrM1XXD4roNcycO
uBlUaX38HlWNlBlwojH1zLcVTTPgmKXQBCJd28wQKA703aMbmhDXvtvyFjL0TUnoiEAeiKsQ1d53
4CTm0qkqWnD7L1vx8zUmHfj+zTpLuBUJRQTtSFjawvEn6jtFoDMaLqzs6jPO2EHzIb2cIivFIeAL
XK5tYlH3RK7tDpvAVFNg5mrGMc4avGrpd5+e2R2XDptTP3cTqgXAduHhWVTUImPKKCLGlyJNMQAc
+3WEI0bJ5KaU0gsGFp2UZf23v7LDFQc0pepMeNImFVvFBA8KtmkEdOyTP4d+zRqkvvsTol6LN0WR
4K0K43ewczREfS69e9LD8VQgsiJ4AyO6DJDMV+suT/72G4fOwSyDP3pvgUwEUqYLt/8HJGkexMSa
MMdKzHR73GbT/diuirntuthMcUux6EodXiAJ1L9zwQEsBGtXMC6iXbJi4H1olNkCZJY3o4DLTyXF
Wts2Q3jEkkjTp7cJRMKTDxYhxCrUZeTyLUtShJjgxOGpdH0Ko3aLLHHrHfnjFBSOm9berM/1G5Bv
d8+wrarM2mcdSa7fzkBGRw20ZtrP3tp8+yOOvEL6k+2Y8hMCXcT40RBnsDg5x1IBAnqOtx2mmSlB
i9QaVRy72v9lgLJmbfdF7e8+bpKxOzuKe0zr+GFRUTPtE40mmYsT7Pndt6DC+rQA7DYkb+sq5aDm
8HFihbdwC0TvtwGXQCEXw0GOoFw1w8ysgm9C8lNaQUaBAtiyAdyw+Ik0iCCzgJrUyyC9w9/3/3L5
phs3j1j3vc++xSYiZpkSS8LG1u1teXPs65hVlUg50xd/6UH1WUgYKgyiZocouP5NNh1pBuoxcsUs
qllGTkmroLY2v7psZ5au6bQImprFeoK7RNsxbkc3tTbC80cIhSF6CwffgWrQmeWHaMbtOIwNDex3
cEZngQbQiq35TOiHEdIjSLdLiOFL9gnu3hNxmXxhk7bIImOPJ951eNLpZoompbNzeuEUqh7ear1y
Ho/T2NymH6t8Fu9K04zZLb+vPb4GjBT1UdJYlUSiFecT1uB7RTfrISO4e39TlywsrsTU5h1L4zbJ
/bHauUyg8L0Di4OHKekOnKn32lIGe2vM/22xjJzIUtF9AURG4iynKsUzZSU1m18qZ9+sGAYKfrWf
oaDLpqdnY+o6xg49w4t2IjrW3h6ZcIEo32qy1nLRkUR+QmtMP2i4Qx7I0raPOtVRQQU8YNc/QqwF
HtpTg6+IK3B9tOimQdrk6R0qJTGyh4Y2GFIbI0FuVEwTmib4qfDwwz9BZpEpUMSd53DHxwtmUHNk
x0mjqlRU32oV4MlSYxCJLOs1j3N8/KlpCQsc2+hipm1z0KkZduBG//ActXp/C1AfYmsiCghFHq2L
SlWAX3mEwDdZAQPGDwJ/0opJ3nFoB5VEwPMbtwLgvfs0PmgBz2MyMn833KYDcaGIGujBRP1Mj1Iz
hSlTHjMYiJqwT1wAb9Lq7whs4UcIJC/OhVQSceUsfiwrZLr1rv3i6xMwRmplkiamOvvfE8Yc9VeY
2WsGi/RwWPoBIA5psfuOgv2FUIiED3OKk8I2pgX4dOgYsPhhHMmVDwaEaDO3ZsrwKdb9jrKuqhE8
9Ksv2b1zRh+b7VGYXtiAbsMb9NEUwUxMy2VfUrIf1ROQFITwfbOxHAn2n7349DNtlASTx8v69o3B
JwOzbkTx916o2FyabJoVQRlk+/i18I3x3Qdkr4Fk85ck0JKI+geooTP8JWSHi3EUIkbW1pb1dHwu
Zri9iRPdfhCTtB1uhSpcb8vxm6Dh986EkybsxufHbLN7PdptgVHro0ckkbwjVGsYOI6dYwwhgQF3
/NH3rdda2OE4z9nYsjTDQfkOd8em3aje5p90YN5xi3V/mBZ98lAnghjaLhPt2m+2Bl148xEEbBRj
BX1Eykeq9tT1OJD+JUt+SpOqU+BKUuk8KVj6omTXEqHHBKY1cm7O2STzqPjqq7FcFoFf7RpTF3m0
iTxGNR8YtLWN7emtRL7LPEJtZyK1PdsQuvb5k54ZWgklYiIJQu1dcv9cq7K3mqKyF7IkSO2YGLoe
NMm3lI0q9McW3BZRcJeUar5aLVzODLMk3ih9cD8rRIrl3xR+weU10PHAxEv+OpSjza7Tbe6v8jV7
w6W3iaTmNA0S+SD64Cy7PphSU8nWYVxaynal6opT3T4eyb5Bi7PitUyh4GYTXfxK+P1NiPTvbAEN
OjyPdi7ZfBMB4FF7Jx7lW3nqGfXg6ILneN8Zp/1xRhs5V1xxjFOG+3nkfmDrsxqDjxMsuMXQBkr6
C3y4MhvMN8huLfavl+Cvj5iJlv7nbFhlntjlvBnvbf6vcMhnrkMR5RKI6GqGnnY5oXfYDm0yPZlN
YBdYVEyrOhWg7m4q+Bf4FzoEG0PNGxjPVQdbQO76l4sEX0x4q3OkCjBES6L94DAjfpMgD67r97i1
9VR8iV64Q9QJAm9X1tgrfKfsn9pSsDnScko7KNuld8L2WBJwsRqYaHC1R1HcedqLVd6k9BILc3kY
2h5vQBI9rrzTtF0G4ZGEbTqzz4yn2dPiP+dNUne4PB04VUNMhJlI5QhYu2Ebo3cx7+y6YjZSrDFr
eKRv/F+fkckSNRC9AhgKcldcvs2XJIttuHjlsN+5i6PPWEZEG233zg51jnyPZW2i/ugASXaFKHFI
3wcxZaNDuBeJHz5htixuZO+zBOpSuFsJ+ns8xTVo/P4a7DsRyxdd23sCAlC3bmyJV++VhgH3mc5U
12Mwk1uZ7D4GiPGM6Z9zcdG6aDiui+/10nSCSnmI4lMRSEualemruAFDQ1W0bp5d8Moi5TKiwT3Z
BFrenkr+JIw/pZu2R5RCLwicfzd7KoCO4APRM5nF5KGDDqbtKK6wQ2YV6yDsh7Uze9uzShcibicM
Aqr6L8JsTViL+1axPq0d363JYnADpY+zHB+MZf1atS1B+j8VCTD96R1BoigCy2JVtyZY95c3gMlN
c8FzpS4pByYb7+rRwdKxgteyvbOHHmBGh7lXCr+9n6VWz4qnfyIaehSxOeG9ArKf4PknnD0L+jV6
+nUR78n1MQ82xdknsFO2suADhAGXkM3Yd6qtaRHn7GJiQyRPJjnX2qMuHpnIwRYksIH0PisFbmEx
gQL9k9leaSbRPgf7eKWon3wr7WFO8OyrlHu/pxXbsBvPXzOTZhj8EapR0X5NV1ETjESlUZqfR2Bh
sXuBhsoeo2R8qOl4G4ZB4jOuq1NnNH9aKAXebDHFxmIqK/oNTnEYBvMMpkrtW6oFqFYViCV9Kx0k
IVxIn9rwidrURKv0Rb9nZfAg5kwgU3jnAFrDi1+ICckTdz10inqDCJxL/uNqUm2Nq5+FztSSHyAm
4sClJ4Znj/hLz5Hju6mD3lGdzWrpjilKCdGWtLt95bgVU/4WRWB2CWCTPnet8ptFeHM2/2nJnY13
Ze1MPVHIlpsrt4VRVQ8FVsgFjxJNq8K1CxT7t0DuPXrU/zv3nb0iNJv+UMFVbMoy7gGiqKkDRcxG
qX13a+KLvgBV9poTtsN5XKK65EwkHtxefvcdxwwATMbxaPHC4LVBmvM7bAX9GCmsaBmOPL6/Lo3Q
ES3lVHsM/ocpd9yo/RO4hrnwDloZW9COOeiD6B7w2XHppHvRZNduZTG2O06bjFcFb7Y7WNI37e9m
DrxJ3deMMSPI4smJXI9/gSA2Kkhh5AwXYdG+2fUNCz+NgsrVIoFhB3Q1Po3f6W7Ocz+Icpzd7NO2
TpKsGRUFO5szo5ugtcZUX6SCoBD2y8AICkrNU4e1g+5QfTGUXdhC3GCacN9PJ/5GAgZMP0HVfJjT
p35G6q7hLfkxqzFdsVbxUYyyepOCgUjTckg0fGAM0uXt+doBrSvlFE3fHIllifgDI2SOS7BwbEi3
sEksl6IW4eWI7aeruWrDykA5ebzvAJ/8I9KfHJ35uznaYmglX0qZKQapZg42RvR3WanXO82LuryZ
7f9DVJWSnAsyDZg58hueGm0ztIugYZoOA5oreYHF7hzuPNEK4J4uGJ32YB4SSVebp4Kr8Je99UlC
VnXtg8QpBIdOCBCYQ+UwTwMACSAjIq8PxOlqrORt1Eb+bOBFzlLrmY+VtS2aNwYDSftiCadDS64j
COrZVKv9011fAidxHKnd2zhYmj9w6DlQgHlfv9F8dyGjdw05/zDd1YsrgCcT4yUEQGUdQ17V7IxK
Bv0VKVOr06zV2bmdlfqtkAZLM9VqnPGqfOkLjFeyw5r73BwutnU/dktlk7YFDqJTFS14L5lt0cWl
irmIH42tvD6fJ0OyqSrM3Kh73K5A5YPDUpv+rsT3L9nJ7lSmt/GGNQprZu5WFDPvXpUnsDY1e49O
98VIZbk1WewlgqQYsKTHvgqshf0BLNloc2quj7DA9RxmjwFBdn2ktCPIZMObwxkbH4rRu7lr0zmL
gxUXsacxzGrxNbQILJWZO1UAEtt2nMl+k0XGk3xGt7Bz0CBNxBxsezgbPAj+CyP0nPEi5MxTXiPG
j4JVXY/+mtFcyp59I5Mcjb/Zzo97HS5t+56XUh+hV9oFmI6WPQEj0Q+4krxBtOWptenCpEFnD0Sv
wBmwVnkFh4XOemzJaPIUn5sjmHhzb/fB1L4ZwFbd99AjmQkTSWP3B2a39qqADCs9JNn2fqt5nhWj
3jIs1JQSOh7zxqTUVDT4ql4u6vIHcvM4add3YXpAgFBBKozPdEopaB6Yb3m82lHHrJ51WRt27NLD
1pxOFQG3CGRS8y55FxG2gTN8q8/AV6uNM5tgmuGJ0e2OFPw73vw5NkYDzM68legtTZJt+zG1ku32
fDCHWElmLFM0+rv+WUo4jIdPheAkErO94F5zkWzSpQmPxlcqtyZaWd17I1PE/kGTcUZVRimSzIRW
2m3rFGHm6/UFe+z5USpbCppla/eQjGPcTLxxNpJCxzwwAA+fVzuHeVGJ7ly2qB66QPEouRrEAH1t
BZAB24+06fG7UU9ZeUfJ50O1P9pBiBAzwcRLwuod4ENUuRyNREXjRQDT0V1ub1XXUbAflQceNlCI
80CIhctjShWBDdFkZqeY9f41y4n1MyGK6i9ItMLUzT/wwD1H+eNngO5vLzRgP1oUYhQx6ZC+nRb/
ddvkCHgSTt4ouJhzKPcea0Zi9kBLwyiL6MgvLFljc6NuG8WMm9ncykVUghz0Pvepze5NkYC7b7Ng
s9qKAeGGZWbXJS8U/T8A4U86E+f5wiWhcir9KpTTM5bRBwd2082XHkBW4OjF47NfOFZwWWpMhPuh
r7l3J4JK0clj9UmU23YZOTR/3NUE0wiqv50bnY/qNZY+NwuN5jkR8JLS7EV8sG2zjvoTLeK9+z/U
Io1Vo0VjClJHUl+9fD7MU3HQY/qjsNOgV0GcVuUUKBbf0H6Sodr4j9YzYy1HOVZ3/aMet78IeXjl
/Lq2SDxhw+hPBzgW4K5q02P7ZGqCn15lOx2QZKzMseRcOcckowo/5Ukn+1ppMYObo5F2JTqU+hCq
4wQAFVF+RuXNSl6VkJaauN/RHNH2QjC0L3N2hHhNboN11aryGCAtsS2IF/u2n4iSzTkVqD9seLFO
0iVmYN7qeoQ7T+ucr3LxFBaic2EHUpCGp3RMtvp4VVjAf8QtHqeo9TrpokIDxvRUPqtBvii9toRz
+RBxxGi6ajmwZcUA9JGyEf1VoGrHgmcWejbnWTJptu4P1c6y9p1qgc/fggpR6Vu2R79EIDcQl5L3
dshUw2NzSKKOOGW0qOHx/XOh5iK2ZxGCx1TqiXxBJ52oipK4jStCj4Zd2TXtm2RwD4j2d4W9+XzF
NyUJ5CfefibD/bujNr2t/H0leZQNhN2vk9+qaJY0Dnn+ivs+VtQAujKUlKq4d8GF+wbzo5KACXyD
BPztAde/Z7mJBi7JPpfDj+g0K/m+/k8Bba5+ylCZmD3vjG0wd6tVehR8smnr8MiKtdFLHDWfZo6a
zZ92oaJ81Zo3B8kodvoAaVb8toZ2auL8+LQh7h1b0vPtwVZrxLBCw4WJHDYFmVN6cN2RDamnRZRn
3pT3d9Yp9iKKf4EzEPvIUCJyezbQdlY1PFFMlN1wBCIClaPkGC5I58bWFjwDlbQAJj7T1k+UVAa9
iY12c7LLGaUiXeEI40aAdTeLc82pQ6+ajD+TCumDzOcWgX0cm5NRjHrRZjkKnw3SDCUty6grDxsF
v63ypu8y6lw7/mPj0vA3hRG5YI7KL79WGTaL/51rOWRQrcpiHsqXDjVTDmYefiACeaQI0p70UzU+
ZBto8ECUxY5Uk1RLulbSLaQvtVgMj4Tkvf+VFvJda6qHGVXToEYSyKAH6bZQEp/zb7hv/U5IjflY
wUjU0OoAGIxA92RhZRWGOS5NucWEaUv7+o/T49854Nr+QBsjPU8NCFyg1GfdmkfZFBRcHRWKspEE
GDV0S1IRdky+QSKJg2LKZvfJYs9TKfD9oKm4fVqN7koWX+CzlOb3Md6ZTkvE+UpB7LaoL5CRa7sL
HgaNY4mJzhZJcgWREA32dak+DSb3AgdMWFwz2H7v87IsbFKmZAF1+9pbTKy0DruXuskIKqzfBpSy
LatdKLOy1lAHiIbZfz7S/YWbGuqyNk21fVEcRmdBrsPeFGSUg5oVp9QMar6Etqi6mbtSLzHIgu8Z
wWboy7FkTw5aVC8ASlGTB9nLXVSbsLQ3/zsVRFffJLzUTKeYUtH36C+Wkmk/+DLgmZo8uR8KVNaS
6hNpeCF7lcxwPBjH1dO+Kzvw2RIdAUW1w0nWCfkjCjj4zIe5V1yTJaA7lMlBA9NTqCwY9C4J6yFR
CGISlCI3rkVPnirPE1StrnvYDDlDO7APN2z2sOx9ZOjO+yALxgIS0N3aXnUDmbjpa5f38kaHVu85
J/1JRQDQWciX0JULVTPIEsB+RmTKF+mNrm4bWaqs+iKUCpVEv47+zs6ASiWdleOSWWQoZ2/j/s9e
wzR3po4eC445+hPge7jtnH7F1BaJVTE5F5W9pi4haOf/uC1qPZtvxb3edKLAOUvNXycL8zU5n7UR
XxvzFIzuJrKk6f7bGKjeCAuXHtryd5Yh7CJmnQNYeS9vj1k/DwTRRhnqB/TzJ6kv4lBCV+WaSJHq
QWOdwTGWGie8akMfpDakA1ptR97uGNlwN4I0ZS/A7K/J+ZKaHavDdFlzJ+n2x83eVAtTl5WZ8eQC
vMuYlDl3c3tSJF8ollfhoN/B0bwGX2lHRWOpLSUtPFqXTNrLYkzOrSkpGNvkyjZG2AUYRqTi+sDg
dWCYaP6Y8il0wLq3k6VY2ab5v/+IYC6XHrljKX+nWr7UYx+9uAnTM7MLV9lMqTIu4h6j6PZdQ/E+
09J9F6rtfMvH+fzuoDsWj1NUYmz/eyQszFTUoHMb2qyxdrez1bMLfbvtw3INsZEV+NFgyxEm42qj
8xGlWkqKKN+6W1yriskhTy11ubJmIX6QDzJPmvZfEnZ2T9zy7sS4EoJKWVc7qG/n5s3DzIf2SIA7
9PjA8joSxzBcvINwTh+tbpChCmi2VljafTvMTldSSwYbQ7nlZJIkKiwuwVZTOEXZ+g/6GBmr55+Z
Gt8taqox/Je2HFkpqGWR9OEvQKPPDkMQpwVhraswgojU6NwWm6H3MyQSjHmMi6yMun2NUFVyJ9+A
oo+LzqEevc8b6pCGtsxaKLbOGzbAZR7GboLDfTuazZzLzcejwf7Qf/E9V834b8rE93W/lmOMixh7
Yea8ZsA3OLPiI5yL2cZAkEb6KDGpOBNoBesKFbhWeKtieSJL93XlLep6UU3Ee+ogLqL1GduOgynu
D3p2sIPehzbxHShi2vWfaV7yfi0BDAIo0pIR1FgfzoI0/a7hhL5tDIeoV03bvNqc6wHDIkftTr09
tJXhFsUKy/lEuMvuEYdjpPQYu2mSGL3e+jZWkIArTtxRTcGdQM/RgIiO21k7OwUhwqIPJnIP/9Nm
uj5bfVoEQ8f+9D8grzhj9cg9v5IAbN53q0jpGmAH0IzgUaiSB9TqqPc/HrgbtiApfMCW/aAs/0If
YlW0RED7VkxQNSNsIv4fZo+plXeLvV2gSYsEfjzJujhw6rc4Dh3g5gnkZZdCHjfhFWdt04k1T7dA
k+NlQ/VWeY01EIZZMt3e6w3Q5ZueovzIaAeIY96BFJWPhABMv8H3Pj7LNUDcqxDg1LhajdUk9Z/M
VarArxj7J4R8FgJWaKbXly9zNTgUJkFd6mX+GtakpiinvRUwfWTen2qBfYc5gM9tMW8m5x3int7Q
7rjpc8y+NhW7aHm9ACTSOgCpBREhV/ZFUXNpZg93TFx99QkB6B0zt9GMIlcTvzMwLNxHxo9uPgAy
nqvUeV5U78RprQ+gzrOqhqkqmaBkIkEXRlNmNzhF3is23uh07MWQc07m+ApZ5Y00+l/8ymmnLiTS
LyB0Rquw3DIEm/xxBRkUFYZfrtZScDaWdSqlYJMF8D+qQ8DoO4TOIhKNlHvX3dysKx/fruXRc7qE
NkB9tU6Pif39qYmA58rENspRiApjA34Js7lDaXpu6Xvd+B7IDph8mO0eJ6hhq5NT3kikuDm17Zqr
i8cmDj3Y9mZWVaFpHI10ueP5zJxpR5QwvRbjbFfvLlhfCuiMD7iZd6jw9bebHBA9GudsnfWqs+Eh
u3zmCNOTaVUjpZOxFm4CK6wofhVPudm1vW/QkwyMPlAKdOGc6v/bmoY+Os67x9ANPA6dHr6MY9Q6
o3rB796oKRk8W/qEYuazfqdsjWO3bHlCJp5zrSgfWV3/kvEmObgJEyxklafgZ7cnafFHrZOmGHon
QJ023YwWHlIVcBnQpVhwoYOyy6fZGX30PNejhS2wuqfEy6DWMqCRrvxW35husIfCsEdJtIth5h6U
Y7mDxcALN6wcti1StmCt7fNTrpIWWBG3E6rV4FnaWjPb13mfQzoBy96dItuo47FQUp3FafCXDdRe
co+lIwkQbNpkXm17fqrdzX0Q5cWNAgEe0TmzTkafsYtASbjQmGRLhXDoL+oC5omQd1kCrx5qWljd
tBItJcFQbe+OZU9M918bQnz8d1nhReuO0optWXmEQO9pTfbbKPAfaTpsSNoD0GM8kHTBLPZP6zht
JC9KDjtT9xJQd6nJspxsdz+FgQnD9KyPXQfc9ktbsD8NS9RLkoFaSU6dba4AUgK2YlO6lWQZ6Uin
mqOT6ZKnAL13HG7RXWKKpZaP0x5rfqVJ9cMzyHp3VxjIzCxsWgidcpc1Xz8Dy5XEx4kKBY3HfmZS
gVyeubjTIs5zV1AxQj7D+voLDfHPY/f1/v/fsaTLwGDi892juLdCgRLLBdpzQ2Kr06GsCs8nHCUh
yWZXp4isc6oZeRM5nZTshgKtZDutHxTsFTOEP/dsCvSnNgp9SZH6RJPUI4vJXecEr3WmAg4xmL49
Xtcs2bveTZk9OZUwSV51XT07hV1pGM2HVcVCUt1GSw81kbgYoS6+TFYjRUjJxs0jAPlX0Z1KDthA
r6krlhEy1u1HiaVCVYejnPto+m5h1XfF9OLsLymy+PdfZfVHmgwQva/yFLCVcPUTqIfv1YQU6wZT
7F7XoEgC13p4A9idO9MJ0u/tY3lF8SVyhbM8cFf+iZX+sloysHv4uZWuBxLFFwY0T/Xw6zxmvh9B
B4YTR8rjUnYONGtKcCHMjvHUeqhAMg+W/ynjKYp/a0b5IKcljH4XVBJ37FlkdmAHvvrTLlr1FjiJ
n0YJCbp6rcFz9Hd4C4w+zzp79tJWXSeBwAhHICOEIL4znPsreHnTGj6ZUwMoiFG1Ddk32IkQdCyS
b7wWT8LcMNVEGIJ5qdrZ/s/8oCjsRruFf4pjGIdEecUGXa1lQ7rNBl46nr1UWMhXxpzJNUgcd9p6
imcInxikYvqKLchpAkBgHADlGNOzFaFvhh1XrUWuy2iWoIuOYjLt40Vx2GXWJMrnhhzdiFiTlwg0
GSA4wpQoC6tSFfVFx9AjiDrlvjRVU+jezXe+IHkbkpToYHWWkoSAPcLga7Nt7+t187msgPCQtcuh
dLR8heobNGqa7Hrt665drjHinenBf9Ea3Z8wBvNiyYydFfeBF8K7TMb8RCUhMKdtFaRIpY5AqOof
3PDRzT/mm8UwO1pEKL1LojP9DIr9+tUI5KQgx+53MG+S8fcIVsroHm9gshMTws1lmTdQzuZJkK5p
1osb68BWr//29v2NZcMFeimEzMbLtiyFfAHIbZSQl1TxzK6PrHk67pEQ33xZsACYa4qGpUzOykct
AO7i8MBWO473SI0iNkJt/0Q5qNDAc5Vz6lQJIkH72n/TklvYiRxFuM4sO68TI2YJ5A2PlhpHFNa7
+deze0Av01U6OBTnaLB0AmpAttvnU9nbCfJF/sxQpNgFVQG8r+5YrOc0ftX36CfxkbCm2LsIO1Sv
FEeuOat0v+r30p2SZTRL+Z0cXJksJwKAPz2OJ3wtFLj2Yws/7m2aKYWlkQ0QNCYbe6B9vfZJrM+i
BT2um1AVHdWzCp3sgkAqaXH0XPF2HE94CutKWggxOhOJoLrbX6n1Tq7/0ucFugVNV+GmV2h6mwVd
1aZ8kiqRD0TTgINe49GE3ujY7477MjA55EX//oAn2Ns9ExeeR+dso95d9J33bbWgkNZr6MDy/WTF
PSxTrX9m5sEB/WVXVJ028tWkKg9w/HfC3dLeuCzxA8Kz4PkrB2JIJ3lIbwhGYSYUc2yxdWF5/AR6
uglmbFSSD63t3r8JP/lBGpeYJQ/u0Ypn1eL0aNNEjes1qSC7/eCMQdbMCTi+1SD4O28413NoCZxC
Y8HYV+uFMst5ej74D2rq7MhlP850mn/KLsD33uS/x3X8oDKeq2xhm6lh9FmQJUP/NmdMtsBrNNYM
5ZGDxMHJLeXgXMewR4msa5rtllAEQ5tBM5ktwPSQH7NJwIuDCuNukWHR4468UY4A09SIVqpxZB/h
YpufuFsiU8q/dXnxCRPD88pSYMDSMAC063uq1ZaOiV1vgWBTMogajZU8O41ahgY/u1K164r0/DHX
E8bcQkx6EJvy/oE7zhhphgDe5JRTNUNcQVF/qFVmMxybaGPXRWe87kqqLg+YT1ZYpRImYATy9Usi
D7RVQYEL7cUkPJOmwz/dx9mETXfkaJd+ZqYpdwsdQB9VDpXF6pr5AdIm0Fphs+KKGkG8wXnZBX+y
nuKJJKsqgwCE0taAKbeJym2Bjiktc8FNNsyKL9iUer4AfOAMSOzwtke/2XHFIT7g0SckpOx4DH5p
CYLFXl8BjKaH1VMA2aKEUoFug7f1STM6OS718c5ExlE8NNJjkE6HcjqbYtgfy8B4NKGpxrcZGjZp
Zow1gGo0QGcTLqqr5OTyGkKoC2H+JGxzgCMlh/K1O/QofYLyvhWG10J6NoLIPH3Xxgic+bN/WUFR
SE9co9qXHDalXqEYa8QIfaYRqQqGSp2AgRPv81/+Ik1MZIOqxM52q09wk6Z6+sBHR40fED0wCHZe
kXLq0F8evg97vpm6WYaCln0Rsv9HktIFXT8XIkOU2Sp81tzl5GKxjouAvwe0bgnAsWSwAOJPOjlf
vDrq7LEJvRdCPfu+UCcFlabQO01Pv75uMlYVAoAcMlwIRuZdLVzHiOjqgdXoYjS8W1UhSLOzrYyH
K9DxVdYRJ453PxGe3UHUwpRZYW10ZY+ppThJ09CuiM4Vn708H/TVrX+800XDE5HDBhJ5kieAUgnh
3iyzDzpgk0ptKKLYfN8FPQoBYB6lXYjBe0RwXk65JKVX8jqyLMO/WzyRa8gz7xQe2YAPXECDqQH0
rayZu1qOMxtxO9Drue6Fqf58FceFOKL+SksMGO+/afAkcgRdZkifr1eeaOtxB0+T/aO6mskXCDQU
8vnPheDn/5T40B3ZUCnx7ylaaA+ZxvE/+GM6HqenDllt79XPG2y3bqul7Zr/ebGm7aCvQd0jNRVR
71fYxI33rl14L7vTGvOgBtErErKxcYuDWTN2wnpAKUL2FBy8X+HphvAqsUJj6okSAtOQ6fsT06yo
E9IMYUzypfUQ2l9JfaGOIW+amKc8rtIhQi+QmEo2qC8aI5lBXV+IKTgNDKBPqFYv1BCBVpYCN17h
zTOYGNq+emZZ0NiRlKHWZlZQ1v1TsgaMPCN+gFVSSJZMH7jQiFoDnoxV+3QTNTo+y7xlRGCEwpAp
JgyCfvvU6tG4mcNu8HDgaoyKYJgDdpgYZ0jHMu+bv5uvtZ2Wrci0oNN4v8s7GIKDjOkS+Yrx6Sjt
zfhk8XxundrZtu3t5KMZs6EnnkDXd7B/kxEPnK/fDjVxR6TMNBTzSDrSNIG4G5ACQxc8RyBkj0EU
89rYCH0EO6HgF/s/NMWzBrTEP61U2NSv5Ei6gr+zsP7YEXaw1HWhN4sgf5ICNPytMFYgIPl1vRS8
g0KbOewfpyS+uKjg3p29ZmnCh4EQq0RYKLowEoMrZcalVHuWEQCSNACAgyrjV0S/a9jIwSz7GYCl
2ar7hpwEIMDZ0DMgVo1SuXXKZ46TTKvUfGaXmx50dMin4Sa2EQdEuYPHSKdK/4RS0tz6Xyb4NLpj
UTilFWHUlG6ct4OoD3eCF+40+8/nzIm7xsFNSB6tY6B/Bnyiu2wSxa3nRCAmTmE5/XEqB1ffd0QU
lW+3ywBPu12Lf/FckYLyXe8Zr2PLAvtVXUnx7fr8xm9Wl5qlHsbpG787KiuuEzlYBNsV7sSmcKFg
tWXwSJSunLekLzKFU6TPQ35eLyZJGMR04zzGzC/bZ4PUMbmIaT0NQBcZJDJoL7uEOD2wjjqxWwaH
NAQxoUUv4tomBafmP+HQtc8FehZpACN16hBkw29okrwQDQsYqwHCKf+Tc3gs/FdB87XH5Zjicygu
8nIk5gMP9I9FW4LfM64u8luN96Q+M5ES+rUhIFVbQQp5maSfntacpGC4580EYzhTOO3AqiI5y2Vz
x2cbvglgPgiaPQQDDH19QZlmg3WwP64HnuQUQfBPVo6DoQ39WS3GLY6LcQKNnGEJIpQu4n4x1MqR
5w4WnlsAPvVPe+0/tu5O9PbnresWnkk9QpbMb8UXuQwhjJOzgBTde+ummrTlo5DAB/LtUr3laglk
KEwlYD8midMDdPbBkhUc55oxFk8cmJNeRaN4Q+qAPm/3ouTNsgEJ7v4AghINd1xPHMBKPUNktvqZ
wiIOC3XX5Beu9Iupqehyzox6BZOiEgEk8/XxH8PztlbnqTTy3DMtsiLUPJL4nUvgy6Ep7XKCXGub
IBcfKCmk3tYD/hmU9sk5MYS1QjyxOg/uTu5zhSrVKfPPONSw8xJzXlt74EVTFtDd2JQN52GfFC8b
gnHA4WEGzY8Wyf06nJmh2MQYBaf2OWInGoNUYkllLMHHOOYET1iIOi3Q3ZlARohH6JcAcpk8MJWu
9GV7CzT+9mWcAI7Y9CiRmDKmxUJVyashY7q/9id8TIf0JojUhalP5EvrNcK9B6bEL/lDgcyVJF5x
1PuoPEPjUDujcGGWlRokMkhF/9Kz+2BSFxTJnEYGRrxgSGlfp0DhPTIa1ONFpoNnz9hkVlhoqxoC
cIhGXZLXOp7h8QRnmzHpwxgTFPkxqe5lLkAcqwZLImW7OCOCIHOdUmerOitRUkhtVsCjSrAotKkG
x6aCPuFpX0xlbcEubiwn9FtkoWBhdY32uLScqGaG0ookmPWcGMX/1fOSPIEm01S/BH7ejxZNkTD4
hEhF/57sdoupOUhfJfLlvH+IODKsTeEx5VLVg8PhkMxx4KkzwVi6v+YjvQtYUzbNq+G2VusPhK4N
7/201LkQxBZFB7N/SC7VLK18s6GVX8anBPi1b/wJ7tCW0wckqeC6YBiwlZu0fa9zS1712EJtogMu
R1xJLWMTJqbSFsrY3XF5Jw9FJCl4je6RIrU/exuQrtqqMKCyZadDDwhND/JCHrHR/lAee6LVPGHr
RFa0XuoUrTqW+uCDXj54YeH1d+glutIE6J8jfBhUt/+A3gemt46Zot7CfxI7732FHWMVCsBu0+wZ
u0k899Eh9og3FU8L7uXxnQV9zKoPT/oVfSNKNMjuhFVUf0yO/5YcGh8s4FpjP9jIk/ndWX+LLaws
q48RmNNpplFQ2iOSwZeK/exmSbejIduvWbKD11hdNIimYNw0bcBJWhPcR846W+Zj5mFebr5mh9Hg
rE/QGkLyHed0gUp7p6uW9qgE51NlngjTkqM03DiY6FAkKUx7nMT94y4bZe5v0UEVvbebit4xF01U
jHmGrwdc2y8aNNzmZylhWe6wb/jW6A+0qm5GJwP+E9myHu9Vc4GsvMP2FD4IPJlbk57xdnnA8mQo
Tw7RQZpfp5p1JMZPdEdkKDlRbgKvHF4Gf94oHcvlVj9b/UxYc3FEmuOt65HI37G2++L2BRWIMYEd
2Jo6uAx8eaOapYs5XqhLU1lN3n780wmMs2BZ4rt6rUe0Wnfm74sL1d6DIZO9TshQ1YNWLYjp5I4a
qox6UQ5VUKHfmw0L8GvGqg3lSxBKsU1mxdz3tKO3sEwkvl1mWYNOR8aGk9sK5bFgdtbaKtpybqOi
R3p5tutkFupLBDyjRe+PowkF5sCZMm79MOIWiGhm4ej/rb2R1SI4335TI5PqylTN8H7UtB2S9Jso
T6nytepGNdcD2r6hrF2uNLEzD12b0GTo/I+6Cu6TW1gtA+/L1Sus7/N7zWb2CrGBAJT76T0UbwnE
MvtDAkGoyLZnV/w8m+eFuShUMBTtktx6BF3AirE5f+/A3YaLyFL7Yxl6jbZ7BXrxXa5EtqzriJaP
nFflrBzB0riixpVcsFnEQVEBqrl0fSptlmjKTxpO+pTUitjWrVOW3xuqUhtnZSq0Vus6wqRyEArZ
vocEgoucZS5aVrG86GJJb/bDN7nPjsp2Hqb9otA9DLgcVsNibKdXF4tPmqfagTpv1OKVR0hbFS5a
da4H/NXscm0tAqhgRN9GQhToxRf+m/Vd0n9vpMhfO4ABTO8y6+hyNJ7RjEpyDmoE5Lujqcpjx+p9
p7+q0dww/Zt72/kaoHMDcVAf1aO0wDCucmXd6o1kWxq+RgXpcIeNfKdkhKI994D5amxBwnX774jm
hg0MwnF7DbgPIPrNA/dMoRfeKxmXLcCVXtVLF6sKseiCbEflrmTS7x6emRPUGlf10G8HOPrPN6hQ
4dprjGc5mGxt8o045LCGfKVFRdqlb635MyDThu10Q2yILrHcoZFjUosAgj5JIPfq76E5ch02vUnV
9sI/bKBRfHtmCNw9MP3WVqku7PmQvcX6PAlkAl40ojc9gX2EyHsWXmxbAfiabT7mSHbZyWfxZqiB
py8AfZMnAeTX+1hpPNRApasJCTLrwwj6EJPl+6iAtYrRK4+kM8pSZ2hwBY13yw8K8RCyzOAAQLIE
5lf+3XUKi8LvcdZRU/x9x56FXb1MgFPo4H6BO3xgnAUW4QnVZ4+lHV+fyq3VOv3Cf/TzhTeVLA0A
0V9KsliNF2U3axJDGNxM/5JN0/uk4KdlhVKijrSVW3uS3Km3BvKz5ft+fkbGEswTltYUf/5GzJfc
tVM4iyweYwyhttor0kYN+3LV//QuhPvNzQx9S1hldNiihRVf8K9D5vqm9ACvS2dHWCs6qaBtRGUG
uR7xEiDZoABfOhTOt7u6Yj9uwViZOKitsaVEbjeMqS4KpT82Z3/X5Je9SKkjAKNJ5bMK1iRng+JJ
XsthUpzXOdjsSbtMZskqbajoEFJaF4yColai6/7GfV+P4V+T2YKhiKKhYRwInxH9L4GNEVpMwPhr
PX/eNpXGDIcxg6x8S4gPjPWApEsWOq06sKk6Zx1UC22wLAlkAXbUVLcjgC22pulhGgDIkHbwK+AP
w2bo+IqOZ8F6/wy3VTA/QzeUROadAUf9aqqkc1eR0tK31txgGnTZhXRfyNA3e0iso0elCZme68J5
KN3DCy/XeyUikJtbjMOQuTvMFPH2vmsomwpRDMhdbIg+OKyJQmRgayw7iEUHNQjhAcnFeS+MB/q/
Fx4ukIlApQIeT80kXit03z3YbErjscfcZ4P5n3a+JaFXVJw6aFRBHQcGhTNV3HnS0BNZEZscVQ0F
famyWKoG1RCwzAxeNs7eZL+S0E2pNeT4Wsq+0FPK6GLUu8GzC7oQL0FhgPdlGGtJG005IkovU2gn
7/1wUMxNf4QOTlFsVR8RSzLdLLgU4reLKe7vDtbeMh+7l0qcCMKC50gFtPJs6p+p72VAblbadmd5
zbZDYR4OSAINtWS5U8EFPX0XBIZEPUOsMOqMrFxdowSHnKR8s5yDkNA9WIWcfUPsYrc+6G0XXEGw
RDGi0d97if4RdQ3tHRZThcfIKgRHdzuc3EqKGJdTr1L0SBTx68bY36vcqZFwY1fjdr9OHiP8Zl6M
WZA7v9ipKd8Bf9zXgpdY7KLBaue0FvLFWa/ND8uLmv+H10N4Rdopi1TX8haFOhxmddJVZ9LW01aw
+MFqE5FujO7l2T6zXapzeRxitHT/ylHzFRnQ/IjBxnTFnrjemT6ZnJuk7T56EC9kFNC3gXDrK/Lu
4a0OE2+QzjCh62Xdu1/CkzppL1/w/aUMbijDcYFr0hccDUl3/H87rOHxkLx8ME+w5BpmqYglARZL
3G/gwZkTq3JgiA00TQuF0vjOaFDsx2SBo1UbLf0bJb9LS3dLSRoSS3tQC9O7Jqqp8PjabYlFdiJu
zP9Tb/tk6xmW4O4v2oMH/S57MNEhpbrCrCSWJUanHWMwAY2XfsuGAo/n9Uxteb5JgCujJBfDXj/z
wKfyId5v0hfcvpkF35u7NosvAFNi0FUTJH0VOW39ebr4sWzK4QXDq3yPFvdx4U3wnytYmlw9dNnY
4QGZ9iAskzxVt+zV0A+WEjW5EMHEv3Rv/5l+v7k2R2p1bGl4R03VTdcrf99d8ABF/rtAkbhNjT5N
msURof9CmO/dPn6a5gQx2OT7kPyC76TKij/NgL+/Q8ZDPYzNxRtwyPbyvwM0PM9rqqZJuEmZyFHU
fJQCMoBW5C++Od6lPAol4VQqxdQsxriveshUDoBmH7bZbiW/lpDp836kQkopCol7ucpHVbT9f8uM
WgRj/u3EdOoCb8kSvdWp74YoVHvA5TnLySLIUTw3MOdHNf0pB1txXu829j1Z4hrowtNks4xHfPRv
r2Kaa77ZMt3r4dVAErxoBPYVXU8NBhxTvuvUsvQiR1R4GckIXECte1Tjj+m8zO4Ydol6Gd0yOnlk
tiyY9jxMTYcyZC7Mkm8jzG2m2lNmiYwxeGfsV7T0ZpHa8hsbCrtdiVEMawMBm5tWF1xIkoSslPaE
/441ydWB6SaSN532t/cI6lPhUIAMa9l436ZZqkGmu3XDY3qYMduUNciZyqGm0HLJNYlU+3H1PCFf
OMbKx8RFeX4sMbVIQFHxQ2tIHdZSEQwvcChZdTKmxbvX2F9S8aQg/lN9AOWOuQe0dvYEUJNOCqii
r4GjbdcJ6R6CDbBoqU2bK5qNlXK1AADKc1HzUspVJIRBF4Yenlkcqpr4mVRhgpdfjhi18k4uElS9
EFjpas/gborkQdxyhklYUubRbSE0RdFQ07dOKpFiESilpuvamiHIVaAG3c0yCu6L+LW0wWkaPvm2
Sa/5JTpXs6TEw0Fd7hOQGdG981UTXpOqgcIYKG0vdgDSyLvlMr0iEJDnYasmD1xWd2deqdQUWkhO
oGsIpKj3ha7hkmnb9xkr3FDWapEedH/YIQ98Fu2PGc2yMgR+duhCaQRtqrPrZPglq0J1+r+2GGCX
jJNbcJMDY1wYTiROY5SQvogw8pu2yjq1548JhVtbG7q4PU6MnJPVqkVWBn0IwukhKOphyV7iyiP2
viuNeTqdryyamkf+vnM025EY7nHFjv2TQopcvGLThxilux69YcwPkpV3E60yKDqAvFSmi4F3+7mm
kOejE4cKiE3Ao4jc85VCpJZkvVRa4/2zlKpStHOzUcuIsJuV22+n3E3oReHBc4JcwE6cjMEhbHFA
mmDqgyRybwQvLANkk0XB2DuIcT9/PUiKMmLOySrUt7PJEuwgdo6JcHqIeqipkmOZJkh/6tKoDg6O
ImP1mEVl7PrtRHC37ohMm8ppQV3D0M/f52s34HCyzz7fEDqPpVCsEjHxJhlxxSuZaVVlZtK5y88s
itS2YswSMgVbuGdpvhswkrHS97xyQZ+VRadfJ8zOE4iXuLPklhAmVxPc1jC4dHaIF/NzRY8cUIwR
QvDCkVWOHLBqsfzmRl69R6n7YYuiEgv1VzjKhFx0LRWy9S4tG7GockOdg+DEk1IvDy9dXjoC4GGI
1EkroF1JJ6mP0N6pSB+azBlAgOz/HRI3wmVMbD9LHi5KBISOc4B0yqcg/nLyrDd6OYA/PIvMmZiD
SmqDt3pUH3yjj6Qa5pKyzzBS89FFz19Ooas4GO6tfKohLm8JeTQsyCh15k/lTC8fzN9kMwvLlgRM
Un3BT8FbRF7sBR8s2cH839Y/0tx5+rNXWvRIg6W+P8v/K1b0NYGQSogxjnP0lWGwIAF5cKpJZwkP
7KNNPFaKcvCmc/jhaosXwNrQ1rTs9CtQHCvRhC8x9mZLk1shyFZNC8Qb0sQGTZcO1VqgV/ZEvgK0
QUJWzlnnR/s4DeojjC6VvT+U1Y4HmTNrZ6vVumsYNG3OWbytDuAnWwL26st16aleFhCu5vi1u7je
/9lHZid+9kqK9FsMyW969sUEIZRjGP/ATFxIdgwn8Nq+5MbXCggD0ee6TT2ULxSCSLQ3fVn8+gFr
X00mCMC4fUnC4HmiXir9/LwR/ZnZDd5f/ZAxRKT0bbZB/+EMUdvGc1YTojWsYd+kYDZ+fxzhR0yi
9UM27xRQQDZdO+x1JzaB5UG8P8BaSO6OuxE1caD/AuXR5EuyU3/2IvmDHw1ALnzTWIqIP9Tef83H
K0mhBsWfotZgA+TSUNb4vgTfozclq6qv6A9lN1lVb9fFwctzQEzVfQ0F7G0i6k2OENlr9yaNkdH+
j0eBEqAnxxtpNqMKM/1abjr7b6stPnADXRY1uEPrULBTE44y6N6/wbVMxt6VdQme1chC0LgdwrSe
3UlDTDmysp97nSIQutYaQ3DNqCbNMvBTCRkssNltyTR99MSTVOcBxK5CkJVxvIN+CukdLO0prF2F
uGGab2w2nIeuVfDZ7fukgb96JX30eeTVp7oSiDHBMEme1z4pF6rrviLIjmevV/yiGqpX+442w6fz
Mn9fBLSnQIKJB9NVB8CDA3zsFcQexyXwctCRqWFZ3gw27JPdkOQEgJkV+SSvxcb3gAOG3CkVI7ml
GiiOinKQdRW8EyoINcCjK/NN4c+HnaSpqpc0QKH762vHsALlqpLyhSwbahlvyZT8HzdAKuvBQNkr
16ga0B/aY9HeOinvrre9q2fmCeuBt3NoOm1IIxm75AfenCzL7oH7BEDpdL1jHzuX+QgOftofXEwO
LPMknEe01bCMW7S9DcruxT4mfBdBQX690H26q8M4WL3MTXWOS5ADD8y2x8vuF9j9KLn7Ob25rKUs
F1ZdQnpO0PcBGHkBK56I/OOrqV3MQzkoJE8Nqd2z5SwDSHI2wPfBzb4dC/Dkj6VUuxtHT07bS+PQ
s4jD+OWfStollJIW5wRcF+9yL9mhMKhiBXbBsH9rdApB6skfuM5ut6dgiDVetH3gh0Dba36yDMzl
/aSEVvkZp74ihYSSvUP/y1Sn9/DVyv9ZrzYzBLKuUR1PuozqfHFj6hgO41Z5JE1Dgke+OBr3HFvG
eU95DG5zqw+mi0rhLU66Xr6Lg1I5z3H9hnA90X78wkThe3kSk8mjiSinNfPp357eZ5rOv/YfSq5G
pgNuoOBXsnkGBqD73CKnnxcMDofdVgbFcKgn3Oa1MyTAYanAS8x+2DMzYZTdjt6i5v2Dpgy3BmcS
GCgOZFwV5LqfuWr56biWrdQwdMY/v1P51TxLvhheM/rFAy0LB+lrs7Kx7iLoNCPe93ZBKYPjOwqi
Blh1OaNwNgqnPSCxOBU6zM02mbiJFpNW5T5Oh2UOYGFjzw6yTrMCv+iNWRGGFvPI+szyqzJYXfYO
lLNoT8YPGq8FjkdZPsTfZ3nwzsDFDH+PmrRChPomv0MUqbkEiM/7ytMtfeAuTtEi2hGeH6HHd+9I
se6P2q0VyeO9MqlLIsYEXtKkUSnIsSoaiSewtRWzHOFuL9qmlBbm3D+AKK07+I+BaaJB9ta7PMfX
/ImjYYkgMEethCbSvfWarWNLAmqxzkjNMjlqaYZ0i4RNZtGgiw5avM+pyxHywvY+NVp2DHarfV6g
NTxwXk4zV7x7tQEW2KemiKAWmm6Cy1qydNN4me0dO4xw4gBpE5hXN/mCzCIhOpPfECfk+myWJ7lS
EUMSxLp7D77c8BJ7kSm3YUfYJ01Cf2DliNC7e8qmg6f7WoRvnegPGKKaaZ8lARaZ4YR0icIr1iMr
eJBuHuh/p32LeQ5lqm82o19kFKPKnm/D7HSd3ITCCRfaiATsfWWjf5NJODAXOP5vN9hPdiAIY2jj
QV+xSwClBaxRozpnySLLTtodcdQ4rBevVVrIsb5NI07+tDsf/dwzaJNurEmit8YWyEjtvNl7YmGK
Ulhby/4DdDtzCHYHd+R/w79wA+bFEHD8hmImJdnW0WSheiHEaMl+TQK08c91PWUlEtxtS8gSzhEq
jMrOlraV6YnPzrCNzqsM20Cs6ileLgfU0oY4RMqvEMn+u2KgC/htpvzsYi8qBEfWkGTPOhWMvIbJ
AV1nSLn/FOdzpoypgUddLzRiB3RaYfXaemPpw6fsWY7RNptK2rdCNsNeIM11OxEGK7xb73GOYM2Z
DWfKbxC8S5SW13a0d61yPtBxg2vWv8drygtjtx/nti2grIzI7cZrgdI82Qws+8h/Z07xUNL1XGcy
rQNmD+YaNyI7/5IvYJkoup0rg9cb2dn+BBDWWOhsH2m6Pt51DvCDGQN8WoDKdNzlvec3+oYwvHFZ
9mvuPPeCQtoa023Ex0SryWDVnTnvK8+QdyhgRz0qeJEigxFfr9xsrUMcVb82waEQZ55WGExHD2l6
E2gt1FZ5eg3xUZy8ckSqBl/Wanavdn/11nuheGuinOftw72Sxo5CNVc5AyekBLJvWoHz84nsp80m
+WNU/t6tfLFmKzu3B3GiaBlWtWFtZYMPS5C2rUJYCwIMszGHqTH7ZqEedN5l9ieP2hQ1cjuiOSIl
BmlNCjWtUW8rwxAa+0qM0UPnldRRgSfZBL7wiECS0ZZ1KKmVcVl86bu1AfvI/1vhDp/Hyo16eBJA
t1A8F99ACkkBpjGo4iMMbaIoEPEDL1cMV6opSxpmo7l3XP/t6UbObmC4if4TQJkYFXsEmDkADhKQ
76UK+7Ejq5Ddb5EphrrJyEcqcNoTby/cnFkubHM8jSb157ZXEWQvCbcB7YCYifoOAhuze89tIWye
0ddQ8pVi7/qz1/ZmvKwzwXADmZvRhRQL+7ZurObIgsvznCKpXR/BdpBfB7V0YoTT+ui225o042Lb
wp9JZoXidH9w8AKK25tGOB5NFl8MdSXnoXd/x4CnjlY1k4d6CCa/htxuQTILZu5rVbW+59KgB2Vw
/uD8l4HCoF+2G0CqptO38Nb/DhNYAmDgqDKsvf+OUABFmfbLIcBWIGmi5myudQ/8IpvyMsW15J1m
o87O+JTEcoWW2HgN8SmXRdqE72wJoq2+ZQZWDRkQ180yf3fZ78kBSsGObVCM/vjoTC/+D6FQYkm2
5ji9L/dd8eGZk6nNSisx/o7K5D2Mt3S7lQq+FDnUNlBhR/aYguseodWuNNMM5VQ5+lyEOVuKncZ5
8cIarmERlwL9sKaRDyZ5vxcEV03+VksgSK0QgP8c08+8qRAdxd457nsNn/JL2f0y7RzxYOFKfgXU
VP04aUwUv5zgiIYONwHPmMO2Iy1BVpAknD6VVkLwkqbEeaPuhOhqfaul2R/2/4XYPIsX2QrcQoGH
tawbp213IJy/dQeEgVaI7nMWLm1kYdst1H7xwaoFKaDuhWqh75g3J0h47AVrd+A8UVdI+I/RX7Fz
B1qN33vTpsXC1+Q7Vkq6DVFLn429Ft7gXkmgHaRtncIVnccVdJT/XjMvNxEdIx37e5Z2GnOviGDO
YDWWywpqSctXZxVvPMDrDEPXWXZ66AkudD9cIYSBJn5Q5sHW/TQ76sk/3sxQ4HtZYUC1Lr2CsuP/
XBmCZGMX/WRHbDYj4apCFcIxSHWNlEoZEwcxMimpx/1vuh0cvR2iGZDBgASb2f1fe2mTXahVYL8z
TY1ECiX3ivW94ARJM+NJlBdjyMaFJ6rGt2cLlT9uAQisvZwhjmTnRAqIQ1OKpq9FIhqLNjO9O2iZ
fYZ25J1cEvfpDJLuGHtibbdxpGVNmsSVwVWwYYpkL2SJQb/d1fXujdpewez2urTWcreLAGEaLaZD
9bZlqES30Ze4zC//NsNER/KOVpep2/so1dX529mzoyA6z+vhSz5iv+qxhbQXWSq0K/RBgGMret53
G/VY5Wm0Tw00zbH7b92PTWLEfpIUESskhetqaU8GrMPnF3oSwmPSIIuXvqCwit6Wr1pvugb2/5Vz
2Da/VM3Cf/1s8BzaIWk4vdYfWuJXMNMW9kgYjxEW7s9WmM8zL8BnUmxK5hua3Ea2p+h0QpEQCyu9
k8Q4l2ySo2iqUioZvSY4ZYlQIMU2rUuBSYaYI8Xy9LgBoYz+9oO2sukzzBd5NEPbBA2bFErmhDVv
r9MHxd/TC31VQTrx3m2nLrPidT4BlUqzBxtP3nS3CoMy4iOHPBYW1wT64MYM7/a5afy+nlokr2Y4
rWjXXLANcqj7ihG2FZjVb9r1WhX4YaLTgyVT12qwcWv7mvcfpeX9d9gu0uwcmvo7k/+AxkfXPnEr
ytUCNKDmurzagPLaQnODdWr0Ls3jtGEdfXoxXw6ap9x20A0+TtRNC66NXpeOCMEQfq6LPx1WjOpg
1UBJ952kJzfrXuUiYm8szy3CRvty6EE824ARqm2IeJoJLowiKK8RlLuEAIJyy0+iZK22O8Kt/HqT
Rac9xEa2jEGUcm7UfY6KjhGS3M/z+yalcvSWQ6VtygIkMc6x2E1z5m5k+842mpjpsP9a3gf2BBqQ
z2OHnkKdm2eIj2jQB46GHSwPCzIS09o6F8K+a/83lfBzkpehEtSHuEAgc/vT2u4z+xXD+LUJi7ZS
sLRtpEBsGMu/IdN94C9ZiUN6ZO1oulTC1nhId1i0mb51aQsPh0nEiUXPARmkznNYv+u3zMZCjdfY
BymJmy6r0YyeqQo75THs5bD+E25YrMIpd2KJwehQ/9sAVAOiTFx651ndqaKy7JE+jA2vKA7m8TCQ
dBsiCDI0WuWhMbxSOGeC6fkMxKAKggFZQ3IN1fcbVVBxFr1DgERxc2INeXTKoyXrCxlX8oJGtbIO
0uj4UxNrFJwQkMEmDvdEgxI6bGxO20Q0Dt+X26Odl2B/PGCuyJm+Z4tgak6erjtsZnvqi7/qCiEd
s5ac0iRAqf6lMdFw6HIwLVzJoH3YQCERUyVjBQKrYnlkX/s2DOjH2ri0taNEToS18X87sJwiggIN
iiOvIrUw2FbFhuQdf69+ttd9XLMdBOISNJplBJy5wOtDIRyS6PF/i9Jy5g2w5COCYDnPKDCezj/i
G4h66zccEa2lWNkot6JZjbbZ5MswmiEXni1vtEM+XRhpaB3alo4sWHknS0jdoLC0+cyZ9Q2S3kRE
MeHrNShlSgqXYhNrJEP+PiqaB6FjiRGQqVgD1lrr9OsMZGF1UgEYBVoiLSw8wlWn1H7Voly3dCTB
Ef1QqT2+7rCFJQIt9hu6jypHjQXuzjVuoGV+70hx6KCCYiOgvEb74dxoTmWJ8zx0T41xtetd8adC
gMD7tFEo6n2T6dimrmASOHpcIbMJn+lwpkZWbEdyXG2joM7+YRtQoefcOb4jcROraHRxhfWmwOh0
QyBWzMTPMesGVdJoLU87Q7O8cqLODt+N1asgXKyFUb1uh/Jf/v1dfd0A547601RVUrGYOJiXRlRK
a8xoe4W/u9w1h72rRI+3tEv9MUoAwnDxVcrpxHkWaAvo9niLbW49xpecuqEAUEu9R9hNYVbClKB5
mlbU1b9dvixyfoOfoqEmB3ofLAyXYykzlzpHjML8C7/asVJaH4MYKLL+GVkCilQt+40vDWb+Kli1
ZxYF2FGtEYDcqbmzrAf+Naf1nCuRP/I0Ed2gJJH+MfrSZYuSiWfSN3ylMa+Hcue9EnJzjLZohpgu
ynR+IcrmYNzN5gy2yCo+904GFQdp9/7jt2qD7jeruYiScJ7SsIdfprmLzlpAfIwjgCgqunlLjaX0
n0ilkg52gM/6tRxWyL4XQj/nFXdn4jVj3YLaas3bfsWrXCnBeNuZlZaOeqE1wdnvxWkqcZBwDsMi
Twa7noCkXTxFrFW65VBy7Rku2YH1fz/VwZ2DINWkww1jGyXodtZMKtkfueD90DNl7P52850SOFL8
ktcWGcjTnCpj7cBknh5SCMacO9xSosG2/v0Kms2o6QZA++us7NrtP2hw81l9KXkNNFdkmkiduPMO
Vl3hkiyC8lX3WnelvmZLm2HXstQY1TA2hnnBs6OjostztcKWJugm1VRLnhnt8cYb2Qske/5i6P5N
TlhURvCkMC1OVfnM4FIHVzKiNZ2uA9GDKdfbbUVT1oZ9dvc8BkZX+W9ZPTyrpVK1Ved5jih4spYC
yAr4M0B11nbbO2cyAeWa0VQRwnjPI1l/NTAXtPJqLDX7fcNofELt5Q7T7bIy48If7W7kKxHPDDYz
sZkk0PB1Qfg97EmSqGejBaUxFJqWs71q/6HQcUWMf9xMc09gBuB3+kDnoJlVzxNGF+S3gXJ45gbG
YmaqWcG/N+hYaZTklsnmBisAMTgvaUUXwKO/dLA3CwEfXA6QfRpFkHE9FgiFas065HblUShYyp4g
p83+D23QZcCdkO6+YEw7pemyqSbPU/9QTj2kYTnMm9W7A+8MccpJQRrrknj9QjMCDwLppsDR4NjG
ETmiAzVEHg8tlbYfYomAM4VP0Cnj0xX2aiUbDoJDK6w1t21aqjd2M5Xv5cN671zMK4OoSuoqP6tR
SgGJ4OVXcrhm6hEOArofhWpMXARKUrVzs0ZWBbM/j5KE33wTHykm67jClsSqKcNncmi9QR5zC29f
AioPsgqqlnyK+Am6n1FCi6nO14i00pHBby//Ow6kt9hIrCBsiEXJghN9qb2Y1R5Z8/AW1ySdOIu+
99pzFU9KEfxxQGfJxD5HqnOebzmlEnLBSCygoyvFf7Q8biw0SyCBzMOvP9c/BFPyyH+Hd6N3E4vp
zbvUP8wm+80lK1arEwThhvbqK87BKqhjCubibghFrrMVenTovKVfqDI/Sj6LwpA1MzlX/9qf/bZ/
57fCGOEKs1lQsoBf/tXkQDoPMA5EJspUeHc3jMA3OSs6jS+cTZgeWasFc7ZhZUaj/btzv1Y1eC6H
P7QZb9OW5y2ctpEe7eeSJequAVHCGLSn5Ihj2GXkIItW+jF3xh6zHI6iRQAd7vbQDyQ874t92JwD
KCpWflAePpnu4GdKMZ9Ep5M5RSXWQPkna4quQX3xZj5qgc9hiAHj9lIBMlFgCm6QAHL7J7HVOwR9
G/knfcG+1hItFss2I2Mp2gfaQ1vdc24VjFU62PgeizsHK8X9kyY1iwPaV/+yEHvrGN0XF6SMhj4m
a9YALBM5tUd4tm52Ski/qo5iIa7LfxpIhQvdo+0+2qQ34WVSoTGd6Um7ON1ahSgL9wSuOGv8sJX+
GuArM57vEZoEdJwuNSwE/zFGoN6cgexLbSAkGAZV+OhuzNO/RlTGURbcb9RFBPwLTGoeDvXj0YJf
YolBZfXeaCtU4SSpxKWGyRORkChUYfLLlOWoA0+E+DqxeKVe3lbG1W+ITq8Z+4BnYtoXfRudoo6+
U43ainzbE6/ySE0MnnctmUWuPo+kQEzDx7KM4uPOMJ/81wkYwIXoQA4gw2Wd5yp832PORY9u7zsg
qpGpH1hYyKjTdJosDabo6NZdvUi1DJC4teruWyKj3MsR3B8F9fiSqwTkmUcbsYeef4vONmKYbPTi
dkNdOYESmajIYZ5qdm2MBWTyo3jrXyGF9C75rxlWfX+krqqgTAOdminitwfoE5H25UV1YCUHNlEy
zM0xsqeNzgZc7gKdoHbEpHrZo2YYQuGHPwZ+gsONQ18CMKxU1dbx6TTchLyjToVARIXO0Aloyxt1
FTEqm/psNYN6Iuo9GECAcqM1gQjMYxRCGEZbmMhSiQMEmUK8Y4EoyaN+ohZdf6VvjdUW0iZdwbl9
BaOrcl8DrDgf1rvK20ho9AzjE4Duspx08fuPrBpSI+vAuQ80n2wUKGgY8yPMgywQU2ZODLp9qMYU
L9t/ArV+PK8MsncxXkTi3vSCf0oxw08vYWzRe2e7i1E2vVC/QkApVAugYsJBodmf0SgIls/cAmH/
eqmZbOc5gvbLjrpr/f63+LeFkl26T4haSKA0uyheW6wwfddUK/fAIDykejhB4o/hedg4Dl1IWJ3Q
fZiVVXGB4+sQJ/w0fsGm3CXWydh4zBZKZrjKGBs6iEIyxY8Ijl59kUIeBPLPxN3FZpGbcKxxc1PL
4rDB7yA4X4hX9O6usUAi02Syde3pU0LhfNIe4q00JtF9v0yqGDK+Eu6p0hDIxrrSGFw5EVexLewZ
F7Ob5Le8vpibGYINct5iP8D/f/gEc02zn/NJAR3d5rnWsL9irYddHUki8K8X53I6tNM7AXhfC3oN
T/JfzpAaP5evkQI9kPFX4RKxa3xxqJRbsN/M9cFubAFErkkDE87JJ1WcnB36rotjuVGOiJQow0dD
GtalcDsgwADX+qhmOUsXDHwEQupmLRVsS0MOxF3bqkmxMZEm6hHDmGqOjiKsPr4fgTwADsWaHZBw
1xiDdNOg9DjOY5QXcXNTT2L3w4xXRgIgwK5YOQLxx61OvO/8mE0V7CmZZbKy8dOCq9lfHzHpYqmw
NLMTnYXhW+D6fe8ip7/3NiW1hkScxRNyizQ1vnTjvLJoTNdvDQxPExGVoRSCt4QJBh1DIdn+LCjy
ATxLZoftvowWSvInOmtMONj7YAfsFstY7xT4EI3omJpayRN+7BQRNLmONtEzyoaD4CglVypW6Xck
JrYfOaWupPCb8J71pt5aVciHhYpKcxAOPNsEncEMtXziVjPnGcsp7MHR+5YPs3ApjFj2xyPVSeak
meiPNsRC6kVH4J8hFEOBWWTzsO2bLT9SjDXsT/pVa+3GMIEhZQia5InVBoXbCY1CjwmsdzAZJLW0
+XyyIqPPiGE4thh8zHX5mxDDZK1uZxz084cmGsdxZLQZYGE5q3doAVx7CZH+c54ALb4F2z4VHzwq
/m6mp2wH7WxGkZ/k/D5b/CtSacbb7abPidBGgeNqU93KCkGWFGfldu/2/o5YlTN0r0PM30PN/awE
g0xEUVHVb6zKtYF0X+92RRniqRhAvfYZwVcuPvVULOMXTk95cuByYFd/aFrJ5XKHPsoBl52EFu2s
Ll7WqigXARUVBERY5Ij+/KlpVtjXmn0YDyVjHsiHkdXghvkbXmGHJZVs13fR54kQ0KlExbEiNO3B
FT9Z46175ShHKKXas9RUq4Q/bNe0X+6uLYcHAxWAabm4ba73Y9iXGD9UEIJ3yDYHU0stoLXqI15H
vuh7IoMURgIMNSr3pvRs/6ZICR2eoD68kVN5YefvN1/i/8CyuWeTFS6+yJLK9klLDuol3nMh5F+E
tBkGGJ2qSHn8eNPIrRn5M8z+wjmRvCDjp4hg3u1KxknWskcK254Zwd9fzKHsbmPyd+ePtdh0Cadi
Vf3J3ZTkqD+D51u+l5liKAtmW6VLL+WsnqFQZDTnefKLJCLo0tD98NYEQVKsXekpDKo4Z9zc6znu
yC060yJBzqfs+Xv+H4XToyxsz9xJQI5OUun3CQOU2IEApNOLEjx20FcH7fr399Pk9dJqWmf2Ogm6
p2iZc0jFRvqZ+Wvza0tsagxSAQGWGnD5TXMmxeo8RGIXwZ9fws8dmpCkLuEtC0s8d3crocFTfRQR
j4oz97UBXf/NkxOwS05qwRu+mxPz9P/gOzo6QO9P0ZyK6VxIYcUprsuq1MYje3wlQ/pwV5NHDAvM
9SF93sduoi4iAEieZwJLv1mHTi4qHDTWsNFOuBM4I1w0n57tmeE7WCpYwhmOkL9Z7Uyisjoz7SE6
CVijcj1Dw7rjcu3TlzIwPkhD+3Xfq9GQp/5Z1bsBhcZLo6ATw+seChGek7tJW+ex9x/qgXydo9Wj
evydkM00XEhqYovozy9f2oRfMqHaVJfIIrLh6A5YSlrAEHl+5yX35fg5w4fABdCjenNng/ziaP0W
yo2pYzkrQeOokLRBWnyRsuR3AUcCq1uPRDlsb73S4dkdoJd8vIDc8QAjwC7WhaXpYTq1qp7cMkIZ
LZgvlgVCAvZLmWwWoIO0JUxBu4MQd4VNX6sIIccCvwZsWBhuDEweuDaYIsV+BWp19oAJYCSOTYZ2
BomN3h4iFCxAAcq1R/6Q/1EKIOCSSTb+HHZO8VxZ+FlZF6NzPLdoQMvl3p1AIN9lJa5ixMVPMiSI
ALPbaZpJSebPxsUcV6wrODB27lFoGGzTscA3KmGe+JcqmEZyH1iHvtc0H45axh9BabHYtxCO945T
L+kCv3aFyscvvWpwTulXN1ockTLN7GCw0lEVf5iT+tlCv7DZR2fa8jz5Y0sB/bHSo0FPA9a5H2Rp
zdz4PuloSavattpO3deSLAKKpiVKEK7SxzkWcvRHuIIgws+MzHXL/HkGij6Cn5NP/x80pxvuQ4wS
XQrbTGFuLrgVcMnG1XmLOZwMH1I0afA9bqUojl090RgNIXnRrI1t98RWmSwmq+tGb2bx3J/grXH2
XXDhNSvsypNKu8fMvtPXDa2FrpVSHjEOYy7l/PAj6F8rNEBqkpblUcS8IinxEeNh996b5GDVlHNJ
SKfKEcChexvBf37RElISRHEoyhvzQvD5zxxv9Pn9bMFc/zuoMxLeA9+QXDfcvS1tHX6oBRiV0dH6
sq3kmDp/GUd9q/WeMuvfugiqDDUPoqwTy3TR3NqV5BJ0Zfb6+FyxLr46WSZBoz6d9gx0r68+jYQF
/q1fyqGKEBfazbhOEsy5gyqI3iQtgld3Z6B19BFC6FLJ3TvbQzWqihc36OGo1yiBUvdRITQOsRp9
8yw+NwFPrNEUqFgKZzfmMXaA1VlWAS4zqW+LnsFrqJUff0XgPdVTa472oeIM1LYowzKAq5c6uErw
y87EU/1IcckXKBr0MwjQVu5WBR2Zsvj5A951MOWrzTvRLGnKEwyTutnOg4QLdr5EJusz93CZ7lFZ
MN9xFrjqneH3tvlNgJOVzyPMWmo1YBPhhKnzr2wxryb+HwZU/w6HMj6QbHLowhQV4OVgnDwYJKxt
PMeKNqyJiwbjN//4xLvazVfmfWKfb4Cu+1Fn0JIQzNnBbeX96xKjNk61lZeHjY19IgrZhUODpbg9
aEOrPoj2WEk7ldK27NhnEN1Hj8Dx3bkRW8E63DGR1toWFCXrMJ29R6E3dfiTTg9ThRBINvvn3F+U
1TJl6G6zE6AXBQaeZUmyk1yUOkf4dcFisE9d8AIqasE3hv4Cffjzf3VMdN2yzvA1F1FFWUeN7hh8
uHOYNYeAjbyviA/2SvmzMsbbXH3htzeKWDcyaU9E3l0WtReqz+iC/MjOOHmdopzGxFEf9kLHDFYv
0X2VBJ30dOStMc5fiZQpdabOzghYGpEyg0Y1TQWUfiAm7KIwzK903Ulh27vl+JIAxP7pVjKjuPpD
Em4T/8FcbALnVsHDbJhmoqFZ3l0zk3WkCTJPXFw3f5IKcraawog3nmg22u/w+IgaKKA6v/eWL0ps
szHQ4s+0Z47jMzkrLSqJp1MLnFbKQfAqG7eIBSt6Z91kWWS1pBs0jp38cFSJ76XKmgT6vtSr/siO
wfN0+OluEm9aSFlbdnwmtV9FDikf2c1UdR39uk+L95xHoFdgxlBhInia8fAzFh2UU6e6B7a0nLi7
4wZPX+JFT9qbG3xueQRj65QcRqhFA3Wo73GCVx96Jm7fXwZj8Dvv3UhuChEagasDVAuYwr3dK9xo
nCvMEUCGUMCjEPtjeWlfldzaA4ONjWv39GwRbdOmdmURxwmJJcskeb9Ld/sb85DDIBGYSDthjrTp
SYKD4G9emWZHDzZjPb6oUQALNdjUDy/sXuyugtFWfdmFDhznTlWZbKhTWb+tWi4N8PWFaSh9BGjG
Lb4Qtwp/p2C5FP/8k7b7oPNXqDvHre63KfPGZYsDm94HblYS2hqvoWfQFDN8RXW7dsARUCp1Nj1F
5JJUcTx3THJ/CuZLoA7aQqVoka8L/kOH8tsX59OUb4TA9/tJ6pozqNI5iMqBixVtmDw5sdWJalpx
CHPrRSQiWekctO3RcE7aMDVkmmnk76NWSOa7qLZnpoF41UCy6mrTIZQ0nVZTeaAyHQ/e2+6HkM+4
vChxnba9wqA1MDotOFwiKEP4tJ6j3qs622S03GAihUYm4fwIuAQcWcyHZbWyt4RQV65SmcC9anN3
85UuqN9O61x+rXh2dLs4Hwmz6JozvsMsKhwMqJQdGSO4KqcscNwFgN0X29AD4U6jyamC3b2Q3tMT
H1qPclmnJqXPgCHD31jkiDVvOD/UNEsha62SwtxaawT6S/CfH21K7ZeSnLBv5yY9JCxXG0kH8Z56
gNtfhug72cdmogj7MU1OyncFgVTvfIlwQ61Do/NrkgSaUFoAtdqbBu6gCVoNlTE3GD8CQYRgrcSb
o4WLX+j0+u/LLGbnKjXxJOozlD8HM2udWJ3/6ZFEq5V/12TU24nsQwMYavyXQJNb0Oi9UYDcu/4P
mQGbzldXMJQtMJDCsRjDMCchAU0Pm7avaM0d3UFSPvF8MkdNsdLyKzeds1TFtrIsL0ZiyKslkAcS
ZG8SUu75uJiH3cP5IQudMATUh03eWsWhjJpUJFHQNcOjfvAenaKFhrC492sPOyGhVIUnEY3vyrF9
iOgtobVZS8oAtxRG9PGLjrNjtBtvcBXzL/KoE/EIMTEN3kMr4CpU0OAsr8Ko9ivosF5BQATXpu8a
yLmzU3BQbExct+McHnFfbljK+IxN4moASswOhNjO7BGKdQu2PcaR5UZrKABc2rG38NNi6Kt1jl4b
nHkgPVI4bCNd2eo8E397rqPgRlZH3iNYCrYZdwGH+BOWgOMApexde+xYqUu8NPj3QpRn5rVadyNJ
W7tw72Ms9NY/vu93j6U6Z/mEWfzZO5Yb8ZTkpeRPhRtxG4uqoYQrPW7ZHt75/HJlxPlHwyPjbNRC
Dnta+y8qdfL2ZsZMDDwFj15H/ze2MS172lcW8ltkm3095eXwGloumHMZoXL+csAWRxO7csAEZDty
NMivxTbUCyezWGbd7KwPjgUh2ICsIw+YRWE7EZ/Gd6vH483CU3ieyl9QDzgBnG12jk6Gls/bPJvj
0f6RTnfc3tgOtSATAcsvVY2K44yzr0v0+GJTVQx/WJE2uBRWITLO31/PLJWUFpDqH5AkvOKLTg6W
8IwdQtr9gRtfHLnd4E+augPHhUHuJrIPmpr8gXF5T6IvPyw57VuW2HvOgPVcgxYJqTYSpyfnl2WF
nO2XsM13fyBRbaJOmsIlffp0rlWOtDR63lTwaJfd95WtV9oB+hcI51/7L2hBHuZJ5FZJfyz0I4tE
4ZWptexzTrwFl0nUfhVmBSVG/I67BW1KUWDwyfsf8xSn9d8TWlSm6DVHvHqnZ4AEb2FCaaxFMOho
YI4bWVsxYdCPDGUv3Z3oszaTo37/YLZKEUk9aT58JE/elZLrn+ZUOkiO+zHX2d5DnmIEtsB4+bw4
TquEqAYNrcBWox8oqRWoJGRTlB85kQtvOqXjRqDzlTqIPVJE/84WjaW84AYzJurEeCEz7HfiYKKc
/nmAQ3qhkz45HC5+l8dXXEwNFiE2qENGpwwdr2JZmwlXTEslioxEKBGBSlFHUIGGhJ+hhigN9MSs
f/b/488yquihLghnQZtDMzr75oiWRPIr/2WRMhWC5e/UU7Cy6Ex+k+J0wnuwbBoR6zWckCybcCvy
bCy03Q/NOby1M7k2Gn0alyCU519djBY3Lm24kkYVOJZpdTph1qlzHJpee1RRL/q7Z7v1ReeL0E6o
5WdwLk7/oKPw4O54++9OfQcTW7SI95BjO0TbLfmFn8vaZZMBIEJLt4H/BmMCQd8DabafBplir8RO
SGNB3KD3IHQTKVaHK6V98qRuJfCdXujdtmtATekv0ygPa6wiMSAcji21j27Uch4w+cyK3kfBicN/
4rWQdbligsJz8jRa8zbfs+tCV9ruEJM97URmw5aV5vKVT3QxBMrJr8Q6u8mT7mJd+J8TmxvO9g6+
QN2sTrGZ7XLXElibtiDm59c2QYN4aYJp+GHEvfkFEPosLU1ArRQY25hJKjyUBqz8I2GZ4iFr19eL
QmxvQ2viAtmLSFlfbAwZW5zIdIZ/sL9Kbji+MRsAk30IYt6LCrAuFHU3GyJa+tKsDUb3cglwpgrK
86UE7jG2YwqoxQSvQjeSrX4DOE5nG70A+J+6/ClUrgj+DT2I8yBN01rJkVeHDfuX17RrPhZdULoY
Mk03HVT+VRzgUea+RPENCEIb+HwpEczlfOmruU1h8T9ZdKt9kpsMzxtDlWJB5pyVb39xWhNPUHal
kdNpr/N5J7tOwpdE7LQAtynv1Rm1SqkxcBPlBzAqwzw4jtlt0DtySXmj4P3MT2+Kwvbv/uoyZadK
ZAJCAnfjf/KsEZb+cHi044wjsXqLhjLcO0OaA7DWbILKvSDCKv1JtfNNAy9zoDuu4jgtx84pJL/2
HwXEJAm/uvcmsBqZBEiOwyfzB70T/jvvNV1DNTmdfYekGr83RcYAKwmhrqzk+dBrI64we2uEIXDA
jjzP0yJPjha5WDgMtiqedaqWmv1/E3S3zxqsvM0Dod/Vrn+zb0yjmhG2jmuv+d67ibaAFuG6D50S
eEpZEj9ryyURyt1OSNegmAQ8TBKoQZOl/lhp2QPxcsZ/gKzf2HmEjfVsA9aBFonLvJsL9b5Int41
/jVJaVgMcKQpJ2jcjsjqRYEnBCOYzNz9Q6uflnY5mtCdhcYhcr60Z9TJpx/BdCc7UHrQdCglYaBa
StdnptRUTWh1SDTYwSJmPUpG6sj+R8htTBQTx8rgb6DOoZffuLBBCvFpEIFjL7rUP5DBKycMK7A5
WNvkC0dxqIT9wLkR7dNS6XnJNtlgpDlO7T0YlRCDVEMWTU2ReFC+jUt78XLHyQUwSIsonW+tbt8V
LKNFHGtVtrvT57tWx/h/rJPNewOwOXYv71uvZbHjLdms4nWjQ0QDChWjLjNl7CPs6vOMqsDaqwDX
MhI3qXA1mB4UMiBF/xchKyOPmHtAyYqiLbNm0OL6AEDfgvLX08/oZX88gI4YO/UomdSq+QctzIov
FQkOqM92XBj3ljJvc3mjPPkuEONHdw1h9TN0c8gm2SrYDJWCaOCNzGY1oR+9LWsHX+TfeFNQYAax
vBGjpuqWis0eywEk4Tz6/+c5bTzwIK00wEL7/DobF0G+a56c0R+B5kzKVOPbkMgdZ8I5+U2daRwf
5H8MnDZElyU2tRxxEE6FuCPnJ6uvh/cdnfS1/Eqq3bvKU5Akwwy7S4qW4RCIpNLmwshvbKcdkkDp
RjJuUALn0/3xE8BVA1mjEXopvgJ3tXRqBoTehhgroYXigK9AEqyHY5WLWTgUrx5EwZoRtrPCWlig
mId1uAu9MtNNCsbk/96cP00Zr6khOCtEYeoVjmYcr8PoMYPnIo7yePPzd29YHJfPKjrBMIfV2kJm
2gPY1QtXJnP4VmOKE90waxolI78xoVL76jFzU0ey7f0bkqKDxxgIHjp18SqDA98rZ0wXfZO9fy3k
tt7YEqmxqei68kqWN/AWuQUiOTk74SKIKYzP7wwqxuH01+2rJy6ZQpC+fMS9hi16dw4WH2Z3KRj9
VZm4N+XSuO0s5F38JyYXCAR37R3xCtcu9ZYldSiI+5OIeteiEUJjeNPu3xfjxiGhwNKObu6xZg1J
nSVeCGyYO97fcNgBcFZEK7VL2ZVFl3z4TX0HUxJluYijQ4eC2/T6X66NeebbRxEHQnRlhDXYnfpL
mz53rz1wUcWnPWb8DNgjSOJFGvfHIcfHkidQOw6n5AGVeryWx/NgEmTHzlAJ7RW9aKMR+mQIe3Cl
CcKLGiwjxH/Vwz54m05QrAWY9mKOvQJ0DM/x2s9/PCxfboOgNOGQ7ndks8clSwYWFo2bhetIJvW3
PpMsuMdCrmdjBGjofSrsX84d95xp6iO2V2GiXhrqo2nFQAJH/azTAqHocPcR5j4WOL5j02uIyUcm
8eWFLiodtKSstD5XcIjVMkEudnQSvh0Ty/R03NB6W7n/3K/iMnpfzGO1UJpeVPoR7RfQW4lsBne0
pt/Qay93kXm0x99b3Ty18TehvO/zf2AmGn5iCqca9l33yn58lnG37Glzki8e5go5KrYsEJnYl7Nr
zJihwIyLj5fNozr/TxA8D5H3wZ4GBqkomKs3k+w8KFTyhfcrvR348nt5qSIZ+7IZpFrsNY80TjJS
eXWs4/5J/z9wUsjVQcp+CRiwcOLdqYw9bt7H/Ho5Ys8y547FxCIYlv+LvlmI/1XxYqD0xF3rJ8t+
QXNsKdl3q96XHHoflyE99gS9t6twdPAd3OgvZmZ6pocZ5PebtJA2tW3EDCOT5Wcpf7mZb2qHwSCE
zqEutwXwekzIu0WRTgEUVCazmFvvrhiDghSRXtnhtYYjqgnZRFzvfwCKC/Zsg6JlL2MgYCwHkmjf
6NClnJyI5LILnXwEfFNUeToBd7F9CUKikJDDqXn2LN/7UNo67MfntA4p0MEJvVW9+27mR7pPatBC
8I/kLd8LoHO0pWeeSrxx9rmTMmBz1hW1e0w0Gyb+cafOAp1vzLzqJbQbhNYC4qr8jYzwz837LiSR
6Y/2p0jPasxtL7+zs1eEtFCkYpVyUDz30djwUw5yFFYzKoWA3mWXMMxJQubQ/OCceSTn3QBJ/1Us
4lOTwt2/a5swUmfMwgClKZ9OZjZ1TwdHiLsi4zXWlCbraUL/7nVsCKbbWgxSnNCqbPmbKaq8X/Dd
S1rDRpeZLPAl24EEcyQP3Lo1hYuMHZ4TUysi7atP3eSoCwF4Fxiu2OPSORHMef1w7fnxnkAR5p02
0tNV4NbaCqTFTGznM2abIL7FDEhYqGRQY37DiWkzM59ElCtFZcM6pPXzcaIrA/mXCBquB6qVb7Py
ow+GoYzBQH96/cDGYbWrpY09SRUBRlIXgDg1H0NiQOtO7Iw/YC3SOJFuMA7JV5Zi4mN/OmQLJu4/
iWuCp58uyM4EGFnTZurqCYdYRtFGLATB6z9qVxx11Rx3sZNO4p6os1v9VYeT/HRg3k8xP+IRv2Np
rZnLoD8xH8b/7RDa1w6Zu3j9EEuz3aRjRq/BJK6kk3mlKAbLkPIdetIWBpxRvngkszZjpPhPZl6D
qifMfg+j1epqvFO0v+0ZMq7ELKrnqIcZ8KPKMWAwHPw1D9gmBbxtsNOgeA0t10a2BbCvZv07Ii12
DbFwwhr/Yj/f/pds6m0ljKhwxaXGPRkMkI7B7Z9NeLgbz6FPa+FivfUdmZnR0DV5ueLdMxgo6MGp
e1BENXEQOMVVUuadJAa8nICSXQEPkrsHCKHXlXBzgOaUzvRrGH6cxgN/xd5d0gFNctNzJyr52sR9
l9bFr4Yd3nDYy9GqpYlgsBGgRRi7fSmu+WddRILtyA7BZmW+PKElEnRMavEg0wdqGiv9kfgYJ8zB
IqTuvOP2WFgV4E8L3trnki1Oy4sghOioC8FOYUnlXL2RsxAZmUGXx12JyXUp+6H8D2b8G2Yk+9vg
quV8OqqttR7LjS3REsIv4nL2txY1YVIhOcPST61DAmneCdGyfA5wLrFBEiHtn7hqeIxtkQ1pJdZO
eHBZZyd7DqtpIvsTWAwdJ04bISSjMTRNDJTCJN0XjCRkVM2Pjfz2Zf6KNR4QiVHVv31upbClUPhh
3WA2bnA+YjxTYehFYeWPsoo3zkK3ZfMuwU0n+WByHWcW9OrDy6k5rsWSBcJmJwsUyeS4b+oxm3EC
HhqVCr3mVuRXQYkhuUhZcSlR0dD7vl/yBOIlXx7rnweKDV4hxq/DNmLud/MVyTEtBTcJaGKZHV6H
tsxXPjBvmp3oqwNP73s2MjGuEG7U4IcYX5aAtVaz81us4PqtdNo8uG2ZYn3A2YWaAGAbI8bGtDrX
7PWG4B4Vmlfo69qVguWsWy3Y4tXaVU7Rz9uzODBcwZS5UWA08TbighEw84VdOh4/WKYpo5mcuaW2
2Q36HhKpK7pWdmfTb311WxYwoscpKOZ8FcuJFuQNX7dPvQUAe0WCH6fBjbl+FGP1Dsfsyrnfciyz
3LE8hv5fcdFB5z4a9h5WuL8lkhkqFB18mwzdiIY8XyzARHaz6y+MYXih7UhVib/73tB8hgP6u2JZ
DZYb7tGEtNNiCWOCz3XFvydsh5CcZ9K7WqTKy+d2xRKmItqEL0o1Q/HEwVQQPbvi0Hu43WFfjIwh
Uz8KU/VdI1nRESxJmQQ+ZdP33aTehO8toVlp/st1AuJP89G8Z3fXxJQRjJTa15BR4lQV6/a+wMmf
T+jMLTBvLuN4+sJSnaHV2FgJyVoMLtH7wyOl7dVxUMb3iGNTw3owseNsFCs2/01Ktjl+/bbXQmfz
WENNqrDqn/PH8g6eq9fEfq6AoZuLQgybq6n1lXNefX9+JGUb0HlKS3Ro5UHU59cirtl5soKvuVXk
mtIr8GubFgTmSlyb2Ibup6w0D/zbJNKfkTTpGREWSWT3ryxi7alYzxnXT5c3sFMYFGF93iccRBsG
1P1VGnmXtlC4e472BeoUPy1slEgIWi1znbiikbeiCpTwxoZBCsqaAVUKS/r5dFo6M+BW75yV8jfe
GZ52YfKXGam0jmAuMPF2Jp523J8zTmSGW8HHzqLoXgAvyG2ojjhnsq1eBVu9sw96zn8JxECQB4z9
L8AS8/zS1D098CU2av9aA8EdUau9Bxa8U/XDGiBQ7VX4odgEfq/DvTxnlaEF2sej0VAsvqOf25mY
Vklf1F86NEvIQa0c2Phuqe+7ifYbYh2h00XObKaCPjXJWVo0DQ8pq1eFLLl4fnpKjnbkz9ab2s44
J7AijJwOYKUKxQSl9gU0MlucM8F90WRqnqpqD1wcn5hf1mxB32c38wBT6GlIwAHQQecaKefZBJNj
YTFFmZ1MdBZQwFbYa4FGmWdL8spkNE5zeIoXYAhP8anzqCoiSNg+k3fyFfBqUEq0kONVtfxZldww
QcJB0Y5r9KS8vZyW5H/3gL8sDdY6zTkYfNPuOPznTRFwngCUQLVaGewy2SHoIT8HkpBp6ffhJVg8
wyyeOtQLH2WSreqgKoBcIaWajU4aiekKLNb46jbBcL8eg1dopEpr5Xld5j/bQT0ife+Oui8jFnp1
t+Jr69t0bV9hKOW8PhwFy6JOqfUtpcgxJq+Hpy3gXUyC+1rk5CDoGvo2TtF8ZYI950rkqCJYJykO
UnfXejOTHll90e6xj8gLuY7ZgtNxf+5PD9ghzFvQcPzJy+xVc03UFpiGtoOZzTO7PA873YBUpSMo
Y4Tt091KCNU51/EjsnoiQiu6dCZocBJ+YKWYTy1w3MmcdZbvqrihvhDjdPzYlkuYxIbDXIY4sbQn
s9Lnb01GMa+F4Qklki8+LDPyGLG2lGAT+oi03ukxKNZaHxotgoGT9Bh5Lf477YBplu9Avk7z3eY9
x59HhV4jPNQVZm9jA5P8jpBxD4Qxw+l5B3TzMmJM24770DLuhVmoFqEyVEQrGwQknulCStV3ZocV
AACzS64LZ+so6d6/2qPX8DqunT6MG6ilDabhOY/KWxyiLuFeFw8icCV3TgPlDdwZ1wDHfE/6xKe8
X4RX0xgha09OC1hfDC/jhqY7PvWfpYCr1RkRqoj0DL7byhgxTR8mL2/diqLzIVWBQvHMm7qYpJJ2
gNMw4iI+dX0P9zlKykrqzYyNcFTcOaSZCQUCQKu+TlWL/4RM9JSXAxF7APu0aTTM/D67q8NYETmH
SWZ6TqArHqMd1jZD/zdPs++f2Yss6pTJAo82dKiwWALhdlpw/mG7RUfHe+62XckHszVfRha+xrEf
Mkuixo+xocrBFKiG9rqW+7VH5mP5OHptC3MmV/SlgvfY38Sk7w0JbHi1XnSSkD9bKfA1pRB32fCD
0id2rw2Mk9V74y0HtqBv+qVnert7iqn4XDCMXlUK823EpywwBEo0efAPqSveOQ1GBQfRqbgFFi5w
49Yf8Fm3tX7i5UZpBGbLUUf/EHAnTymrdAgZIVo0+w+WmDw+HGy1rYH/xfDTlBGqGRd3xsN5jVsz
QpH2ueGIX3/b2tcgW5L5H8svh3JWNJQnSRu3+dbXJoGZGaXeUpd+xYI+GMna18FUzkYNwFS721+2
leNMe2EN6KkOokxmFIVVIHjzQAOLUblpAfaErv2EmCHK/6H5AzsXRxDu0x63SzRKjwA89c+iZZQc
fd4y0NKRwGdhYeHqvurFFGqxC5LD0HBKGANYTrOKRnt6jakqFq7ioJdkPhx2wD+pEnqfKe4ULcwk
fZQEKBj7IwgGiLPqMk8+T9G58WiZ/8y0xpQbUAibrYkDmTFJJ3JRDV16Q1ScwtRjdJTRw/VIXzmz
GV7YAFVN1BHnTowdU1MSi99R3EjK1j7jwiu3Xk2Cxy043gcAKjIdil7a9dXgCoJaUQ7h1nDLompG
nm2Lg3QTS1wesu75C0v+tJ/Ue4g37/SFguC9dfc9l0x0PjkXXoaq0KtiO/Vt3uZ5t1VF3PdElHTM
XlilXwO9TcBZ/l4+DcRp2zvnLx+LqDxo/1tkpGD7RBzzJ1wxJOJFC88AWyWk63h7K7kTmWf8pBpC
phlYFXALoM+kdkBeiAYlCjBhYaXWmy00Qf77o+KrNOqnksRzIt11XWpqocnBi5UQjOuUMCYc4JhR
FkUATkHy9OpvInfFz/TWamPlvZ6eYb8ayaM5X5lfC7yxsV1XuEOQVBDaxy148bsGNu8Abpwt4UmO
dvqZOOZ3UjqlPmT4Ig0EJMXaleYj9jRCKuArgbrcKb+h2QUoY/deX9pwV2zx8pYy16FRd0QpWA8f
8ANftMzQk5dj/vuGkdWCrVXrNdBPheuX0K9Rozm3RjhvpQ+GpEJGRO3mTuJcfz7lckKjCGg7TUNR
f7XtwzZSt669qY3dXTqX9kxKGjAaefQzG4aKC//tXyJI3jyTteDeBGqJ0g7Cdwvklgs0Dwas3h+m
Y5X+QrCSu1tefjIcT/8Ko20xoN3qX2GaY7R57H93COo0DF0ngZrFEier7mofee+GGkIYyBN3qn0K
Eoj7GYBRCeANV+Uvm/Z/QYQwpGvj++Dsfq8GlKl4P8zZ+CR34CD2Lh7tJQqkTxPcvlS6lZedbKxF
InmpVqPM1HSq+NslX6qLU2jXxeotVvbni388MdoOMt+YRZv5bT1x1INTwQzZn5XaqZ/D49FzosV8
12oFpHyGymAQAcLAmjwSYyl1Bn46Doj1treopPawj85ckXpnF2rSwArjDwNhvFq+M3eqk6GbVNmi
3y2Q0n1zpz67K3iu+kp/A/N7wQYJl1W5dIAC9CpUB2QfCOdR81NqNvODxxtz7w6DIzwT9bXv/z3A
9Aa69/cGzJOVsKk91mQi2oJKS+/zNtrbloblJhEzX4eUjV8Om3Fq1kyABBFyt7N6FyU3dHkpwCrt
FH8bd4yWIrdPFoWg8ph6ORdMqagOt+mZR6onxub5onk/bJVSW1/T566beIo2fgQTUvdjp0cXHVpr
Rp0smOmmz+MmjNdezvuP67iJJlSvYMYMohmRmzh74gORa0/VU1vSig0jzU6MUq5Yt3srsRvpv1m1
uMgCaAokWcfrcsuGGCZ58DH9/OFQZ/24bmJ0FZqZ7LHj7Mp71U7LE0rIJzwdaKyLxQNoTGLhIPI1
3+AYt7x0RvZlYFo8V/drzgxmxaSZTHGOmXWGmAbDmAeZtY+PPG6SKp0MQtV/So8GC6yqtmEwYgRi
k7BHQnm8fT+Gxz1pXDDeTMRqZY5+z1yJrbSbO6G6wdfcw4QJiUkBwkKAYWrOQ69OZG1zB4hitt/p
P4gut8jFi4B4LuBoazzbkG8W+4cTJrSxP6ipFFZsbi+WSR0KH1lTcIwpM8Q7FuhHRFZ4An3T6wMT
LrCE8fPcnL3mCiv1CutOInut+r+ksnv5QOCxX4zR40aYGiNObCcnfwUboDps+4mZ/TygjluUhxsm
UoWl5wz/mjLPUdbs1SyFGIsfWiiX4HupwBlUCXlf19CYsVqml4isEg1IwBkml1uzYBOhuKMzW74u
uh+FULufqcESENO/InyWpejUydZSslL10HXyK+ZsUn6RChE/2XkjEZuPIE64eql6Hg0rkEnRNxjm
ko/tDDi9wfUy+h6zWbkv8DQapdUKChODYfEFANZVARW8WSLqmYpDVr1NwRQOojL18/ZZI5ahuPHd
i9O8DSYMe7oIacLyMs9J2NNfLkxgteQtvAs/ajrlFL6EmVM3wxvY5JClPidflzilml86mMhqKetD
5VVZWZQUK/uqFeFU9fmIaxODYkutBWggqM3E4X8vlH6VjsTipa1PWIFIflV3Bg/a5yE7dSxQqwnZ
DvtIUOKHefUluKwsqE4UqpzL2nj7sCBJrZNb5OHTLPouuiU27auPGM93WCQcCzd13DN6BhrN80mr
p0xWQMpzM28C6GbUpErea0L+DTGDUHwWWyDf/POt2ICFf0SsJbaKKcK8Fjji7oZ+YwFxKUak3Xmf
dkYSyz8cqDZ3Iz1kGRqPXa0mC792YVhXySknxPLuo1UxM0p1AsOIHgEW4bNDBqIr9QCt+JFJMsrl
pX/xMHoISBclvc8+ZFfCioVeiQ26YE7gTdigZOzBDt6F4TEXKDGvALixL67XhG9o/vJzTVy83h+b
NQpqQWQfiDvCPVupJDoNWC/5/6KH+YFr+DQVXNMw5MYVqtQbnaMysCMYopzXw7iWIqAA/60gxD+R
O6Aj37P4ci8/3gBTOaufFnonRgUN/TZOY7pR+XaGqJiHDOvLN5fd0SbNmTnw7Zjr3Z7ji1SCOwsz
asjWikzJsAj/iX+5NIdFP2goHZ8XEXrhkIxKPTrYDx94DDaSLm4uF9INmPtpWlvnrgz1t73gfkY9
G2ydV5xx3hi8hMuUHVYdsUDG2FNO83rjkDN6lqh7/NihHOSvcPd7t81M2/7YhlGsTAp/94uC86RK
Yz8Rlb04ryr+9wiBJ/jslNoIBWOm7q8XNrTjnrkts18/QYYDsrqsGGnwJQtYGPl1mJ2qErySr2ni
MT4SxviK8HcB8WZDiHCCrGSi62Cjbwtr6Du0XnGUi45VusKGWL1dZ5V02bMNeY4BH+bydGC8vvgN
4GyvVrMl6v00CiiFja9uSmoDJOdy+uaeaamxwbzsQJjigFu0y8LwOK6lsi/geelqXyrjWaCGX5e4
tIDgSM88xIASDpgToB1c7L63Xxi1/697dGvEoUqIeerde/1hTbtR8P2dlb5YhT4vHDHYI80CZ+qb
xpUkWxvDs6LVnKGd8GAID8P/pVla3jv1FZJbF8NWiEAMa1d0ZpGCH3Jt8JeTP5Nthh3EoQqzObNZ
/Vk8vBqJutJHKDeV4W237rryLwNVi37LCLata/sb/RSd30MfhBUeFQhr32gQlSAhuEvLyAIQ7o43
kpAwy2siixj4VuioqBJjDrIRYrcua2DIIouHIK1kBzUYBR6mvNtR58/WATpot7JzEp7cv012rVys
KAhMq3y/n004/H6oegNyMMd14LAawVITOhlpE+1JsSzFIs0FhLaSEOg4UKqg74zOZz9p+WUHdeHR
c+mhenLNB5RGtT/nDdzsh2EPRwsSX0V5qA62oIqvMigx4CUkpnzAn84LtQ5VjkRrr/TRPqQrhxyd
ENrXAu4NYbHQ3p8xv4FTkzukPdLJ2VR4iPAd1kxI5D+IxjbjISKZBIDxB/TJin+IGX89ufUXDJ4v
jbrc1i5Y1kgxMQB3O72VBxwJ0RpQANJy7HQ/c6IlL5/ScV/+bN/l15/dvNs8K4tJ4G7MlRiEu9Xp
d49D0BZhGGbbs0euHOEn0Rl/C9o9HGyqPE+eHFQu8gA4d8IgkPsXRzoni//OHWsrM8/hKuu4fISJ
zvDMFkF5pY3M4uWw6hefCE4R5sRqWWYQ1zuNijDEc5/NVqmUKO8ty3FLC52XKOmKD2GirIwpXxq0
O/asq2z+0f3CZYHxJUhh+GvmmvSg7brHjo1C9L+/GTC81QwRNexZUyausb7fkAvilN5x5uTcwkIi
CmUhzTjdybDyWhflzTsii/nDwu3vqt4PnGYnSfez/bOcc35Cx2Jx9YSX4hlhZzfY3Wi/S6Fc3ybh
XDHVfypILGSr5uDCjLCwFiNsTaksEp3HiU9LpFubZmutIlTu7ay9u2ipeuuf6ADXB1oKLD5O2Zr/
6ml05VwCjv2+rC04uuZQaqiwuMrIvgfdYIRQzEwQQB0268NRMickFEOb+GRa8TKD5sP5D9YgRupT
gN3u2mJFMnXUOlEVudFV+ZgqRs6s0V0JYEmuCHcvRo7/hObtv3AOkMGB4M0nfl8BIVqj+QAAqSS4
VEnYkK2DM0zDRkUyhZIBpwFrG670U3060Dpf7vmwmaBHizjhYSasD+k4/0HMVVnm6zxmKPxoinju
EzyIY75pXX84P84/qpiLEBF173wg2Ok6QOx6NuoJTfnQnMQtIP/WTDwhciIbHBYG7WbuCrDvZ4j8
h94UURLCTYoFHO7WcMDIxHM78g6orBOKONwmxhuUazqry+WgrgSTBcwpCbs2vQ33chsK8HABwCl+
aU7ndT0uacSR4B1CuJEKw0bmEEkj6Xm6cKCioLryo+FT/zPjk+2HcfruKOGu4pzkNa2bKhE5jLhm
qcxC+VvQe2HEZOsZPxPNb/+PIXxjhmYlCEYh5Phdexok2uZjWER0tWsxwVPxS4CgIS0HE+gAanP7
JYIDGfhWwj+g3hmoW2pvzrBNGtIlADtKMHGgsq7adY16B/dzamSro2GyYI/VgrCwRH/ChVZMR8zu
CGQq6GgXD7OLUljbEx2N5IBwv63bynxhRkmZKJ2Zo+YSR4rDDdnQCVdFhpbYUS7iE7vpr/HX+Qd8
2HCjEYzc5ti1x3C+MCwsFnvhYNKrm+cWUOlbU6q+J43ElSAlFj33SIALr4s581viB2ylgDR3fT3H
AKVN8EoSaxYfk19i0FukNTmhhnnkhZZ1HiPCl1P9HJSLaUiJOvL4QP1vT8Hh1EIJXHwTkyk0b6Wk
k3z6BdmqF/0CgZRWAiPLRwqT7sW1pTbFfP9Q9AHi+ph/Dl+A/4twpDQIM0qcoCEidZuH3roy3yub
ij1XIS7wb5Ju6B/AFthcadqn7YjJSHD1twJlBXgDISR3u8YulSYg5iTXAS5ZF9jk81c9uRaeihdo
95ZRAXki6i/iNslCXiFxSe8fJ5rRo7Pl5NbgMhvp5hN6LCKTwL73ucQ5HcbCRImrt6SUH92l1KPK
eb6txg3Zazp5NbiLOeDPhYuHIylfrFF5GV3xV4JhXec/UbpTUdL2GzOxsLIRuty1PKxQmVDQ0Yqw
jtoYnYw4Jj7radlvn01bqTFvb9i1DnTvc0eAYts5tqJNw6BMR7oFc7ok776DcBxopIi3Wg9Cm6N2
6vx8WYIGGoGvbCfRnCRMAXd9j90fjonDQkYmly462LM9c1BLMUx/r/WueeEMyl9p47YuK2xKHZCg
+zDial49kdKLXc3MHNmcn6zMyFGXDQfBrrd0yW197pu0Nrzj8nL32ZqKId4mHSXDTu1GXwE8omcL
rPZzbV8ridyNs22qg+eadZ2HkNu0l4DhbY3Y1e8nn0PRAa6uW7oVt0kmrqid6IvwfCzuvffxkkmc
ypN/rFTb2gtrRM2Qm7I97xHKYPvt+zlG4w+LA4+rSKoKVQlaFQVVKBZhWc/39aXjHxSJ59yl7C0k
cLJlxuSBlooncGyt3Un/WqVlOFFx5bL0isl6LCDqnjX8HlddcEXFHT2Oea2CI92n6t3lfkxrhuvM
hCmVhho6wp3Mlk6ICQ+6FeLdgj5Uv4fO9qH0cNEtjVP/pcimeegzGLnoKYjWkvZCWOVe0UEqAVSp
8J38C3zh/RpV6bVeM0uY09Kj/18lAiuPKRBuJuPIVswwdz8s8jrZ1bw6fAPFa+uv+WpMpRBveexK
WvI0wz4aWVbk5Ir2reWFHSkaZIb8RCCahPKTwAtTfmAMMSZ8SrF6ce8nv/RiaC7yDw9Ptd19npbE
46MgcX7LI0eUeZVeMTvymZF4gdQGCjKZNOXYsVxYUj8OMev4Ed80BYnnEC73ykOL3aoxHEPEw2k4
M0m2HXugnYGVyU7ztQz8oaUbbzhpPAffi3s17L1Lx82thF/f+2erVqFXEpnrVce60yrO24v0yg59
SfXez7L+D+yEU5VA6mEAPjiSWiZtbGCcao+7IqwkDkVK1V975hq7zplBO+1LDEjKT8ZvmsM0svO6
KGsRAPGRGpUWbr27Yd7oQOz+I7Zw6rb687UpAmCzh51Y9b+r5N+BlxyZMKzMJEHw1297EJtwGByV
I6BxGhe2R3M/cL9Iu434lZR8W6Ygqq7S4989zc5WIoKYBDsIPRMS8Xm7Zu8Tciosb0kcQi5UWqyV
dxVmWPFWQX2WlfpiDzGGGc0Tmo3b9zjg070LdRAxsJmHBlEWZvTtlSdz5imbyD+xN20CbNpxf6YH
W5HnOiBnaVOi3Gq7aLx5HkSqISiVgcVBGg0Wpbw11t03aQyrrxK9BJy1LPuCh65QaXBNj4R06/WQ
erYPJDq1LLRZxz7uLpjxaPPYVAWhedxntFuz6+rz+NDL7kRHyPm1Pk/XhrVGy5ep6RgtVSskovxd
QwXtkOOMOAUZhwPsaIMeDbm16GYNe9TUFiVX/p0KjpME1cv6Xo+vQZDL0Iom5A5s1HrDYkM9bBo1
TwOiw5ChPg9sFNqV3XHmcLnjCnYgMjw0tVfRGYMcQZl4d8fdmk4bJQqsFBUv+Zif4VOqWW69kAIE
tKuHNZ58Op83X07b747VYVtZ5Xkvs/IxOJe/JM30muh9aPQAbfY2WqhoTay5L1A/bF4MHb9ebikn
sqNASjUajExBoz/ceQ7iZnMxOLABAggUEgs0FVy8uusFpjGA2wHsFwkjKrme6PA+RyC09PvUv0KC
DduHTXawJ/q6D4CWKg6nZUvYd9YTpP+xmzbmDQHhT9zeZoN0JAv2B7TPr+68ZKNW6AhFYGxFgRwL
EBjyL6lePE/Z7qk3XjZidBic9Bglq4rAao/A/D95EQGB6DMnZOwgHeNohTyEx8HKqSD3vyEqnGHR
1uyW6N/lGDw9g+ZWCBSHOz5eBWwMVtPoQZ0dJhndmuwTYd3H/QylZ5T9HQVN8yqehCYsdOxvQ2B+
VRljGWMNpFk9WbbAGJrZBTBPKwUjUCJeLaWooe/qNTw6TEmsakOWXhxCcB4iWHnJaqpswvEBrQf8
zIgUwxPLHAhnzhI/NdTsoza9T9j7e3cWqUg0QhOZiWawdrv3tIYwEWGYSiHTszIbljGo7n5OMu07
qhsaP/vPEjkuwyJMZJPHp4NagYwbF7zvfFixvty8/F9iuy6T5bknOBkFrK9CGQhhn4UdEaOUgKeZ
lvHfXPc/xRfXsg+4lI4XRIAxm3qyQmlDqSo+I4P2eGSaTZCIMvinhZykWA19k+idMzoGBAIigNXB
95shLAAZHLFdXRPVbBw9WXpyTCfj5fAB0lrUGQ65FXhF4x08Zy3CKX8barLMjAheAv7Tgx4IsBaH
XXly+ihSWWsFVaTn3Uc7JZEn5XKt0MUGy//KmsZH7gDvTTddWQbhob+vOe4QfCcS8atbPM+cA4jZ
HbNbWrluVq0uNWBBY8YRVSaNxwSbULINmtnvGgmmcoYnPOZgZz3cRl1O2cwbg42PwVAYYbSHXDEW
eQpeo7CRkUnM+ICwKAVKkf7ehHzbBHywOxfFmdBzkLUhqIUTCIAqk8XdjhDeYxI9yfTBAVjfTDfN
V6A9CEQ7XFkeMPU+7EG7k8Ly1MAYkWwzpBNwNqfk6E8P+nwqE6LKsWjCp4nwJuybxDYSyEIqmLCT
aYEiO8RfcIyqFIVel8Ff7h3nkQ+0yo9GwIFCdoVZ3jaNqZ4xKXP7+8tbCE8E6wAHMja81R4YvUiK
auggsqfiGWtOb1ykmatbSwpnogTdoJ4Dmn94eOQGQ9ze1OTxbO2mMAdXEK1Ijjv4LsSSUg+YEMpo
JmRw72Rllwt242vTiGYsOTuYTuCZX8W9Q/O1BAOEL+Vpv6ewzRynPVEltimRWa/MWYZWvXmkIjFl
L8Z/hS94Gro2qHQcs19e/7/5WOtX4BDKzAoI4W+X++9NOietQO7AutMASs3RXtwzei5j3TfkrVAU
xD0hBJiHihG9b00qBPbnSrkhja5w22Sp8eWz98oGgQoy3AE+yf3T2mPwfOT0K5UVU9Oc7PLai8qi
uMIgaLRvA7L07olE1WqclZqp3FmubUZ/qXmWyQTyIFMNdeBCmzqfDx8pUqCjXGUN9g7zSP+vF4um
ZMo3Y1aJpH3e1n4YA9IXwvU2gmjNddz64sqyFfJSd/nHV/4hqBRRuA+34OtCrwt7s5Ph85f7hwt1
c527V3EBkrvjiTYS26+2IdHp7voecKrbD625SYXcqzyFBKcb1SN/JwWVN71BeNBsbVgCW6PSCuZD
PlysbFByWm++cWmNXN7ckLew0Gt4R3C88GLukMvvtTe+0sjA9cV88/hD52R92K0cV3DpPitwluvJ
0YplDjNRfvNGybFKuNF3b4h9hYmfOvV3eKprZds4KsWdXlj776JHvu3GnZwZFXY5w2DfOD08WIIO
UHHDDgWPXrfAqMaZfeHY/UdxgJ3M1Y8OUpgbYcfRM0T/KgM/aDq72O7303zf7ulYowlKcAZrA1cy
HFX1jcz0g359XLptWfsdKF2dKtaUXi8wdL8cpBxgl1gzJwpQFGBtMgHR4Hct8lqTrVyeEswS5+Ow
xhU69yb7L0w2WVkxAGW6VpZxJOiAl49aJtwrcOn0EIzX3AHwYTfVAfIRoFKYXwPqdBCykMvGgNWY
iyAzj2LoJhFKQv5F/YKisZnZJ7bxOaEyRaKsISwzHaSyogN/zE+SFobX6gr7OZbzCLF4bE+8RwJj
0dn+FeGjRUeiz621LP4cP/adZhqgX2ik7m6GiTsaQ+pUN7AL32EUN4XqOs/YktXeJuXgOwW50IZp
jKnpr+3/X11uP19ZyU4QKBaJrzDS4oAUvdN5yvBkqUOk16bpCzcYCvDY59yXWDo083U5k8a77K3w
UuL3GRAvE59xjGaWuvFTGQQjZWlitkbKSxwMIGm7oloAFe/GsS1d2nvosSbka3UptUyqcmsQQOr3
k7IE2DuohKqk4uXSBjQ5UUoGf2VFYkdSLEno5ClMvqKN+dYmLjBTx5KB2ZnuF7irUNLKCAGOC09i
ij4a4GYde5Xc6CY0b7Z/uiQJuSOUGAKjgMP2owgJ7LYizH5XbqbCJ9neYIkYUPT8tc5LOAwJrEms
yM7i1HPPTyHXKvIfIsu0xsTbx9sBb9spgjwtpwYI9S2TYehnbe/VOB4aT0zuJ+AX9XLy3F9mc5PB
KQMjJa9A+G4m5zjpnoTWQkYPQ+zhoW7sCHdVZWvvK3CukGJBmRqSic74kWtTSBIB9mMca1wSFyE5
3mQgfc6uYqD5QSEhd1giOfpPuT+bdQ6fUaVXTP6BJ5RdTMVG8gAr9JqxK0JxJGI2cZ/oZDl4d9C1
pXgOJqsXLdMLf9iRbix33B0Jz9NB9pIlu2qXZePxtVrGy4PV5WqPNlBptWIgwF4V9hVyqAaADRuX
ZQtkKYzQR3Eu7jFk4iI4rwrftTBM0bHB5xSXEbw6Dv7lYpjhsXDjiRFRk7wqbEz02wK43rCrCgEl
A7w2+Xv/S5YPOS0wdlLQUMhU3yDHadMbAZ43hggf2iJ/+HyKxPlJvUJvWRtfT0EJe0QwOKhYPqED
1RvjWHdzMHKnQzEK9/qoSnaesZZCVANxzz6+2jSdznWipCE4/w1LO+SUO7TO5gjM+ivYz1VJUGi9
uKir8SsTMFBI4c37WybI3I7cLZQoPnuEYiCIyI1qHmLdpjADjE/OlJi+BDih8SVGKr51F8Mq2ZJ/
qzNIvyWbvr6iCvgCACDDV/DPy9ainrGvxLoPe2ds2ryMuADsUrSXybZWpI8mCrtPv26ALDZCaOmy
ndmgYw7A7tbyDATm0/fbKluZ2PFStXHAAKB3ONGRqReHey50AHFrVhG3dyQrmVnvpeRazeIX7m9K
vrHhA+s4lEjIef9/Xuhz+RJcLoQl0wgbn3XJmAtfw6+uXPEz6cB8VmlXAmUg6Y2nYNxXl0AkKkpU
Okl+rSXonxAFyW24hzC8kb18/ap5ubt+VcbqXOfYDHBGxteKzU9W+a2w5yDIFrZ0hhBMJEIbImkV
N0f487459k+dsVpbf0ary5N6VuAKnX3mIaVj2QioOQ4CVzncko8Vmq6E55MdYY6G/2zDgGPWn73a
oYrUTNwQiD/iKh/gDYZWoOVLd3Hl/ZjJvky1DTZJUdCeAQYqS2X50Hgu9m5q97JWmFkNqIP74KzO
IjLC5bp9X3Y+RT56AsilIV1JY+/aKF6rPoCaOnMNwmtb4tsfE6ZEjh/S/TMqogBj6MprH0Cs2EIe
Qhb00I/5jAIGFLv0XlgqqQbH5tr4ZH5jdy3spSkdZESeFKNvR5H7stQq55SZgrgVCvlcR/yMoyVT
ntXOv9u++a5CaZ80SCFQ/bslGEG/k1VKtl2RfFbjf2tDMt0DerBErFU2mHbOGJsZjRmFn55r1OiL
F5UlDgxZkuPx4xgkt/cqptPV4mMrli8p1O6tSpXU9MR6BJKwmrWdWCvlXWLVYMPXOj++SULXbexG
Z4bhPgTrSC9vARZ7iJJ1okmXUWSh9N8WbydcuDjmqKYCmSxamc6pbJP2sQsWhmvilApR/LOdkx97
wSUV0w+TH1r1UmJomkLFUUb+UUt2VeXX2GtXtaTh1i6g4K3jH6iC76AdpVTl5+Bos3Vs3zJJgBgA
IQzdgXtS2D1NKM+7NNS8V6wExiLmRk10QFEYUCartTWJVSFgAyVEyMzlajBT2eozQLmoh1d0I4xX
t6ceUzQEhTOo2hEKdbGKSmgjkN8lI8AEBv47uxwthrCMFjh3fmZJPRj8olY++E73ZnNwk5JCgaKI
XbMSnRsEp68LSk9ATcotw/cHC7VkwBGknmTgO5dU8O0dKg+qBWL6Hpvnu+ELJ/xwWXdSch+2G6ED
VgbtbsO1bgQ/sp195IabqSlGtKQ4wvH4eYs2PuO/IuL/X5QOzWz3zJTd+vlyGYwJatbzdNVeNxIs
sSCLFNRFTb1RfW/L1wP0PINSapDefx6f+J+oPg89ZZPcnodvuOzmQrmUTPrUDCcs46BEUl29nh6V
aFfl0FsBsdJpE20UyhC/3co0jsF3f9uXftjJ2S3tG8Z8GkptpSmKxcaUOoxmHRFF5vrx2F0ad5ni
emHcZJVxpOYKbtLH5/6GtUeASxvipfHehY6YDGj28HEp4rLaz9cLLH/s5a1JPj+gl+r/KX9UIULW
NEWpn+DA4YnteTAGcJtnLziz5aX465DFRzK8TeKriW5IdIHbSVMwrVNPLIYrVFaiVcEEbFQ1A6FP
8CUSCeaRatF7QoASlOHfHfcRKiSNEA7RmC+Qos8QBXkIlItBYCArY7GypGT1DQlaCGR4u85dq7mc
TcQsZHiVmreH8bNdGeKpRofstn+X/jb5UZ1qnqFSn+aErZWJFUkefKydsZwe3qikdRLgFGbFCAkR
9zQ6gIIA5snxBy9CTfAqokNlki4BKXn1R19SbIbjbUlcKH0ixEXwj+8FkLQrlnfBhlYSBYzqSq88
fQ3lXRba2O+v1qQdQHN4U6Tk4G6v13b9m6QVOUb4aZ2GT0LNT9GqPZONTOYnQdlhCGxaB9ZyyHI4
gGmjRpS5rLCuchPF0BX/1v6Fw1p90LZYZ+zqkz/HnVGZ2ZRB04sWOtGMHdbM0jlQLzI8kI10/Csf
UYTFzNGZmKNcKGPKvgFLUzu0B4rDyHPKGz5/P1F4I31hO83SZGGMEj9vszxXWL5chp2hC1Czspai
qAj+EShPjd5kT1iepNVUt1B8j46nt/3Zgvdmwyselqu0nmxHFDVFjTyQSj4fh3xiirAUrwxH3+G1
t9u+BdMi7BdfR91CpqWYAd4ZG8WhIJkcXadT308azuMsvSPfXJjMNt3oN54qe0h9nqSSIBFwsxRN
ozbWj1ns0fGW4xgxo2wNjuNhcDug8bq50GtzgsrTUaDWK7A08EBdkEdiFyUw2cnQREq9dM3FclSg
U0eKBexQXTyXHlH59C/Wf0Q3SQM0MmuTlbFlkpzVFPoaIL3mrtFDhiA47W8rA0X09KH4p0TovfwB
CPd7/wlb1mXm7xdTEAAl09xPJReHqptaCjdqcjKeu3jHIEd6O6XalAbwJIhWW+4Q4sdj38UvY7Gj
nbhxYS6hDwlrbx6wL8JRwdBplHpKZaObQ1i07LFn94W9ffwoRNMImkU+Zodk5kQOCCWlhBZ/TNHs
lKOT1cgKk/EKiyUZWzLGxilXFYvSOFuThLqbydXfDaqtQIu8Up7c1qorVd8lnDAGAXe2MhatAo2D
xYWvq0pYyRFGWPklJqWGv4qKKmnV8mnDeM6+Q2qtGj6l5wSw8gMup4XaaP+XnK6NZ2oT4WUD2FMv
ZIl+/YqLgGld8fTEOGiPiysOM+I250MT4JCHyn2FT+M4ygJUDGLFi/gV0zrsBls1kFpq8PLuw+RV
B+W6agmIOO1BNWpY3dJFXPiCtuHb3Wsm4oK5M0MjEBl0/T5m1pfhxhxy3IOtDojXAks599ck1Kva
+ySCmDbFZKjYh/y4o99Rofx3Zr7+tC4APlGWLARUQ1cM5IE9hc+9ZYmKtbExRpp8W35wb3rmUht1
kzsKHLhW25gppnW/D14ZbTzQVN0hHchSSaWm5IQoPzzJ7LLIEBvOA3uyHRmlKAjFV+DddlFWrAYm
sNYVRuC5Dq0kaTe3G+0KlImx7EAclpHImaKvpmXpAN6vwV85s2vrk6IxCqGfxc69AWZnEAkrUVrd
rENN1+/hhrbuYf6GEuFPVFoRWaknKPHUdrSeYRO1Hz1q4K8UJlMe5vn8Vuk3wBprajLxxWWpi+z8
HHGaJognNZH2uhAqp9Ycgj9/tD0Of4r6qr5GhSn1v581qg5kgfFEnv9X2/rURICrYuuUfyXaNJoO
05xukecCpwQVs6d98x+H5JwjTioUEyRfJbjyXlbpFMcOBs7e6Jdwx6IbD0L1PE+sfUtT5cD7EqYO
W2tBsJ/c+iZ33/b8lS/9IXz4n1HC5V1YX+fIR8wW/EH80Rq7vU5UCwcC59MWlO6ERcQN+7Pknufl
dIyDS4F1n3wbgpLFAlpkSccfkoEWafgwETAov+io34vMG+yrdoSAx2OZun/d2FRhTKD17smK6oc2
RPf1vDR2ujOQ9RkD6g6l2toqahu97Q60dvmeXYZQKTE3cAy9ySbtpqZLpDCYTTFiKDpZqWJ21lbD
gdRHDH2gUg9F4PDvBCja6jeF7pMsU4Sn2EQwT5tZwPoyCEnFaUXULAsr1+8la+n43DdXphXiUiM0
HAZAJMa1nlMmj07xUISDty0K2DFL2WmA6SkdVZ8Z3xOhzN6NlcN0cTFXh85baSF1yWBxLChn0dko
diT3O4GIi5nU7Rduv/icbba4OCfA51GVQRjjY5BXVhEUBVaB39wrlg2OVdZPiLhkmHv9s30+LPyE
lzH+25CCPPqGXomBMOPlV+4VuXKJ2+XKtDHbNwVHluuBf6B0mkW0LG1Iq7WokO2Xhns/axemlcfg
t2CbnucMMG3oB6q0jsjF/fsriWxvImsFb0yj1VadQHcEwyktFmd1gjJkzPhjIDTjHeC2Y5QvNNih
Y4FSXCeCeVQ+K0NZh3jDxT3AYjmHcqu/foQDAeO2kIwG4fe4/WOjjCcnH+vjCoMEb0BoQQJIOs0O
WOCcJ7xCt3VpJQrcByrdiZbbKOkB4HoayPMTh1HdLcKTKDQgalUN6QFN6ETTZLdkiVirC/3aavHm
l9nQT/DShNIwqFQ1Fh+LEgVnmCdYG03DBWCmk4Wtr5M6/k6QHIU2+1cDjlCcANZHnJ+OEWFeDaHJ
xL8tjucy/CPy8t7/uliE4YPoAS2ByM05LqnetbFvGW3SEyw4D5UPMaCENAMKE/iMS5A7KJUFqL9M
Nm8y5tc9nwRNkalk0jkYOnJES4SDJslMzicFWZAYezw8ohFHlJPpwn2HNVk1PumsD1kcaQ/pYjrx
I2tBXPM0Q4oBN6q4pIKmHzAuGCeJlihyBANVohrft+CEZZGIndsyQBjTsgLkYfkuN1RS3XQdj/ZM
LCjqboyIj3uom9XZuoMijZ2/LxNtjMoeswq/vbdm8w6DALxDPLeAqV+MMmH9EgrDaoAXeWDlKoK/
qX2zS4qfZxFDNIJ4bWHCLtdn/OtqR+VG2AyNUd+KjJ4hPoP6MX+5aoiUgs6S/J23M/moCB6Ad+ZM
DHJWZUqaozrVxwyUQPD/pULU/VTkN+QuR9J4MGnPrNinUSoh12oD1nHjktHbglAzuK22auCXcZEF
ntGmN5mta4TUeYVG/6EXKUbceu0/i5cUFOO+CC8+MQSwtJAmr3AHz/K/UB5SZpUyJUw9EXCUcyTd
uhP0bIN7gIaDlnUq6WOpjmI8Q+igmIp6jhh77jHKYZtXrPzpnRjbiglhdXQC97Auc6z/xV/pP+x0
LYErSUoTvrfcojEmgDVPWs97z9CyKmgfFhc8OQIreS8fGHJqlS3jnVGBoce7aYtWWfTlrwe69FNf
ugZGgQgIsNTxh4CAJd8rTbGwDgRPa5DHUB34FXY0lcNqPOUUEgEqESVgUcYV48Cr2XYi0w3DsjN+
TzxkFHjsv+30kR9mtK/MM5RfrzpOx71bxkRFK50mcu0ACYhBmIWtYS2BHNwpaj+02XiH3/ebWHGM
t+fjWUfo9TI/YyKZTfKKyl5jEYlsuB+0vYL+nXDtNa7XL8BhUfmir5ZLbznqfg7+bqBPcq9uuFK4
WkO2VyaQUzreov6fzGksxu9ChxlbZydMz6KxgkpW0lXaBpQESzvR1/qERWbehV3WiHAQuN6KSdOZ
nUyRca9nr1gDhiBEhUjPRaGkO4r2PJKwNeuInrIcbIbOk+OG6B4a3iAgfQEPUs2TXKVNyg0ze86H
K/hCNcp86ss5egnIUrnOIcu41HQR6CKmBVRtSJvE0oeMqFcMzRTc1hhgpsQxM3QiS+8wDxalC8Ol
i0FNuVo0zDkdZ/tiPbRu75OE39ezi1YDOmsqMCs2DuKZFQWHYfCdB418f2lItb35jfS8Zov0uZfI
74M+jbT3dh5WgfDnumigN+I2mnj41m+7f24qBPTly1laZPtHCdzI7IQKVvUflWiZ1OXqxA909aca
2cghj5GP0ubude2THTADUqNWuNsX1cLRhDEqd9pAQ4ITrmvRnDewWW3c2JHp2CfV7FcP4JMfWgvV
3xIy02wpwH+WJ7XbAqJxw15A5jZxVRzEMUBXQ0htPuTcmbKyq9jBy573q8DHug4ISaseD2+X93M/
X9cYhJMKPDtimS4MMDHKlGAiOu854caIlRDuuh3OBMYJ5EwAZo7TlMHSvlI+kBqXFuUi3lYmFTg4
kYJHcrrUAhHIeSqNcZp7iZbTXoIpGcl5G+lkAL2PEDz2RyZ986HpESnoYkmA0oR9FAbmvFegJOC6
gux47QJ2BBi++xdFHzi+0LBL7QG09274p3g1Hq3BAN7kZnG+NZ1/gx7sWPluY5kkrTGgFErN/mnt
zXa4r+LHLgl8SDceM6fPhFpmFTKBfcEW4JkenjLuLVqyDW9fJ/C4LxEl0vGRoIOcZS74cWxMRJnD
KRQcf2+kxeQQ2XScl8Y3/4c+HNsuta6CcpqjQ+a7jAEV377fQplmrDomzNPG6yBa6Pu87X5pON8T
DixPuPeSkuCfnWtPjOTUtjvRn+EnygIn3vB3Ufz4Me1bF1WLZ+o/8H2OKwSFCXAjFU1WZnH/CqlD
GVcoLtS9hRUWoKyWxlDRAZF9q7hOp139MYlB6AedjUebnp/WF8JH3z5dwvw43TTYZoaMd8sdQjr+
6r9KI7bB81UrMHENsksadspGlhmH53mg6VWg8/SXzBUIcHaNykxI1VhCT5IRTganhh4LZZezbUAB
uj+f/HlG/kK+l+KtqqqNZYPihve2CzlLZnWJZzky30Is5gihFh8SMyJgt3O5hk1EZM1lmo1R4zyS
nozMvljDHIToag/8E/tNw6VSTOT+VAEfWY8bZl0SXN2m60fTgHQ+U0bA1h9eL4+IIJfxY0DHXVXf
dPmbdNroDOD7J2bGCDNiWDW8cZYgxknV7mq3CQHUwiBt2uIP63+euQnpHhQh8w9jjn3vgEjALUF7
h7OR75H2orWGqpxNHTNJngPUn/0eBKgPv7qyHNN6WJEkjspPmuM2vKt0BNnS9xr6RafvCmdKFF0W
7Vc2xNSB3Yqzii1ktMJ7q6sQoNG4amSqzjEoZyyjqxE9TXS1wAtCBm+FPl4AeqlactBXgmbIpktL
vZKobgaLOfFA/UpJYh6hGiH+vlEpfcPVPC3ERMKa6PDCmX2mr/7ee0HbJS5t+f7sizZJ0pu4xbFt
nN0P/7ARXzM4+C6qeZ975VqafR0pryQ5kkV0eLh0/HkOKyQdxtKtqsnVkXnV3VZHR3jJtUbot4C/
sAs42DU4JO4jCFbAslqQggln2ziBwZlDUM/DRh9YfGWocJ1/Ej6B4zjPJEhUsf0rrJ+8y8xLo9lv
pR3Njq3LLPJ7bRMZna9BjS/E4brBysgER+mz1rzhX+QV69YT6aL4nGxB9YL1k853jbUr08BmqQOe
dyrM7Q/GcjAybWAzPd2HCFd3RVabkVN0IhMsxgbonDjukE+Ogf1gsMBTYa3oDfyuL8YuTSFq47A3
S/qrNf01a0oUQuMlzhtFjmaBoorruCup30ntV8L4sWGSjgqFFzMasPJnzJfUIPpUNc7BrN1Pk/6c
WejsZAtaqe7EmtSPGU6NzPQ3WQ5fUU6RJ0Nu6CEgASRYvhi7gz/tvcWlyFItplCFDqIq1Cz7akQn
RmGmZBR4NABNzfFO7B1vIRlRD9+xD/EakEdsQkoZvVvZco4pLFhkr5Rqu3NoYpRT4sKuiXah9Kx7
7Z6aBZGoyjuLJIX0lZlY/sNkNxEEbs9xD6xSY3xIUpqkBjBxNQZr3bM5uf1w7YkEEh8O2uwFXsh2
dwwggQRV8EznESB/03jZw5eDHu0ViHzwI50fcIZc85uJcjpCp1Zn/zy9k7fnhffNwseYRmsEi6iL
B4GLxT1L4/QTIBJEM1P88ZpmJGvTMQbB+6+mprDkGmXmryQ/Mey2qLGUn4wx3MY0CzU4oBggV27O
BhdfukHGhy+8mnWn5cHb6AcsxByS3dop70XqpDqtufV8Yn9jOyMtAQoJwJgYrKf01n0wZAgl93FN
kl0rhixfNhKtidE7wvNBm8svVPPUlPLVPlYXb5v59gbH3VaaeO/kTvLbBOQxRPsR5JCUWVR1llzA
EIrigoE257q0gfQUVFe1jBKZPZiXekxc6hI2r8j9A3Fb31YmcUVbj90KjCatedXMCbfj/LfynL1/
JcrilgWeSKMY7RDnL+T0kdVkLYLBBureA3/Ko64n3SPQf3wALPyjHESHOh4rfAjt6xXka7Rs4jcS
XSRv99Foqia35rKXaql69t6XUuTpjAOAO4bvkdlZbU2L/u7womwVxOp3hgceFbHzy7gytWD3WVzc
zdETtabswcKFS2RFfXGaf70pQMdevFpyFVm7s0oXUqIqRP9Vo6N0d9ygWS7Ey3HIBX456yXQBn7H
dsMeSc3LTAa6wI7KZO7ezCCGSStedxxwRLEZUg48SwYrHGhNlpYFAVcDhvPhcXgeNF5QzXhbsBs5
MLufVAHkmoQvCEOYUVfkAE397Ll1I5NJkn2I2JTM6UTtVPpMB+ODnbSiKD/UOIew7uZgB4CYB3WH
lD9qtrwWeCt7f19HBUzJWSdGJWBtyZLCHjYWW549DhHdT3V/o4yZJ4x2WXNk572wDLsNd6gSXxc/
HCxakVtQoJEiPs1DqlMoxgTEw2IByiS+yd1gZ2M24QjWc8VPpLGFgM67dQVXMKyOzn2T45CMeDPz
80ZRJApwY+P5AIQNz0iVfhkTY4/E7wiozKcMT2XacTxP78rk6SUNR9Yu51ZVowRecWBtjllbAFkW
7B+w0pgH8Fimym8IxDPgVucsqQabqDQTsoZxNrfcXW2voYslfaWSQLdCMICqRbtLKDr9twpcMTbb
q5EEOCs7LD/5jB8sKnSCn+M0QLDjqY3JQ/CM5E/see+2773kS5TScqXbFfbFo7PI1BOJ0mDv7LcY
vIsydFY7PIEE4VaSzRFkHOmideNw4c5390aVW5z3TxJ5XXv9DQ/+4cTzWlNg3i7ZBDw5Vt9OyK1c
WaVAGHRjJVfVlGBwDmpESrqxwXG7SU7BJuYw6HDP22w+Skwes3Q+SsBeFRSUQR0L5Crw4HmiVPij
dIaLjedtQF0nF75UcKkkTGxOGTtxmqPxhMevDzyc+1iSodk7jTjLLK6lryovSjUdVJ+LpRt6jBdz
PZLE96KIaikGH7xWVNynN3u1/wwX9mWbhI11hR6+axCUHvuXAJl2vJ1sRWqAxE/Wd+34qznhCF1k
dOHrJ8M76AN+3pCGRFHGi1DGjwujkjhIW9dqXbI+I4kDFPbfdodohe7alc3FgWe3dNIKt/b5baoD
8SteSsAB8ag2cpe3feF+fj+6SZnEn+nPbZjbO90uUDIeIwdvYpj+edPXMnqlMq/xD3p9rIAyJ9RU
dpGSnGfCFjSo6htUBB2CFQT8/PBpJ/NRvjg3knBrh3PclOkFTQXD1sR5eTwhLsm4A6iI7Gd9CNt+
Irra9BsTv+/0mkLNdxL7oXGgrwp+GTvMA4AQD0DGjMI+5ynYy8t4ytdZ8aznGXEODHIwiIh82Lnc
OOlZJF6lpcGpWF+Jd1c0qora7nAHkswIIuxa9IelGbSlPUBo2kIsN6mgNE9Y9mgmvAyP8GDXhsKd
2Dw7PuPLWjEu21RxRqE6tgShwe8wTDHezd+95yqE/7qCQZUQ+38c/IDhxwtFmlV3EDTlTozH0TEd
B9VDOvVKX4VTnVxffMfDjk53DNAUg5Hm89mKbGodvyuttd2zQJkJnT2YsRoGlOv3xDJWpQpVNWyh
5tQ73mAz64M8M0jFjtdunwgchuwoyxwxCuUSpb6JBQ7bsOJW0fyNVIp1Z2Dd89qjP1EN3NDDNTWi
Ix0eG0t3mg0Js5TInB9AE9+YHePJqHG5LOin2b5BIeyokkyyl/K2hQ5go1rJxALtDI4Klan4dxDN
Y4uElB4lDrJuUlE2M62cxgfLxplHzanSXAapn4W3KUAWlI2+kjKEdoymwnkiL38NyFXl9d/weBon
Skk2eaczJ5f1Ecq35h302ydo73eRBovJNLcxuEpo68w+5Jg9wdzT5H4MpjHlHex6OTnvuQUF0g8q
mwbtg27ElqLTyh/dWBsTrhTbGpHhnpV8jrIpU2hxQWfytK5Yvn9/rny5qDkYcTTNq/9HyB7PWtSG
azGq5V+VVwH+OTBL9f4BYWRCxT6x8FK+0el9GbGETQOPBUY9r4/r7VfI8sPXzELIrZ8CjOV+B//+
7hal/4DlBHJi9bKcgE07g8brPs42OuQcjnkKfDE9C6VWhmsnc0zewW3Z58aQmvEhZoJBwsqBX4P5
ZcoLzoaMsPYbpnb64HgkhGWeVvmsEX0edFQ3RpWMbJ5ju82XTQLiXtip9jRd7Wfo2TMYrYNfZsBB
Hy1yS3O0Z9+kMHfPZVXlnwBxzyt4IwDxuymYiEsp72XvY1t2s4Q1XXTXYFASqY37RdssnBMp+yOA
Bh3Cwyk6tyK3jckDycGPWVHQXG4uftUuAFgZNZ5uGfDnWN5qQRnh4lFEikm3k+VRK/hZmLpBsnYZ
z1TQ9nryKoH+dhqbd69hw8/6xkvA+Ir5w2a7U0mCkXH9Oj1FsTVvyArmtv/NBJALVG6XwNS2ALu/
rtb0UKCOMxxrIeclmv3aF7HAfU+0nxeF89pDaeojjOmh0xY7n5eFH5SKe/5HOtpgnop2aF5kchbC
N3HK3i/T0yNpaIXtp0ugug3AN54hOWjyUMUiY3gPq2hN8jEQQ4ppb2fsVI/I/Frnl/tTIg3w3dvw
3M4RZCyDcIXuuKNGjKFnG5miYnl9xrzhjzKcXaOrJzGNYhaNT0HFsMZEp2ZgnXGBSC7wAqslbd/K
8fePXfkPipfquM9QfUYpjS/W4RNL42Kwxw5C4w5jiM6XZ8rjw77G0qO/DaAMGmurOry2k1AWWIYK
RrC/KDbNjlL9dh0E+2JlOTqEMBC+ViX9brLRfRRbcd7818QyW37+jarrNh76QhYdPe/wIzerXzLV
G8Ndzc6A/hkc77Gb9BeLeqESRYmJcSG4hNmWeRJ9MM04dmj/u3zagt+O5MW0FX54bzOA9z0CqSwJ
DsznN+JbpwfiPft4alb/vTzju6cmHOJWW+5yEdSUyg5D5cdN8J2So+086Q1td2F49P9h8zHWaT/O
gvZSnUJmjPK3aCIIoZw0lXolruK6vrzDJZDOvt6ldPz8IkRwiynl4LcrDh2FCLefijv6A9VGLgk7
/bpFnhQO+SrrPgQW1adbRY5DKwinfSedUGE+8b+LrGGlEcizpKloh3faOLfCqKy3UF7UPxcePYMk
JBZgZSWOJ+ZnFF1Xb+oegStxfCf9fX5RvHCrLAir2bMFD3zMOoQ7nraDTXQlQy90Og9D1R2SlHgq
JWCqkyCi/mobqHx61/V9oCPMmOPH0j31fcHaWvNAlCISVbP5cZHymq47itz7pggelho6GBETA5uK
ckNkNPjv5IYixOkILVzK+sFOZoUAOMiZsQbpPUoRTIIIyWGqx6dzZviIbL+1rxAjsKMKoJpjiz3e
rAsDtJLTD56am0pxpjX68lo3PoQubmKKhMglWg7KLm9rLM0k4iJ1j+NhBHCFynX7POyN5X6PC5S5
na/7/A4cpxntt2/y61uJflsSpw6ehh9EKfRe/S2LoTX/Z/QzldeTGfnB+qd/RQHpN/ORwrUw3pfc
BQ78YKdBUO/3nivvugqPgbfBdr9qCmTriW2Xe7naI2S2AWUaMjaikT7oe8y7ssac9ToSIagqJcyO
1z+eH8g5dBrSa/YiUAPTJj6bi4M4UkBkbuyZQYctdbcn3+Sc7HjpawjvOU2zB/6b4YUpXU8xbe82
hybDNvsoeONrGCKEOOS/tsZRcE+ctzMcBRfDYM2To7asaSxqY6jwjDbGKBqQH5RQVS+Ru4f7rW4P
oHUnoNXEWQLk30Eif/YqXYp2tCOxtIF4t7vLuma0YVgyCZM0pdeSONU8Djt7CG2cO1oR8t1/DxzE
ueuN59oSsuLDbOyOdxQfMP4veYQ2oRHtb/9yA/gXTpAP1AFFSIHao+YfA2k13zfFWY/Pvnmt+STh
Duy1WuuhtGl5CWo3SKIw2t1SRR3ZQKmOIp6l39FOmsErnOpbaBLVgqALNhvvjnLmukhH8IIdNotT
xcCzLtvzQdI4QkWrVmbiZpBCbmgifUU9zF5dEUiM187uvtkHqLD6Jt7yhR+YkNJmi9h8BfEmvQHg
ocKACcBTEIk8HAgH+DdWch4uYWBCkDb160sVRj4xsYhYZYIPSXUwZuWsmjNgFNbYkQbhqPJTowCz
/q145dvoxMZsbRM5O6WQCnfE9jtBt3GoVOoh6ICNSzOlZJs9JLUimDDh4U0dqk0BX4ADelstlS1Y
IS8Yk/qzCsChngbjEpwu/2tQYmJzHhp0vlxj4yko4vnPdARdD9nhFpKwS0g6Bep1p314XKgwRvce
PZNTdro/E57diJjMhS/t2X6uk6stKbLHUYQ8N+JcVELEL6I1i8Lxa+luiL2j+fiQOJ43s0A9/3y0
dQQ/lVs2W735DM3bo3OeS8k0JmFUTFPHxvmuFU6wKZR/Nt1OFSYKjjNhjwKZ6xGViX9tKqx20ZwX
qkc9YeLvoU/5dP1rRHMCRkg3jf+L4rmFWjC/yhrkrJ/hvOp60s2BKLu8xQiHtW56qEqyBAvZme4S
02O+GU2j9Fvbqi6d+flqQhtQLjJZTLEkXrFYROzX0pW1i0WuCe5OX0rzKn7fdaHJ3Z7mPl9d4rcN
zaStniTGih+MXGDlczvHXEoJf0ZRBvIbKTrQVpWVs5vQof5GMnuaA12riV95XdyIUOlTZpjzGxEO
7yP0sNdMbEib9B7AFbJC+GaMbsEQ2hoTqkVV4flqGBAePt9qxMphbaxf6hG9A7cxK3zjPBiVjnBy
ll5m4f0dZkdI4yCLPRxswKa2esa5zbIsF0ZyIIn7Tg3jtcgutfCTCjLn1IAAh8utflIrk0MmAIiX
sgXoMHw8K4qfpjvGqaRhMKyeVmow2fo6rkZ9yLc4G9DBFs7W0T0ZAQlLxdqupeh3jQINp2EVQWUB
WkzvnLoV4JJv2Xozb7hkmZP/nMfbkoXbNKyQ+vC7gN2Zx2PfAaxO4AyQ8YljjGQJ788IZdEOuo7M
90APsW2+ndSBiAwGpAoRrF0DdEwwwGDPDstVoMxY2OgPshFb/HXhPx4v8RVWH3WENOxn/Rh0UBrI
Njspc4IhLitqZVh8MO8GO1Gs9absCRj3q72Zpyvp6ZDJ8AqSZLN9DzpEs0+BLd+ixeB9mkmaGkPX
laZlaChMjtY5RHHjgIIArlHxVm/8Xna+0TaxI2dHm+K79GKcS2F0lkOkRuJRBWWr0z2RHJXT2H4g
v6gslkqp9rxqL6dalSg4t6Nz4AyGY0Or6HcAK/Rfx0wcWwU3y3SaucNZJs4wJBcUtV+HGQhS+O7m
pOuYupBoRxq8bQze8AaobVO2mnIDAdJbUCSBT2Nbj6nj48EiYe0ULqikIe1oC02WUQkO5yfC+UHH
NZSlQXxneUyxINq+//u8FJNEjsh4vZBYtJKOKeT/wjRVr02ht8+A4nLz+Wl5ZYAdpMAv7mK/dBQ3
lSoTVUI2s/sIzfKdnZkgg/14q4dHnFD646m6Ey9kTM68s+C+ZW/6h1zRL+d07O9QUuAph4ToFTTW
Oyi438JbvmGF7zp4Y1IF4wS7P0dffAZCadXndGaISYKG1YfD9W8XhcLwD397VQ2J6dF45Oz2xvwF
q/w/YLz2kBzk2kfKEgEDLUsBQlysSd83edMveQsZMnDv/4U4iGDMTE/AIsAiniLRLFJ5EXrtjl3n
6sjlk0noTXtEBFwvfpZYWp0/z0e+g9YPeKUrb6kLgxc+peVqryBIGcdzAjvZkRt00K3tIoBOOar4
n1aG4UsEo5/S5W/JxI6suK6lDolWVdG7291EDRtCIHqFNicsjdFxN294Q/4IAoQ4Vzbkl5uu9Zh5
zUqeKbwdDEFpNAvMyy9yNfULcjwsVWrfT84msQsfjQM3HjIF1yNS6VcmZCErvQQOc0oWdHC3A8b6
d4MsHDYS0LfWM/fp3DztnVxnnaCaXhLMeF66IaFC2qpTy0qNPhYKxgwXNT5aCPlB/ovhDiMrgXYA
QW9bz2KJUhg7BI29RmGeG8X3SU5x6k5gku6nJ+W3hV1gy35e0U+dyvA4SJwn2gI2DlN8+eqKrdW6
WnsdxiAt2HPuroplQNkEyfQb3uMT5yOYbPw2/wowP+P+7THnL5r23f9L5/aDWJZNLnAug6u7TnWH
CKP//FOfn7peEWjDth0Iwevh+YK/yhtoF1DWnUA6+yQMiSLGtRt9wVCZt+FOL8CC7UTqeDtXH3pI
YTd0HnutrkbDs28GmLHG7r6GpSOdg2OqyXKlZz+FL4bGN8vj5/fhYlwUtTjNonEoJ4PpoCrr1ipw
Ou/Td4fOjU8cMWOVFdGpcDZiI4d0Z2KoFiJ8KY9gHpe1vXStSKViDd8KYKUWLfkJbn5dGi17mw/K
51hclVmiHefcSFFN3e+TonvLMT/Uh+f3Qe+j8IcpKoaOQ2HflbQ1wPFGrCQ3kno6s/2qPjxMjIro
FgC3QCQ+tAPs3wmt1iZkhTIOeZZ5N5E/6uja3NVt3lEG3LPCNtRlNTgkVi8Ks7QfC0zRpgIFYADm
XnPQ4jkkNZl6mMte80AsU8Lp8794+hsDkw1LGC7Ox+2J3TGO8uHCq5didanciO03eIcV+ImmOL3x
VaPbJuge1lbAYBHybu/oYYX8lOgwE7UQhBoIJ1Gu8YzHCtvUpNtTkdagIL365mxv6aCsXZXy7NKb
QhkZaNtoAQHtUCcz6VLOZ+HcTTBMeogBanzmlOLLFTkwahqI5LTjCk4U45q+5NFVUfLEZJEqQLXs
OFQekE6/8VryaV6BEnR6lisUkcCKxfEFKNIFxXciq5+V4ck80nDOTtwLWuHs0KHwTVP2Vm2UcjtL
rTWiNhN1Gihus+3HxcrxeSG2fAe9XrVUkYAugFWz5F5FiLzu3crlKIUmnTUsbsSSxxw7fWMjGN5/
6gR5dVeygtIGBUcu/zLZyJCAfIEINrbG+U1UXUfddl9gUuOFTYcwFLC86qky/jVYrCBNXECyYK2c
w9gNKe5HzQwvnX3/R9rXVpSyN0iHITAkgr/CLWmvjAGaGSi4Z5E7E1cCPE3igPn0Z2/tB7e/u0yL
fZM1CNTvpcCI3V43Aid7Yy2F9M6UM1DXrgVZUIXFmLlZ8Oc2NDJ7ue3VypkzoLgEu27j6r0IrOj+
xyDsoq9U91kYCZFdFpFgS3+uzSpuiknRCWGcTQsof7WlIkkhqFG8PXwc9qHI9bFkfNyKtRZBMOhS
2SpnlUfJDLvq2Qn/p/ZkwgHQt81RC47TeqsvLu6VCmtzvmJhb4q+kOELCqdefWbaTnk/QtaYvHhB
1pwCpMtYdjt95w4OuicPIRKmuboXmZeoLUZ6AvHMpZCIGmi8rKccqJZiaUFTh9ylsmSqTPkB+ExL
jwJW8Assw4Swr2um0g4b5NSkSxjC/pB1wvQGRTGoA9cdBXAFSzoevNgxAkDz5d2xjB731b/A5Hqb
+0c3TciloeNgHizmow9vtyenD7LVcz4lJpny3D8hOZ1rZFXqyatvQ9dSpnRw718X0r5r1g9dZS5p
zse5eIPCtW5ZTGB1jUord2iQj00yUAbsdrigrhjCXvdUCguDaha1uzJ8FQULekYb8RlfVFfFb2bz
7q9EbTFUNoULGxl254Qc4T9K1g3TcaCfpbdVU/3HHOqk/tZfi7J9Au8eDfI5BMPEd+zXype4nB8A
/R36UIuyWBPG+7P6nh4qo/0ubBnyJjhUn/Ws0ESg6b0NbzP0sXEvq+jhI4FGn0PAepG9L9ocsqK9
zBNyDPcVd9zom7gPCtfuW8LjgsEt8ylW5p/gOScVShVDNOu0Q0XXJO2coZ2/Lk0hLB30DU7fkHEh
nK3pCFb9Jjv3q+t53BFYSsttUhB4FhpKNhF7AVr6b2Gm9AF6dCls3SJYMsBfSk70VL0kObQAUZAC
j+YRsTiGlHTQ0ufEwTrF3CBZ75BLuUzTjwTR35oxSlaPehLbC/WExYBI39+IlCXptantH8ktzkrV
NNfnpuM2OAoTi0AoelwBvwOsu80DaneJy8WoF39h6WzenvT60nx1p5D5MHhvD7wWaMuG5IEDrpQt
/3JlYCXstDwhSxE0HViCrnNu4jTJUTT+SNgWzn1sMDfq+GFiOmGb2jj3dtmNX5S2SU32qxTrRQGC
WWopo5oEQ6WUpliS+xuONi7vugzr7xSFmXIk8UQoRAUlL5H3bVa2s+XZyEm91DIS+RbyZhA3VjQj
vbu9Am5PoMeuQkriQLifu9MJ3S0ia5mKSGHA0vazCyupPttU9f+eWhryb7UpvvEDFZsVGrZvfBZR
O9Q7EKvo4CTeq+OoPSahVjpB2TpWQTjS9P2pl/p0nn9EpNTX94f7h3GnlUsXyTNMoXidnyJl2J2B
7oHgoOIMC+Ol7rq6/uH9zOVCSZxgtAwJZmFoPy8Mid5npFe1HFiUX1se4vydbXTZQkb94dmDPIN0
+fsDQaunqe7/ZY480fHlezSGNeDC1oPfT3A6lwax5/6Vv+mflwpjZy59hh9Ju3nuRKLrwNdJhM7X
7t1e4/+pHsVLzh7baJEsgNm/jXPUkn7Ve1gydMgYxH+Yrv2TDtir0eXkCo6EAjnazAIViHpAgFkH
yxUwSgzZ8SgvNrG1A36m95PRMPXBRsYZO9e5iRu3fJ2jDqc4IZ4ZqdHEL5B3aOnKmttiAqlHrUdh
vjjQYLq4XfU5hN2K7kE/afoRgDp6U3VhtvFhFYu1/EVjXANsruuxwtoFcUJrxLlfxwEWAJaMo+rc
utYDOknoSrBVutCdVPdDkjgamhWUyLuskrKiuJNsqcFi1m7hrYEy8OVkGdnjXIUAEaJapiCGX5VF
clEQVJEdhKNRAjaDneCHiwO0/fuI+jLFZSSrs8PfEU7BwDJM/H7EP2G/KLpW4DYkfGlNXHOf7k4K
zjzrSb+i0bCC4pVNfMwS1/Spz6iwIe6vP78sSWRdRpS/YkiMvA5fxPygfAK5Ydk1PGc0MJ0fvvgU
Bs/rnZ/3593cLN32T6AcdSADQkMRpZea6XnqPZcrMnClnQ3KMrens70PWL6YqCBbXNp6qoCREN9e
iOPbQv77xhQaTCYAOkG6gVqH7lHH5Rj7nsHMa/a+9JjkYdNRKM6QFzi0JBWwIrQBM6HgRPq3yakb
PmX5STQuYLTZCn2G3q74OvEEwjdTMgn+c4WbXuS4fezth+tbNfZaxH7v9rKm4EBlDKSRcddZ1FbH
FhgiwhrxZ7LkJQ4/yOzNEzN/R+Zja17uvh3X/JpyuNohQlHPnlYg2QeDqya5AJ7SxbviEzenlSI0
cS1BxOuoB4uJDojnACJJNf0x+VaVfy8QO0CW/dKR4sZLuD4WskWM9RWsbBamgN0XLq55oRaKiulT
HXR9ukUu0xr8uuxIo6JfJ4R4Z6uJNxgtsab0HM/H9G2c8ZQNzQMqSG/pdZ+ZmA5yjwOqmXT5O3KJ
b7cJxnmXiJcAPAGk19J5I4DEqbfx+31GawcRxsnFFawkdHRr9gtw9zxvj/kkWsVJJeV+4sLBz0La
JWUP8mXSJoMgE5TSweKF9YSpeOqFpULutmqvqVNY4pB77TPUzE1maz+B+bNyl0UeVWEgZMNU5jaT
l5JUWvuv5ubfOBcqcRnGihaQg/LcJygq23+6Gsjm6jwbbgQuEoJcyQjAxm8iB9ST+600XRK+e9Fu
QVImgcL1RYx7RwAiyn0lkZOntCW5MlS9PV6tkRHEACTAHwP9KRzPRBgOx2D6+YhUMs/1RtrMQu/S
KxzXLHTmGPdfdR50IJhouKaNQVmqDhuVEG1RwV9BO72j5VgcFP4okHJiEuG0fei5QuQdUPWBtQnh
60lGTqmYB495Zz9fW0n6fHG+PnG2BU/2h/OeuaRK7IL2YuYOGQKDdFbvJzGR4xkJ1Csjqbp4WugC
ZJ/0oYd6iuWCiM/t5hNdvVlziOpf6yPSwBWxV7JxRdLlZwHFt5nreEsmVXA7Y77gp6DJ0ddE1vEh
b1TzqaYj3KfesW92B+2sjFVB+0NtYkEjxkdZNx/SxroJyYlb34p2eWBOFRC7Zgj7fpzxTtwbmFhV
wppSUJOOUF9OiBh46VkXopjfsGYPJsY/I1ajm/4NtsVNBSAthUjYIpEILWmxNhTHIsBV9eT3yPD+
LaOTVV+1QigP4kRGkIsD6zxJw4SpVVXoSunEzX/Todpy7ltyDaPsVX9RZCdW7FvGW3R2o0zjYo6T
yTREvxmAakA+KBFSwP7u1MIpBaDnb4zq9jj7AGJnns/m66yxUqiOfDQ71DYivDlP2Ed5zOgP6ccD
qaGzqlftQB42lN3LzNamXzmIBQbs6pdcwTmZBmpUor1p4xeVo5w2aL+iGzlLnJ7Qm6czoV/9pZ0c
x+grp3aXF5OU0mXaekJjWxV5GQlZEShYq8g0HgBXXrtkL7eTUdfU413cePmTVqry3xrtbW5pBD/C
5LqX1A5vNZUHZcojR+6Q6n2n/eVaK0+hCUeUBAFreAmhH0Tmz6h3xarGJW9Ef5+C4e1lVs9obSSm
iwMMT93D8hZYsBCM8Um2shvgM1e9dPyK5xWP8pqQ/MeTVtVQwCWG4VY7S2FqXJyd9PVAg1Vv4vQQ
cK85zSK41JzMx7UpRl48iJw8QNg6U7P652wNsNKFkYV2g/kE6XQQYWuGoDMLd4fOJwG8n8IrNaj1
1RK06wlRBsfamLzqebE4mipK1UwBhqS5pcz8KOiADrVn/KbB2R6sYbzAplgaOVYz4sSOuzgo+/ha
V5cxa86LVR7IlU6AfEzBhD+aP8+Zf6KBzS6GnBToUQyTnjrRJ1KaGgXeg5duASZV6Kq9ULohIzlj
BwQjwv/Mz2IMpl24whqccHqfnH7zIgLUvL/l8slGFEuO4MHCAXz5t3RbMbd8gqqMopqk3qMCwLAl
fyr1HcYGjFWsjnE1xVxouawBfi1o16tHy1Y/tNQag6OrKQ73ujE6qMYVgRMYsFIaryi2fG+qTHPf
0dCL8NHtGv+qDNqB71vCIfRKYMIrgf6Mxe7oYSTzSfDUnUzHJG0ZQBmSfKDIjyS0vsnFFH2Xu5jD
C/X76N2kFyGYJ6h6SjJ4I6yCJA8w+24SO1qwbWWjyHcmIxDoKchP1CAkjjJ20izIHhE69MM/7IFI
BrPDVic7/WCUKM9bolSl7D6gYKbQGB3DzddaQYZUEnce2c1Wev0Sa0VkjbLNw4tpZ53LtN9csOks
1ivBeLbU+5RDqAQVsLBc856jZIFoW7SNoWHgcin8KYIwART9H084GrLe1DrHEZC9c1pK1MACpg0C
vCK1+ChG86+yI38vfanEfqC10Xo4g8gwgXJrU6tfaDfIZe2nyi91z2B+/iITW/p7R0l2PGapMXTv
8QtImydoe6ovvwLjGpapfc2L/r7RcFWhh/YFCeAXEgBPDzGLCxVHKjUwkLFIIVZmiFy+QtwaU1oq
n/psPWGnCxcwvGcKbFKqa4OUk0vuotSGJ9zV7o2PFE+eXWTQRIvU8T2rOmnwhjWMLw0QCUXVhgz+
VdTocKmKrtuGXGx6mr6w5Ng79OakXXTbe/2QhcQjCnIlh4iggnl0cNKaCAB7pv7WJLlltaTAItyn
2+C+GUd5t2H0e5jCfkQHw5osbXnpVjDAlI5UIWT+7VJyo8zCM95JcrN9xGm+BSwe1BwIu0dmbZVJ
xnCJVQW+2arVDJn2PK146bADUq0YaryzgJffDlbS/Tpwt69ZcO60fTQXCK+MvC6w9Ql6Zbs9AK9p
BDQ64KISsb9roAdlFrP38By0qnaslPQNgQiKY9/vYCmxCMuo2vu4sVxaE/W/RK1+0kFTe4X+JZH9
+YR+PN2xoPoTb27Rftss3HJGNwF6b47GPpcTPhaQoVUNu+0yggmAPtj9RqIKT5pJwNnV0kabsh9x
TS5ycmrenfIrFA+G1HMt8UpQugR1FuXvw8e9CiJpij8JVhal/Rh0tnssJ3Bk+Cffx6rpS+HGde81
P5t2D0GbV7qjIb+a4w2TXP8UNc6QBpXr3XuVaWhKLzSHRrLhurxf/GKXtrVouwMFLvgSUYND5CUx
dVEnSOf9BQ9k/K7G1yX7I0cC4mEeEPSEim+hizp6lVDc/+cacY+YaFjTW1InywYMMmhOnyQUfiTf
wrAjzSCVAsofinAMK2y3Pmk7TDND7jkHgnk7jlbxZwdCkZJPmunKbxHeAbzhqsywftyboYl5KPz6
E403BLGdxK2J+mQxB78AlOr9b07exx03yE7LD+q64mC6Rvxe7YtBBOXsPSU9z72NkB6Qho4fNXRN
zbYLGxzY7wB/eFDMNw7raxPNq6TVYL9zgGycK270SDpgR41qXrT2eIL8zuVPteW8qlTXzr7H8gk6
CKHnCSDTb0qpPLDN6KZhi/EvL1DhPM2AlheU8FONu8MeOXL/zMliXMaALpONRaJpqW75lEub0qKZ
vvwg4oN3OhsUK8Bc8p4qg0dUJKDkRfNDcO7UYjSJ6t73Gki8jxDemNka1zi8Wgfs1w2NfXyPo6fo
DET6SFYlPGh8mWPYRXcArSJ9AvEju9DXRt840caSQr5dSD0XWzEl3XcOE1NbJFwdACr+kHHYflVJ
KfLFrWXOxvaXQp0xiW1nEKyef/AmE1gsIzPLOR9gAvR5yShxnF6v5bk5OXXe3GFbIEnKMEswhcG5
LjFEcxHGZUT5jX+qUC6LN2L/OZPieWV8xaSYDBQhR9ZJNLEZrSCHpmMQpkpwZJhyW6UrabFPXddJ
0WQpkR6W+hxWjcyuFLTO3rI0wKt7Kc+APFwELcC5oGIENNoJtmlO6tlBdsWWQOZ2YJVHmGlxxPyY
o7c+jQh07+g6jri8dEWA9URFcYTOQooPX3rllxM0eLRJYRr7f0CMTMFpFaLG0HSNxmJ4/IVuvAg/
5dngIPe8/c7Vou1gx2OqgeE24In5JlBX9wWYOP2SocIYkfcIiLspDF/JYeh/eOb48MYY9fBJm19H
wwF/XHrPlvX3Xs8COID2NDfytmlf5ktOLkJHl0njgVBrKRKipA02+SCsVQY3zLduKq4KuRuk+ysj
CBO/jOYKxFE6p4vJPMtKggbww6VlHhZPEKqLFhMajrtt3VDe9wrfg6y3ET47/tNBFCHYwszYGu3k
6bfCjW+nvrfxgKBWfOUeOQCb5PE2LivvMjNuwoR57qjpq9mHbhD6wMEaYAPaI8ZMIZ3LoLXhqHsE
xgOBDUWSqMM3CMb7jr8damQhik8NaY88uWYFDZ9j2HMkMmGh1NqxD9izhqIgxDlXFI6cOVin1s+7
IIBMrW8w4EEtZuhEE3ipSAZD2EhsPkpuMaZCI+AGaZzk0WmQb+PlHcMwztVdJ4vFvSufZ3kKeP1e
hPYyKFPzDBAFo2FrnbflvYf9DTSx8ybI4QK5HmssZwar9V7mO9Vi6Rd+5SXYKHOEFAlB5QDmsj0/
kglDvl535CaQB6pelSrIWE1rU7dtw+FwpVbJ18jXeW7m0hJtuI9pL8N44oykeiiRzzGlnOH4fuz2
9KKJT/co6mxr+5Uwt44DrucR0o4p4UFX+0mClBXrrrpt60rzi6FrL4M+FZYHasaB9QEIZqDjJfTO
c+Eidxmv58bKm96aQ32jTvzD22xEKw/F9iI4bQEnHjhFi4HVGkUEuqOQY5UcfIMNDRh/yytU12+t
K4l+lYbqzZEiGXLvsQKZUHeyGbVtV6GO41LFGBljToU23oIIrpHSNHydyaqO36/K2wTFdHSsgu8p
2ciWGy86CcpFEDVVWUyYfHsLlNwomQM5CWD9EzR+Z20wKFMOVYHVUW1kZ1//3M/A2rSNlmDj3H8m
lR24qD8rdiiUPi6uQvK6GYY7JQ3T6wesaSD6y1W7XaVRXlLx+I9wKF4CjJQRDmUf0Eh1MovZD0RA
+utiz3/ad7hB55W4w1OK9YXsvAbb1B0P/wvzKbGsnGzw9ToeWVjHb6p5N2buX3ntE/Te2U8lchmW
zxN4sBhCmKUnA3psll8d6OLJ4HT4kHQ3zF/59R0BklR0YRtuv8hvr0gUFJHRXAMJS391l2b/+ZGA
LcXg/y2HwFE5mvf8467t/842KDoAkqWHESzuCmHJS05wsmsJD+OCVrTlcJ5NYoUiFLYJFQcFqNNm
2qewst+AtNaP7Pq5V8ULXxSXqHihhAdX0AjkB6NdQTEzZDD3WrOgVBUjUb6sECVZXxnif+YHfHdJ
wGO0DiHzdA6WWAsr3zkkKdtBSHL29eM9PlrEqWUW/cxw9IXGnXTt0eo2Ibl13l1jR3QQ2pr1otz5
Opsooz9aAde/EdztIzlenYmGHNsFxlqj2DDwBUIYDNMGP+gELhFBHNS/mNaWOgaSnjPOfh4ysGMD
w0aFi9ds6Ob150f2B/skyXAyhLkHer0y/4v2VT5QiaS1fYbh56s3Ms8MULQan2UEX/azn2DzkO59
L6DtGSn1Dil6gJMAoVYO/64NyIHQRpX68pzkVantzkRVRgPaDLphM4zJ/O7kBY/Ci5Qbzgig7eeL
4SrKKHxxByDrVMzWNF8RzuBBy2mnvmxaMqHVH9lDRJW+pi7lO0LQTbohNAyfK3mIWh6Pyms8tE0h
Ach3NS2wURyOd5JkdkNadsyIc0/roqpzoE3NXjtqBm40lxP2FjcrS6hqofPcMGvfiDnJ/fbgdjSP
buT2xsMhzzTON9nHwdY8atqAhmAN4JnkPmEHLgdr84+m+h8gZLx1GFpy56X5V5qCM3U2NaG1b1eS
q9fcig6ZWx/dHY8OxWmHY8Q3cAUWWnqFaWfT1iIJ5ewpyhtz8RvIzvVA24ZJlvcTB0pkuRCW9oYz
DDgFBUTH1EbVTlzQ15hdsis/Ui1q6GI0oHwUnrkQwDnxAHDnesibTFTgV8i43zvCK7hOv87GWH6K
FjOxYCxJXPBJV/N7idBXhUVvVcb1BvL5Ch4OGjl3SCcch0oMic0Royl9G4zUB/0hDl8BqXJQfDvH
VNI8dmhEejwMa0jEGsT+LbH0I2/bnwnR4fFEM79H1wz7gAyfEvBHJuYakIfAra21m2/+IIvV1qN+
0/oOqwVE7sNIreC1alqPJgN3CRJ/z0pWIVxbfzrSeTzRraFY5xJXmFn3M/RtnMnutDjYrAd1oAzL
OWrDLaB/3btw44Z0hHfSa5F7VisNH4xlZ1kyASRnUoAzE7ZHya1eJH6BjTHLW9STEKc6fcvAVdkN
vrC7SU1PbETr8Hg3EZtIdqeimG1M7TdGbvQA0MeofHHo5GZ4z5YZe7IVrUbucnc3ALq36qPvK7ml
vRco5EXmf4NOWZy+cIvUPRVF3fSnovBm9en6UISp0iyLL6to4OPu4Cn9k9DupDGJ/x8h6rwJVuxF
5SgeJQvaTIX3H4tix7ik9bsv9WCVkKklsf5C0UGMgEddfdL3DTMVFXjAtNenQJWCvEF5ChWZB6ey
LUakNtpBWz0NYqt6gweXInNeEhyd+sf3WmLubJUQmbsKYM4Ys+mM4Y3uqJScbrWLhTlfr5yjic7V
DMHlgsDGLWcxVASZtiKMYIZ4Z2aUflXXbBwJQUyr4QpK9mnPzsOVZG95s1dbJV1hCqY5oNuZTOFm
3+Rrx7KJbz97DB4gJFiyrKBWcOSa1HBodO6LwrUQ00Fm2bWenLs9h7np6FujpS4Oob6Fdn+vU7Rz
vT0pehqwfhWS4WG3YR+6pAwelVuKYDJicVItRzX3IyJBOwGcIIjbafLN8NG8BnJD0vbJtaefD5Aw
85Ns2gS+qwBxLzlGDj2KL94hzrSccUSxfyGPoRN1ltORRpOv4xjBKNYQDvKYuyYMimactQe46F0p
MtUICUUbwjtgTSP7gNdoOWJRTDq0auFJl03XLC/Id5F90iPpHBNZV4ZzMgodOQ2W/UnbsOtH99uk
IANujc2ONA8eFguJv8SrKXEowIbqADHcugVmBAcGhpXI3BbVWZd6TBMjaCA/mAuEPlHbYkDK++b+
W2DqHnec0RBOqYaLvOYtdhdi9PTBuueWSLtiPFD/F+thlHwLl5OQvU6ijnWtr0hDDg+UWkzig+E5
y7cePuPLaowdd1JZucZ5KcUnwVki4/Bd+k4NHotnax5wlMDm8IGt9dGPeLLh1sDkl0bvnaG9iick
CapLa3mnD47An0iipMq3E1+0UeIofQE5nWyb3hDPYgS7tkLG6cdjeEd9MrpKZ+3yJMBh6c6B165D
VJ7EGevnVdbD0C6bTBC0BQr2n31Nwx6BEyb0H+qnYsoh4+MSzJEAzZe/ymI1bxhFF7NUZNb/9PAb
Lly3QqFdBSlyV68fAOYFv37htEESSvufuIwEIMCALfAp4W0qA54t1ZCfI1y/VoIVAHbwSYrI2A4X
DJ4/48GR5W/0pkm2RkBYkdNBvoelGj9Cnmaaj5BaNufkJiBKfv91HCRyaBwDCtjS4D5osmNyFKAb
Y9pOABACRqQGB3YEuv/zDK34eY2BLHWmkcp3SWcazPoqmXS7aHYt9fnK35zvSH0nv392N5JIQUkf
zvLVeWEI4lUX+gbqwdPKVU7D/8mAUTcYMdGJ7bZG65csdO7zFalK1JvkF0ODJ20cB0xTPUfv3fPe
Ro8lnzjc/dO76Zt54gdrKSWBu1P0SOBxXEOvg5BOslkmAQiYGEnVqGChfz0tJ99YefaUzOmdaZjK
nvuE2rYKk0rukSqp8G0+MevR+IE9UUNUcQH+gpQqjzFkV3/dMiyAZNrwO3W+oPC6STftPfdD8Qux
bpqc3Zz0JEaUblSWPuVTK957gxEeoGnoMwNsCOYTN2ItFjn9iPK8I4eSZi1BI+ma6L8AvxGmVJsF
1y3RJWAolZiLKD6ygybdMWHcmuunvnWhCTrdULu0uaUise6uzSXjAuE6Diobee8DWlcA7gBJc6G5
K/+xivG82hGGRllNvPr17YGGrNX8KhccD0okmechkmxJntWde3hWpgbGN+dULCYC37+Il7YStBsE
DI+XS11/2fEOK5Yvh1f5VD3F8ZQr2kgGbDfpboFH+g5l2fz7dKyxdz8Kv534s8S3d/AZ/6VeoBop
4vU037A5yJVXayL1XVYd1jC7VHD8xezDeMe4EqP4hI9CbKXtBZpkgiMkgfYBPiTw84Fgws0gvKLE
xooUqYvybD7k/A7dOeNwfRT28Vb5F0TlwBoGHL3FZTZsGz+lwISymKqE7uieSqihhGFwcfermQeH
9ijBV2atPKlmYjO7+I23YtqQMzsxBYzbvlgVgvG56nbQL7j17B5pmjuQDKGUii9UeIOis3MDTP4t
RqcRC/w2ItRCTHecuSYqEcjTixYfuWiX5Lrj6l+WNECiUYoR8I8hJo+SQs8dDlBGHl6MJaIMUiTj
TMWkcj7YWf4+BWA86fXQDdBaIwMzE2+G9VI3PYgKQyON7bcGRRGvtnoLhazVxjNRBCGDzBp9diCP
DUhjV2KHa9wfon6JHALmxV1b+q5mxyBPWEiAsvAVQ2tIidBr1fZyzR72nFnJALQx1Vy6LDrJ/uc5
hYPnpXcku2pZ7rzLfmfmW5fyDiqjkVWqfSA5saLm60gf7938t/RWQn13Awz78TsjWo/KmG5OKG0Y
eCsfavoFUi77R1337JjEWRrZgVXN4DZE/4no8nn8v0heGrSf2jdNaFAmomQN8qzAz87mV+aKsyfC
smxZJCuzjY5zjDx4UFaxrS1tUdaPdMSTJU9WM8CuhEid7janvD2GTpyfvVJdnUgjX6lWG50AyfFh
Q4VUPZLLMsArznjntnxjZ5f7DeSLymHqqoT+w3PvntfT5s2SJhfTleL5ErUKl2jgZM7TteEn0jZM
8pjk+wX1TCrk0nY6Gttr39RNRIgNKAltMIr+p8TUBeLar57R6tNjhILldRjhEZ1R3p7mOnOXtj71
EQ5Zm7q0jEUQYjSsGUu6S9vHFy9WKTy1UIeXIxYO/X7CUed8XQAfu63+kKHshiar3BFyJPSITu5T
lmYltiW1uabJXh2AZJkcvWKEuPBnKc5Wkc+v5xYQw5Q0+aEx5AzMdmi9AMHiI0QLH1Q0ZF5IKhdb
5V7bkSOHwvhe8/S0S1vfw2o45uMqbPDoOBhltB/frNNpQvd3ipZAvM+LclrLd9cjW6anwPvPXyH+
WZGCCHF5oFUODo8O4vYkGqczmMlLSoubEiOe1P/sDFcwH0jp/qnnqS5V1hPnZq0Z3+aRqaXX1ASu
WgkLAmA9Wa5NaudfKQLSKcAI4PDaHE08s5AiIehVyQLk2koYm9CpeAlw9LopC5Hc1JLX/TiB54Pg
6HiE01LEHLLvsGk7MD3I+Jh377358DcWYji2mYVyeDZH72wujXRLqIMLreT+vy7XcTkxxwSvp0U9
01BF1xzJloD58+xArgLObCfxlM74Bb2DYqUhbDbtGCM16rvlETTCj2XtVnp32Mci15jq0Ho5puDv
aRf25EzE4CXL+DC6BA1pQv6y8VniszUHPc1hfo9cfwpEdE6SMdSflo1dvQHPj7YcWotuJ9p7BGok
k0CCVGK4CHN5CK9csO6E+SI1mGDhe3+X9P5p+RoRAmmrvoO/GVXD2kOpvrn+JqaiV7jT8CwkhC2b
OUNcn8fBH/TkpEJIX+LGqcbWBejS35Z4WNCJGtTLC+WO0reHgrmoGXoL0q50CtaXCB/72pKVirDL
TWX1OKoZo5IYf/m4Pu5N9FE89HBVWUy/AQkzlYL6IajPdmj3BmP2vAGlgmKqK0iEYsaMuJ7h8SvN
y6g+mRmoUd3i+Z2mP8VnZ1EG0GySBG+TqEr8yCq7l6nSEJTJ2OiFmM7XE3vZj00u+hNxk9icrFDx
tkRIKpmb7JetVho3wy8jCidjlhIqoa3frHKORSuifOHgqeV92g6zD8GoGgJb9QNb5ihOgHasUt1i
EK6+79bd8sQ65pVaqs2BW7uZqE6YGzR/ud25HuSaadj1jpVgkfcz5goCLLH4ruMFG5g7fekZmH03
CTwdFTc2uieg5XweFS+usWMG/95p4NYTrwwlSLQbyzPYlVfkyxrJUhKsUnK+y9xGJG6KAlc+5TUO
5cWHHwO1GjqpQYOVqabPehAWpjldO/WQnKMGWd7RFGQoYOJ29ftMu6aSVqkvic+Zlmc/Kh4uoiJO
sH4Rr9HYWCUg2FXy1CymXsoZmutjtPibHo7Ux44JHWysla/r9G5XCYrfOqy0b9UDvzwc2Du6M0+B
vLbAOM6buAoFrizDDdJMXwBdayFwQc15wI0XSQjW7tmMsEgWST81Hcrlk10Xjj7NwHnGHvnj9KhW
Hhb5r9M/FFYu+I42hV7VG+MeUeY5wOeHJjOKYwxuWLClbZ5GlSB1QDI8WLYPAOBWjNS1x3fEVLkU
jlY7F7ABFS/+otiP32tgSzFhOscNfFfeaCmMP48cXIuC0Ne+jJpKFx5xjGujqMyN8KLH6SyfBbB3
6fZY/Bf/dHal9eFhrNJyN2Wl1XzDJ2D/uno8AHnWUjz6T/FpiN4AMceJS5vnDHwbFYnkYtNL2zpI
HWASWHKjiFKmxjOtKGgJWXrO0BEGt9En2rtp3GnjN+NwltJhXTNAld5O/lExA47wl8VVI1Gq4mri
hOO8tCVinJS+MyeHU+IMSoZtsg3QR2PKaaZOxTEkwWJGWGv+oBgrOwnEtl1gp4U1oNBhEH+SO72a
fI/3Z+NDuqYlvc9h2CyFyJ/04oh7aLIqzVeOedYZg459wX6Y3P6XMJNYtNeeJjaon0fbLqm4YhWm
Scj0HFAeSDtrqE69fCtIr9k6UcvSs3DOLcVXbdwfdoHGfZuMYZUuzRETz5kNcbunLkKDrSILT11k
IACzwSwZTmO5psxneYDLp36YS1swziulAYGgEY2Zyk1E+UQ+y7IAguSiQ9vNZ+XQP6rlVVQqM8Vt
ARXHdP3jEmaDmTkmTTTlOKR/qOa0azGp04ZsNDy4X0Q8/LN3W0Zg/b0OJAYDNY58V79Nx+kE8QZk
VMPrRQSOmeDVKDc4+AavgaKT2GGOOX4D86SHI7Zsthhv9kFzwVUHX3Q+/rOGo1V7/iXRV8VDKqNT
p5J+el8C2oEFVzC1RdoEtaPqyFWsesO506kaeWSlzAv2hmAMdD0kVbYq4gs6fIrsBYfmD0bufmbt
4524yojL8/h0XiHemfkUkrvVQUmj3Uukw59I3JG+fIqS55i1BHNmqWQlEsTQHEQLoBohcNT/XqiA
kDxoE+/WMU0kxdalKjfCEt1c0ngGaYT1XiVTtetdydo7ijJKo4fhcLoi4Hp02zwke/HaLq1zprr6
qqw0BHnLWQDfbDuXHXKp6lHOK0cgjYjRaojCToVRnazBX5m7nnPng8FoY4uAbQbEr7c7ZdUVMqb/
AaCNImSbYhukxtfhD+yOQWMJFoRuyx3bXB3gYRjGOiX+inat5LzYp4Xa1Eh32H5qzPEeXXu1BAnx
4x+nD3xfYCbzqehtJAymMN/CcyKoH/pcQnB8fwLG2sC/VJi1dP2zBc5V5vv6H8mThhX1qq6DB5jM
b5eyV/sg/jEnfbz7DUNymwa3ydF151Yw1lC5dZuX1MQ+9B+65x/NyljSYsW2TRqoy/A3y3OSzwB7
pcy8S+V+yDZPvt1Iyv3ydVuU8BwZywT29xQd9vv/H1BjSfxVh217JiWIlli5HRJRlWKvR1sH5rFP
4R2XMn4IIYASZq2lHQDrsR74hSFPXXnPutqSP/lQsGl/xVqAperBV7Vvy7l+gX1EVzDzxVPXSo57
X+0ngTd+IoP8B9OKnijH4zsmcTn8PGEU7A02Wl4IcXs9pnrcIme4I7zxfdVCoJGjrr9IP1XQkPCf
Q6pYM0BhGWHhpfrliOHYdpeMaedJ9A9BBsVSY3Lerr/uekgKYlfQZtSgTTTg/Yi8J2qaBokweviV
dAvEbNpfKfTCBaiCwV57SnJxQRujaAL2exz8J9ouaGSkE21UPv2y3ToUDPpY+q5bTiBAOAuI682N
7ReeDUKcOZYv3sj9BFcWllqkLvKfGoL4fd1uC1UnjFsIs7hic6ZVZYx3m34Bqt8Rr8UbIf5Yti7v
ZZ2SUtBE2jBYJRnOOsAiWlzaapk+ZKwiaoGgOV2NLQ1EeWFKBWr5cH1NYw4fzjRdGTdkwBXdZYZ/
D9V1dNkUUaM9tOM8WX0oojrO4Vaocmamzotu6F4mbuCr9dM+UFdl4b5/ZSRMo5F9cryWlDQAChpV
va8x5Bqba92JANhsIj/VdLAzjjNdZIpFbVPfsrinyooBz2Y8h8lVoFqw43+zqvvAub71GFR/UF3c
Eha4DNBQWHQlH5RZufMxnuyxYwruR3JosUu1G0PxK4GXoyn12SU+BLheVzAz8rVTmeKDnv8fBY0N
6sxCvFVrR4zZS9dlPkbl53rn+rhWUtuQL1QnE9KIdt/Z8nXngg/MWT2weZsqFz2tiaecBeTpDY/d
eCcrTCyoVkdxoo9u4P6vaP3s+sKWVIlnhzJ1ViZCpp6YElme8uS/VkFuUEBFk9p2J1cj+6IUOBKw
EmSYsDgdZU6f73n0brWbEBCfDNrnDSCjX7Ipmfeaqm9xEJuhcmXOQ/AcXM0rVDh5JfpScDmDdMK1
Lf1Y7urkWLbGkPagX5gpFH1hL9ehkBtrfA4XFvG8gXv0ps0qAFQD31K94g2uB8/oG7+gRcWifMlI
fPvNcse/nEAZMNM73LAjHcJdhyms+IwdO7tbl5CzcEUi2kSfY3xe/8hB609ZND+tYtAbus0OdGgo
QywgUBjpY1qCfnPQYiTzDmxeAfTvOhOLna5mJ6pOsNAZhdqR8csN08JpjhTYTSbWgy/PyJLFqOzh
GwlR8wbSXN29cnIWr3pEYjMLgCr0iQlcEw/MvWl058qLWTN5+NilPoKcAluP7BDo/1ED5yISi5PW
DiuSS5ORZXELLe/b0IaiInlMN/xnLNJVYjELJ7lZ7QZh2JIvBB0SI6TuE4l+0LIaY/DMhsKs/sXV
qGr+eaIS6+bmsU/CAzbKkNvxsmCBseJ9gxhpNG7bn6/LNapDsLY5BApM9J1ale9gEtqTGolM4rlx
A5Rh7vO7tD+ie8rN1RulEUVXKaIn6fHGJpeLHUPGPUIUJ00gPNvh5zf3Z9s1+EDBk0LuU4tmEQBL
Y66xhSU0BZf9y5h8XIUPrKska8VJNTOunw5MYUJCXShWWK9wwsMt7J4NcFSAJ4FJZXFfXRI0DFqp
C6PELCIk2uxj8x+dvmZOdOdUrGMnHitWR1dgl69rnh4Ds0ZRhda2+8TQULRkrabOZ9CVdeSwrAXx
TVaCabOI8CLXhe55GpMDeFbSUltAoOu09Ur+yzCc/Ajv8eKu7NNPRkSIrZBS7E94lcO4vk5NbHi1
JKWENQ9S/yBZEjBhGd3oTPSNQ2ot7D02vyl2nwmvZD4sbgJp+BiuZyzRU9YSsqbOSr27V0yA+koJ
TyPyFsjTShIzme2mDe2GWwZmbK2uiZ4MD3LZ4ocGi//cC0oD/rREkR4THgZYxXvyq4y0jft9Mitt
FQT6UB2KKSPgfXlxTXmYoSrSBwH0l8i9ls6SBbm3BLifbOSbwE5LUqWClOcr/1OvK/972LlPF2ip
bVsJPihnkEYxrHK5jN4rl8ATBFwTi2I+1/gzB4HlN21TTVoqoVVbz/+UHM8QbCCH/7OMYln8bDaO
RQj/rRHORpEvKz0W/IHpjQkSDmTbOoZMQJGjrzyBpKNzgjIcw7isMhQP3exj7+SF2IQjUZc3nUnf
WXOj4Nw3mqIh8hQpf9JpJzaZec2g4SosMsi7wgywwPCOC/RXA+5CBsSjGK3AIrhAASy7aXv9rFUU
emkUlwgRzO9VCiCUY3vfIaWzzJsemfvfHvXs+4PvVSICWo9WIwtBOO5O2R7FEz/1d7DCPiTNDinv
iOqfWNvLaBYcro7cP6Cm6TgDvGe/GdfIC2DmY0mKqpP44DHNsti1ZBymvRfyXuqcXsTuM9IxAwWK
NZgt+Keo31oAb+IGiIxAa3fU4BA+hGyDrqJNMylA3E8/c1JmB5VGOvSX906QX/TMOkW0S656RlsP
sNbn5mlTMRnJe7So+TgVtL8LC+YMsTi7VtotAKTrKxCUO9xXZQ2a5mhbwRGMLHe0/CFwgQZtVJVf
szLxSjp74KCIxr0Lvm6xLq63Sk53Zt4onUpJ6MP69kxti3DdDzJwTfet7eQVsZ6DrVcvO9yUCvCt
sIQ44H0bVmh2xEtO1LxyMYiwxTG+gYgXz5Zy8xJGEk75xpHUxxcHd0a5fiRyTTc9Y66eTl9IXndF
eAiIgkrjdFP/wxXk1iZP0QTxYuIbLewDuEhbUH8mC/UMehm7r9OtQeTEhNdOtxLzuoYm41DeDxtL
18FL4n8leq76aW84QPZgCAHu+TXUQVSDN9N32SyFlOH5a0oFjMLp6HIZbQY3QiBd+hiyTMKFt/jG
gg6haODQu2ed2C1RdtNCSupi/xvpzPpRoW9sIAcCjtUNfxl2egmc+eYF8wv48IkZO5XJDzV50oqa
LZ1+EPeQRRWfMSaeHep4Hw5tCErH33gwqgwqx9b/TA1jZQj37LSbY3uYuxPODaOPG9uirjPLSpU6
EWOzp7EEKRPrhUBGooNDrnjJyTUzydxDAxFivqcWQVO8wHKY13lv9Qpm1SKzpgFTUX5KcGjZ7qPY
cGDY5DgSjLtgSR29zSKTXwUVIZWU4iCWqhEEoYKW7hShKtiam3ZyI0dAzWRN89cWCctIw7XzuRNs
3ctxUAkweqbybnXKT3Nx9ezFyLGQ6Ee+g22H+D8ubK9VqH3UWjT/qKV4SPyBUoObdh19B2exMf3T
00RV0UdHjT+wS9UxIwVpC0W3+x9OCItBbsm6EK8ka0+ylqNBanJfVMcNWqQD9y2KjSz9Dr2+ALiU
FG4IaLeOvLGAUyn2r+C+dhzvJxc2AwH3YpoI5kTexo7EtYahs6BuPyog1Pe16MU+DYRjwG6udoiE
q2WeDJrTAwLdQ4ZnuVqgwxjNQjwBiQ5Dkb8KFI4sv+PTIffRgLeFyVneNsoFZp75EiVyxuX1KIcx
I15dZDrBZ0rdPWCzlUZtlQm4AptRqWVMT41qk/tvZMrsCTPGIPMmc/syCiwki1ClKJGcYKHVuYDt
Q0MU04Ju4rC+8Qd55xsthIL0OoA4EGnCdkRoIxQ+jRMv9TT3VscQmiyMHEG6fxYhTalST7GfyfsM
b/okd2CbeDZssozxcSCJeGlGY9z5wXiPOkeSDjF1bkXvL3JTxRlaZxLxcudDKqhJS1T2MB8hR7Ol
49Ely96DFWxLQDWzJXiWAxvv7zkXO3PeerBW3KNowXBHsiWoE3WMsEnnKgGQJ1GF/JPAmSQ/4Inz
Dx9+021525KKtBI7PeSEI05a2NXZNVCidUIHVi3elmkJlB0LCZ+urB/Jua8lyW1wHCzZ/ipZSkkQ
Y1wkEEaM6DUVul1G20CDJKfQFj1u6AY14aq9A5vmWufZrAoak8AfkiLb5FFCEdRWMZlE3ZLWxtFt
cXS9NRfWIDjmvjPGNdE4ydsMaCfz3R1O7UGXexzxbEOJN1rdW7jOyP+j/vTw5nlIL8DCdrFTy6Nv
338t8UcAfyR/f/WJsYoJ3sMi1clX40O3KVOFVL+ZGR1YI8zlmmtq5M7SvoyzHvXkCOSH0KR6IYr2
wblfAx2n3Z6ZBsQQiqGLBrs9FYl9Fmg9QJesghWyaVhmzkyAQr1n0mLDz3i/jgJctayWWmesM0au
3r8SuRBetXkVZlEUJ2buA6gcuRApnJekRq//gMlTLYRcqsPoF2yg42skLy9/SS+5yZCZ73jeTtbt
kR/0GZjD+PD6ZlT50/z2tGKmcaag4bG9pNU4g84HOyWUUiWsIpF4GGqaQzMYaTlbSYcRn87XqeTs
vp1NuqgOYnpHi3i4QyCIKh+T6+ahdcv6qb52fgU7bcYVG+0Ag6LG7qqVQV3BgdOCjFoROPlfn8Su
ZlTK2QHM4RG3v0cBOEoizAFnNH+xXySsVDlrfGzt1FVpQVIs/c1n1Ow2piYzPhPdGDO/9MKcnSc2
gxdA3MVrOPCQEyvPbQCpXoVlhYJMom7IzEY1+oBhjni5ax+kNp8gdPu1teGgrDeTcMunA9Jlu/QR
gA67hQvDxSfuyuWmOmNjuMMj6e1dfOClRcKEDbSsKNm999njaSEG0/biNxHFYeORrTX0TdMmbl+I
2wLvUqkRj1bZK2FG3WcoWx6BJ2VVsRrHaEvm0L/weEwGNHFp08KBJTpqTtPI8fi9bQ1ulNICWOMF
o2a35j1aU6HwUEEPSYPYiixJvJBNLEC8Hh8T/VvJPmyEFLFgDESsz8mU6+JqfdnhLApy8VOqwPkm
iZXkxVyQmNrMPsZfqFBtDrdpyNrDURZwQmnv39DLojNAYjNuWOkWIuUZ8tMSIdRkVZAKWw8YXnne
2Gesi9XEQZvmY80F+MrbkTPqkhKT3FZSxZIWO1tGormyljVGDZ4XyuqHQWt2BHbOzKTVZUi+JryP
ES7spQLNisPbROShyluvKzuqyEiCKpt8zx4r2cFKaZHacUNmiAkpTumC8XbDQ/dFWUQgiPGJgtaQ
dBcSbPIrn06liWB/L7msWXuh2LeZpa0/0qqPKtDFTSWP1qXviAUPKRsLHJCAbIDicyU6ccZvTNIh
pUgqiqwRVock5KQbCtqs+iFxUjpYgoyRiKNwBmJzhTwbA2eemR/c1ZdW+lTmD1+ZfjFsjfBJl9y+
QvvHsVeUL39zXCJK+UPa6G7dQWXhlPyvN+QTjRRiAhuO2ZlxVQDQtAJTwIG9Lx/0MtOCmhh3Goxf
7Vn5wGzgRk2uKWaLJAaCzmIVzSxt/m62D53vEIUYxj+eKRPAi+5ih9XwGsRK0JACmOBqUs2BWL5Y
Ax/6xkw6l0P17UGnK7PAr2gQSYlp8D2mLQrg6J9uV4Bh1lOq3dlV4RTRO1lh6sq3BnbnjV5zJtDW
iPR8uPjMYE1Fj8wXH548cdozKRw0mP14/IQ2W3zJ2DPUsOvPuryJxfRfZfjsznNjr0ydeI1Zfm1o
J6438Wv5J1t2/gpnTDaLQKxBmOCsBlltWPAKNKBlxXO/q6TFfCaJVti4IGlhr2hB6osr1jUf/JDr
6jaW+sFEfU+HAsWiPdzvpdm5eRpVtHC7HlAi0XKlrafaIhIEGQYFMn2UaVsydyvX/C5AqKclLml6
rS1Bd1vMJezgAMoWcxVEyczZFHYCdMOtSHzHPogCGSiVI0v0Ym0YwouxGs9EvVMYGUkwJ6Ydbhao
IpkVPEUl938VRtVGy20QkIvlyywan8RRN5k2DcvP6CgGJVhAtN8pDSQqDNHVWjvONiIjkMHiiHEG
uZ0AnJwNIEhhVrMI1iNa9g5WkfNX39BW5dc0HbhlIAIcmaennsG2O7q+e8vo1t2YOrLACekZNXPd
pld+Y9eI4TKFZbjy7gETM3zGG7TE7oNAkkCIf1Ga0c4aMO3AifRfKsIC+M5U71l3Ns2GZWFl6bXH
XXP/03zDj4hWiGd/8MRYQ1BnX8BDx1sD7//tnRJ2yp8Z+ofR1dzkflKfKbwrLPIURq71Nzn+7y6L
RYJVaRtLiuYffLExjtebAtWJy5NdHRyPwooKYpd1ZWY+0L3ViL2nSP3dW62U4eLS8NafBDEtjhBM
Uf3cvNQ9MUHz812247kL6G/b0t0J7pIEXnP1BS3gqJ1BXGjmiKTZk06m75EKZCg8Dkg8ws/jPuH9
K09Trpt7E6vcRNSk94ko76G3CL25OtQc5bUfuOv2yXzP8z6DciFpmTxbMxir5ew7Ga7I2Unvrc0o
+WlGcJtIDe9jt1UD3FwiP+p6TEM3s6xDLV4DngKhsxKV+EWwgAzfbPx/klj/elnjrY5IC13mmq7W
eV0U80hNYXWQP9dIb8iA3Nway38LDDbW2glksk+ok+B4Ln3UCQVhsB0CoeHjI6BfaDxyKMV3sBGM
qBigixeV9Jg2lqotsvOgNWa3LzK2mUm5X3/TeClfrJJhT07uX3v5yXtJlDiAHj77jVEJocN6VEmX
rq6ae0BtYWgqHgeO3aPgoi9QY7SeNIJQN4b9j9mRd5Vl+c+eru3ADSoki2n04etsImBzCg1KNKL5
EHHZ3f7lIlow7xvOGyxumNRh/UHChDkc9Mdf//0c0r6NXzbRz2WcyZ9w6XE1qMDwQPWlv2bcjBb3
5zq/PMs7e/uvVTk4yxft1irGpch+ZhVwznW5smKRGWPitg9bcDaVOfA/SXNV6w0tDIGeA3rQlLhj
iPl6kZJaH1oTC+0ab2onTcic8H2PX5rYULtUcnZX9Lqpo0jtg5XY0K9saKjzCTeG9ddIv93PBK18
Iwjmf95JJRlUIIRA9GfsSBZJcsU0nZu0zRio5QRMCDkVy8yVJdeFhxMTzGcHwgLJBThgWEcYuvpL
QAzltesCbMNUxH4OiCQ6+mC+8rfJka0S8wnDF6dmyY/aWZa1EDxyXpPsiZBRUZ8+rOYboePtm7vr
/Ar+fErx2z0IzwEE6UtLvlT8jh+/7RGR9Oks6QBmFqUPS5c5FOAS/0j67RGL5MijD/9p0EfD3R0m
5HTOebushxE/FmmHuoaeDgFpXSkDYiVqU0gRRTlOS99aYQZbVWHwwfNBOkqtirUJB2KL4p2yuehu
rxaGuRzvqeKEg44uNWRdDh5tPbbvoxv9Pzyydr8V2bokgpaa2z+MU1YX8MstiwdePobsP3O/Wqim
JEqPBIqfDI4QMCBtNCoSm4S1vbDTn/Di9rqh4a5I62uqNTiPAsCL2YyFmv0XEv8l9QdbokWeHnJ/
/S+3TPFxsB660DuYoQLLVEb+7N3SL7nAgx2I5lrdv/9AT/i73EB9WktpeIVaBE7e7TSZtmPZ03VU
UJBsuvYpkQOifyVdRvI/iq4kr8KyTTN+R2PlRXSvz/W6/UOFmLZKf5P8t+mlbkZcagM2jPNR8Lyz
p4+h4tu9DZ+cqqj0enhx2GOoGHg9Jp8D5g25kVbC4WFl1+xVs7MPLoeJ44J9fc39WUkYzWPB30xc
awlzN361mZrnoo4aUyhmNWHdjN5fuqJCd/dtPm9PISkTbOAc59s/ghwNMfnNxVo6GinHQXpXg512
cBZ6f3ZVmR807zZlTmxLW/KibNJsQVPbgZoaEcrhw4B5RY2J1kYxMauYcvx+30nJ3XHileITDH36
+JWnIpcAeAwsn96wXbHdbCoh1MUhLQvSjyAG37CpYlDE0H/W+wIN/ggHUxBXvj94Jj8gYFt+3yrk
g6O9h/P42BOixI8/7YuugTRQId3O3m22cIA5/c+LWxI41c1SUohwVAF+161ZVHUTGO4UmxVUoc0P
Y+UOuoJwYTH1Jfmk8VzAZ/XpWM4009uSg0GQlWv3mHtQz4kyAkwepebp1K9gAYyLW0QMAMjmf5Xw
Fob2Kv+PuWcJ3rvhSQQgCOWxQOVaOk03Mih719gsk6kv5WRHrrWOPNxapGnoOp78y8vYmvq/jd+z
ZQTpXMXRsKbBUtZ9u19qsKvEUkXGctuqfVdMmqsaSe4YZwxHZkeAXlK5wsr4r3DCf3lurIsvJSA3
5kN9g1O+n8+/eOqkPifSaUmIogHk+6ez1En/eNEGsha3D30nV8TxGXTff5ySR4jOJWWI74DQLBI0
irOdO37iqGSW1Hi1AGSR4Fk6ck6rl8tsCTJ+oUuIHQLox+eM0HGC11VyFR/QKkevTjQ8DFeJpjXu
CxiXD7PE4JeK0P1dK4w7sF9H/tG4n/ZIAKtEUH8aq7wze0EXBue/U88HUHIIxQ6fexMneAEIZFj9
twUChXMjxBoRzcrDXXQBjO6sOLRfUu3s/is6uuNnKcNvkAlfUUHi5G6N1TfqAgJfRR4xdneuGr22
uwwmkLT/5TEbRHs4/Q9C9hRp+YEpnPqTP4oF2XiWlmogL6JLQTaQicqhkPap6ghOuTe3naru8ClC
uWsk1LNBNxIrQzQ/R48j1QsC/iqX2MZiDHPBZhg8tR379hhmL6oWj1oyHKpTI9wE+1XW7d8iTMGA
+tE0yY/PVBEEztwBToaw68aKDpG4nqxLMjQKcITjDkmlk3a+sBd319E+HpOJazzcSUsGuShBsXeI
svgYQbN6nD9UGuGDY1CRXf2a6XqVzqx0PAEVDAk8iqNasCb6s+OiWDBPOeOMneATgmZNzeuaqb12
hqu+dGdI2Ce7hP0aE58FWu/m3H6qt8Dz7but7siVT3CaPym/35jtIoBU8a6YnxX9peY73rld8BW5
yewmGZCrDqc0exI0IXNTkTzjQeUgXSsiACoJuGWP7fqZ5JWHd9q+8cN5GjVnbIQ7Mvfyfl7Ox5c6
kWFIDzsXNPHlcANPqtEMaQky8nSz8iPBPWOk9hY/WvcZ8uqyiGYPeTFCS74M5hw1p2z3u+iYk92D
3NJgco/MRHUmoyk7PuR9UcoONa4AofmN46ZmoWyX9Y721fS1veHagy1u3zZmArQu8FgoiZcGrJSb
ZACC+excM208AN2MfVq4KfhFZZ8o2CDbXp5H6txG0x9ulk7ptFJRLoGkemzz494TuPUq4mNqnSWt
c/LY/JmL9alGJL9bIWZpl46uqcgUY15ZPVNL2b7TJ553UzFF9wjCBfu8RtMlKYnBAxkhF8XQXQ2z
aYNQ234ixexcjoUXdC1hbXHeeUd+v3+ALQGyGcnk3vaMPzSvQ/hrSK15Fu9gwfU+GE6AUR96crJW
NdOCJESBNVRwl9agIhj3WBapZV5NwvSV2nC8tKutt7NK/LVl+KPv5yS0LznhPOJqJistUEzG1STn
BaARCKu7lG/nxvrj91YP+O4L3uMBpgHxHhumZoBdsfUJxxDAoMMZ2uO3z17yK/UIC1RvqLGO4HhZ
sJ4RS/APJHYrfdmdz6cLvAvl7NmRTWN73qfZJhG4gimWFpQSPx8J8t1oIOscZisDhUQtkXM02jT1
r08OAQvWEH1TtTT+EpUs6C+1iO2Ia+1YeAlgC03BxCYXxSiut2BwnurtTdfw4aZv4AvkqmfKCTVJ
UF1wJyQLOGZ+5Esnuav8Yz2EtBuyP41WpGUXeito/DNQijDZbFxKqimg1whZmrxNbjazD3japeVq
niVpuY88lfowzYlAFmqEaSM8nO3YdervEc1c90m5i/2m8KWaXNN9m99JPGUbJ0a1xq+o82E2RQ0p
VzvV7LA2KwcZKvifZnkaDTEGMs5DB+asTnBf8+VDKbv8fs+hHScnpkEtK7qY6UbiU4BGWGyCKVCX
/20RA+ZEhnh5V21QluB9df3yWishAWe5gTt/I0JDE1HCChLLYAFxT0MjLDtPdSzMFGGe0T+24hir
fl1EFzYWqC6c+qX5y9DxGJdyc0Xg2upQyK30z3rsWVnaC7HLL/jDoc3YrQMq36Z0SCDdqhj+JXYV
6OPAiQuoIUynZN6FC4XDGx5L2/ohOfsWON5uN4wF0hOuV65qNptS8p3iutsUUcv4UzIRi5EDkoAM
qBSkm7w+h3I0WrTvmvmq9orIOgJq6xgf8oz8nVxtLDa/LoGSDMdkdpkfqZOE8CCxce1Kfy0Wxisc
7Ls/gZxmibFk7Z46ou82MbIT5B+ejNpNDsWPh09GPkGiMS5UAv2wE4ldI/ogJH3Mtp40wEKZDWVi
tQ0iPQUlFWZhvA29tOACORhgJ6R7HgNp5Pm6Xc12kyVP+q0LFldanC9Y5bpwFCj9DUQ8rrqNZX41
wS8qdSvcL3bkILQycufmF409eNXFmiw+iNzNePHEqCUe9eQ2zYyr2BuOHguXu+k7tRrvL5dsCleg
0bOeEIJ7gN35G4zjfSyP35vnKmd8VtcwFASoIeS8qB8xr2s4gcPee9SCQSlFqXniqtGsGI8Zw1OQ
dYRivA7q1PuFJ4OwDS3/hZzAp/U8V8Vt6iKkHcY9XZbXs66pZbqf3Awsq3J+gxhtRpT6WLe0Q9DM
DQSLADGG34Zm4nkU/Y9Kua2rUMtrFRpojozGzdha2FD9jhJ+ZM0NysS8Woug1lAa3YcVzEMv2x3h
Vz/wjZ/SQqPOcpfn0k4XlxeDQlldJlWaB9SMKyEdbIGUv23n3mb96HO8OA0qXNGTW7RaaLfq+Fqm
CTEi3QBCACrzauZY0mZBtesMkV4b2cOaitxfJIxDl7IK5AX/GfMpp2PT3zk2vCJI0anz52p0M5xA
qAJvIWuSPc4hkMegVMLNnH/Pn0I2mXe7FK0scEqi7cUKPhdZrAexUavc8U8jhdeyeRyp+Pz9cFbl
C7HpRq7TK/NlQdXeiZsdU6cH40NGAVJUEBxJcIeFwi8b7vo0xA+55fzKyFg0DExZxjyFObP6ZADh
eFUTPHiKeQlRI4a65KJkAx4i6vdnocQbwD0rAkgw4f3JsH/XaPf2EdvjSTSmePCv5ut7hcTUyCAe
CQm/qWtj9S3QvSQdtldsM/KzpW+xIFWI3EtiLbhDtfdsWmMS+IsR5zPjbzRtA0xtf9C9xhGzxNwb
e1W1TK3XQflfdt7NMyUxih0zVIyhWoIGk+IYuOXHGZCsfkpFBQ50rd7OebWSM74dqo1oAunHMXFl
zE2lzOugYDL4QXuYIkCrxwvI6WL0dMqg9AECZr6W4Vbn/tMoCp00xiGG9RWNKIYcCCo6KjRD4vdk
H2Kwav180c84mTFvmpdXkRds4rO3HpA5oAg06q/iIcHdtInMNafkeMpUKlauYZgRzTfusUvS0Wua
VPyV0gOhw6epxgpeInlgKx6Q5ahfuLC4Vtezhnabi82rrghKVVw0AQ2nWUO99RXqthZa2QC1wuML
HoxAFqF5b4xYzR4KXsR1vHsMVQ5D1uKFPctTHUDlWNLOKJBBsHCDsIV7mTxW5Sjikf0DTd5ABZhQ
yF5LbnrTe7Q+dFAFdhrU6qYzgKKaSAr2KRRDHtgDP1vR/f379Y5YuP/VUiAvkRnWMTupqLaYGBR7
D4N1H2su6BRvqdT/4JCd71LOegHGzIuBmgtMfGKCOroQeLvKLYLkwyYDVmMdg4Sg4DfBQOqUnLaK
tuDi9T75QjSvY7AnezSMcTMLo4ayrOo0U8f0FSEDCS4Jwpp0QszJ6QzfRdc1Sl7geK44dyZNfHVt
ohgPjRyPUO7F7D746dT1AYVx7Fq7SXTcIRRiXXM3QY9Y0IWqyFSI0cxip0eZRwvYScmIOk9emWcR
Utx2TwamQw15aVfUQaMKkasAfPcuI3/Ipx+fNDuUxHhB4LFat5OHabdyVNm7Gi25u2BLFgPBVgYq
cmuCpyTbJvgGMc6bCKyRUL1mBgQiZYty5fgsQDpvm6ozHfw2c6Gacx8XhVTZiKLzGPp7eWNhvFVx
25wVo+D8+Tz/ZO5j4KZ6642EJYVsHJUeDOWU/7uBfRs82BtoyhtBnjExMu8A5CrI6wggvMk3GPjH
r8Um+WAcxKzo1Fnkz3FCrHXGiDR/H96jymbzTw3N/BjubF+m+p1ApIpryAPeRE1+Bd8fuWkCtTux
vuHFA5yJofzzP8vFhuGexJElPAwO8dyCJxoFbIQTPk2PtU2ypixxCJB3Fs07ALAu3I/MpfJYJyvV
wvQkmdF62PJK5FE6qZ1k2/URPz+qzWJ6yz7CJ5UyQUC2p5Iy458PxQ9/4/hAG9Wk7ggAzS5PvOJv
5wdAG7dfiCO64hX9Ks4Pn0iWMAdqh0tcdCjIUpXT61ArIZE8c1aKWkfKyCcOp+vlpi4w4l3g+YnS
kVLI6HmZOxjN4giBHzTNUwOChK8B3bC/Y7iKM6eMhRg+85id2rTi4sm75dxNyZiGta2WGNiUj2mT
C3mt/f3WnUxS8IqH3DZht3lYt0PWCV1z3wDfAbzXWRVUkk1tWS84f/UHdwFn+kTcb0wi40gY+aK8
ZVcY9pHWidkzB3xKOqOfNKr4YVECxc+J4qjUggIGA2f5GzVY1xFuhZFtXZJuwI1H6gCtFvlWvyFG
uUEqxji57GAg+zJ0auILhBOyU0hUgscvqdp3OAtGbc/vTCzPFx6aYGF4DcIQVO6xOQBuqWsqWOOp
Md1+YDawfgqgvqhhW8zIwVIUaGPkZigetWOBL8XMn5bYml0CC3FkShYqQ1NAylI5HKvALLywPMCr
xmO1mjnGie8szP+s4AR8gFEnk1qkSOethgFpb/e29KzP34eMyg5dyeEGWA+nx0PzY4Lz/djs1Gto
EB7ujusHIJa6vlNrRKyT1k+y8AECQyg0558cMx1iXRNI7MExiviiAXcRaWYAN/cqPdYsLsirI3LQ
5s0ttOFy2Vlaar+lU7d83/U25oR2HacHo7/k6skFUnSjZNOrQy6Wn+l0qvpmNUmmi/Mi0+tfRukt
umPR+axuPb3frv+7i9+8CUOj6IYG+tJxDsTbeWWV5fv3tdHvGqQ54MYGJeNer1f82nwnZ7IbrkFY
2V9lBuHLnz0znNZT7ce5lmp+SasH3U5mbvlGau3urxCGQ+KaKoB6rKeVnMqwlxipwJGbgJaYoNS2
62/t7pm+rbq2f3cytr7oy1CSEUxs4cqU3knVD3XIom4fclqOrOt6zZH5SuNJ6Z7N0CvsSpcV4Stb
uSPdv6YT4VSYHiVIDXhheGm32q+KFWjpoWJbYkAkmvIji3OsfkoSdgEm0jmU8zZd5NPDow0Tvz2D
FDuu7BMS+azufEFOflmh8hDqrmBju5EPToed6cQ8fBLGdJzstoqf/swH0VbQQ5BfigITR+bpF8FI
rzEIgdtXwtZ15cVxH9OBZn7ciOoJ5COfcu8GME8SEBnT2pbRmsnFC/f0rAaIzAlTBU2OQFh7Uus3
8aB/lzD1IqSIaDMdjyWlnkzDSAYXRV3qOS2SU/PYZ+iLCxtV8+w1MRqpf5ia2lUVrRbcqDHRVjLK
cJGgN1GzTHTOP/xdn9fF5yrVtOojhrO51qpjA5B7dfE68+wBal2ykj3MJubrJWw7Hcdmz4yhvna3
aVIZiHXFQ+wInBTtNvAXE/tCqsBkNk5+ZR+wr1wxBld0Dwhlyi9cbqeSImUaN0dZfFJBNGgSfDSU
VK8oY7XYo3eGa4soJ+s3b9IcZWuWSgjSPgZIsi0ZZojdfaLY1OpjOrOGUdUuUuoJ2lFCmhyr/eel
mD9pTZE8DgVLzwwslNvUqTR1HbG8yB1qrftfSZw/tz20L46DA2mzg86+qX/kVcJkt3YmFjAZkR1C
COm9B4+D9IX3aQj+q9n9OxNP2UNEaS5dYCUUKuynd95DfRtKqG67yMSPmaiVAamT6ZPcvgAC7Own
oDZGsQ4P6xUrpkywoUzBVcrxCkV6rybEACz/nYLzSlZJb1tU67FRJ+Pzf0fJ/haOkX1WHg0nY9xZ
ITqDkt4PmBJb5kItyZARPkandklSAt7XHd6+BFBMy0FEhKvrC+Unhxr5yKl7U4cTauFsY1YeL3qg
9wh8wKEJqKjwWtEOzSXu3+q6e2Gd0AZBZzKykXLPJM6hQKRp7I/x04u7eUzVJO7/Qykk1PPWsM5/
J6jo8cCqeRRqZTLo1TaKJ5rvLuq48KRDoiWhwQ3NOSp8bwivWvX8TceRyaMwx26PDA4QM5oO1JwP
ZVMHyweZploOP1pFU5XkfjESBDUSl6wHmx8gPEDaUQ+IGE6bMkxzQFQub2BYEHrYLDm9CnAJI0YM
6e01CvfVBRHoSFVH9rh3IuKwPfxRfnsCzvexfmW6fNVzrVZXOtKJTcpsxjsS30RtCjes2AaYDopZ
5X/ldVFMqb1DClZuF66H/Hc16TpoeQQZz001dQHzRtXN9WPGrKbWzMUZMk3I/9NATfbjtsouuv3Z
bo4QYJ1v54TP35cgHiG0WCXsSw9muj+ziZVcuA4U8nHhMq3L8oMELIMVawqto3ddidFz2mIUuw1g
hshqmdewknOvGPoE9X8Ck8c5Vcsrf9rAftRE38tygtDwtYLxDdhrxNxFRtBGzuMZyakehxMHhAlu
BxR6+KolpxbnO/19V6ttL8q+DpVeprHy3U6mtFWqj8WFu8QysFb7xQjEy30NVQWCvyqts5mlKJW9
6GsORmzdVZG8HZQ1BhljfSsUixHkEpYsTfoYMKmb8YN41OH2RABAOmOwVrK8F8IfVUdbaAs89Qau
xekfmKHlPW6NhsBrgtrSLNqllBqVLNii+4PipXvEQJ/muBVfrdWvhiih3V1X6dGwOldoGmUuZmZ7
t6AzAxClIEEtuXV5yeAwbfubbbpnUS2rl2eDdIpXYFzu+U/FXTojq8O/kxJ+hp8IJPvNvdXI5HjV
w0EhLEJ8ognfvne1O/PrGmTV3GJEOUXfqeKNhJSPGJZD9WRMDrSN/Lt3IzGovhIoPIzS5Ve4PPJ5
73gmTHjMdVM1c6EBOMCRmxm3gEZbuYRJanJjBdmdjoS+omFME/U/bILSBnGR0szKBzILChjnqmtV
ISK56pDxaqx2aXrtWd4/2A887ox551KxhDwquTEZMb/WSMtC1Pho0dvLXWUshrqK1Ehkx+9737ZJ
lWDgUSPp+1OQAuOzMVSf+wz3xROHTYLdGwtcHhfChPPGsIOkWuJyWsYeJti8/eMN6Kd47LG4gl4H
odIzVjfxmrU6yPApvbeOrVlpCXHQ1nKnzyL/2FvRQJ4HJ1ZeVi1Jv2UctuB4xvQKdPwZTqeHxzh5
UCcSp2MjKMm5httg4czBqQDOW8v2eRW4rrrQRUC6snPlXcct9j7SlSh1nthfj5U1heCaMgGTzcCk
KsMEOzKpMq8sX4n/+1ThC3xO9sAKw0SbWJiuavPbgymKrNUMCw7OcEGITTyhjTE2W9eGf3U5yJc1
5jLwhAdmPZ3uCNaxmW9ihmo6nLWSAN4aDwiDgxpS/ppUy5xOk0AypuTjgHfPVgdX2wCg6MYCLKy+
E4SDOnmfP61AsMxolhuAn46CFNfHmEeESTlIYTCYtTHiN9D0f3WMjTIKwBA9vW80Ze9QhcFPdoK7
0WxOQfbfAf+sd8d6fOgThDjxT1MmVuP/xeJr6Wwb//ZcLeq2AaAci2CUHzs21c8q1F9GJSKpCGhr
1k+Xgpm4xGtju9KeuvS3UqL+++OhDOs9uYNMuwiYrxVg88Oye9POWQluiNtOmcEbC2iOvqms8Hyt
MF4KCdP6Tc7ANYBzVMLQc6XlDuYRcwcY/r4h3HT8uwJF3yhI3O641bbG47YRyOBUiV7v4So/P/uo
w0GHVFpxmnZ9P9NMM7y8QFu7Luszal38FYbbOxDdC6uhAzfAKDR8mhZXvCK7zFNj4Od78rRwNGD8
q+7US16iQKaGUEOzYJc8U9BhwDzh5R8IjYyrNN/gd9am8tCRxmstMV+sYUjzaE/1VgkYr6tfMhHF
I2XYWFz8iyE7jxUotBlnN/YsDgNVmuI7QqXquE1HfLmXYThCGiEctt9YZoi92YicJgc3v2Y6rpwW
Egq9S8SzSt+eZU4u4mFx3A4ob0BZO5Md5U9O5QSKAgBxfBiHFrfud5mHc0sx4EhORKFEqRlyzJpF
FKpsbWd6QKcW4qiCyssg5DSOCD4T1BCcrL53TMN+fFGKha91y+z28GlloFdLV0LOGaLiydgaAztX
sB9YGwOloi/IvmycpO87LWkfG3B2mE+UTxdLQOPJtIg27C0Fs3q7Yl/7yhVDhGzzojBqnuBV0vT8
CvV0y7LCBChVgPs65q2NxIzXYIbrmto5lWreRGCe8bHBlUiwPKDhW4Ey8J69GoN/wuD61cOcKGj2
lRpWNO6GR9VWHTEAEKCxjar1/3jyn0wKs/inACW096GpjRWkEAU//bJY3m/V4WpWI06hvkTcA0UG
KM8XqcrlwxeXZrJokJ3EQZPmvallkAYSvjYSumlPYQRB7svgFx7Nb+hR/4ix+GheYuUq63SK46sW
7EgVTzZU0zej11dAztv5zGNDLaz3wBBZkcel1MG0fEi6BLoo7zBB+61gxFIVhyBnMUKfdCtl2zF0
T/iEdU0s/m/u4+i6UynoEYPaaV6UUesiucpuAbQP7cRO294AYGJT7d5scjqtvWrB0VGmfQKQnbzW
kdgW3jBVIn3iUhAKXqHZleoEQBtKe0lLzFsMLZBd8pkZ13HGpQltZnT0OwtnKaT2ipzsNtbMky39
JeeWE16JP+a68dVG0Ea96pLrH1yVvFr7eCXS6XdyY+YQgeSQMQqew/1sGNiVjIkXWcrVJZbFN133
r2wFdowajjwCl/Pbd9ss+5HkmNs30iNhS6Jdlhhjr+SBMvDwWww9UPoLSWQx0KwZYOJJjBzEDnTe
KI7EpMk8fZG/+gwKtcC7FWjuBpGb16fM/aTVNJPdmM/+9e7QXkN/d1LUJ10+Okl4GYPgrZ56+wv9
hBaK7sDHOM1ItAPnM2YlmuzIACsNg6NPdpuBWCE2jeyLp+T2HdAVgSTV/0bbR1kfd+ZSb/7zd0Z3
ulRPQOCNup4/F+Vzn41sz5lxhBU7Nkk423dc45eKQ3jgv0PJNEf+tlJ02bjnA4pAQ8CZ6v5H3gP7
0FhNx24RiFMdSAn5KMvtCVa5leWHhQ8s/4dl0NCwu0nFZEQUjfw8LT8Y9QuHpzG8XbcCSy6q8RYz
Mbgvw/powft6Tnhu9BZ/8Qbq0ar7bB01/UAMt0Y9I+YX70ogwghPamQumbgqMw3OGybf9bEPbkr+
r8X23U3tTk6ZnoCmsTzfhclpFztAyN1FjJL5J7NI1QHP+A8NL4FPVvtVYe1JE8zBu2P3S2DDIwo3
48Dd4EZ13DWw/mKkJ+iTymgdLxVq8erBZ1k8uapQT7KEeOqj1ATHjln0FkoCfqUFL01WX1Qr6+TC
YsOXZ3xxocMOZDEuRKKTa4pHm3lFK9DyJEn+ZlipsJK3ftiKADaLkHa0vCEQ9xY6IS3tnQVs2Kh9
S9yYCHCRFF/+0QD9ENsezn+nc//FZz2HWHqswfXKaj7MAkB6gyBne4WBRah+CMPEvB6kL3HpB75c
ztvzXPKGpViohPQzcRH8wjl6xSAOmAu/YIcninVsmqlRLXXzvsUNk/QZ/v9RhirmpY7L/ZgQCISh
e3umK1EqnEoFvwsawRXX2+WGe2HPqx50GmV0jU+ifhSio6H8aP2nSAH3PZRErv7GClOcGKXVV+uU
614OigbVaoma+sfDuXxROmb0c5yr5jfiFxy2ouyhs4OW2E84Iw/1vV4XS8V06Rz9sF6v7TrAc3Xi
FgwGbYfADXDMKgK+fNFhJlTa7m5WlNnKmMSKV//jC/7bScQiDV4j9cjGh22Q4QHu6O5F9m78vPXI
fc12S+qLJ/H5R6mDF+kz/kj8GHBRYwuQm9huUNsb6vpNSNfkPbSp/rOjm/Pu8W/cyjs0QbGJHNI7
+Yy30VQpOpI9bK//rmn7CkaIzKNAGai9DEURPgmN39gdB2xr0yuVY+PKFs/QvzSbmnIS/5pvjZ58
yA7q1hh++RemSOgQzycq2P6IlFn/tno+SZAkuEqqLlZrlA5KYLuEMyz43FYg5mCqZvm7kDxbWb3b
U7SMdzXKWn6CGTWtgPsp7BSzZ4hnc0qBILu4EEjYYoZGSWMzYYQfmvY8KJ6UQHn2fQcPkp+2LRz2
Cr6Onr/KncJN1/xpkraFUZ0BZ23tH1P3ks+ETR8tizV5mUF/qIkM+X4eCZX66CEsuch3fseNE83N
/jOr/3YFRwk/sdVZd4gZI7ItZtxxoClrlUlzzzSzb0Q4BIyOuLjbZgWO/jBbjuGI+litZ/+1BnW2
GnMt0tofP3xVTveQbM/tL0YZD2AcAo0OawERt+vgWMdqWZ01E737stKa301+ofrhFO6ukW+3ONQs
WeVki6V+Vtf0IpL00n7lAMU3NGbtPRBSgWN3YPPU5NwtF4ecNkxqg6jqGujvh8uPthKtAKbIf1i7
3D9PShrs6T5iMtWcepkd9iIrTUEnYl/oy/7LL4+iZVpqJ2AfRJ1WlevusoTf9tgEza9uF+2/ylk3
O6mT7cvPDjIs8Gxw6hWPGH8xIFanpymxD94fHwtninLMpwrffU+qTxdFffdVMFv0WRY4aIcsdgwW
8djnkblPE522dnxlK2OTP8HFxOUlY1PfjMHf+lgwwrFrKSuqMklka/0EzIVs2QD26uDYxOjfVQPK
sSPTs/yN1WP7Jq5twuz6jxmkt8KsvOhnISFWtdDFiFmPbPgqSVtlzZvWIsojVtLLKCcAt9A44PHk
sJ8CVnz5qvICaEHhU+6ZfQ8s78dX7u3p8sNtG3+HKPeij5AUZWKg7P/QSnvVwxJkbynY+D1aWSRP
Kk0hmnly/qo0o+oqiQEewVpyX2EAd2swccWUzqvrmKrCJe23YR5Lq+g+1f1pd59Nx+5Im2QjFyXW
qzoKeJ143DBsT6IxC3vRgKqDyUPeCd0rkAsAQuILshlOUKQ6naB6rZw//JVtO8EHrNOyRXzaejzo
+Y59wUZlFEmGHV1nNlG9KiP8AwMG1EoNxZbmoHr/joNrYjPKBAXkI+KwHFlx7QhSHm54kz9LvYOi
shoN4ZkTdDHkAm/zwtYo9czutJRk2Y8zD+pZE1d4NXZBBqrDBoSK0oAL3LX5iRKRcPQvpZBXOuWK
POV8GRVGSl3bpFsDNjXfn84pTKZD8Dk6Rseo9fUzXDybvF2o6f53lcfwBXZvsozJ/jrgd+i8re+u
jhNFhJVaiRTS/mu4IjEX8U/FgBekfj/ITUxEOM9rTZR8kow6i9urVRFhX3HCXPXcGeQxDIV2z709
qsDy1/ikw3nfqmr0DpwsT8X76qcYJO7GFzY9Z4fBdwbYLjtADEyKEx0NyNkV1gYXsWfL5wYrjQ/5
MeultV05t/lncGG8QH+JBWJOUdeXXBZ1BuF9kf5LYxC12N8UxesNaIhS7GgOHH3hE5DpI+8m0J/6
66un15BzGFm1ieZYQBNlo2qQIvfRZF2mzBfI8lfm5fbUP3mgKR4lct6wjac8iVRyUBeZ3ockvi10
qX08GtIM3FA7oznwnkUvttoE69ynhziiOdgWQx1XrZXjh4TLFQ4Vv0mKqhKhjjn2v2GYb/wRsJX9
10yfd9VI+arj1wR/hovdc/D9X3+AQjoYtPhugSD4CQTdbzP05GCRGWFyoFGyL4szNy6Sb81QTkhc
R62naDaWx8gCQIS11+Jk4kBaxxtw8tCtLYTz8xq18yOz7UQ3HNS21Yt87wtTlBsY6CBa9GyYdxwm
nVTu7bR8mNGAgw/rZkbOvSV042hbVvXh/komFBF16rMKDS6iXTOgKqooehgeDUojypuqu/H1FVix
A7vNYB4Ti7tNi7G272rmje8zfp2dLwske0xjFocGfMwdEpqRmkuh8HS8r4WQdgcbw+cGJ6y+WedU
VaVy/Kqugy8KP1vSVfzeo3bbULid9BWB4yZqOcS3Wev838UUUEKAJBmB6Hup0W93A8WNH/ZjmHtw
ylOJhJ6glL98xS+Qi/rrfBOgeHbvICMZCyPPk7B7ejn+u73ymG9gLqKGqX0GSH3GwpwZg1Kc3p1O
N6xGUbrj7nXaohIOfKhWgboUsTQT2YefF4Nh3bBgMPzIHKk/vHFXxmzMXq3qq0EZsW43dxNSIVb2
LfSJ252MKPVkyBf+IHUiJO+IpH1HRQb8cHZRlswI825CGTzAnEyJspr0K8FR1mevSBADnKHwDUes
TtKE5GyxrrAdR3b9nEur5m6XUFlYrHwuuYlQvfkYy2EZXPWbRucQvbEYUTOQBD52C5strwHGhRbQ
DlDnZoOX4cO3hR/nzaj/pRwwT1AFTtT6J+mO8nXHVjdNR9/kcethNIYqVQ4JX5sQ+C0rdeh3XyTX
FJwpHRoQ/wRN3vilKEqRnk7ts7mSlpkVJWhSSJ0D41ZR7WS2cBTDf/5aoXhk8GMAWa9ozaELqTus
OL4F6HGJZHHb7TIcq8ZBO14ZeQ5veRSuKHdBK/oFFtxboGw+OABoixqxpJf34jJBDWEHHI6sksOl
AQl4Xrf0AGlh23zVeKusK9nonKfX4feQOc6EhgfaLye6rybaXP7XHgrS5pJLFrOBy2Ko87J2Fa9P
lRKVruO0uAlo0zZIa4M5liwJGgkZkD3hxgBeTHwJMpD+VH9btTsmGqLLUn0+1+zr8edJn3Qp5xvE
TNhfGZC9JRoc5DLeffBlOjS5zXexIhKwWufM7VBXSj34P+7zV/20fLJ2p9MTK+bBG63VxMw5I8w8
0+azkaFVqeY+5lqcgWwZw37eMpdpCyJe/fnKKbJJz+C2LlQuwqG+M3k1Ej+DuMQpXYKd+4sg8uOO
2lgAXArQHnwqTc+19x+nVyo9690Hsbl0APUDhHUryI52lolrh3+gISGwAszn+hqkAg7k4WOUmIuF
8D4zcfZg27BlpnwVAJebOEwSHE3UENS6tyYj6CyeQf5OxaS3MstDNm7uHciCU9XkDH2KiVAvaRj9
EZajILuPm4WC4xJ7oxf43RKAvQrQe/kWnA+0HcgnE2vE+Ny+slTWVP2wQwOzDOE84znU0VYA32bV
NCEMnn/i1ZTUC3cBGTlS/3XRJYukEEmUTbdAqJF1jht/jpkukHMMB1W1TFcMuNKMH8d3/t4PoMEJ
FvBzH5He1Uht0t+dfmEHE5rj6cH9VpUcBgjlFh/7/RYsY+z6mG6iIcsxNtOcs/jZU2UjQLAWjLmQ
4wHfSW1RJWtEncHCIRqAxg63f3mBud2C8lzyyS79RPpV2c6HcfKp09tsyD1LiVwmmFXMMJiiWVCz
11z/HKpWUijf3qaqZSz+VXW1AT8sDvX8todRFyo7FVxC4g4355vm47VN0YkKusCqCIucM0izxD/6
OGMW8bm9DAteLUKyxVVoLamx9LgK4lzu54bd5nIQFhmmhCy246ahGkWZMtmofXXzOfLhzklyPwrd
5NaAjvESp8ULfMdDW+HME/9u3aGIlaOVtN3MrYOAFKa33BOQniqzYPShlCGRjQ22V1f4D07Y8gyw
F3T4grgbWxzJt98ekxdEiuBWRZeN7DMrlMDV3NPH9XVLUJDOHhBhjgG8J7H+McQmJ1jgIMSd0EQh
PaQINiquMIgubHedUJV9EMbrOlIpCuWlwX7R57OmqDnRmCxxxprNUZYW7ZTK7s+MFmbhrQeUpdy0
14YDVcWGmDvcgPEanxi+TcjhqOyZrsAHsCLTdBRQIq/7jua95YpxQrwZXbR41qX+5gel8jwvSnkF
nHlRphoOAfLt2/J4u3fp3hFPJ71H/HKFZcIgHlUcTFdERP/c5gAV+z/VXGm/lIHj2gbV1Z6tYtsI
sh+MrQAgkn9ZpVnXqtz5mqkLefZIQb0m0CRHRz7O98dnCgt5noQMLnXikRWJ5S4mLv6R2OrGcwpV
ZqDK0wP5ABK3ipqlEadsAnxRtOQY0St/88cOxeDmFSszJgGmiV5HwHAD+NUb/pSv1manqIwcBiwb
3NT/6074Fuo4B0eurd0K/o3b55uP2VSwPAjErtdJ4i5vPNnKQnHzGVL+VlaJ6PzRMxLcCdHdyaCH
b6IbWvpRd4vmg0l2OQF+JAIP55XByKnpSgLgdUq/uFIIaEofvbk4qMxQ74AXqt3dZVizRkmL5v3N
kzgirLjUENszJazQpOm0n8IvXf/wsNjNkG9fErEDK+DO5TJAx4Upi/ksFPsP9T6m7GzS3/L0Q9Jy
tf/5+SQrdTO0kv2FK5OJIYfeVnglIXY1A/dj3qiP2fx9q1OhByXDM3OS0TPB9hjq4+c0mSyqBUpt
JCeSwXknRgsfZPEBxUEgK1FgMACMCkW1hUJRLP1UfenBw2qdZJd4PLD5Y78vYs3WgkIqiMo/Qu9j
AtADdpFzTSQrEXZdHUDdLEc9kB4vMCiMqYJQhI6EKL0ZqcqxtYkNl/KIWvWOM7UP1LiMvjI8ndVn
JVnBTf/yAJaMZHhIXFh5hiEVEqwKkP9AZVBk+WhBWnQRGmG+szSvGe3tyHl5pO/NN1Mfl1qAUt9v
sPzMHq/nqBJHjel3jZHFPGAwNsUOaAfWZT9p/7DP4t+yW+kJx7xu2Lxbew8RulipVjmzVtvvD0iG
upU5dSXHIzblMekSrkVDB95Dv674nZxmPDjgh46nAb1J4j+8gbQ+xkUOGQGqGbdW755C6tAteae0
kx2E+yMW4Nt2BtpQy5fmBTMycjc/bC85TUFdBx2PAAi/S/Qx2/iRVs6RnJ8903ThgN46kgJtaqXG
XqxGMwS1M1L9P0Ncg+25/mE5BMoSeYx/42/zwxTtLBu/ZWxbST81DrrWrMrnh+fQTn9pWfKkMUPf
LIcMHYH6mfwRHlswd/BbKvzntArG4mbYdoG/WrYUXyl7fLMzedrnsr97zDDvSPJ5JSC8xe8QOZXS
ZTSITV4mxnmDRaOKG5jCjQGpZ6WEfIFUIhxRsWn4WsCmeeefUX/qczUTsSvNjaSTza0GAGiFFigN
mIp/hZ1A3u3tzYMBs7vpghafpA8TQmjQvrWcueTmDeK5ijFDd34F8KKm6r9nAgjdC8T/VH8PiMPw
df9q8+f81Zwl0xFS95EpPobLYWSXFnnTr0b/KVt0V4njV4jK1dSFE6OaMrL43AVurZimLBSuvd9h
s/seRy1NyBHvTUbMcn2SOCSdLyV3IFJPcxHWmpSDu5lNPySOvIid8Z/iiqi7GOv0bTd4LlBrAm3O
LF80Isimp9MK8EcNihEw2ca73IKvEaisUSGBUMOxcPNycbmHpiVyZXgljTB57EUAq8aEcPex2IDb
1rfo5ghS0VmX/QKcfvwNafk/ED+KxjXcKmvbhNQ9QRJo2mWDYYMVqTgsguo31NfVUL9nz4dKOWmZ
roKPIXVp3Q/vngD8xeLeDWBiUil7Zs9uK87wR5gqCpvYqTjXsBrdyd5DSgBZQdKcIp8aO0PC0E/8
g71k+dIyrmwaQMLLrxGdeTnjQ0cfUn7OF1kQYrqLbkQqKpAMIlL3iFXhQFGV2lxQT4Bi7SByrKgZ
GmxDBHTSm0QZE8oUbE93F7/67DACbzTHPyaGXNrULh/ni5rzuY5riRocJD9JODtmXRK5aYSrylHX
L/DbeP4O68VsAMcU7/XH6rjxm1N3eHK3/3gxv6T9FxKaTbbB9g8EEbuMjPipY8f6+KQ4i5P1T730
+TlsEo/jit3QW5XZmk+j1IitTaXXDNMFqfti5TfY4YH3RuNHbkw2G2LtuEfUGy9lDaWsPKUqEA6/
SALQ4iA5YL1u0vAcag7vseSzTP1IlThHxiBY0vbIIlOTfgnjSR8v2HJ1llYBJKAqwpeqHGea32Dx
61Lx3BtkQ4nK+lam0CUraQqWEY06PZsNjUdXos9wK3MEfLlneOKx84zJyoKNwxOK2Hbd11aByHvW
pWDc2RfbJLSW9Vg6x3T0YhgBUjWbjqvntiUkGI/lX6sJ3iCvnRTiwIZswNptD0RHGSB15oTjZb5A
QdbnUKm0+utIo9guE/SSkHiPv44gn81r517dRzR+lMmR4YLAiZSkT0ehfjE0zLWlApHupWLyLB4v
IKHjPdRG61NOOY1Lc1iPuS3t3eRuGMs1KK2z02uvmBbd7ClH6S+opdn5ZtU2qzZvOLWWDo1Nd5AN
Dl/MC/QQPmI5aYK1fwmrMzD6TnBZy4tNATQpmQ5w9B0M4qzeXTjxj/r2RfYwaqEsYrTg7HqMn7pV
UWQatgC12Wu+o54NBiZvjJRk3YF7Gc9J5vm4nn4/oS27fk87kzgBfHyefv8uTxR88iXAqsVsVC8m
DNhVuMbXAe6MJ5aRt0RNuNs1SEICoA1B+4bFCg9wAoXmUI6/6XHmtstqgQbO1YOwGG/wPrPImMLu
l5MtgAXn7psvYdpTqV2Hw0ZxZq58bvELmhTbtcampWifY9XKZB6EA97Qls3ZH0KRulVC8gGKRJ3m
/VhIfcSvuIGIRDlEw2oTRXDidPhPKoisrXB+QNqrptYwswoFLlRDbu34df/kCJ0wCQBFHePtrqbc
5qtMFn88ChnkD0yXyhxicuWRfXsAMqc1Bno3WPUNXXiUfeXkqrfzRXEEIaPsW228udn0blp18dOX
BmpSe5CJEYurFlkNhQixNtVztrMywzmQG64P8SjvICQCpcIuyYYVgl9w8nv1suDo794QyJ1E0zRZ
EGimyzXS7OQxuXJXjbxJfKDw4BY1LZK6MlPKTH9v2DDrUomLERNDmaoto2DnVfS/pCjPB3DcIdpF
clVzpddjqLclx3uLlCxI/ykCpGom4yXVve5uOlAjR/nTlTuYqTuhKvkmMWSkypa5gZ3Yc8J0kq0H
/7mmdcik3q/Sz7aopC+uTktBSw89vMzWDwjFpyfBvdqf7wUVa834lNhrQC3ihsUpuQ2VzrUYyduw
rngCtXaZP5GL4vlysITWx5W+/8sY0E2y9Kk6iJse1X4kPPmTFgmCTbwfHQqOmIQVUxmRKoWz7CCT
bkWhXFgeTjGjg0ETtzY02eIrcR87yCBX0yB6FzcMTFRPJQLtpT+If/2b8LUt4uvs1zkrHKHf/FbA
QpVa1tvNiYXdhwYYXfeCo8xdDBgfAT1u70iwQUzrGckMEoYDW/UI69fHKURXb67yLQtKIZvi2Up0
fjy6G/C9czTEk5w6MBSupfprSDaIP8eK1BvtSLVdyyHeBow2iG4o892h6ISx5Cg1hIEedFX8obn8
/ECyg3lGSqL3Ts3/ICCRBScI66o+SePcX+BertnZZMV7YB6O0MxYBv1/ab/19Kg3y6aa7gl0aT/+
gzhJbkhfZt8Dy9SW1gxV/nW2q/9B+H0Aqw6AxP0YJ+1rM7C4h6JG/OBWEdj6f108OnbnA7I2pwuU
6tkPb/+XlUUr6tMJbQTfxfQS4UpGLmfeS9POpAr6KxNDrBXVQu/c3Ho8rEHUN8KEDYNl64pfiRpY
URH65p4IfmrbKL+1e5zAgU0h4R0QjZnOaqzQBAawqqviUYdtjPpWzXSqKsQLCK8pi3tlLWA7dBa0
m/XFn4k8kkfpq5DUmbgDeG1bG0brpMASX0+FtvsgCYpz5LpiIGG9ru/Wgk2yDFEGGP4uSiulAEhu
F/0bP+JOznYE6y4b6qJSJVl9wOWOcFY0r1Di0GfCZD8s6WjUUkAPTfXpQotDvFdF2VKzvlowxqa9
bBE9yPo6yLCdFH+snzgbd4ipvO5j2rx9EnNQrjoB/ExcfJHM/FwwFAZrnj8F6Yaw0dfaek4CAAXk
9heWtgoqhi8qXEdxfGou6LGQ4pCylKSY368BwFxNS+cZvXcnh6h/RxOJLc6V1WWjAheMUwWtXkfp
as5KdRtPZiyDtt0ao3r3fcANlUXx3kLTQ7qIU+HviEgGlpDaSoBEF/bZmKx9e1EaIZPUl5Bojro5
ioPARi64sK2ZOdV6H4SBkRWgwSXRWM6ANKvPpiA33BpBD0lGQ8S4d+99NIuq6katJ8m+sy1fGcLU
SwC/y8zzSXxK3BUirWMTQgF7ZgRVcsJLR/HSGoNBb+szjjGNLRX+OTbWJdk71e8fAv+c/cFxREFS
Zx9SMKBUsFKSx8aD3KTXwX3emM3M3CMkhs4WmEMg/AhBx0K5S2guHtwJVBPIMkib4waH0aAH9RrP
kKO6++/PKn0AOEExmOIMv+kJSm6EFBvyWo/G5b/oc5dDrvfNA7Ob+TZvUjOYid9Tj4j0e4scyCn0
pFHTE5MzRRRNcu2gM5I5s4HjTTFzDgVLoFgrzVPlH5Hgzwcu7Wgtko59JfJxVPDHG5A4WpXTGugu
0oh2bxhsF5ODKHqjau1tSaGCArGsFeM33XKEE7EraNwwCTofdo62oCv4qrrQqsNgLzzw4ETIE46s
tNJMlRY64l1xG9HGOlW28caJO1MRCSav1qo6GAWrR8YqWvd+2acqQjA8bchsKg4zJiev2OB8NKcY
N9aT/wECuxV2T4ROuHLFD7duSvcoGYPI+bTbQUzHIQturVlhyak3wTmiEOMJ6R5TKxW/R5htfHWc
9uTpK+hz/8IHQsxDX0EHMLD1I4GtB0K31YG84elhNk9S4YexCyYaeazc6qO4sC35tqv8zhjVar/l
0QT8WEF6MPxClT4l11F5SfjkkCupc3LJgzRFapuYFCiD4EQQMQj5D7FQ4CzbXBFz7HxaZFffpey3
zAAnVV6vTAw40NyupNv/gHYV2f5nj0zBuGUa1HRko6mFQp9fX2IplJcn7HTSEbvU+lYUKiVaP9q5
GKQDnkQurCCZ1NgVlr1Cwvv7K9uZ5h9z1lU7JE8w9EPzFUxdWJ88Rmrh2OxJ+WAeBBIYxKwC8GPV
KuCFIM6poH2zxaDpRQG5+F1o3wC2cGNfrLRJJ/DxaMAkTcQBt2fU3vVj1is1ltCEWaMoKOFMRazg
CDk+1A+YX0m9p+W2VYhdO+tUm/YwZhTvKT62U8KQfT8H8mRtydsKuVjAcV2SEsUtJjiHDwClUuVk
H2bDSuF5VvOQAqSIZaCeqjJEUooP+O0GG6yragf20oFEe6C/bov5SsbCSPnQy4oxc6KFbUSKGokC
+WJgnAx/HIU49QLfQLaz3VXfHfzZT5gJKGO+cLY78iwKrjZ/McXmyjqX9x6ZFtp6Ay5pQl5JpwAE
XRmBmoHEGOk5gOOWZG7+r81QDRVDnLg+eRmUSADNdb8+VS3+waN5BpadSzhkrz3h5whSBSjURjea
RMXNmvesgHAVODx/ZWw+gClE/BjcmJoeJRvhluuwcOm27vGWpf4GIBTIE+JwwE3OggJMcKR/Y7LG
/iZwddoGoNyGxIj+e/o+2av/rYvQG5fgBQ7NP5jxpjqAdkGUcrPnDvoFHObrt0f+38rJ9aW7Yq+B
aMR9UlOR4BqamLBZoDkUQMrwQuUZvngvCzxhUZWx97+lA0hK6fpWyWKoty3fy+z2A/UlCoQ7KbON
Wku23CuoiShUPeSdZHP3sr1ZpvgHQ28dMju8+MR6+g5EutNSEDUJL9C9Bz5tbZdyDR3CnxR5ByfW
gtwFtQs0vXN0qW3+ep7AlYztLZVUpDPJFYjc8IEwON7NwazBel9SwImEBYenJcherz/UfqRwXWLu
QiC9u/0MZKXA0Z8iZKDWIjiCi64u5EDwYzMpVIVoGwmeefvqwhVgo8GmhUz8XqtDo0ij44VstLgS
Z/12sb0Fd1Y4PbL6sg3TF0fkyQYtcDXGv47OZeBWtG+622mVyDIkTe/5u5H91WWg41FI2AnkBh9C
SLrCabwj5aIX/pznd0vXDOiOTH8orhhkaMSPDKFBC7iyBIx5jo80tX1aJ+TnJu8/Y6l3U9ct4pak
Su5NlOreHc6q38RnVaI7/IMCXjLdD3uRRtTYZQ8une9Z6/B3nRhmIMK2Pv9tqrl7zSGLZ/X72msh
oYD7+De6zLg5C9RzmOT9mnhttQO9mJLtgazz6bxB8iUmp2e4v9G2QsEVDf1yzK91MTAZeVv/egk6
xA36kIVjM30mbQsuxqNwaQWZja/stHdMXvgO8T6DOfnbHWhX1hyrWEpfTUs75FmVMYb1xuZy3fsp
PGUQr9dp4wg+i4fgee5VPzC7SFYtImZIQ7SpD9jPvhaUFZgLOLqdsuRAjCra623hcJjfPExF3lKs
ldOnYiWA0GhV8yKIgE6svgv5pln+ym1DnG3pJXOoDnA/1AcNl0Xp5rT2buVga06G23Puk1XuYJa6
qxKTXLHND8eKMl3i6eClR7jwYu4kSn7MIMLdfATSiChjGZde9EnxhfQ2W7jfOXb/jahbh1mb6TmG
JXSg8/1xTrZwLlzW+6niK9OznKtK+tVXEtzrUtyHMwSVpFMPbsxT3jiM6UgyxjSIOxZL5oKtQAR8
ZY8LzW2XvmCbQ0KlLH8Tm2FlHQpwKnEY/zrLv4mx5y5qS/aHW3p/NJP3jJYocfJjaqMbPj4oMnDP
wpkIMYQICyrojSsx3RVhGMZZVSDP4jArisaZf5Lu718kusTwnxL3JaY307VAij3DLQ8Oh6PkavdC
yIuvca6g27kMYD4futzXhgzZPeRuRcC6eyCAZS0DbkOASPjdstyeidFQM3oRvUq946VW5CD6a6b+
QR2R5N6Aq84suiIy56nBBI9l5Z2xkhy0bfL/Bq8zMmuWE0e6Q971t7cJGfJhbyfuBurd706wfhx5
B3kjN/wlX4RtFbbY2Sq5S3yhFjsx2NDWV0Xjha6o04oFts8nfe0eABmOZq6ka+jSntTMPm9Ah9wP
0kbV4+hiZf+ho5hO+H6PZgbXa9zw9Hg4oqjXva6/olxBFUbFR4LEvMDDLK0WPMhrN1u5mReTCFLg
3WFt7AxgUyT1A6bVzcL16EM67cpBZjIQa5uYQ0Xn1wybzY8gaNzvND2vkGvEThK2q3pdziixN2Vr
Rmn8EZxDFpfwcsEYfuuaMF5n0toucothpCmQJtjOyIlll1ZlhTxAxrEUiRBaWOrJjtXPlwPQFaW2
tr8FICOimQNg5/SMwPkLI1caFR0zbobow0NtKUtsVZ2EZEoLZDppdsfABnTiU9NdGdd3oRq6JmBK
kzfg+pHXW7vkRal8CU+At7Zm834GV8lXGnjX/mZqV4lpPRcBFZG9vgX3xhA9ADTPtRYQhIQW7UzM
rib5NxK25DsT9J468qVbd5U+eQTc+f/sDRrtTA21Bt51Noi0wE1ikjV2r3oHMUcXwYvBzFG+X8oN
6rRYrkulTSGUKt0bTCZbmwzSYunfIHxuGCuujVNVwebcb8TEBDfYbppF9dvZswBmED1JNsmQXPBo
XVKA+JOH03CefR+RYJoCyQ+smPC2pFlCH6wVMjaOvACiXPVwrFMypu9nw1ufL/SMfmSAIJ8cWIMp
4m9aEskFMMN1K0+vfDKv8I2+9Wnee+VPVmX35nq7I6dwpLVQznXpsB3XYC3PPrIg7qdAKcMC3PSS
mLlA1kosQHMvOpnYYG36owt3+4bLXpHl/Pc0CpzJHeCjcr8GHsDxUjQw36aTqI0CxvHHVJXbCjCP
nglZJ9rXWfJM6Zz1JPXGFQVc+PpdF25w49getod4ijNm0Uwr196T1zHD2tTabDyEkdvLvkTNBQUg
l+xAuaWNlbC8WHutfu9bTJfQF05XoJfCvuu8kcobSCGsX6OtcJxUGT8OFZUJFokw762j+wMvqbUA
NEESbBrorS1ltLMBx2Qaf2/KtorAO/LCR3IV+SPiEg9FNT8EELBUSRtaNdVjbk1qDC2u9e2K2amu
XtAqvQav6BGlLHo/PMCsU9P4PZQ5JsoaLXThUKpdQBFrr+r2FJUl7Nn6vgnySLYUbD2pnTp4Ly9/
daGfr4J3LmsggRAsBopBQmnutW6i/zplpwLRI3Ml2aY9KxvWmFUydhql3r7LDpvurcNqiYxlcmob
14bwZIPsi3rEKpLLipaHIRPMo9kOXGxfMPGmhWLDXDMeQySh8KqWpmmYFeCgSKbfg7hKSesknff7
3yBu/QYWRW9DEq0U0o3JV/9u73df4tXyiQKN+BUU8EiqSjVyNVTGKggYyGnhZkGsAyoLSW8jaMCc
6ImqrAlmvp9dyUrTk9Aql5ek+h0Dj0uAZSW5j2+SGLs7zdvYX9PBgV5qMP8wx5vQufFreeCXdhgc
H3USMGR3a+BEPipG8P99YamoS4/cmsI6BsdzfQGoMILSIljY4J/GMUwBHTlWXWJm/QQfnPf7o3C7
8xBX6Q1SYHq4zag2jRCCqsaB8PSaD2Y/zyI44wV3sPDyixkEg1/TUOg/CPlfyikua+DWxauUOFK7
LflY/yBuIK0qooMxXPkFtwstcJgce0Rxxq1COeYPjQhLejLZGCvwLAAwVYDAGpFHFqJOWsn5TFon
XGZpjdcMgAqUT7ZpDEe6CspmJiCHzZafLMHDlK4DyKgC5s0nwPnuzPQnTGYkK2in8Y5/Q5RMQdnB
xZEuXeFs6bF0LreEeBE1/Vlg77N11LEQWajodOytxfTkc22UNZ1PgbqJK22unr1vs/BpjGjhQE5l
d13mgc95HMSWGtQjg7KKOL7qRcJMDaj+sMJ4rXbso/VryHuwOLRiYzgxWKh7vCN91MZila398ii5
YJIHS/pqZVFwvU6KTcKPoS57cvqQALwp+7W6cCbYbXX9I/bYeIcQ45NEq6GGn4jK95p263oT7gFn
DheAR7gvSqP3UsiLki8HfsmXZsF9r1v/JV2Sv2qw+b+QX2GQQobr/31j+6C0QaAoNYW3naMukqzj
5ExYVaiFowWFRiI6pO5TOULxwzwx7XyZDhTp6iE5XhICeUDAlHRVIlugNfERcAOORYS4KVfFGrSg
dATp/dnaq5zC6LsE+Yeuqial6Zj+zF8KkuD6n3UBn/z5XMMDgqhjTzuGpq7I4uOW5f9WtLGxZ1na
IHQU2PIqlZPUPrZqTqvTsaUQDQgVUmUV7+0m+u1xZr+3YA6QtrYIHOaMxdLlgvkQRWvxEKL3LJGf
jC04+y/youe5UaqiJyf8aJ6fjdFE1qv43theoLjWwNaENGidERaAvW9fmBvn/d/zHdKTobqCXQxR
IGA4IRVkb9e48bOrc+tonCOHxByPSVHDMW5j8AIl3BIwLOFq+kGoRRav+aZuXcsU4U8ZLoT7neJO
IyS9tMFFiPUccx7UStGCnmoSXDlcQ7Nf+gndfuECudgIWREU7Vbla9SOR0QdjwRvCwQwAeAxedSd
VGWEzCK1Se3aLXZQIs50q58gKoBmZs97NxNSUL+bmEuCUT4tfNFaEAayyhmQomGy+h6CCJUCdpEV
i7Rqn3Ne0mZa6AkF8eL+XOrv7+5+nfsAYIrVMGM62R6lTkV0sMMJK0ScKQp9Exl9QUOF6sHgPxds
Hqf7XYfWmXGHQuSVQOklj+AZtvA40hDSaQsiLbdOgOB4U1tHRFZe1WTeDtjOrxPEXfqgv7t9XwBe
ubz4WWCC5WZ0hVXUccHfdjrGKasUsicgWrYnSThMtdvvD6wtBkODd3igkdhHmvZv3boyqLJOrPYL
1UwnVIu64Dqc1WD5bBF09IARwlwz4CDd0ke5lnIpyzCgjVekVWJhI/BpU2R/CZrYjZeKWIJ8e70+
8FzWO20Fn/EB1Gvn+UfHdsd4Za12GzrcNEz/Whgwt03Ow9J2iiseJe3DylMJosjJLSOkgD7xI93w
kN81SKPwLjJwa8qlJIaoLe+zrLGxo4wtbZLPn+ZQnWs+haXvmiHucRY7GV9O5roErwMadUE9bNsB
cy+3nPRViW6FblGDa0IMtXgcWzbsDcVmHhGBOmH/Be4u2gtua714dQucX9KpTjU8euyunEeMJMXq
96khHfeZqqY8XqPr4SBF6JBSugazCKkkbw9feFAM33ERGGq9wwlTozE0J00NKTBvrZE+YTsZyBx0
WtknaP68DzNuC9K2LxpbcCVQb5gTdGiu1d6LftJM1LAFgtAeNLnvbjQ0T+L3koKYHTkh9v3yG/tn
XCb6bnsf5VyB6Q4prmwukgn+Rojb6HZSef3wA9Y8QEHOcnKGsNd+3NsHtxevYuKgjul7NbbXBceE
8yBqeQGcKkcgZ/uKLqzEa6zHva2lEPk+jC5orwBGJ9ejPdIdsr5+ChKSZOWswrgQegEBsWRsZU1O
8zPqurcdlI3cMK+Rnk9wGqA9PdwhXNBYBtQqj+vni0GPnPXu9JKv/P66ZQGJ02Cc/oTbST5Zics8
iGJJ8u6UaUNOyK7Hh2+HsUF73v0Xs0yNjSywMVnTS5269CAKa8gSJ7Vdhg6zj5UuhlS5yaz6IEC5
WvH7q/gFWkPYGXjRChkEAPJVdfwUKpxYr6yHomnXvqusuVO6GVanna48eQ5VvNT+gA3IBnnplZZM
QCXSLMJCj0CTFs6Za3nC9Iy+JvfPP0bic0ACO8q3E5QeCKJ6iQStt5U+voPfTTKbe3UXN09kpWS5
3+5L+Zh3/IUH5+kjjImwSu0tdDfZoQQsaGiT1KAYADfDLvUADaVLyJxrlVOnQQQaRguCyOhDkHow
V3j/1ERbCLej/YiyePrFw+5wzvKeV11fKyD1BA9D38C1pVZiSFJZl46WoH5P4LAatr5bianBKOyB
1geQRhgk9I47dukYAZNl/Hd2TpK6Tbmdf1iTiMm37vNdRfXrm4QLUcQpFQ0R7ETDGlWpGFsSRpvM
qyhVvxuTppgi2VVGOLKnGwXnj9Bitdb+r7jAN5x+orFri/50AZnLYYh1Zv64Dl9lorbUM/qQLmA2
49Dm5Ed1ZHUcpV/how4qaLL8ZzoOjU6M7aKxDMKRtvVqJHL+ZHUCzcV8XUMOomeCVFkHBanQh2fO
QTe7jPmVce9dOjutVxf6I+PRuCpM8zhVAnpzFOq2IjGz1Z2P7DTwrmlFUpVSXYSdBlkB/OKa9+q/
iG5LKM1oG92WSAgXpmH5VRA7aYt/VbkFNcPlMSci01xUrOlZ8dkRlv+8os82v+bpKvABPGBNba0z
DDfula0VfhZpKuwlRGENLiPfr/vo0fr67rfY2b2TLt4lCR0cJOq8/908Bp0paVfWixDe4XSvEzKY
y59Y5mEeA2KThBQwEg2+6xRqfjXrUFdCU8nSxilFGzoI/p19ZHswHVnpKBT0nCEFZDrSz8K06d4v
ZTl0hzdxOyfNQzehDbSCHsQCksFlaPZX3I3nf6Vdz9odVV4SfYeBgIgVWSvbaYVMYUd5fnUIQb0c
224J/iW0d5JektjscWSLJuIS9RHTQP6HxIkRFLzYt60QIFwbghGwngqIYoHtKnYv8/Ui2MoFRjLG
77XudlmRjpY9r4GuFwjmSOESAaV4v1/ssaPdWvneCxhaDxc7YwrRSnLWsRc/Q36xXSqyOddo9mX+
rjZWgT+ZVj9EeYxBkTc/8/WSFwuqaq7FyS7Y8OElCbS6xBJCLkSkAYiDEOk+H3Ud70ND5xlqoKOW
cq7kDdtje1+wIlGER3htrtcYAbQ6EEBd9FLAqaJkR5+Kr8MloFrYc2wVbB/f179H36fA0O38Pgmt
u400gxuHKNTiPs7qbAPhH+xtC1WoXRxI1uk1Xx5Q0NC/GuoeIDLyzZCC0iBQ/WTrliKSRSQ0atTx
DVQAG7ANB2bXXOXbudtN9Ae5oDBG4nPUc7zzIkVwxQ+y3X0CrfjhWwky1h+iXWddzwaVag+Uo+2N
FiCJyqj2YvG4Eo23ZD1kUN1wfe4GEQctzbOHy3chU5FnmT8GfoGG4w7K9Y3X8hp0pQkRUw1aE2Lr
2Vj8VE/yw77rfr2T1NfLKdCXp3fNIyCBpFd/AwJvZi8Q/k1ykODFqtEHWUpt2vqe0h/yv0aZddTE
2D7HGZuuV2OSMSMqI5PJb4NE763QlfYCYEpovjpgLdDahbeF09RPxQvuGXmW8glZcNVfk9KpdGKS
PVmgLOlKEkhD56OklA7ZhntOwDeIGnfTPKdMrHzBAnk+qSPZjf2msGCW/JRVbOLAEGjMqWqEKYPL
ZVGCWxWyOTCP9G0/zBLAEoyhTtFXQPOhCVju6CUC2l/gO3foxPuOyFtQXlAHuCJ1BFlk7w5bG7HS
QOwKd2Sa7HWy/Yi1Cz+pxUd4kOhBMgmbHw5p4yyHEMk8bw6K9uPPbeF4QuqSCnUdUKz/roPptKWY
6j7TkjspzdLVrrriQ7ghEEFXWyrdA0j8jOeE2pqEszMUgEWhjMSBPobFBfAu/P/6LYVKyoAeGYTc
Ky4thHQCClxGkAKN/Rp6O4kpvPzmRvmLdEoZVyMCSD/o6Gj9I6mOt4u2XV3ZhRFbaEQVIa1+SZGy
/4umA1XD7/8K1qFYCSY+SZftqHDxyXphYOVbCzw11kJCXe6Jtlf3NJhfogpv/dZ59nj3HVjvnxgU
qyoYfhYpSGaGojRB8oSv8/leAI1sdu7xZ1a8LXN7rifVyMvDfocYyIZvbs0CDN5zsAyGpb4xCeLV
37UKs/e4kDRczfFyH3b2xoAWo1KeyPkNpGt+iVgn+0RIgjJtcfvK948TlN8zthPaHHAEWnHVKA9G
McNjdqQmFC8FSjSJqV24GfBruUz5APT0Fcv3uP9lYYIwXem/WpZ6DveaoKlOZ/rP0mymWiiiXrvK
hTgviENmOQBAUTrrABrnlA491WSr9csdGlzjJ4Ghu9GGXZqTEW5CVvxptTAh5DK9aUsQlJr1dz+j
ptyeAl3QsAxS7kNnX3a4NKyiAm5kBdCUrIKdfGeAXB6yr3Oce/hOzX5fnp6pBTUcCgw3XNsJ1o6M
pwGF0Mvga+pwXzx0ClAfssm90cNIn4VgmJjfBiY6qs7GuJj2vqWgyVv9sDmxVgQjAwpmLYcyj98L
BFpVLmbBcZL7FCPBN4dh/VjaGYEXv2o5VuxLVFHQEd1mWmfB+czRYVI1rh0R1Hbuy2v4HVbRshu0
mtR+pBQCxlhxDm3PqxA8prrRFyhl34KzhKDcYcHRhTVWz3OTON65Cw7+Z1UZmPdqtcxq4gjfh+8e
i3q+f9+a/OnkSDiBIFA690QFv5DVwlOTyynw6GtJfWeVu8KURIgu4Ee0rA0H5oPnezfY61Y6oXRM
QKUDT2+XaBbiefaSU14iQU9wleNkZo4Muya09bv/pbnPDg+HCczu5pLcc2dYczgdvExvSWIMDIB+
QuGRf6POi1EJyA+8K9N5Ac4H/lf5fMpTD0raKA6DzeUN1Zn7PdUc+CGMvTnsFqKp7goZsUzSVUUK
oJHQSgijnz4FzN2Xwq2Iatqq1yuqtIaELYnGZ0hi6z/iKg8Z/y+w96BV/hdjpNCn6mqGFRV8wgkd
+38s3puy/Jl3pMCHSX/ZTuW8RxG+BjCi1hYJauxwhgjuQRR7GLiWcB8MznLXfatlTMPE0Pat20NP
45DLeZVpFv4CGfpMx+tEpH/hCuGVhBSAZKDJJz7NzTiY2VkljpwTJGeLyW8bYpyCWvvLVH2AEe1f
RYpPKCNX/3DJ0cyIO1ZAQmt2BBisFwyTH64neyQlW60mJt1JCplV6Cahn01dQ4yFKegyxpR+4LbK
H7gWuPoRBJickx5MqWP8WSay/GFwX0svD36hkHawu/AUOxeKgMux4I3RDnLtuutIAEHZvr9twslo
QA6UwTSYAPLLHQn2Oua9RUCHJNVzRrncDaDsUu1jGvlyiI/ffUO0B8pnKCIbDZNPSH9Fwb2b9M9l
zldK38cgrZq6B9AThzdVrRHHnR6eY7j4kMQWu9HHTEXtQbBQcxtIMWkM+eJsPi2VQ04eA0DjY6Pg
Ei5J32FVrQ725YcvBBXmdTvZpexySEmfGX76VIe348sXDFU4KRYU5gYyKTt37iXac5oO2l1Yrytj
wU+iI/PYKo0WIpU2s+CXCJ7BLz+ezLN1KvHhyTEOw1jFwJXc9R5XS3AWlq/tO4WZO0dPJ1RhNZuw
sxXeyRz3h1SzQWzKg3hIXXSo14KqrWbOBeegjMdrW5KL2vWJDpCtoqnImeZYe1LnS7Hf61Uous/W
Wc+8RcpssBHar4a4J8TpqnKUC0xabmS5bGkg0kt2rX7Tk+TLtbwqps7/pb+aBgzJVj/hCfqNNDyA
WzE1+iWqxf7o9B+eHRaLh/doU5dNPahTHjYPl3uz6uU3wqevssUT4hDFAmpYqReDwt6BfNzo0ASJ
klGrZr9NlQo+ETj08ErCANGvvCeZrrh6O6EKHgstgdaE81ix0mRIbccUgpLkd2iMncV4mJFjWNxh
pU8eu1jf5NhMjKTTA6zxHnIGpWfG6a+VI+4oaH95/qoq8Sf2lumasjGzZKsf8Vz/19rTN7j9JV5Z
ZsFUJaQNrhtpVylIJPVL3a3/960mKYuS1D3hXLRIExTuoV5BvaIqp8hRZk6fNtRCmtxcE5Edmjcl
kJ2m/shazA2QIgELA1cvRh2NqYj5npvghPiedxbXkNNwf1F7cuIL+J9IIhusmveaE9sSG0h2/BnN
ESibActPBEUJ1nl4PYpyyHsiULoCXgYiQxkj3vSrclz+IqmQsKTV0LzPZKwOIDZp5X9ZidsWHknN
orlpw18yLNDXfXRWoAofPzoVaDIDci2yeVeRGoFizNTmmDqYKVLDhWua7vwUnC4+3WCcgq9ZLjqi
ulZJeXxKSFcysUpz4zRvLBb/xIUSi5WdEiZlt25eu7lvmBHR8fBRUP68sGuqqmZDkP5PNxArR7oY
mgrvh//CqZoxQPF1EueVK456sDESLMepCHTEsaLUdo/lGiIDLlL6mhAs/Q92KCKLgkA/CiOBvwBB
NN9ziLs0PzBH+mn3IyIPyoC+MfKUKR1dG80/D+ryLJn0MANCsOjB++aK1C+raP7mSb13q41BzHnd
lay/zctpsmwdTYrqQ+gYyBkd7KqNotAVVFDY0Yzfttr1irHXP/iAGhIPsnF9Q1lSwg9DBHdwVZDp
dQRuP91N6JbDGYYoNtd8j8YdC0tKfxHkOYCPG2toOTVVi6vbzpw+0UwkWM4GdCZhW0RPyFsp0dDe
zAP3uGH70ucp0RdJ9/EP324xcw60A7s37VIlgkRPMc3d/wB1bpHKwqJ/L8jEb084uTjvNb/o6jEU
7DwRLrom35AtA03+E4t2zTovD42ZBuiyZknfPC8TarWCV09DIJj5in/l+AKbkhRWj/B17WjC15U2
kd07FrxuXIlax13LTQEUVt52L7dAapznM8Inv7gpm1jf0I52lzWaqoVQC+sfFfivtTzgllz+CaVF
bxxuOJd5gZ9yQWqi91k4ux/KDjbWC8Q2l/I1mQzkTSJ/KrvrhorV5kil2dCWf2UBBWCt7XOPq3ZJ
Mr7FJIfvoi1QqyrkhseO9+UAwMpDGZbCN+MPmflImXULZuNSnIkOWExY4LdCZHZZ+YRc3ERjslEy
/Ba8yaGdCul69SM0FnzLXhoUKsNDzx3clTNfm48AfjAzJXT1bbeXl3P8Pi5vRaZ2fWxZbKKeMJhU
kkU7/wNud8b2La97PD1XCTtRfKrUeVjcekxDRpEg2foxTqraKe4FbHlgxgNIzrswxnGRDxF9UB3g
hvBMH1JAKGEvv6eHlBlI0bV15KrWG3RyLUPkgvga/6WbBKD3XAQhZTEbUJP81b7cnnhzjWBWLyxH
fZswSRQuyMpDDtkLl5rNZOZZ1T8qWmzLZ0cZpo6mqD14FO4jDcSOZ1K86sQhmx7OfWgbH7fSGwy9
R6o75r7F+I6jIbfkvT9eqG1T75/Y5nLSCtuad9iknlck8KXZ0QKI7UkGTXGyCvW8MITih24px5n3
vfupjDpIF7nGybGb6PLdfWtlWc58oJFn6/O6DgbVnwO16hJh77oMZdtC9OWlQh8dRGfKqDH7rtjN
A5QnTZwingtQGNX9ZpSxH8RtYPH7uxE7UUsRJdnMUjI5BkK/bxrsfd0hND0sczQ3mmuTpdBFBDXD
6m8gSe/Aj1NDgCZmB1BW2a/czzeQXjl7+fdq/iobkf1Y48HPzrWygKABIir0GL2kqElJUuvh2NEz
eyUif7AMzaOkyOVrzGddKgfmIvHGbXdH7lBsEt24DZd7XBmGDug9dzianV7JlPmDRazr+Y6o1+5N
lJFlOm05QYZpebw2gcHCbXNlw7YxBlPQbeycS4sIRKG5rd4X7cSmaYgRpIJu3uie8K0RtAwz96b/
Se8PISkQw5K6/gnHvfBmCid89s0bzh7+MprHgSOlJrg+penhTSJxBq6pixw5Dk3oIX/SH3Gwuc12
T+odFDaoSL+EpKnQ6A+zHiudM2M+bzJ7SKZTUCTn6UAggzIY7lULKj4LdVCZzb638FljJExyDLsP
NXWV9cSZ2L89T1dd8F9ohykJGpH8OVaVZrws2A+P+Ml6Gt3hDBBbcW9mgzpuFoAeOfSuKQcrQTwY
0pHm5Y3ojLRnvcvQYdSbuAKwQXTtUiETW/nfgc4rz8ZTnNuxW+066AWJ047v+Xswmy5UHFK0aFWk
DCzenXQRgiEmSB3TMa3l+sAvIdh9klMiBPJEVSQ3NohXSCpt5TNjDqaP6bixqSrMVPgHol0GUHmE
auiGzTnxK8uqz717ggVYYZacSqblqpY3KKHzt48gOpitv6Fudtec9aCUt3SmnHyf1MteGzXQFFIN
Yt5bdV0Gc5lsBU2ucn5szlmV47fNiQGgrO4KVxNCGVyLSAqQmYOtvJBDspa7ZytYLGTiXjcuGkHe
nFhs1tmoA4TksjnCeiL4bjerTI8gcWX+8zUT6svf1I0zyeEUbGZ6G61L1739hSTp2Nvw2TlLHp7M
J30tvrafI4eF/Tnyw42aZuUQtGLAFB56HMeF4IXdfh8TxU8cNvZ7RasVF9Mw1sfkviyc2McJS3AC
YBbg+LoQE6+hvQ+FOhA6qA++f22kCYW9qjrS8p9EP/j+NtVkuEgyMXnOZfYzptJCr0D5gwEfGGkj
DcZUV2dZDAkgCFyf0a636V2RwhySY+riNtjpJ83yjUkwHWGXUdm3hPH4q90EsTPndjMaOnptdmwK
uA5VgGEp6L4J6FMmJHFbp3JYGDdo4Kgdmij8J8FcXFL3N7sYa5osiI854r9tsJC0/ik3cO7bSeBt
o23H4DY9fB3sxgj91NO3/heAW2qX0IDJO6U2kJvVnlv1aPqg1aBiduF/OlS+9Sajsv1gdMfLps1Z
CX/IQizazL7k+NLAw7ySf7Dzj9w3t2w0+PdcxMS2ln7LmT1B43b7YwPUeh2hCskn1aUiEatCHGyB
0FnrdWTdlOMcbWjkinD3BS5e3f0FcAxrusifLfV8DGcWnPV7flBO28ZI8xH6GjNE5YkExFjesN77
ms6nDtz2HCV28iC3NoHt+cPqpBbZ1iUgeJ+mS7Qx2LTBqRfDx2qplVcKnYf4ONvGCRo42Mcg9RQD
BwJaAV1HKCca0r4x6sryuwyba15eJ3gR2xPrWLH9+5JLCyMs1l4sAfeRuLGL4Y0gNbXT80056NRJ
3GsbdwJAc8/boKBaS3zHRPwPQRnN07XonFx6lVf+m0xgIRh7w0JggLfVntq33ae36dtRV0j2Bzni
UfEUH88nVTQu9ZyL76CR2BcgrVrhxx4y6nk41OOmUqrnzbkzkwkY10gIP21Hr/wRoStyrqltEV7j
vy1FTRtRf+CcExynry2/DaOO8G0IQX87cdm4IyXtFe/+SL+PamfMx8YN8bzRTnmZ8leq4tAAWfhd
P9yVZaBq0z0tdKyT5sJV/mICLerRti+ytYWtKEU41DrQbUP0u7UhcxoOkyMnA3MjDXzqwU6u7r0F
c6xP+pZmHJaGGzgeMOTWkkbYhZTOx45sh+ROqjA0ig9yEimwD4qyhKKRvq4BrK8zuoS/XpvGQBac
Jd8sMz8qAPB/G/AhGY5R82SdAlnlC8huJuVchOEbG8NhJIKvkqLn+1ljrtukZXp+ZxJpQtIuxHzp
We/FWjHp1e373VJ9Q4NP9ZvNvujv2R1mBmk7kh4DJATUDW0x1SPuoywF4OS7yHG4+mZTN3zKTwz4
HGe46gCSLE36eOgTY/bW8RAOS8FLbV+ojm6P8WmufHv6CA63EglEAOb6wXvdJkvnYR8sd0V28eRw
B5vwpoFGeKTfp+c2ygMlw9fktihbonkQ0D2lsr7CUGnJVOD1a534HpY/Gs6vLQE5WHeeK+lA2hwz
w8TKr/lQ0+rXg7s7on6e20gq3qqnnBnOM2OYEd1U3BqjZ5n0QSP5u+zsB5QN/4EwhP9ixPJQ4hmg
0SW4JE6jVoZfO/DpIt78kELOfSdlZY8JA2qZyFWKIUTW6XY5DP6n9dJ27H4aud5o9tWbo1/q5wsV
eAPUp/b2Qx+pkLv54dKBzLM63qllSYY1j9RazIpBJp1/Xn5fbzlkc65fMFFgRwGg9u7lh+x3dTcU
4mOyhOtxxu0/ankaIFqqOC8ZpRNr2NiHYgrGujeh/0Fe6I3vzrGQyJMNKXVeXx51QT+oqyReUrUE
dDmryYenh71zSNWiMmdu6u5LQKuXpPooBOR5j0Aj3Q9q3O1sDsyW7oqjcghkoWTVB6Ssoo7a73SA
RGIexPb8HdLCi1u4V2qtzsbQTp/b5238/67B0dmcIifiicclioK25mBsKCjA+oUlbavZOVkw458g
KDboGlYh9cbJwojRjc3WySNPjUpg13rw8IupJ+0t/AybFbzoC0/XZRS96aglQKbTMnC3lzoTQwDx
wKD57El/irLXEIpIy5sTI5QqvihphBq7PNvFcRu5IyuTvPSY6DHndqNdeko1S0Y/G/D/y+Kx09YQ
FNGhOYPxOFCOzFRD76RF7Pel0Gd3bGjkiRcOhWmkyTQenxIb/yRdx+OpnHDkc2YxEkcVeMJik02m
zYrAc2nENRoTBeSL1oAsZg49NjzF0ClyxZUCOuElrcAuHJ0kk1VIVouLqxYNlJaF71T1yd8BnCJm
OgW/4Ytsc/j1dP9GwU4o53WGxqg5M7HEh9gQ1WT4+yVuvvccGUobb+Du/krZwC7zWph4mEsBO5qH
VaoJSnTlMEevDIVS435YBnTh3Km3SKdmY35VAzDkCQGrTFOP+fXJofc7b+v9dtjnwuxxpuRmKTbA
jb5J2EERCteSjk4NR7erdNGxLyhKFrNwtWEqYvoVV036B4HMuw6N9g6zDwK05zKA8JLjN7vq7U17
4Bxm7H7o6/ZsWV7k+XNJG2A8JRbqrKEra4FO955ci6oa2zwgnPZy4ysH90VtxvQcrb5h0pbjaOzh
r79UD++0fBeeIFXN1SyvAtvERFT6nDLqxzXdT3laaL19F+U3Ryauwz6FK+mqsMNF2RWu5MMgR9+L
4N3pAfGtsXs7Wjo8ACX5EJBg/Rtj2J/xWRPOMLoW5Wt6srqRkdWCN9FmJ0EnvXfgj9KaLRw/e4nr
51K0ZyoHblUFBHF9ATm1aby0KAqr4WNWzzsLCB1ssxx4FqKi11a2fvsRARZdC3qHkFhSlwcSvIhS
Ip1ItmKzsShRISG3BMSk9HYt1UH8CN5nOJlI9Fz+KaLKay7CocWAJ3kEuV5pEMB+ftZqpcEQtXgT
4FUtVr0mcn1m7XbLlgbYGPPo7cNfy0YRL5hMzAAQk2mBOTEJZVUcdBpgpcXFzRdt/TzZEqLZM/Tv
Jo1RoAbPiH8vPoDhk+4QZaX4STU/YC9P/swGVOKY/kXqcT1obWztNqz6oBIjFwblJJ0kmVmcaQc6
cgwM4yFIPpO26/NhkmdLGo15QkbQxnyw1Bcd88ppp09GsJ05jbY81vm+7lvN6x53kcFznw7axzMS
ZKDob5syhA0g2Oo8+Jmn7pDs/MtaY8PriDwMuILu7mGvNZ9n+dGTyoyluEKs26fZGiQV1Uul3U/5
k/xGKwHR9CBT35fqREzJycVV2n57A/OI5y898VERn7+Y36oi0uXKfAGOAuwhyMyqOsx0nZMImccA
sSUDpDTDjiyQxveXWoq9W0lQf051xMc/15dTolzUvGBNd1zspYd88pnZcLcKY305tFiaTg2WmhGu
eOZTueLndIGTWxZ6qgwQsgohQW9+R0U+l8wTgNTOB/AsTJzh4b/wQXkTmb0HIvy7dzbfOefYoUwy
zUDMtAEA0vywGa0LcnX4q4wByWRceekFWjnRHEgHGS/DOL6O1Xa3zESsfmUb2bCM+wu6WpJNyPTy
thgrMUdLuib2jT+Qjk0O70w+M3u10ewsm4E0lQ9fn1ZZIwo9PpodXGvTCZfL/R9fT0AcoRR3vfzv
ci+zd9Z6Epkqsawlbrrp94jzQM90PeRbK13PK8c9W2wjzON8CewltJ2Bo92owJRX+0NGfDydmF6J
1kYqXLEzWvV/3xUW7/E6f9fS+kNXGDX26MaH+7XzOgj9U8/nY0DuUfWQi12c6+2IZMOJcIgwKCaa
blFutZEUik/MaN/j0sGbHAW7sL+b2xumMm2ccKwx2++oclcQ22BPE7hfb+FgXpNCgbA1cpKPmB3m
ywpaTvaT0nJxzo86MF0BBGQUWxMt5tzsqj47vnklkx4UBrEXt/EFmqt7fbAx+zOJf9Sm1WAu3JJ7
UU1Hw7RA6OD1bJLM+BB1ax7dUw+gBakIOtVorPqF1dAAYKKB/xaHchtry0Ot35vGoMbU5BLuX3Tn
s8wjnx1Pq0KJV/rErTrPYv2B0ZxG8hf7xLOQ+l2xCsZkcUXryRaOJVIKeSdxTy0lvOZ5/laeiO1g
+sIo+Ah7hHZ9VU0gV0HbaRZ2TvNnQ2AQAft+mdgRGRDUTpfkGqoszE33fV0EdA627wOcavPNr4rd
PYUCFIa5/Rg6wskh7K/HQwUnIgZkeylgz+uY3uW3DrmD6QpnvMrMNFuB3SwRRRoyQsZ7fSiwzUXo
LOMV7pgrvyup9EmDw7cSL89xX5im0Nvkdipdpo9YWIYswhPOSeG4TGyWYbP89Qb1gmX8kUrzBehs
Z/rSe61w6eQXG4uOvisUXcROyhDjKZZFz439yP0+cPUK0rquXlEKDlIc78rXOn9GYP4P524yirge
TSG7K4hUzhFKuvlGd4bYuoNkaxOgTsBF1qerKVplJYIOfqU2DKf2Ez681ttDlzoXxI8T7nSIuS1i
nlxBfEStdKmF1hX7vyoWFOOS18eV7D+pu4cKUEtLx9mTKTGbKZZa6Mkh1NPKAbg/e7vv2kTPemN+
6eyoBJ8E4ank6DzO2C4xLtkFmcdUVIhJSOlZLGW3TvdtriiZ5jcQxRdUzQYYZDwE9TW63sXAxHCM
T/3AOtXL46b+fymPqHfEGPm1YrGOG066areWS27yzJCdO+zKclUZnNEXRnJrmfhj+QRtjpspxTR/
0i4VygfKPj6NzKwT+xkS2yRb9ulVdJPVo9NoAZ1k5YdT4a34Z+WGDPMISDQC9QRwih71qdLLzOK+
mBIgaYQfHFt2WoufwKkluU6v2ohcsnzU8h4LAUiwEKw0Htyzu5A3QDIKfUPsMjGpabi0Sq0ayUWi
M5Jxz+xYpIMM/cUIZ3oBCaARdHAeuBt9nGNuYtM04jb4sOLqkajnLqeUuFKYkFBP5FmkOEMqcvrR
hBJKfhvT0IdwGJaU+PvhJSOEqB8Xa8WyBQMlXhdhumxzY+HkXG5MrS3g1T3zlgwQRBItIot9/oRh
k6X5mrwfY91CMamK7UPqqcN07bvNTg6o5KgXLgMX2t736XWt7M9DqhlRXPoC3zZP5Dgt1qAROPpv
XryE0FCykmKu8qDztlnkEJW0/OGl2Wdvl4OdHdNLlWunLnqIACwILEOHdgv2gDxmtH+R8wEIOzTe
SAwfJeMPhBMiLIIhb+BcWskD9XrGje2OmOXl1pt5uFGTdFO0RQW63Lr5PuNK0VTO5cR7ZlnvdADH
TKBpCWdQYxv1+EG/yWB/kGPndLOHeg+KUFWjA1P7+esrHwt5ux6s+LOtM+4wCcJwB2netrsOzQ+1
PY/DcdRHCgBVw7DmNtnAz8iSo/j7pjxU1XHrgM6FCY3fINQGCM4fXX+SOLsLHZIe5JftVvH0wxTp
jt+eq+vIOYPpfatTxf1c6bgv8ziZVkwQ5Q/XbXlqjPzdM9pX3UFGRCl6jWsTM+iAONQeTtMBfMvL
XOnTiJuU/6YlIFz6HHreUvv/MHId7gR8/PJ7XwBdYQE4MFl1ao3NEWq1FPypmaIbOetEPzaJXolw
CIgaufDWx+R879cTixtM2Y376/VHs9p4sOvFzVJKC6F8/nMhjLRUDsMqG9zVmGlXiK+WiRPWnJ5c
Zk3FAbwPpzAxapfO2fe6A/fNnmrwhLJ1o7QoyfrNkmlg0g3r5SYGdeCZz5J85+FdxAWGzoFuOSkn
mc6P3XS1ec63KF5dUfHbOgEe/0XlxL9/FM87SXcEIcC0CSGsOrQiKbKm8pKUOJIM69F/wcjskl26
WwKFViilOxv/G2zenwGr4LuZsZogSHdDV+kuISgykSIALLj9yFxjaQImwZDuJac8sUeOZbpENLFt
Mjl8tm+LaLdcHLEPglDe9XkoSQZk881kP66kZSWZn9YhQ+NOXsFB2KPS1xEEy1dTWwWfYIE5OLR5
kbAW+Ba42LFbJwYAS6LKh3uEe/DL25I7SKLStanGYHb5f/hY+5ZlGwn+Q0xztGBQnCU64mgLv28E
/IuPs5khLdCeTY95wVsGAVL7/7znM4hrU3RSaweQsNvb5vsC/85Edce1abj9WXi3P0E19aYh2MFI
6Z3CoRhkEHWU3uuc7WCzA/Iko/M6KGdXpfaT4erpLw6pfNsyXfDsUHRQ/i3ZXfJ6Mmn69MYKZMCU
yvs23Dnzm3x/BpIgy5Wt7zUACO38P0WQUG9CkcKpigiib+BHd2Yuf6bhyo/DRK6J2HNzwHPcTW9I
3Ir7A6GHAuSVdgy41lUP79cO1tMu1kiojljBtzD+VKsfaiA7e83SBA0uoA+GEFaNJVLBbhDmsS5Z
TgufSUB3LrLptQ08NYkav7+0Rp5Aiki0jVsjY4IwX/OqjnYEh/0z/eQ9Scs6TKKrCDDhDmCkelCA
gh7H0N6NGUGVFu0CAwZRuq2KrSMjjW6Eyo3Ra7vGXNbiJTe9NQ7eABCiVNTi9NsddjnI9o9/UqGC
A4T5RVSInrhm0uYpL2YJcEkKJKRMQhcIcH6lQCNlu11ItDme8oFfdERddF5WYVY8cZHdB71j6v9A
ZdQiP9e5sk0Bh3YvdVaOMAx4131rBuM5BKt4WR7JJTFCscKNNQRzsHfVg5Y6Z0910Qnihmdq8FLu
pWIjArjNyvrHTm0nUNe5UDAG48ros1QolMxUuneD1WCY1sPcZbSglPw+pmrblM/kVGTJQU9Nv5CX
2W91Xqc84vrr0D2hrtkzH+rVagaMjOEkv6dQ+7TZDG6v/WCQh0ShAf01G0G82I2Cz2dV3k2TRuHA
4FZywNe006qlX0CUJAZqq9Is81PwGRnoGP39dWv6yamPgobvlgZRynGfOih8hkfJb/IrtfN02i0K
HL8BwhVraPu7gr9Jp7X47bHmOzPa/I3wZdaXsWh/FmNzxsyfjvg0hZbnAoMWvNoReeAhk2ii/rbf
QBZFnUdq5GqfVPT5ah1S1RTfTw0EoUGp0NXf+D2opdGlQZuRX4cn39yE2d+QV2KSuvF13eBGJV8y
fDiOYenFkP7U9+6bT8bWw/09mAcdQBJaBEZ0idKx2sJFcPv7blcqrUeZu79t8bR/5Qyk0BcKAuwy
YhZfEcE8jLZXavf2BY9i6fSJQ+zGx0Ib6v5gGbsbM5MxWs0yxURH4OHntUUjQanMgMqac3GpEMjy
bUEJdesVUWoTnoIJI7Jh30DTcAB8+PXNovOWXwljVrXl4R8pO66iMaNwZs/9D6jX9NfxRMOz3jXr
kL0Cc/w7og3FH59/aVx0dAuNGaKnJ8GYxTzwYZa0C0/X9Wm3CTU9XChXWyzJ25tb9EupygN/+PHj
hoSmG2DScZpkPdi+jWeE7UI92h9xTQTSCkxUSI0yzU9+awiViG1pAk6Yocgk+jv0wrntAAS79xjX
YfXSk/7/Q8wW6xdpLFo2W4WnJy4DGPj6vkQHBDZ2uS+MSCZlyDnmSA9fuZSG1sI3CR3FlC8mqSaQ
hCpoz9rP7llQhQQTFcTqojLtRvyYTBDRN7DoBkt75UMuZZ4Q7wnSleo4XM60/Tq7t13b+ckqYwiV
apUbfOryliNXbo1UfMYs+V9ie9LwUE/Gl8s8nt0XZg3mEECdFMTutdMVZkKZWSAJPRefI0S53U1Y
tCsworvkm3AiDOKPOYPvPaKiLufPJUDjtooujh/6eTVgjZUxwb8HBo+m8T8ryUzbQ9chjKcC4dnG
7c70EMFH9z/+Tp94L1/VjLOzJYIDsVsxEb8WPd/yu1HT3gyzOWh+jHjrJhf/RXOAJu/d/ClhZ7vk
JMGXSuw25e6S0CPzgW6EW8/YEfbeyC2NVoOKdvDkmC+CtUtPWcvx78e76/yuOarSpqlfdxLFwjrS
2r+QXtPKThIgg7Wvs57Sc7LJeHbE9UCHXf0DIbMnW4s416zxGJVeN6Ips8/Z69jMUgCGM98fsyZQ
zQYjV0sbseaozNadlWW5dX01J59bkjFX5PBXmQwtiGt0kq8caQVwToVAIoiZS9Ph8dRGKO8Sc7qi
sS47BOUWg/xyeQ01ToH4ubP2FuHPsDXrPdIxiWq/mag7jpp37SSeMyFEC9yz0Xznaox9DHb8Ctok
Vd6HHJ6eEVVp+s2ddL0TDkljmUEQhZ20FSPZzlOhpy6NrHLDywCeO/pGhXFOByHaCjGXNSzKP+4K
DIPWIagIXrJPdEstRMD5zDCd5F6MI/N4AHujM+04SKOHBCj/PrkXItg3m/zJvsJrF9x3l2MC25rL
ikKb59wT+D4htm73RF1Liae8IBCVDbGtY7LvlgGvVuwYbU86cQ6ucuhRHdC4Zv7bLb2IddhRIzor
GLp/edS3OKm9p+DOj3rk5jtp+5ZHxOwBD1i9jrwp2/oVUHMm8J+3xBMZKFlEEaslJThJ8vfhbesL
BtZvH92WGHQDE+CwE+60SGxTitmPB7ioMw/lQHG/7zJpop2gIrtf8gKcVAZD9Czongc11EqFIU2I
ncxxKyElZwb/JftjGR6kIm8c5t2jqWJWgHPIcBlPOeVi7lfQgnuw8Kn4E05EqAIKHVioBfabOr0z
CN7STSGyPTUwxYHmLN3Q9R43H62pmnZX8xj0gw1TDwASjQ1gMHKF0AYXMKcw2jpZuWI6Ncbc6iI2
aj+p4MayGTLtp5gLRJc0LUMNXSqe7fvEQvguQ72cg3bZn67GvexIPvZXsv4HEJ9pLOXLuDikwEif
Hpv+XIGWgKlMHKel4W+Zng/Kv7B2ym2n5w1P0L/PUHS6gLz1YbgvsGoGmD07IYR7MxnstR+YPwSN
574uhTRJjT2vUm+qTOHaVL2GCBr4/6rteNJHzdelHTN9IahqC6YWa89hUEnNd70svSSC9IaxFg2a
SGOO/8aPEmSbckSXnNpd9x+K+SBdAV5N1ZzYuWzT4Oic5Gwx/tEjvS21Oo2VbCGURcXlDuMKyvYv
akng1j0l05fd8AGvRuLeYPbKADvBpdrEB+vDlLm6+Xz28p1U+xDDyVAUIM6cEME7fPZyZf6wtggc
rjRqHUidYtzuO9z8QUX/+0O+do5ORm5GR5DO1kA6C8DOosgnp8QiUvyng4ecPpLnwoaluVS5qkxD
rr3nNdYlM/4TZIHflz1XEWVvLgihG2mR6eI9LI9Sfoj4NPnB+uk7tk7d3yfkSQBsSvZATJ8x8ecf
J92mDaW0liCjstwAVvrFBPH3ttUJOlHiSxIpk11x5JtGWRGUC6iGdDHjd2A6fOq4DiKD3VGKD6uG
F8K7Od92eGIIwnaPSnBJtcA1rxi0jgwGX87xBOZT4XqFRsDqDBlC8HvSfIXVCCVY84fmBmMThUov
tTNmNoYJHV499Z2jus1Pvien2TH1giLKYU/a9nRIDEZ2qdVFq1DkvaNsu6n1+JsRv0arDv5vDQem
dLVf2JcnWXMNLVRzva0UYIqhCD74LglRur4TD6EUgn3GiYKGKNSeJYODO5JALCeMz/UxWvuNp2vy
NSAu4aYPSxRHcszHMzUdUV27IPI+qNYgDXOxb8FjvzxtUWbwzQiwzqK+A1El2UZ8EuJPgoed0MMf
JnVsESf0sPVPucucckRMOecGeNeaj4BnIYHkBnK5iraVu3sOdBG9ZVdRniruGgWqmcXaUrBxr9i7
yQ9EwecGWIlJRfbIlT5bI5pajBuKOp4wV8st9ZxLWN3WSYTRCjlTF/dLbwn45aVoSZD0vnmXMRW3
fBIWs5ymEXUkYtkI60/UCEXcjcWicdosdskgyyPt4N6AopzNrwSSvMEGqcg+LP/eqqJJNBd5bMD/
A7N+EGfeRMd53lAtowOyrs6CGH+qFg2U10xjt2SkxSg4g63c4ltup6yK+0vhAmIMNOq2da7WTEnH
BkEigZxHMZQgSXIeiF2Q9n5dqH5/vI7o4ScLzYUST307hqvH2LT4YfPjwZlcvA1G3ji3R9Gu0sh5
VsDtcRGiqQZt5AWsxq/1kqOilzFnnnQbFhqSmETvyNq/SvWXiInA9QjClpfs0MV0uxp200lTvsLZ
YyqDZgnraGQc3iKxCIiXnGvZYd/r4kMPqRWx7xDPAdh2544OqdOVrKK5K+iCY716FWk5iODGwzL8
Busfx88wbvQq3YBp9tICMGjB+KQFJ8THDejAvpy8V95wQKPVrf7E8bk0UrlYbD6k4YYwEHjAVolz
LSbPHez3LTBPSWXeIoeBvb+yKtxgV9H9KiofS5gzy3j1QfGcrMvh80bhxCsRq9hg+U0rmX32eIxE
YBcGleLAeN1TEnc+3Lqeiqe3fGT6/1NKyw+gb/ljHviUgrR6YgzdvaNFQl2zGuLB67TrD3xjERQh
3R8RCk4O9fN3mJrdBAw/qX9LrY9rJc2CirfJdRjjMxYTaNWkF+sLvjAD65m7OgnPEu9XbIfK/4Pk
rf7NWsp10ZP3WAOEPGeH/+RzhUqtxTFCrVpSlw38EjuiszI5woTr97/ZeOtTUeQI0dHO3gr/nxa/
u0jlez9yg9yybqb/yRLQZeMIHVKofkoma/1ape2tfwp6P8lyGnXXlu/+nsR6X30MysToKptvRqPI
Fea2r7u7ba2+RmclkJliqUAa38b+ZLq2aycMtuXq1+/JnxqO2mPGrQRvIPbty+HIDkSkmEcYIGXo
eKKaGzOE8BToeVo3Z8TuAumbBJqayG/X4BryHKntu4AlRV6n4vs7V8YtElv/vyPvniFjzfdN44bX
VkWeksIiHY+om2tUmUOxNnoTc39NyT4oKjM7qiGny8Ibzqnfc987iZo4L//3x0qNeAM07hwOY0s0
hUdJHWgI/cSDDhhrK2ftswTy14wk3cw1H+5W85qfRsO4ozRpXDmbtUtb+F3wYvIGf7NKG4MtTd7J
hn1MuVtQrKWcT9MC++iNrRNlXtIoPOfVUtHctMUmRtUXPGkalr/UCGhio/+JOlLKfapJ82ZNojPc
jDED0nV3UqqYDKkeEEU43gS/683fSUHlWWb9AhOfWD0ahJAemPXnaGIhKyHE3Z7vVPLdIuO/UO2T
0nrg1EOUE+G1dAkIQQcujwelLVFVsLfZvfXUJDyj27Xxj7SIta70/eOO6/B3snQthvkgbF8118LK
mVh9Cg+4rlFg9ZkxK/NkRpfN0c2OaPzpAYqzUplOlyKsraun18z+TALDP5gZSIEb1jyVfyP5Ih1r
POSO76X5W2oBN3ef5E7EIYk6LMCMbwvasLnCHYxzivHWhJLti2L0MGKBPLOL0+9oVJ8auJqIeglY
iw8Puh1sfua1IU308tdux5oR3VE7H5OophVUxPbdFJCfWEH+H1Q5l2b5DtDQV1N8vQ9uluznN83P
SVXAo1A80z3Br7CObKfnx6grcJzneDJJQV2X8aKlIfdtuoebpAMEeASrHQYtYN4IGbY1RiaosRJb
p6QdAvy7qIiGp2ObDqI3ZNSezJcVQMgsdGbK1mnaO3TA0koCBZrW6lX9rUrQ5uOxcfbc4ohPnX9J
ChxRu8QuhyIfp6H+3HbUW3QgnG1bHi/3aqLOYxGq5nD3bZBL/jXOCzfMHBFGoisPrL95YjQi44Bh
FffrKi6y26dK4/SqM1bvseuesNXAYCmGvr6lTCnS5xE+MNL07nk4nZmmJqJO8VSsPi+T2YpyrRWi
iHXr2TC8O99Yqg6yo1jnaR/yz5sptptn4qGpiZyBxReb+ulbM5RjoNmreRJQNQu7LcjE+qpHHcYV
WZlMgVmm4hXYxfW7k6nX2DDTOi6SQSZvhB3i99CBclxSVGFHNj2IkXOZb45S/ngusxHOtDp9psZ+
b/ou/VBprsCEXz1uUQe6C75dtKRVflwuaEf8QpBIEDl3lCy9MZyJpf1Znx2zeAjQo3tXRmyKRIop
5T3iCEQASw9K31Qc/Mc9MzWqyEBf7eyEWr70lVewpWXnqu4Ykdqk1+fuuQ/P4t/uNJsVJhkGFXkA
3lMPIUVJjNS/nFAHpJEuwvGnGj0WySu9FRbtR7oPKGO078DhrZXmUXW9g0xAy23NvZKnTx32FmKH
uEenx/pMdYjIYs7izlLdUVGpmNgNo9si9LwXDD6v7jgeD4tYYTQy2nJN2lH1NHw/WK3DaM5p2tgy
y5cUTIV9COr9iLBMWLMBkt9/UinQ6aIA01xB8AueS59RClmnQETiqJ/9YxQ5DmQR+Oc9U4yoQTS1
bv30aXmxLqRv20S8L8lA74qiWUTxSF8VnvtPowXrEMjh1a3Wm92Pwe4mrzSchunez4Z+iDnpLyoQ
7nXgvbU0CnH55LLIWMa3oPVcZLxzEbqMYpJYAETuefAionW9oRV43PsxHm8yBvG8+tqIJf2kEfAw
5E66JIa9sc1hl2ZREiU3y++yGgBnYsXymAqSKRkJ/8+fZbSmwEcrXJTmdV4pj/t/CrquVXYSVOBf
kbAadf/tDdKDoS9NM7IgQeYk0/Z57RKYWZIjS9PfxjlvZgC6FWTsWd+luqqEvQOuEZzu+hYCCL0V
+evwL+qt1VsN+bzqfSctqQPIwroULK6vQjs7LheZmjah5JjyLlH9VekizUSGI7L42gGsTsIGO0qk
6HRwGDus/QnI1Y2sIxxi04fvhZvSLSZozMyjX4ahtaRvt5RcWYnFydlT4iIcb5oWoGJcjQfmKI46
FQAL4ULIDr4SjroljnPKoUJHISuh7+DKAZaZGdIjpaV0rgGJr5lQTLJdvLfvjurdE6tD0mfHKM83
FctJajQ/MavmeVsIuDDOSL51FQZCSu6EXBfhZXF1aA2xuF1ZMpc7L6uTbeT3Iqmdccd3fKDzHlXb
V0+yAnCqlUDV3dCPEs8cZCOBtXgE+hWzjd6rXJt11iua9h9UCwW8hWuXGpFKD0Mogdnq4bx//u2Y
lzIjSiR3YF25SUGzaSS06HVNub2uY/mrkQ7ydaDo+/2pUsX7iHsE8PGowauILZQrzKv0U4u991Wr
HShQV60+ift4dUmroP0T84INEpvHiywzRzsrdarT7ZYjsHn7kcx6lvhmiRTDXkKk3mN8vRMgnZ/Z
GiT/rI8Mv2hS1yF/KFjYGsCDrMDagAkeIwwjQ2lYa4EF7V+oTFMpDQz//Om26NWNi0FbyhYSS+Pb
VsP4bHlLfBDIUR20nB4/sqKVxpX++l8ntyPDrFeeHE+qJj/qIdZ8PGAzAJxUJuwWI445DFTT0Q66
TgGOPY8dKAjIbdQk/9mBkLCdMTS3QjFVvhUd3+mzHCfIwUOPEnMCv9nvMwDoRLm1mT5nWTfqm9id
dNt5PY9vY9BwKSSnkD72b5tU1tmyR22st40on4L5c9HYwO+KgMS2vHEvSxWXD5XKjSa+qYla3DBm
u96AOOrI1yWr29q8O8AlidnnN7+usO1AwHvdYeVeBae1iPg/QLy2FlXd+OpCfOBKpVXnO2BAwCQe
OAAq/IcXaIbTF26kkrPuHsRCsdU+zn34brNlcYFXEZbHSwg3OfUSrePHG98ZHkqOP9ZFmCF9eube
cGkYEP9mX7qYnw5+MMFwrmZ4vBcaxyw5ZMJRMlGWi+tqlBBj/i63hsjGfDYIzK9h1A7gaQS969we
PPeeflD67xvSnEeFlzIDaXfPm6yKzaY9YNQU2NP6ksGQEhWCxPglVfXAwaDsQiFmkLpyRzeIAumI
8hk49WVIgodmB4DbfgqQIhvEDtLBvu3HBXXUS9wg0zIbtpCGTQGAK0PeDMkxQhMnwAA9dDWmBcN+
BiO2LYYDd1m4CLoUCWil7zat7SZ6O1pABba5tCNBJeH5f80B7sE8loHymsR28VMwRYaMDtEnaBOW
AXw9tfD8/UbVuGzC2/VSmK8YDIIXnHqumr28opofNLqIm5d7ZxZ/EGcda2un8PyIbc0A/EF4KbLP
Umq+yuDgMXq0mNCsmx8zSeuhGW/oq4ogzwvrF29fnnK1piqxUEWACoTEHkkptUOtQ7eLq1cGlV+D
shBhmPlTpQ6Q5M48tmqHKjkuuKeoXctblry1SwQwSvDS4A9FzWpZn7Om60e0QYiGLoM3uelRquoQ
PG9lE2MTIAM92/YOOIRwdoZnSh3B3nt4kypZC5kGm9c98iW2F4mNZMyr6WSb5dQ/CaCwGSXjt1nZ
BE4dZz5o9vqosqG5q+hpg63uIdpL0LMlAzSaFq2IQwBHDlR+8kgNw7jOzb8my2/g1udyhBHVKSvU
IOK4C+YaKK0FG+Vq8JZt9SYOMw1kHXjyBSrL/o2byFdp6eqgwX4M38WWFpYZK053B1aJCUo1vHbI
D+cl8mXD5GwTULxMKpTStx0DpotGRvbYgTJXC8xz5QTyusSJMZ8n16BUsCaHXUiH7ZNHKChzm5GB
uvE+UdjWYe+hkxjTpkPpofQfpIO1uImNe8bPgOpf4isIYrd+LwsuR71OJ1cmrCF6Jwl1cJq5klkr
KbPyDjgN3szin/qWa1vP+f4ffNhhv97UnVM5L2zoIOUsJdAjAbWdB9VHUgu3zOxn5h3fi6OQbjOA
sq4Y++IhDsYgxa7E10Q1uXZa3/vOCuhuvJ8ZMWurYJVxocQ9ckS4bJdt95Gd48Yha//kSgDw5j9r
cWqm78yz9LecYMNv5FxcWf6eEIpLRu3IjDPYgz003ea/NaQHRB3XQIgkMl5X1F5KF8dM03wCWXGW
+9HR6j2k75u7z+qP1cXrJRd4pLYUVn9PwvgW1MeoGpCJy+5rCY0AlA0C4aBab8r3Nh1COXgSbfHf
gAYXEPMJned38iU2f6cGRZsMn99e/SGfIfAoMYJivmlT6u9Zc2LOWNEjDzAniX3X9gpXMfLVaqzj
6v6zmLO87E0RcO08c16HKbPLZGL2dqN+S5utJOYIHso0mWtwJO1ppiz2zZhz80Bl4yvkThQH8mpT
oy0I9nfwWHWfwVF0irvSM9BTDX3OZ6ZZqRvu4nrpV7YSq52+i0KaxSZ0NaMDtF9WAOdX+zhm/gaA
U6vyY2hOFR87wGcMszrhMvS4vN9MKXCHJD89GEEWyE3Ln4+WHeh/ZxyhjlhM0EKGLHivv515HmPO
eEExw4yBt6DjuTZPGc9G1UFNaxjA8BDUYSHChfQ/OlaYUf4xROnqHiCzao2kNrG/COHEPQhu3Eik
rMbgYK7+aTeRIk+V66TH/fxDrivg0RlTIeWoSSN9ZiMJv5hQHlhmOeJcb6fY1vvdmy4lEppBoSRA
fEq4RuEUU7jiQasRNnk/lXTRxS8cFILnTCmIYcXvLtPTALhGkI62IQ8RfoaX+wkke/3RDYVzDT2H
PC8lK+wAalIL6M2MfNQMtnjuvhhv/IDTQ0hi4OTfzOS7gyBDUglrdlndlr+jJUCIwo55nImTAZAW
FMQRLCqnqFvo1rIdWihq99rOuFdKzf+YJ/Fw4ZX/XspKvA64GnygZqUHqmL0D/gaSWjqO90tR3eW
ypgnD8bYpnwKGXP7CGFMCJ4ZKztNctIGIIPdNHnmgYsnEsZzz63Am9G2utkk8sJdtZIq4SQSmwJW
i3MqXQVOt9ddM5Y1+6xy1j4w3j0MicL+Ka+5HiN9Uvo6o1+iPTbUZsRmdCZD8LB7f0ObhF0wgjyG
e6nQSMCEPOHBLnToSFbAffjdpXe6835aVn5ApFpuA5c4Qv2aYwFxOJtoAjNWoNzvP1TC9RriLObR
IykICZJBZOwjb22P51JWXqZcoGnbRsyGq/DuuX4Rt+swjBnoseAfMId56srfAMbb4Bqx1iOULYqh
NLd0hbtCKbX8gRtyKfPUIvl6bcBIq8dskKe6ltUdTCT/r/DA8PYL+nFG6kK+NkkB+PQk5DdJaqzc
kkK0cn5q8EpozWsDtxC88nXpdEc1Wm2ng5S+hkGOOVOkcrEAgnhSl7h+UNVnT1afc95rT3JuTU1c
C9w4v3trsK2DfSPGZrSF8oh5jjEFmWu47Ce5KiPZG2edpkVlhdhQ3DABDLK/ioRHHgAPDxq4VtSs
h+uzdmC4vdm/Gyy8QpYZb0C0iuY6h8MfHz4eJw74Lr0gxic43ipUe3eygwu4OSAH2osdkr4Vlxns
AwKAQiNQrFfWHH9ok1gLF+ipnViBocDIpmM02RRUUpRI0vP6o5hZvZVK7ijK91kE3pXqDZfV7B95
WtRytlBNPlKFRGVZaV7sLSJyumDCUG/BALKWSz9jgirTgk6x5BFC+Ee8ZWUdk+gZA22c96XPh1Xv
gcRBeqlTrG3iG0XtHes4UQt363h+ukvbhmjKsvpsN19kECylgS+mS4NuZEJsTBstEROOaKk616Uf
EanjCzKCCmxp7YSyK90xd7CfquS2c8FGiinDHc5iFzhPb+LI5pThZNziaZ8VCZkyOPQX5L9m+Oek
2b+Z+WxDE4mvaqxrZ73U/M6FCk9nZuit6Xw9UkTDj0NICHDggqOQJsDe3hKveJqbiMOb3tmsnMt4
GIihrQkkYZJ77vo1PzSx3kCRmkx0mpPWjTPYwBbnC7MVSkEaziJczuij6YLDpRi7Wm4+txi92Iqq
kYTpxgJl7stxXmUDMzjTlz08s54m5gom3pnkrBnvrzc8RNF4zKLiIR8GRpzosLRfvUNyJiDvt8xl
WciueW4vdwq7DCZhX6JYJEwxMCMUA1MOFC9Rh465NMwAKy76hWAwI+UXGR82bmiofUdDsyXs8k2l
mQmKtaaiGLsQ3KGMAurkfWQatLtFY7KNB1XEpg36tTTHCO6zCb+BxtYSRb5hryQScpGiW3rBvhTB
Yo9k4W848/hhzd8JGin7y4v/fUqevNIts9ud/rZ1lFDVSB0MUfhGEC0nDxKw2cWPLbgLIf8l7bHM
j9zlp/AkahNGy2uISs5KOjYY2WjRedyDZnF+dfBY50vJIMIPUMEYYNn7CjdL/e8ILTILnmngKvg/
3klrHjjvRUzYb7wFZy1pNw3vmS5BC9GQuWWkqYJZ4tnCt3Bbi/de76E7bcF76XO3lUm/yds3mXwb
VS309iG4PdRTCx/D0N0d8L78A7o7Zd77/qGfbIu0UjWxnbFZ3DdLhxS7LMXLJYtQcfh16bkelSTt
uOev399c76IUgAE8NhC4ftQYIpNASUGp5noFmqk+g1R5vbpdm1B56lhx9ssBX3WJRxYgL8XVeOXj
65c8vDELhnbXQ5VqD7gplmM4qkKt7FLKyPXUoVqKS4FrCx42MUY3R9ki3OQaSkZ14E+X3WrGx6tE
OdGHl4SOsjy61lJAVT7NSBEYtIFHY6WXOJ/eyrbHRM3I7J03q+4Puxziubcc9ekDQfzHACV6wO/e
S8WeUyEBW2D1h7+flXGth17cY0DUT01LOW6jmaQ2NJBlymekZGQN2HFfNvRtKDkR0rZsyF9zRBDX
C+P2R4RUxA6Z4XSaVSYcdChteFdF+wQY2NSnvAPu+qBa2Ep6/UJdszdiOOno4pcw9y0ehNDWztgW
jZv0S9h7J8V+Ipwuvz+pJOb+p/1YZxJRyi/fSJSmKpwVY+KTzTszB2NgIdiqtaUEBpoodOvVR6S8
7p+Do+98UzqTk2Gzu7akaq441xF3saOASyAi2rHjC0D5QSy3V9sWAUDuSNoTia1p9ApN+TpfXxSM
wkwgu6euKqeHLpIfiOklCcBlyOUxLhvLBFgL/SNvAMXARYKEH0qXpBGGu8yanLeHSvPc9eHJqLl2
S0b9g2ledFktUXSMo2jM3mQyeEdEJhLBW7xpwn6hChjLU81QrpOUobj7YpKnXElMoc8ZqCxl16TE
0J76M7EnLqX89vbYBPeNWKN6kwEUf3qb5fb6bwq2NoPmhCX+aENm5yuek+/44jYQFnSPoPF2Wwy5
9ry2lgMQP567C1LeY/aa6/J/glPRaAeJzmohpDeHCvJZF/2aLuYqHTnPWM3qqXOpZuPR8OZjBtMM
TzuhW54ocXV5WftIKryGKDXyzTk6dKIf1/ipYOfFhVOUXblJu37VUUpJ0F4V8ICNSqFHLf4Bx2mW
kEeG+EkDMJ3mULvH60Agf8DfC0Iv39v3uW2pIFGhvLvUY6hCKMr8yujUR6oWmehRZN6Jr6rjtRmc
uN26Hprl/+Tck+jyQXZK++gTrO6lweilw2j+MslPr2GkNjbZNdIbCgGAQtahoNM2zzeCV94gZl/P
6lT9fZ3ufz2Ljd2efOHCesrH7ULh1EELQg3u8MP/PfxQEyIJC4x8RSS4DUrfW4KUgrb99uyQiIZS
Nz/tv+BX5uj/E6FoqR3DTOdPc29ibWzPCAudcLpdqtZmpqzxjzl2IW42yYue4IlUSwRHO/uFEgWN
q5DKCqhqSqnpzlxIMOBQihK33lBvDml+ZxAffPojxERkvisFK5rLQgrhspxzzpJVLQ5l3TveynrJ
XeUnWIwvRZbde97wUzKmfbKW8qaEFnIealIE/JRH+0WWSXUhexn7goXJMBGE1s9hdP7GKOZHbrSG
WsWIXnX0qEimvcKE8nBIXmXimqloVM9rWkjs6oQrn6VMgnDJKLr8DPX+VpO2JR3AZyPeTLk+OLAZ
9GLYqzQcYio5KZqBbCVlDtfR4I05Yi49O4IWLkVkoOXNBTlLf+qtya6s7WNiipCwm3mv/ECHkMEu
8t6Wut0I1TFIWaNgc3sNljpvsdIVLKPn9FCs7zkzb31yJIUX9J3pjopzKxW9+ojCrvK9my7+NZ0S
xpnZsIGckJedT+YkoKRxkxB4qg9Jzc+m27h6fTHN++EpCIBp1paz+ILVYovL6bbpW6D4PTK2DNRY
4ofxQW3IQIwWHwdVQUo6VR8njkOKATsJRCS97ektxeKAFPSxlHOWSbD3+qspgAD8GPFUT4v6WFYI
yotAhj7/g+rTE6O7MULlRW7P69LZ+vO3JDdSmaSem0DIuWBiRv/c7OBQ1G2vgEhRfYp1oZhZ/4UT
YbUctwmur+5ixjxojZNe6LfPmhvs9Jy/CTcDMiD4ZntmQ+tluDrSiv+FtjZq1LwWN4cqjvQXhOro
/hVWdzmDc8+Rw40rRjNPTrWihH2JSNh6i9Ro7laAMZ6mf5xdkyEkyXpEuHqTrxorxu+ooLAihW/u
UNBDdjBbBRRoIaZJDXnWmgyZi1x6Dww5+J5KcOy9icdfxdCnilKRYMINOsLhgfFdeD0AZcPXc9pw
hajFZa4EfBFWHC/Rj8D8LIc0WJG/WD38h5U5M54W144u1Pv1moD92Vp8Z5uypmgYtrvJM1jnPPCP
hItLqfOb2Qgs2dCv1+VxL0yJ+g/eKeMtN6wu9Q41Tp6vby6FrmV2tvbH7GcSm0/zkyfoLJN906xE
eH/T6RP7hoBPCms7kGn7rgHEFsA5d0pQOJW47H4KBgHhrhuzTUUQs8h+lJhAfDrRez23TFmQ7/NX
A0Juuu6IfJEn+1WD1G25hezKV+wqrTMrlZEVDFuYo2J6daq/dKagWG8DQogZQ+fcuLvukbauRU9X
Yu3BsHY0/0hsS6BYXvrNZlmdylS35LSQFUkxWdnpJH7dM2+pJz8Xe6iZaTmX9HVRCQIH3nuEqVat
4yPDE1+WH+qL/LOKMAr2oQlr/leEv4d9DvDdcIv5556FF2EzVrMnmLiGWlKNEUeHApQ34pxZEYJV
M8c7ilV+u3hY2J+8k2IQp9ghHHIX/8W07VjQdQWIrItatziZgY4j+EHdnvy4jAtj8SWv0tSAADD+
HAFNonDHTVsQmwAxh+E/WzLImKK+Bi04YPOHk4E0X8fveQeoSDCfGzKiNlLxxwnyWUjbKnMSyxJe
GyLotxFQgyblvQn+j9l3qjP0SWq8d3i15NrL3AGhwwXvrpLQSkJ/KWj0u5ZBJVKL1K247pPK+AY/
KA39fftFcjVJ5B7K+UF+NrE+Wamgmbh7Ur255OKIAs6LcgKMXj+ZQsgMEPIJRmYyfZWbgqohfOvS
z3mEDDJfbJ2/biSVPG3YlMaMWijKYnCrZicfph12vTAGTTSicYIWSrQwDOnF/G0ladOWQy4Wwks7
VHCThOZ7xJNbe4rka05skSvmkUIjGTuC/n+HBIqeMT2szF4WKDNuzeK58/9mTnthm4AsjRkaugok
+LzGAz0b5b6oFq3arfjcb3qqLa4L06slYEtcyCmeks53daQoyH/cFIFmRTW30Fp6jS4ApFR3VpIe
EqD/wclBBrHbtiN1UrPYzwWcnWwUfDYsDwdRoW2MZ5ZEoVryAnSUdtGYp12zwo40+qZyhyTE6whl
j0ehk371vI2vJwoBM3SfFwHBPb7ihoYR6uTU8NC/QPYDZLyOLR9KqUsykabBP7zpWCV01Wm1OYn8
gSyE89Xl2LT1mGb+4TtT5SJ4dkuMJXLx/0zPjoqhbPxruO+9974XXIrZHftY3ivd/lRxQ4voshhj
Q/GygAzqyue7/kbiMhOGASNY7r7G71izc7fZtPsxmGHd8vkcC+oyRJKlNa87sqE0YZLcYadb3yjG
/0nFQx6YcTwaWTkjgjImusS3y/0JBRiEqEcWjxLyJB0rtm4n7OpjPtZys9VGMUSDMeQ4BxKRQmwx
S636j6SE49Hc4Qz3gY3fqwZpzQ1xsfWa1qeKAakNPlqm/VU52gww2DbwFfs31l7DHpox6AyFN3PX
mlk9ZVeasnyXcoUuSciSCU9t0sElgTDncjKzgasNgiUlTxizChF4Ls4QpIcTgYr1sxVansykIxl0
bQ5DvoWxA4GxzM7KuNEJRsbof7BiwNn4jaWfJlg47Kaj6LXoAG9pwDe9U/sfUnlaqtFCnJPfjMlj
aEjEsLDsEL7PWdUSiwFI2SttAmdKlxBV0nVK8yawERn27WJxaUw7D+Jl29SfOkm9yWMMIARlkj8/
cfJ3Lpe9Qj//PggweEXHg+m5f6RpE+eMMRl30aN+U2HjDjWe4vkya3EosQ1ONHAyQ7qhKTq9otgK
hdQHwpd7FEXQ72hI/V2v4yl0Nw4le5w2na9bf9uGflbohgJ4R8xKkrcX6XtlCM6TpNymYD2UqcjU
GK7h8mhwLEJnEvWVyQwt2OdDkKKrmgXVr5TmpO/tCkP9jukzrUgPO7VyHAfGzdhwxUKi2wiIIufI
TBrBZ/AMjDfT5rBTtoeYaqSdm6HyQoN7fHoSOafrcqCkAJ7yleZg3crgTx2hVWe3k9hY6LUHuSSD
KETegGEth51lw0x2VgYoW9THaA6UpdXL37keANp6OzMjf/9zL9z4IMGkmGMERejEHhf2gzbACE2P
OdLcYsyG6iQfqo91L0pKxXve5i7AwI9VV7znSWet2xYgzaVNPjbpSm/88dM9s2zRZWW0E/QjyCtI
e1OXE8ndYVmQ7WKBZNG+j8q8FG8XO1XVGtAc+NoxxAqGHkh7gHZXpZNb5XbdfFDrq8xOx8DXe/yC
908w6caKVcXOPPNrjGz5wd3o0gs82rwKdirUc6zj6hLjpXfv6wZOVmz6gXsQmxA2JZGrBbrGLIAf
1thN11k9M25KjFbqciqXBP3533IuzuO7LNuVIwuZ2vndtbRsqII4oRfat99GTzha0GmCpgY5LrET
MefQJuJOZqP1O2vqCFCZK2hKNiK7EgEGGWqklaxTLu7iQE5eNl202goMOWwKpClb4Q29KBflBUsh
ZerjG1f3xi/snQDDIH+CewZjfFFpqFnjaY6xaT0Q0JG/qLadbHVloFiJOIDW1zRHQOiebxW0ls/y
Oce1xxZQCItz2gxozJgZY0tPbDmW2wl/W2mni9ZOHmZ7AH2907No+Za4sfqpzbXSjUhbjM8dEngU
082fTR/658QsTjokEIwscSV8fH9xFpClTYSqF20+tFThgGURTo1qEQO5jD32fIXhsGBx2JTT6Tqj
S4f9b6y940EB3gNDnFsflfzmWKtDb1I/fFsYxc8J4H4VC3y7Px42aZ2d4syQjmafYkM5nHUpeSTp
cYH2YdkIo++siRlxU9rt6QNPf/NI+FjxuednX9Bh7Z9MnqsDJcjuVF3oNy7+2YgZr7/qo1KYQwWs
Sq2ArDR/fNwB2ooIKfHLZ/fEPvsTnDD3PigEYhvx/odFUwfQQZEPljjaMoaEUZM6nEG7gXe8w0IY
KKnqMsMgYJ5DNb0iuTBfavQ8I12XGXVnram/UEkeYTrueCixjLtgixKwy87OqN0SY/P9FHovBBrF
drFAmOlunkNc/5eq2HhALmrQD/sSSOoevutmKSdnorujmo66wSQrvWrKcTY3QKHgYhgzcsARl3Bo
dRBrpG4iSFbtoeaYbuTWGRsU772CzIIqd34xHh93v/VkyoM2tUFB/QvJdTNktvbKe5BX3s5SXFCy
Td3mQQD0LRKi4xQiWrofx1Pddiqe3HBA/axenNMFjvDCYz9PM8Y+aSrlzp9pdoV+MCGG9GEpmQ4P
5V/llX0dApwvPjX8j8z6m4z1uLzOnk/RC/7hn0YKKfqBxvWnu3DS8cxpEl/34HoVu6arYRsJ5hHf
dOBARrelP/j838vo9j2zDUawBwLmzixvzsBWH0ScYYZLB+l9lgjADa5mD9SPxQMUauodz7AJ00p/
7O3YzD9cK2pn4uV+kFzc+Uvw8n/lOzeXmAgENk57+lO1b7O4c13rTWjYagEJ3lN3C5Gk2+yJIt9w
kTG4NQPEj1a8gI6FZpuQbFxSRDcQ8997CW++lQQuS+dH51RzAKqTwxeT0XWeaIXP/C7vXqQKGLs2
NVlHXK7Hk3zgq1yAGdFbTXusAKmDOrzzCnXCJ/xLvJk8lboEGXPA3XbxB6KhGQ0jxp2wT8M23xLh
Cy14aeVTZ+GghmafGWVHbamMfVpsgsjPWrqUXzoVDoD0a7W7VPD/cxiJYkwcGWmZT6wGvounNzg1
allSllgMwU9qI3QKdjKS3mJmNM7i/aT6ze/6Ds5YlFM4Mdro27lgDgYlr66bbYkeT8VOQ+e4tBjz
emH7zuUX8Zxkx3O0pJ2SoU4K+byrqS2bhV6bCvh0UPpg7G4CCez9u8sWHHC5k059C73qHszVepHX
udQozNuuGelyVCJkYtlj/BQgvXhT5YnHTMgl7xpJTqM1jd+SbKoc8hylVsDZooK/YWzQYpKkkZTt
rL8RtvRQ5kdmajtGvjro8Dkw+QEQEGSHW6Z9y+/4TaPNjgDPusNLYyOoPcaGcPL6kasnng/cDQzk
KchFfzrCvxs21P+je4tDxZ2zRgo2kFgqLBriNHUD64j71KhUsdx2qnDlghWCqgv8x7eJWEuKqO5o
THlWX60K6M6oUR18YIu4bliwd3/vfvPgYU7UseFrAgZdsXpLEE5ZH4yoH0Fak10u0L+Ynfddi+pV
6pwKn8Kgnd9S1RetQaez361XnBmuhANVFfMB6O37qYtamHF758K0rc8zAW8zU8KKIQ/sI1eJhdAn
M4udrbQEQlf0u/dR7NSt+LmNvTJ/N4YOHU04STDSc2Lr/eHwen39SigsI3uekv8XYPuhegitAeLz
2idNNufkmaFGp43nyYo3FoIJRtSnjSYXVtqw5/gl3b6KYc2cHXTJF2iuJQD7s29Wzn1Jz1cTDOVR
WKTA6y2yC/Yu1eVDVqpIjDdwhTIYSBW6DWt/hBuOpEsdMFkgGIN1755P4yEuA2CSrW4jwerQpjeI
VatsdFAIPqlT9wK7eB8E653WcGz1vCleqX8YNi6nVef5xdXND4y/i4w6u+GGr7clWkIOYYjYkbzu
M6yoVhAPQjUNr4Ooguqr2p36iJg8y74KdsSB8EzwImZSLoOuJU91xNuONx9OHh2PQZWcQfB2KnsP
c6DH4A/fUYnf50225B30MB0KPmfsN2+GTL1yd8lSllKR/1yT9ATIEntAi70mTdVYiden4v0GEQGB
C106THN3vF/dTe5kDBPTT6HAZ0ltg7af6i8FOh4wuIV7/EnVYYQqpYBNNL+0uclbv4+MLgUh/+5j
BkDDEerwE4+JZrhWmqQOo3JIHAHiQnGZoUiulhyTmnF9tCjP+LrtKhf+x2ujpb1dNbhmDqg8nX6T
8AgPYzBImmAT252hvjthurr6PD7Fpr5jsZKLOaCartmnTrAqEqzOISk/eEkUA/sg9uYVyLHcCW47
oWRwaZXM4Es3oow+R1ijZ7M19Du36BnwHJXxwZ8XXw5rkw8g9FBcX53dUMXWyKdrG/iNc5gCjyF7
sgLQFY9AUZ+eysrKPoyKE49kvc2RhL0jTnrkZBy7tYtL/tPeb0S2z3FvxXMlxbG1DMHl2e3TUvhT
h9bAJCZp+EB6JDByF9Ega/jjG2Fk89tOltyBSUhI+Ms+WikP0/K06UI2b6ymk2uKtUEnYPEE615S
S3IDvymBMxpoQ18aWkw0i2WHfHQLIZ1oi64lBy12q5UPItcBA7ae7uzlyi/V+JIO96K0HrclGdht
YLNss7EVdhOx+fjKzvmlznh4upn8eQj6IvpeEoZ6dUViX+3a8PDIm0O00/pk5EMveOG8xRXe5rEf
wxXyFXOsloHneXd+bizKUAVPT4JA5xFue7E2IoWbvVgJqrJL1mgbwuepoZrJfSm0di6Ztd/xWfYN
+wHSFjfZiGSiZMMVl3jpxoZFrTkQtV7wQx4nrsHPjBeUbpvIE6CZ919mja9rzstcCcIZsmIR5Xuw
kQChyUI5CyX0P/C6J6WUYg2PfjVC4SBog1dgys6JFoLZEthwDlHw5mthJ3w3u1R07UdnpxR8QEVE
9tu780yoZT/uHoHjpmW0wbMxUVcYNiYmvGaPwzmwHHPfyv+qusTOMUvYtpX9j7rzPqucFHPZMoTt
zKOE+nWO3Ey5uKUibzbSlUcQpJgOaXVvLBu35GXxeexRHeYxwiK1bESTH4ylPU4XspeW+isrGqmT
rB5kdaakl1LpxSSPqklgb3ezb3uiXEBVZgIb0j7PXSrx6uGgHZv1bMb5QgXv5KBsHX5W+XqBLOuj
+2eV/88NCDFZCmKvB77bLvnL42kDsoDmJbITyBRoFEZE5U3e8hkiA/gIj8fwSqonDkTLVJ6z9+TC
0ixg4fkpZ3q1psia2OBOZmF7dLMFoApnxqy8ePPaYOHpm0UwMS+L1NNkm+zEpw0VQ2d4vzo81Uqv
lOB9jsbVwvo/59Of1BIssnNX9aUskdC9XZjSpXcIBg9UNAqCFbaaOCAb6zH0rGQoDeM+lGC90ZaW
n6i3mHwDmdaNq/iK5dUTbZiYW+p/bq+t4tZGQLMX1WlkLKRMeaU7ODoYmeJ4d+46pqOHK3zdO7eG
3CwdAtmKIPZD7u7g4EJ3LhJv4plZ5HD3gjXtDzgEaUmJCyQ5Wl42uK/Mfctt/lxS0TJEvw+0fAsY
zdoWIxoMclaXp+YgGELtykuNqrFrByCaBtEPJ4VYWetYURLaE2tCVtqnVvRxPSkGIPvImnj7GqIn
lgfFHhaJsImXBJ/9+R3v+W6XP6Zf3EpS98pGahiLjrs//W4oyq/4WJvsFt28slT/GbtNmDX5OL0i
+r4XUXlywrMoZPlWKmILulNoNF7OBTLHxLHex0/JGP5jV6q7CNL/0WzM+1u/2Hhqm1xHy3E4MmlP
8yHl2Rsgqg7suKdCeCDhRupWzC99QWfOHdS1kSX3DiQvVjbJlb097o1lWHZUw1fDLIayRR1GZceo
QH7ii6R5T42VCPWk65ELGdw7vo50E4+X7DmHpeiLjLCBjbbrTlwCrKsURez0pnPnE0Xt04JEVtzg
yK8VcIDCHHfxbvwI7G+XO7qmVNOJdb98aWuSXjFK36dDdDznzjKTAa2tqByiTaVxVrVrtivq2XnV
nvdg8YNmPTQXFF91eTwWQR0Bw/oP/JUYqZFFrKamk4rqBbOsssVU6X47qB2QXf/S9lTeCsQcfRKN
oqAdZAuBtocsLg16hp5RlJD8Ix76HVNqf7qLlThbiT54g9FHnYNT+RLNpeDYlLrYHdL1Af8rOh7v
VYuVveKHkTG0s+Xue5vsNbMbOEKssJBvopfkew7DuA+q3Yh0LQGqE6wSoSmxxsZGUweFkNt4me0T
e7gFaNffBFFjrL/0DLMrFh4wxuiZlEAOHpLu2tJqaOEyAS0jGnLcFKa27j85uQHSCqjHk05HG/lX
txXwhr6c8PgaVbRWybEPZT6gf+htMxYLgZEfLZ6VDdGuTy7jzQhkdvuuBGccjNOAoTcrBrfJ6PCN
35Qe2gLK3W7OaGW+NiMu9v0AWkrBUTYvP7bH5bMidAJcYOUBTa1I8KjoMU+IQMqJz9zgLtTBdhF3
cO47etaE+XirfcAeJeDm1EO3N28wdC6eVUUaEQKQK5uzHIxSRIriLj3PiXkqYxBtZf5N19C4ccq/
XjzpdRRAjA8dWp2375XxUrp5smFNbpBtcH3aj4eggOMZlxsw8C8oGO/9Wu7qX+8PdoyZj6HVBpB0
1dGd5soQosxWxOtr9w0mc8P0V068VykvQPsWRTj+axZSxoX1QR/fxCeOcMyAR1+C6WJnwAQBf7Rh
jBiPC/RRYpddibqR8mAWIA9b+ixq3QFIcPftEZX1FVAiijHp7Poyrc5K5GpyQWfAqxKHZHSu1iZQ
GMGddFyaIkhBHPrw/EUiRkVoUUKB5cYj6zTt+Zd9YmSqLc81dFQ+jeh7O2TPROuM7IkIVGQ86pSQ
4xoLawbxMwk+p8N8T5xMOReH9qf2aRg4XOnUCz1h3mQfBGrO/WJMZg6Ato+7tjlVRIXKYcYGB2H2
npIBYABaCwpfzGZYF94zzHIk0OS/5XtcP89NZ3qen4gL60tJdPRYPXpr9gcv1xK+lttpmqZ/CNL5
L7qVagIm6XnN7iFbw/P2ou8canDzGLoAWWYCg+lIlCizG4YkytkG4m9MyxuKsP02bS6yW6L6m0pT
tklEYKqKAmUjiorph1xIc7IIpkMJthsZ6O0IkU9fBf2Vp3LQ04KnrKWVLWeg6yc3RVuhDbZpK5pm
WEdCR+qpwAdEmsGpjIH0alQ4rNERV2qjXJfbOD7pnxee5r7CbwtmStf75I3b+wdHTsmIZ1d3ynQ2
XYEpukmuBWHW4cM3L69Jm3BtodWKC4fpKqiAh8bCc64gw0TfnHZCsrRCXxvvqGSvfdLxUwn91Amv
j8zqUo70A029j7iD7VchifCVVGN7UAZI7FBI+Gt566p1zSsvL2CvEMNXJwqebgJI08tLjMQFi9aL
dQxXL7MmSgetL+RCMoi/+nB71VMgkes1v8z07h1j925Ty+LxpdXk/Ak1tlP5ftjl/aGu3ZYVgSdJ
Onwi/rIwoidpJYsQGKcombm4CuN2U7iXCPHHX/9K/uHbJCnSlcHGwlydALyWmp/xLVCKKeyW5d+f
KQMhm7zrnaG/AEElgi8QIzUQfmt7FpwYhEN9raEd3cJcYEzUNWF2R3oktnFcR/uIvdYhkWV/MZfo
E0+tYpOOrshT+UBOEwArNTexUzaVzWLv377tjDBEvc5aW4IDNWbLfG1QO7tDRsHxpoE/L2E0k7s7
cMLA+zmcSKx6Y+BDokXoWm5Y0eLlyfZVrKQn1LEJqsIrnzQmCmPmhMsUDDQoo1BiEuAb0QrKgSSP
DzOtN4VKy5BmGgk912WuS+A3+6knCYWCakYD0YrfhB07BzbCECB1iNZOafVtpEajmCGSX5PvL9LL
z7Z4xyTkFHG55FaYiWZNyUScnf0T9sNp0dqes14hDwZAiH9y7OfLfZlyKAGVG2spPYl3WEl8bGZX
R+GsCxt7934OLHXKQnTUG8XqexvNvufLz5dHCaOegPDkafAkWlG8/Vwvae7eIe6Yvz3a+ez6K0T+
lv0rP0v15oOVevpz/kyv+0C3/1DYsmpbzX77awN7eDM0d9D0d0agpWwB3KLkZL6ybpr+2aAPCNAt
nhHP6mLb9EFmzHzyTszGf4TJohJsan/HpEno9/bH+YjJehYor8KohZK7Re9C8eJCBpo5ZAEqRAPr
ZQyqhrCZDETpttMp8TFiDML8UIsLZmun/f7dhVED6vEhi7g0J2/G3CAqH2G7PSLjfMYo0VUkfC45
G6Zpzkdnu34+s+ASsXYJztjK4fb5Xy9RfrSLSx/TjKdIYQzE2fQDXGjzqdO1Rcs3maOLIWXt6R/G
gIYzY19YTh2JaufIfHwikT8sLGhFeCr7sqG/S9zHucOtyYG/v33Nm3mzHMVIOVokEGu7NrNJth+s
ax2raVFv/TsXHCEdTSr+Z60upRShAMk3H9bQ4nhWWX+nOdXbRWtB4CgFbtu0ZSog5n01tlB23+aF
QqojxfPmIsx5tZYDlbD6zqdha+jUFk7Ymv4QbMHDauRniFoLwCR2dsyZUL9Azxy4127pPiG2Y8En
94urAP4w+Iv+7K5If+RK72J47AWz3BGOBKN6WyOtcJNKmmne3wab+ERXcSRaa2wEiZnd4RjyXDPI
02S314soznTjGEdp+kIdorpnsiSqzTU5dABO1dRRDryT9uC9nYEY8xBLKvxxFCrT2xc9dzje3UHg
nZb2Owa2906XWq+OqMlmQH2k0b8lJo5tNc+w83BQfNpND4hi41BjNWgoUbOClQ0Vsq2WuRbVA31V
iqpi1t512x9bToxA0vns9ozd3oDVnKhbnsrEA2EBMda1i1nTz/J1cAHuUsPwBfCvvSTCBiIB6u/Z
jY7Qa80uFf8EtP8SEvTp0aP3Y1jPsAuYsl1H4i2CdGaC2FgSf6k7KnO2rtnNgWDFly0MtGAhsfVH
b/6GteNEATooXJq2CmHkKo6h4tYwhqY23HPVQbDN4UmAdj9qLqx9ql1rOrRGPr1R7peR178usp+N
gGZECfs4USRNXc7ChUbnbE7QricCIV8bqJAyK1HoOIO9cuCGStgmcoj/JSFjfgE6UkwFog5UdK4t
KOxld2Xq6AcLHtr+nkgtG5Z1Iu5vheYlFEo/4RJxHPqtvcjILbONIziZT8FuNCkp+m4UK3/61t8z
91pVZ2dTLGB3GnUZ26m8d8fPG21PjBuy8tHvTh4wXrv8VUgw2CZFkkrprT8+43eLmcAXPTiRSy7P
ERb1oXwcrrvYNOMKQMA5w8/DgMrTCyCDzW+/q4zCOEmg+agv0RNagwBtmTT7WPKkvB0KbRB4jkHu
iDwfG7ma/Uj8bSnFZicA6B8OZbXNkAuLh7sBu16wFFfwq2zvDmtiJnT6RMockjaHdy0fcoY+JQ62
oDfG1qgtIIoUKwM51znRdefwU6eYaO3zkGSh1ybYn18xI/jKbv7JDzwvT4R0EGx9jR9InGdlLRkf
un6eDswMDS8UyQSqisqNdmHL4MPAOs3B6QcpYUjYhY3kWHHR8CWaAsANIyTBKr1y90/PZX957FM3
xYydffUHnd5ae3GYWpdH+zb1pmYZAAYpakvlq5zhNgoBchJcsQVZwf+5vCZoS7DVrtv3ljZ6Q1Zg
e0FNGZAZFD7Isd8ScmL3IQ/lUqVn0n38xA/UCuEM62GZ6DPA4XXtFlGWqK4GhdO3DDr4Q7SoXrCf
+xyIAMfiRQgu6rAZ8NaNIPvNFBEdYaXmJFyNJ0zAfBHFGh3kqI3hGTBIFWaqZpSZ8CGhOeH5wB77
nAbJAVP5b6gb1G/ZRtSEwsNSTZMKZncA9ZcAaKecMEDr3kbh+nAe0SfxlURyhk+7cWPwljvl9k3c
u+uJhQYCruQJUzH5j9Dt96DtJmMgNYKPn3xnGf7kccnT7iYBqtarx4laMXyuQu23fO+5l8xLe3h7
Q3jwNI1Z+1bfi4X1cg9wq4KY1ifd6Il+iAnBm8NtxSEV4hp3lDw9uoRVXOkH3xglPDlqEHB0BPc0
A4GMJfWFuEQuiTo2fvpcVdLURAyGNMGUKh5+26V8xFuhFTI1Osm454h03/zrQd/7GRfrib6ZFvvp
t+N/Oh+nfStT9arFbVFIkpwIZBLKukUb/k4UwGuFZ/wivJ99wOMkULamK5bhDqAg3tfZA7kbjfBk
1oBjaGqTpVAP0WAnYVeUha+xcRCZxD91BcUVSfJjZ1B/TNepT/yLiHf7bFmP2ZPHx+axluQRYljo
w5hbe+6Bv57NByJE/U3drJWZ3w3xxaZJz6W5YUO3pPKh1l7GKYrDFcdArNU5O6bLLI6M2vR7savf
OzcVOWRwk+AZZ7/VBZ/AY/FHnMN0CnwKlx+DK26IE8Po068I6UDEpLAG5vdNKjqmIHnZgY/97f4u
9Cf0QzUQq1d47JKBCyUjyK7Osln5/5E+UyA1pu7UU9L0ucM+s6OKObL88HFcsTQO+BSooAB35de4
P8wAKF9afrwwO8AyygssSQcHDJOy4kjGwvuavwK5c5TDZ9yFDchB3xMImvczkT2b2niHcvUuvKje
VsNDx/s56faKB20oW+m8qpAqcYkad7Y2dg5thOkwR//fkXb0DgjsK5WcUA74u3nuiBvpeXzVhZ7k
1bQYFx5As1SFSuzXjArhvn15D+6+aKVmC8p23DB3NXVSKsd3FiX84iLgN2SwjLF2t6qmrZBPWLcI
3YtTUoi1McKY2auMlfgYzvAtrO/+ifnPZq5XW0tzf866DGMxQgbuEGSeIQPFhH0iDHoGWkc7VdNA
/KFJpVCUPBWGgZtxidIi8hxKREOdtZuWDHWozSmc4G0U67notEAfBp9mDvXCsNb1lHqwHAGMgDcQ
43Gi2uCfOI3VZgc6+DpGJkrwWeGO29I3PfyT6Wic71q9rQpuIwfZxjRazGyt7Y+/fftMXa9HBaMz
Nqq+ADo1Ds5sxoqnAGHlT4WDvzbGOmQXJrxe2v7myBYmrcdvlvYznU4FGRLx64peTTWhVjABG2qk
oTqJG/oohcQmjPOeBUtlEj40B0b+2YneyuNPsYO0JVQboTnY1AN5oLfgSEWm5jlRHPa17GlVUvxI
3yTsAm2JvbH00XrtKOJNLMCTYG1YLbsmZdrYalEjySNWIC/gvviZfRfmVxpOeG0QT/fqdGJ3HjXb
kzl/Qnp9ZOAUywmwgCBl8Qp35zBaSTcJ/TdPWtKlAF9Oo0d1y/4Hk/Q89RMMy3K9mkzmrbJ9TGSk
wgfXMy9NssXi11yS8Es04/fncPJuvGbwwRlwT2+eAqLpHRKZ5KGMC0oA914Bbu5nMcORT19xMYaJ
r5jD2WWO7JFMiHm0Qrqeyy/Y/8eKXzJbqGkK32aAh+nrJxug54pOycU6UH3hMOtnc1lA0Wg5jJQO
oRI2X6HHPNvk5SdiVzFb/u77ny+oLGucZ55GUN31OSFtkAyK4QZu/iKoiTqAM1+VpPqFF6c08exq
VzYGL/ngdlbYRn9vX+GrHQT7eDseqLbGHsXrHntSTJ0IOLE2zBWjJrLhTTHHvFbh3pi0LiEaxiTp
nNwV3uO106/NR/+Wx8S15s+9edXb6iKNgMMvLYuUFV/MrjCe91Rv5/aPRq7Gy7f0yQh65GcmPHDh
0/fqUOFjsjSXokPneXgPT7stVUXIEqsTVhG/ELU47V9sfQ0KT8VXgGIJpfB6H1vO1spn0zt03hmG
Z24pgsH4/zKGgQEvrmbOnLoGFbXRG/sKAhBglD6+efff73oVUAgIdMmdwpPoM342D1b0jYSyjMPM
JdNtEg3FLXycdBTzCgUDUQ8iTzjQWyRS8xgjXsbozI+BvpKlp7p1LYa9vQZouTojbqiaO3kIYb8l
NsPZTcsiFobcxy46wrq0OYEh6cgiooCEtzpvFvqWQnGW7PW/LmKY6KSQIOzsdCTo/gRwhQTGA5Uq
Yg46HZF4szpUjTgiuiNiKpYAwSvR+18psrz2Tj+ksWjAOK5NWKrYZGq5adueVunAvSei8dZ75EdV
k4/yZYNG9ohOyOaoxv4oFoM51dpVFDILmv9h2+2u3Z2fprrcIWyXOhN1/MDrbbJNFjAf7BIY6srF
XRlu7xcsA1iSCfpHUqiUwLGx1WFmgVBz5Gw7W7+EKo9pz6dBGmTQa/lAeno6DkhGdzPc3ulPsCAD
thDvPLTF94mw/NzhOpflPh5w/7E1cMyqB2HiTDfWZtQh9cm1Ockj/kq16mBCAy37CwI7GbUJz7r3
ea9ieBGrXKDExbQAAuAxuURECUwWYC+GlZqE6A8OjiWwJUK/AO7jBTzbSSL0gk424/WQbI8pYKJQ
NLPG1JTufO72KH1inzIQ9kkKMchTmBjtMJ23oOsz7z43BTsJszkJcj59RO2SLBuL1x5WE6ntve8b
nj8lj/kcKLIbKJHTblif8voTfi4R9HU296eNPBT1gJDxKOMD02lFaFDO9JRSO3Ia4uF71ql1B3L/
nPQ+2xXbaerpTrCQCistfHImU4b6A0UzlQbwcZ61lBUC1dw2ECB+ostjwyTFvoEj7LtCHphmxq+6
Cp+wqIrX6z9wpSx0qYhuKFWp8bECsoiZl3q2sawbnI5emoKAthMoBSaN+EQLtQjPkBIQOjueDh6/
vPO18G/dxcgqJ8EwMLJ3ELGYuyo3Za9EYvluiBdG2TDOYaqPiKC10jZ/wqko5/BtudLbvRr6Yybx
s5HR68L4afEjQvFS96dlhL1EQWVffxHgHsajo5IGcJJsadvFqZUYMIUC4TB14hmSshQ3yNCLxwOE
skHekeQw/WmNOBPyg/qGVDj4lAmZz+tTxfz0xviEn6sjZYd3bGDhsYTbhUavJUUeiZHqBFWSzVc4
9GI44tw8UzRuxwZ0POfjKFPgwIkesR2JM/ULkGxltQhDdbB9aqS1CCyjdk9z96gqPi+Qp42L/Eas
OYgXvnwmcGedIym+Xtu+sF52oHkq2CJY2LVnLgA6UD7bvL7k7S/STc1ehKLli1mxxlnVFvca+eDt
bVS9WR3jZyGinOyX9K9uHAi7YpfseAFURBJw3dnIa4SRLMBhkIpYy/zNZOh+HCgc+e9vTixB4uTt
mkL1nNtEAjFbvmtty+RiMR3jN/6wIsFk+XqpTZQQjWJFcKIv4gAT4Yrn3NMtIA10+GNzWFhjwNpL
Wh2s1hGSzaaRthDytxr4Wzx+eOwGbzNRP74FmwlJDhajbO30RvrmujPjCjKdYrKICrGKFmUXhE2w
2Z+UpbQ7GycW+ln2uRyUOy6oPBzNy2rR9NYgcd3l5J8ApWIh63tZQLzY3Tk1yz5pdtG5Myw6xtbk
lPWTmSXmaHvDtv3zQlj/F45OGvRfWUdTXjnDq4rRPWsC1negH+DIXCXNfqA/k997QQTbQx+U+7gh
tD3QlW55E92NY8p77wTsUTn3nqL3IYip4VpLgHq52w/9w5/eih8kCXQfyb0ZE0RdWpxgwhodagE2
Fgd2zn922rkYMgFQCiJfFuJO+9ZBRV2NPeLkv5VmPu6zHxxOsn0kj+R75cmz4cpCK+q8mICTkWwX
OCI45RZYZTdBH+F7j1lkdXNCN0g44C6aycBirrMnqJzw4TwevcI+ItncLX4vaybWCeTaI1Z7Q8GY
9pUCK3ziNk+bnOPuGfX7xfGC8XnwWJO68C+dg+uFde3xqfnqMdvJsIVSku91cqrOXQffOrtSOO3f
zqPZbqvok68QYe6pBYV86oNGQmJVg6Kk12BI87w4AeUD9EDaIkW4v9RqzkoU7itOr/NRSnmKR/av
JxiAMjHqE9pFMc9Sd9EotVYXSAjLzRGlIBhTwoJy4+MHodoDxWYhdTQG3+CIej+83fWY34UsJ5tb
qN+3Nc+TGgctcOg3+X0btA+v58ohEMMYYvSy6DqijBs1+cXjHxuslK0EDbQDTFqNacMxZzzpXAeD
0tixfPBDQtEBHN8WASRHfcyr1D9aRddfZO0Ajh6zzxirVh7Qffj20H80wK/12UAZdVZONKgfk26v
9cUDqiB0lkWhx8clNUi93jrKN5rsxTPxlql7ha86EyCXQL99VuqoEH8q959VYR2rcWXiZFM9PqgZ
NHqH84WlIX3r88MhtvIlutwshUgHl1nNq2XnDmOhjwcN+He8VBCjK3K/BollMHyaFnEJjegUWoFU
vdCG4A9NRZNhrdL2yx+FjbB90bvMRbz2UnBwt0xlpu9L2lsLzDDHDWM/dHtNmGO1Lec9uXzhMeS0
zHUviLuigyvptGMgB+MpCWhpE6/5hyPS2XQ7Fb6JfCWmn8i7Ri2JvbJUriTVuVbjqcjs+X4fWgGl
XYp3+z+Ay5XDanWTP+yCCPHARumXiHCFoqt6qsRITyu9VHER2AmbgWbygcjie3pIflCUXZyaYjrO
b3rNxL9bp/9PVEVcbLN6ByVwt0Feo/yEFWZlnSwAp6wA12zuJxED7nFKpBbGMY0CgUpYy+f3+TPq
Mv6qF+rtbmW0GoWIVWKLhNqLOzWGH54iMZcorbD3ii1WkVsSfFrEk566P77sO8wHO6X69+DSkOin
KqNMt5u+67RkN65ln3sT725UD6iXw9QXVTgTTw3eUHLlHCNnX60a3pU/lf2b6szy6oLllwqYv5N4
qXdBDTwYnzmWd0ldMy8z5kzaImq8g7lY5AU4SpU1j82QKbHT2QgcYCZcNqWNgCRtFVpj5GXLrSAJ
ggbHLrKkR2BJ6mcAL/inHN1qsurH13S0E3aLmBUTI0y/q2Ca8jxpnqr7d87+Q4XZXSHaSqg5PJtt
9cv+NigN0blIn70FdWjKq42TDxtWx4+6Ktqr8C3HFMeT61S5lVSOvSZ6zIiEzlGnc3cok0x/Pl/q
T9OrveBBTekvj7Sk/UYTwT6d7czl8oD9siVxoKmr+cyJv1RlRuOsAuiEnAabD307Gz59+K+4kJ0N
fpSFDQkjAPbqR26Xs6p/zcCY4q6trM3q/MzhYq5xtE+qocz/H8QdMNBPlzwOIQOKAcDHtS4yWZ6H
7LJHrosOiPdDCmpFMTpAlttb+mX9qu3SvAa+Xj5KZ2QRrJFfAD7koV04Igscg7ukN+Fk11bm1nAT
7f89J6CpUPh2f7lrO2O48eSkxCzIjCpj+a4JIhCRw9x/p28iMEDDgpFqkw0WTSEguKh2YOQbV90A
6yQTR2clGKLkykHyMr9F3g0j3i8UKEh+xfCApa6ePRBcHBSvUyTdbVyFHTgZIla1jO+jh8CnuEtR
/DyngKUK2ClFEcfBKmVbN4iw5acOCuj//EU/aspXk/I8KSGrxa6wsVTJ6gPFjsAZJyFCkFY60rP0
cyawJbXyHtz/qcZbXtsmgMrh9ESgVzjGS3Re1Zi87awe6to8dQ7L0RTKnjaNh/QgAHINX8DCSY8d
zKoHFJv8ecWLE8bttRGYJGBfgnlwsfDnhfv2QIzKXtL36zsE1UuEp62MwIXuuvRGBkTMBd8+uglR
HCbkrVomA1evnDMiGYr8OBS91rES2keRf98hRD/ouRpOT2hb45XUmDOWIAtRRx3ybxhM2ojE914/
AlsS6KgZkzHuofbCsdgWak1fkvihYwp8w4duxMSl+tGazg3NzX64EJ811cugPxbNZswKFPh6NDEC
nH53aPqOVzxajv0X32roqEE3BIam5KaELcMGq/gIoGNIRLyhFcuv1uS20HZEI2RTT7TWtJSeErM4
++whw8nVsJ8JwvPinmm6lvlXir3HEtBMIEJvErXNKNKEMyJxL6Ta2pfpuvCUzscRwCvTAE4eT+vT
Vkv9B10s6Jd2jQUatLeE+u6jmxPNPYVtMWkPTls8yruSXra1c4kL8ELVRyGxLY+nhcm2Rri53F6U
feiqAhsU1Ij45z4obhdQ7stRlumGp0YxB7+HnT9YExBJGnl06S8reJqmC0Ne9EyrUYhIpFkkANOq
wasx9pO4f+Je0XW+T7A6fCncJexVaBOfF7aSW8HF843OFBZithC2zn0EE9oSbmIO5IwHPtxTMv1m
aX2BCOENzgtNFNWSTQTem3snMN6Xq0RSTh1Vyq04REWua6yqYkrU2gCJQfF9clzifbOEW/OJQdhq
EZiOrcv19KrThyxEeiwf/1ua0lxEdpzpQ/HAHIICbQ7kq0K63j9NtgqT1PvsLu0TFq2KKki3yQg9
VqyittPA5VWA6Z3ce264LY0rUE0x77hSMnJ+2DUEBB+M0DVHZwXtrJFv1jRwiYaG4hlvooCfJt3a
AuuT4bFwLZ7oKyAOjls/qqrfHPgrHoDE482R8PlasC8yYjgCGVUrBvCCkNkz+YmqubQMoaFzmGG4
PpbJbZPZ5NJOS+vpTpuS4l6WuKw5tVw38S0cmv7AyXrTwTHW0InSlW/AMrGQsLpbAlSFr0M4DukJ
KEzfe2aDlR9whJXxDtNBSTGNNzgrghLTPuQyventbDUx/v3l+aZgwQqmcaeGMps/JQZ9LUVAzyXV
p0bz3c+Gf9w3Xsop+LDflRd8bmMDAD+6STHzT0KjE5u/VGtGbjIfIoXZEtjltvjtjLIGurd4susS
lT6kv6HwNgUlKLA8CKbpkAf5qsAsmNZM5d0R3c5BuGjsmIdue8m4f/2uwMBvrFKlxce+yzRf7gXD
DPoVn8QFf2a3FGDN4FngtZ/yHl8NxCDNPKviMBgAPYmTWeAZX/JIH9fRGEYUD8gyba/+bt9lleUd
/Mc100RDxYdO8DXE5BVhbNyfkNNJQbObrm4vjitQZIq6FIkNQZSht9UcNXfZKxFaPy30nhdQA7Bi
aDgrTL81wHeETKhuSdCV9ZwEQx5gwxzN45kEO5WQg/uPub6TmfziU+d2i6MjGHSrmiRHq87/PLd+
T3Hu84WIwLmHVk9zRbMQikV96ap8aluMtNHlvQIFh7HhnBrczWqlF5clW28EnQ1ioXp9iOLAHBJT
TiXfAMHaWzYl0QJHkk4qMaZ4tddGKHwsNljCyH6kxn9kCAhEcpLD3KAxVWmV0KSXbr5FSWze/2s9
e1L6gHYi2r0A9R+ZFDb3kyMFNQ1Pe3gqZNoAOH7ITohMDFKuJZ5g5oMfbOAwCfAOYl4M8p/G8K0s
ppYDRyulyJGDTeHiHugpWM41fFJRUruhjRu6IVeMt4Zbcmzomds6WJyquAvoChHA3QSEa1+0Hf5U
CiNYQR4S6iRTPMguHPvEGXGZF1b2GfEIhVJlTkRF0QxjR9kh0eFyM44Q/E298KzTmOCl4wqxLJDb
Sh/tGoGLa+KL3tWsJggicoSko5Q5M8YhGotMpt3xqoAO8k9RPrCLUe4ZVc/7Hy4mlptbG8cg2VqT
7KjE1g8hLMN6nRZEbCYo6LR3gxSKX9/qkIrLEwQo/CiZLuXhk6+5E1OGdT1NfqzpeAWcC4EH2PgZ
Na/hW8fzy6vOAGfZuAqqbEDuFUDSibLQOSsTxpD+Xcg7d949l/9Po3E+rz6QPZql2XEzC7wozkSS
AbcZJFjfi3IZRIGNRaauUll4NqMCtgfp0kyagMlwAx48fMr5SnOXeu+2gZlRJ+41mSCBKGMnjur5
sakbXCfkB/d0CIlYlSY1yYbAP7KVUp6Pfn2GHWE4FYASxsvW5FHIpKUy1KzxzHNGtDGSqI2YJA5Z
lkLEbIQlg4bvgRxx5GMQFS8uaxJJY5bbJYcOPHuezdhhrUBc2zs1lTBEFs45rM6DztG8k7w4r/xH
vhC70/K+0VYDQav3bT3jhp/OvCz0oXBwktDjWzUdnCE979Oa+WRltOw+kYGQ3BHIqO6paFDNNE/P
C/mr23GdjbIrjK5FD+ZHJ26fEVjfsLJQkkAc6hNNmkJQPA3RpFXtyHXjIWwJicHtBdbOKdzybmF9
IAx29+NMvcmpF8sXzs9rXsZaeo4Zl0OVTnCGskZAGHtoz8QZCHegYv7XuPm02ugZKurcneDNL/mt
UOeMgF71W5key7RZL9fCKSm3tjhHdDKCUsTdfvgtxqMZuMhMP9jv08kA18enyf8fvqblZx4eaXWo
OreWOIsqx+fUpAzJBi1Yp5tY2En7Rh0zPPv1atLII9mZwV29iw0GEMCcmSHFKgMr4Fo7jDOWFD7Q
YQ9rTZ8Nf0b+BTMkjBAYBxXRWYhL50nxIQ9yysc8++/M7+j/yswoyYALAuVcdQ20p7dGj8S++Gea
KQ7JjdPthE8ha2BssQd7i5fdUhd5h1BbeE6T7gktmSJexqRszaBDvetEU51WonUVVKtzkh6+klH+
4v7hxaOxJEfwomSiCHxxXMlj88pzu4y4B+r15x85cOLsThvbarlOuiEO6L1MQ22/uJrImxsFF+SU
wT9SHUtJPzWhmwrJLO6IgHZ+vEEqwqbN97eAhgG4kgz5B13bxz6I69/nYBKJYtcnFYEM1i3S8Xt8
vu9eA4bfjuCNf8Fjpw1jX+qzFWf7Qe72G3EVU6bDEiyt8U5Fh/TcF0NQFzHGammSn+mwMvWtq7RM
ZEs1hJwhePFy6Jw+CIdz4InYT68QaacWn1CPvqHA8dRpuB7SjUm6uWkRBlTZbv/v5Sy+XgTAA/Fy
4HIm0K3V+muRShTAMoToio2jN3yAXZFdEFiBIRnO2iKiWilMvup6qO//EtSJGGB0a7rrRe8n1Q0O
jmZe+UMMflQ6KHYJXAPsOPxS9ZdbarbP9p/QDU/s3Kb1kbm153WqFUTYChuDIyh/zuaThF8bnQhn
MJ0O9TkByLim+gAjDKDL7a3vP3/vK5OqYvSg4oa7qM+uxeSFQeelDn09EIBIldYR+WaB5ZVaeoy8
QaScN5nj4HdJRNlvKd6nUvKaY+egv8OfR6Qg9s+PYC5dzMgXocevC539LKSQmMUn0c674MissH5b
TtmSPEPOjfv98NYCFO9QUgl+3iN6NDbJnCz17awFEG0Q6WDqRot9aSfGnEYOojmzZggWzEGazsMB
KgDf0t+yKsnHZVDbEZtrNLfnBOAE1NWx62fwEQJ6Imrd81VTTJG1bU/X8Etnp1Vo7tZwzbkMaNyW
pGBO9I+8OWz61Igx7xgAM8+xX9BxHwy5ybUZ5o7wBhWPwvP+L3fDOukggvhN+ZPpJ5Vw8yTthadq
8hOz3si/BsVpcWx1F6Bn+Dmojzz6dQUWTqxffu42krwGMkRt834/NJpAPPuytbk3SzOurA2LRS6z
71nkkVHETO3CvMhPrs4vTHioU48KagHUu2uFjQh6srC75odTXiBGil+w5i9siyrj1EVTOP2KCJcM
1ye5bBQQedj3ADD/kyT5HqB7VIDLOg2mM8XCEpjKQm+6/uZgF9tI7YaimXRIFoAqE++QcwvdDaxz
rupjFJyqza+Vgnk6ZD0rfxDfP+beqI8Srer5tBKV5gSYOP2cyTuouoDQ+nZFcsfYS/YyjHODE95g
Nqe+6SM99GlGvKDS16Xrp5kwBf53eKvOUemEOwGuyUOaMy7PcrzIONlJYfhj2GqVe4V91CmtT4G0
fTrDlLsWkCGOFZjD3hNGbw9tycYLqykk7BsonKaXTlL1i7h02OJttGSmrhhUZv9SZNYVrFXdmqg/
c+DTeLdmX1AwxA/bsakyAks+o7MUXzhmu+JPVgCt86VI11Yr1SfKfGudXLiilKnowgQ9uxP47AvD
BQJ2DdN19w/sDJZ9TAYDhYGI/S0GL7y50kYb57KFmQ4bKPSojM3XxiF4wJSGVMB8xSKlp8HfIMF1
l+Unfq7kD5Wdi5TVGkTmyv5Zk85h9xuoCDRQdJFuFbf9suAJw6/xtChDbG9fdFA5xMT2kDp5YPq6
Ds2FjlkYLAVIpvv+W7r+uK0TXB9yr/SqyeYFIbs4DfgR+vovgpy8lHqCcFauQ4r4dLG423xq1sIG
h11pMwTPitwakw/SaLXwYx/CjanQYJJ9wXf9bcwoqPI4BBWy9lmDXQkxjTb+zenZhCeP/QQYzG+d
aDB5Er3+TocEF4O5inRbLWbuD6xYPymxaTt5TB85//658+kr8Gu8wTe4pPbsTd1/HkkXz3u9gg5V
XIiwSDUNCQI5y6QpwFtYz5Gw4pUeBjma24bEe7RSxrO7mi1/iO5T2hlPX4TQ9L+O7Y8ehySRK6gs
4t+015zjAgi7xeWJEqrWfk60Iwbg1D9ZEdTY2Us+2BSeAEsKVV3hYSbUxV11VJHA95Ycv3ndETTz
CH5TtBQ01gPyg02usdUQgaaj42khFs1NkPJoLaKRPazmLIXGr8eVdcwE1c5uYw3LNoKSlKMMfhf+
Novo+cv2+aycuAljWWtrzXe+f+nazvDyBV1vJVC7vpaZorHD/4I/OsmvP6j/2BhtBLo+KDcxvBmh
by/Kn0XDMlMezjA16yUNHelo7flykF5bxHp31wJXRESsW7OIgnjeARW1HU3LvBvcPEzM4dbmqhd9
Q4P44II5Rz07R3qUdlfbIMrQHVgdsSVk3ad86kt22QVYsrhdUivYbszw2jnT7i1MCrE8H6ig5XtX
M4AT7K+zX4USvmC7epqH7gl5bA4bruufB4+i26+g8DjeI5CwzE47N0tjd4MjYOqyNsbUfWXjtGU7
1ylpMGa/8QEPHvMI77SKk/8hHuekUTC7mirEQI/JVSuEYRw2cF1Veid30RQA6bzt3yBCg0raI8X1
TU8C0Dyo6VMg0RG/dErWaG1vwgBAyB5eXkXS03Ri564aexbLkhzIXVJBPZdX02e1b2Z1g1kukGMQ
uFX1cZ8evDed4HOo6NGFqyolEsXAZ6glCmxFRahJh+h2aNQ03It4hE8qFi4aL1PM2cjc28BT5uxX
O5zidIObfNlsadQVpPdl9y8tQzHnxABsQkBppt+Nliqvl3SnJAsgO4f6liSWQA2w6QG9aAhFJslW
fwMVzPvh++wc1Uy6DEOHcJ9g7NlXBuen8o5NXQ+jIWUAcB4jNzJIwbdb0SABeDHyNmqOj72vWlDp
bFCEXgSH0oM4EKjXqTYdugmrUCtZxZtu71m7R2klopCxsTVddtp7ISC47fekeKwRn/odkjLsrpTz
0oVs8MtRsIs/NfHah/+zcT4wkMAC59r95iht3WYMHcnfKzwEBET3cjtTR4ZVUoQKUj/+PbCMz+yp
6d3d0dmzxfyVc5j9PnMmKwLgJ9KD5pvaPt3IoUZg2dG7feonOREP3g6HXPOfFm5x6OiNAjm1ULZX
7SHlQ/xBSMAMlP+6Ha/QedE0eCbYUUMRS6xO6dm/vZSWdZ3M0Ob+i2utr500BngnrOMuND6EqFyo
+ZZvu0BfxhLOC6DIHsWLEdKGfvueXP7wNLsu2jeYcIlULRnV1LsuENq7EA7h0oOOkKnBZsoSMJdh
Ok3M7unK1M0hm5Ecl2f0htWoa14HR/uxBf8r3KN9VDtKVTGqf/Whau8Z120ZhE2dwRzYRLEt1Aa2
hBFe2w8jZYJVPewCl3YYMmGZ4wNBlVaRsXeeCsRE6aGdIDbhI30vjbavsx+ib7NmdrHwC/yt7fBm
2Uck7rqITnTf8wszyKw52l/gRZA2CxUk68YHEHQ8eLm7M6GPlfiTPpdFIiKDJIkxJO3++3oJf+vE
dfVJLsYUJyQkIo6/C+ZOvFiAkNlwFJEJUblyzUxsuwITXB6i4RRXR2TjumF27w7RF4P2MOYboP/3
pK9YeTHLoX5DEr2bM9PxFtP/gRkqqR8N+tpmIKD4Tky/aOYbfxo4tkfqPLzPXVZPv+HP7ro0LBk6
RNwTQ5JbSjRVZedi632Xo7P2woTlGZZf995JPpLaTBnUsOrdf7YvdhpVb8NzsVyFKyuYBSV9X6xf
09BbyvSF6hTZ2i11a6NX6Q+Qxnjlp7YuAydoXvBrZoyKiCfuBTQ5YB7mYXLiXSyytbfyP3mDz/W8
FxedGzeg7y4sxTjGm9CgjTNEZaWgteR3sWmS6FEBMpQDw5n1PjS4qlyMOzcMIxWxj11YsZvR3tQw
HjScucZOmdy+rbMvfzx8dV/DWj5DLEmcWeEW9mcOg8soRgKiijxMLzFkcMiIRtcn5zNTAOCrrDd0
2wlKaMuIj8Qx3/kj+cSnWOOWFkor9l9Eb0rIwGO/o/5hesrl4HRDRHcE3SYjantQHMHtFsPnFnn8
GUR8eqbYbCXKBHosXzTepSagPW8aqCXFdCDag+2XEkFFk5p1Oie9zddaKA4IgtNnQhVypSyfKFeo
jburLvo4+7gNYASua3d8whqbVsr+iKfes7DEJpGGrqzdWnUsge/yU/E/TTJR77HOoeIrVkrj2DGT
bzGBOx6i7EdcXnVdza+QdljWPyeu2q63pD57beTCFPT6/QCTpSS4yYfKzJM+ooBQPCrLBUQqL7mC
XPWzWhhkC5FqhFHAKvNEsbin20NT+nniamDg2cswbxH6pOXs2JpRS6pqARNpcbRCMJAk3vVuU2BN
G4lrsSCaSibIopnh9gcF2MGJH9/nIXcAguiwNOi9Rkz6G7Oj3adZANmEcxwx/nh6mwlhWvt997NX
9UhzJhTTKwOd1Nv+ktf1sj9382y5Y9StYIhKuzDTpJtrWhAh6nc3A7J/lVvv9Ngi2nal8dNm/emg
mo9epjlc9yX10blDJTKm0Ons4V8K6w+nOqvjH/9m+zxQMCnm/+X5LxQ5hr8ROC64XX1LicKRp4Y6
pUGwoZlWx+G+CZ3Sb9oGeAfo613EGwnCKKtF4asrppCKailkAVclNdQgaizrl7sEk1rtaL4TzId+
V35WeEx2Kuv5JmTA6un3VQbXSI+M84M02n3pFFgaaHvFy/GmpPDmU2hs78HCqEoczsvte2nw64bo
/DKS3geVbpAiGSoTmKM+5tHZZBDyRJNxKlnO2EBpcFXRpZkqQNtm5wtiK7vUeI5bXZ8T35CCY9nH
qAGJnb4Towx/Rj06F1WJbknne0jnlv8D/zKOvllf4SmbbJtWDS+J6joLMmkP/IU/NHexDomzxZhw
/Zqn0NXH5hhJm/wQZniI4/ZkVFr28GnFhiSFay5hZ4XHHY0Pxc+EVk1vb9uzMy6T7pRoaloMloeH
tcxeCiEvXDytkCGmjK0jcwDvcqRxb4V9rFuxrBbRVPYbs8p4MtUvDckIJZKpTh3aQnqYQRO7uWKl
hNw9zUpORSoqJJDNKsSqtb+x7EgWlntL6Gtvy1rlTNGAh+D3IbdQNH5twz71dv+wpWsqHijWKrNV
9zAcd/39GLH7N/aina3cbKtULJslUFWHCAWoAVig5Yq8qvzSn2R71ZgVd+nWLsYMOyHRw9OszjhA
UGhgDpFvCF4n9SqLLoyL1e0rtqfllq/egBF7jI4uTI4nBdeNaad6L/XU195zJrtj5wZi0iiWIpN4
wsGKOOQt+rgiSCMRW6KC5FLYF08Xsfek1QGs/R1ccSF0F90mJFArzn0PbemItaJQndrZqgTcWt1q
afCl4w6MVFWnqNrjIB/tUSBsdkOrvll2/pJhSBXK+Igm7cd01F/2ul6HiqOy9knOQlxAevKuggj1
i6qRuJdTcn6Xuytn6koMNa9J1iloybaE//Urqn/PJuWyX2/qZX9heCuD1ixVm7ZKVTg1S3lOad5h
1qllWgy+ImkWH3TNuGUVhW3npyV48d6yPbHGVcg2ma73899zWIaH4CSrRE7Y/vjw0w0CqcDfw/Mn
udXS2ecuIx8t4cpjpQVlNT5ggu5HN8WXihujEqDwDiwOZHOIpOwRcQvwiYWXSZPMntZBj5FOJa/g
g3RSg1MXbzVLZcGDnB5t8v3CAvL0t+j4S431Pkq9g/H+GMb59922aX59jzzQMZqX3oKC9zxOIwSF
LIqjN6arLAN4L0CyPVOkklr4ajdqE3sc7FDxZp29bWQHYDSkxXmjn2h28QzKyPxLlOGuJQQAZMUI
c8C+JR4fEbM610HOWMNnOw6XIiHkq0IkI5y+bf/x+lbvyUYXvxVk0nijtE4/cNI3JUt8fpamL6w1
shjCW+YsM74SW76hUDvN/M3FfxqghDufqYRkxEHmhkUyERXseHK0nPiMcGeruFksWpN7mLQ4IjlC
g0XHp5AcjvnoYIq6cP+LxcoKyp6CGuZK+ClFFI0KlZCG2Gi5kUcPc3BW5tpklLukW2uS461D2WL9
NKWEm+J7iHEkk0ET6ITSOBpDpr3JzvDI8xelteDrnmgLPQPR5mDFfCC7WX62yp5t+aKUPFNhTyFE
w4VUiIq2YX4fPSfz5qHhMykLw4m7U52PAdWlvIjhULqumK/REb6/+GKJgASWCkibowxdDsMkz+ph
X8yxudz3MoAURUkhQ2BE1R6TG4c4Pk4tfB/i9tKERkS3N6hNUxvfamUJNVsj7/OiwuGErA63tQg2
tn7B+TS5pEIXRVh/Sf+MTjByL8azFoxEeNbrxKPRNqyE6CENOEfZlDU9hV220H3gu/4x2QEpBO07
cITOwm9WZc0bALpKzBcsApgrXwKLfHjw63QX89Dg0hzqyKz0+EYN2IequuhvjDQDpW290U5JvwEE
vfiTf9X1s8lpB8dK969roxIxGK2uuYyOChsu7ih9BINARTyuxDdPQGOw+i2paLKdiFWHoNWTt/6g
zMW8BG5rHCctqTxTHr9/fTurW6qcLJHFqvnt7s6uf/aB0BbK7+X7r/pkuRJsWu/VJNdBxHLMQIwE
ImLWA1Rlor41khCNbsaWhDkEvtG4+wYOHjfwz83L1XUfvUGfUB1YQlBDpkFIJDQbWEsdcQiAPKj0
rmvO1dyEokZq5X9N7Jq+gtocBWMMsQoxx5YusA0gG5luwVGVw/mVb+BrE44OBW1nyRzunm6yV4Pi
4ByW72LOw9nOV9QBIsk7AHWQ713ohAW2kSWCIEMsPF406MiCOiXJECXKJOUEu4E7AqTCr1qZp6zr
7CZ9Z9s/K4TgRpE+Aplx+6n8Liny+wLq18gU8YTp8Es9w1PyMSF0AguJlFs7S5+6GPVZaacc4dLG
9w0OGSxrbZ3RrHdYHFFdZtkxtpOwj80lnWWOKwzGYVPGsry6PS4aajKPpi1kGsXW0M3g7zSBDzLS
1l5QbKql2ndmIbig/uRsW0Kas7GTI4RYiX3Yc69L3t3tdajfQLbIj45JqiBZ9mi5Rq1LxpnSptFY
aerUzqOb5Ifchhw1RoFfmcHccjzTZ8Kqdq86JW8Q+aeyzpQUezWE4ws56uEuAZbIgXqoNJMAsez2
hcbGbDGOmZnLgUa8U8yNPj9+LhJJFi546MeWgBoLR9A0scZcMlxDMTEKRKUbJdigWNFphJZCrtUz
YaDp33E1qaGbAUnDFuSCYVR08yudPI5aad9cLy2SwqCGkPOb9x4yX3qm9bnBaHVUzWl+vhLrHJGc
Qz10YMugbfkg2zyxX/4pv1QC9NMHTIG95SDVT86gNywnyihTSWyDUd1m+4QEKJq9fOtUPpu1M/x3
cN7VqkZ9NMtfxDKNGOzaW9bQ77MsjF9SUEKZD9IMA5ZanEtnEF0soxV+FbTsiPWEZdoBtjorqDfu
UxBOCSBuwuI+6jJk13nUCOlGGgZrpnhuwH+sqYjIKPBC/7BXk1YgKptkl4f4EOFXrP3m9K7RL0vv
TxITcCyTYToS6j4APa92Pr+fmUhwdRPe71pojYgkLfD4yrYvoeJcWVnT83VI1CqEUR9SNc4ClpR6
MuQADKtlTttU8LJ+BggUYMiXEJ/seEgU4D+tJBSnoDqLlcsCT261eZiyEIFaQipebKqdxaJsurBT
O10ujsfwW8DFpCaa98tf+NSt0bEUdbAI+JPpAvaxtnsafZNt9R/9R1hLESq49n7ANkdz5PFlhH2k
iT+IrVjLM0/kaRuO+fxUJCIgbNyzJ6Z3fTrOuWjVhIbTLouDb0d+4apMIOIHQTg7JrmtrUu5ecTa
phzABb3baVTS1GyhtNedYsfxtBOdERDE9Of8QdTYW78KXzcEMkqxFvgoJsYB9K6icWr+crUxoZ5L
GSChG2l/DZIFEYQ7iBnJXaJxQ95OjwakAOnfo5WA1PxuU/3AzRw8OUoQlytqWjs+ho5eFWnYA5Oc
zGXYRpSt0yD3VM1dLQT8FB414lamMOlk9DcLeBaxaivJ4mjN9F0r9LWxMRMloUNdbm3JgRDq0QBu
JBRwFZ+MnWcLnrrrOMyz1d2KcpNoWB2DUX6SN3qAmwS9lefq8kZeM+gwP+OKu3Rf3U6GeEeoOgDB
YHnFIx2fsZ5uuYU5/nDnIhWUqqufH/Iccrlj6/YcbygNtmzvPiQKOddEvuVZ91ie+ogx7wcqXuGo
mc+Xao6TwlpOGM3hTrIpwpqcTO3Fp20CMoCya3rwYWZXnpFEh8ig24I6SryAwIdSlSaVkyMaEVY9
M9AA978YDW+MR1Dv5BZ2qFDqt9x8vmN0EX4ZQyImw7scbAnpCMEw7HGjdDbhHHa04LuMeLt872Wb
xpxpqWPzu/NRg2Fj7OUSc+cuszL2CjPmImDalSfah8T3X9b/dEHBVPVELJTiKSaahqIEHePmeYwm
bdYy1V1AFETyF2v2kWy4PpKY2ikHKBdJX8Oqdtto6Hp1bmXct1VEyavyEzPLHcbwD+wPaaU37nWd
htoNCMiDi4zv5D90iuv2z8yIHnzkP3IetM1Bw4iLIfkXp+TfMrDCf0uiu2nA/M5kO1mPfbEvM6WN
NKiuEYJPOxuas746Skh6YrXgd4Py2RBrIzfDqOPOrlQBK5d2hjsNowxcNM7ajtk0eU7cTY1XOowa
iQRpj4kmALq1bWosDRq/5pnl26Q5JPyu/eGgMScqnVqopjn1/jkZ3x1wp2pW+xvLCheyR37S0CBh
r/9axsOcTdeLdHK4RK4CAR0KIs9cokJuO8Kn+/X7oc1Vz5h6OK3Sk12C+VQO1AqNOxt8ptmEw9TW
gRHDKVpjkcISjD3JMMKkiQbkrknVh8s1JHfwC6CRmFnAeMFsdmVWA+ITngH9WHj/z9NvolK8w4na
zAL3Mb58Mqtmf5tBbWN1kH385GF17M1SpCZDSNykYh18vWdunP+ZQxKNUFinkNcyIQh4S0k0GzXE
c3/sDAnTjle1X1l9aOA7j6qrllzCO8NViDrD+IzZjMuc9PLS9vbya0R4XBLuz4RqdVJbjaXn4C+h
N1+Xp3oMV2AEQXCE+1Lskt+QdRCTbt+lNuXdclRbfGVjKw55Akn2ihmtIGwNenkwOjaYXD5tBsoX
57vdV6FQBD+YrykqTMRnaRqhqJd3ESAjzDp2xzx9B781zEsJq6IILkwtM6BRkruiZ6LuD0fyPdn1
ohV8eI2OrG7x9ErtmmTNfv+0+S9P+sRxbp0CrTeHpk0RPc4r8L/ARl+8EjoDT423C6sx3HIPFxRV
t2nQl+jI459ucecjl1gU5FdKNgmBOPrVYmkU6vLHwB+/Yk3Az6BvkoW/gsoV8hteRtT9EuIHeGXC
jQwcAdkeIjzYWkFCam4vsRFGa2U+17BW6OXtTyO2XbWxc8+C4YY5gKKvs/tsgkx/wrBQdB6p6T3s
9ou7yOMnlDvqkF6RYCUy/zQWDtlDxj1PH2CLXGMIJhoNwaLUrCGpMC7CDps/aLQxwDnYNRHhcS05
1IFoBC/4+7hfde2QcNFht8x7pbxcCuhkpYEmY0nmzoIndJhRJoTfT9UTeArBTj9siY7yOonjSsHX
vyhaQYcS43bcdk61lz8uHw/hWQgC46htoliMirwDpo5wXmmr/7vwhz8y+uExNXxkfGOwXPCdFlM2
01I+ow5KeLcnWHC2OAwl+f+0KqC4ITFD2ZxJqrFFoxCxQtbISA5icYo32HsTAv3a/xIouM7FGiXq
iVaHGUofFc0R5MspI1clBYmdYcLRLwAxtrn/HKjKj/6lRzAszAYsZX2Cl72/Tb0+jreiRWw+5mWv
5wcNMpoQFqq4DpfE9savmF3rFsx1Ugxc/kyK0LLB6Wr2Bf5fEnx7Q0bSPDYNEJYcAUvE7Me+bbTN
Ou7udDrMpkxjlIF7mXxjncjHhmrPQpAQzPmYvgv/zvq0jF2+MwkkQI18Akk6+BNBIUZKPYOUaASz
8oln7nbSv2E4+SsB/nJzBWhMLLaLLj0C1RxHjs6oUvTEVeIooSfSlFm7+C8VNGZMfxWc49WTOdVI
EgvUo0ajiAssniy9LCKVnZpsXtPFd3nuak1lkVpPBG/LCR8Ojdza1cNQB/SldVVjad83rek9P27Y
CY+PK5kFnR//VHMTkKM4tQfk3Vh+QeAhdio7BFnl8N94K98Ktj9XBggy1JmFduDCuYQY73rOVVXb
qPyxQxhEiDDsiKk+2zSGRfH3aB9bQ5Z0IGlHcS5Qllp5GaBXOmo4b/w8pRJhu3RMYo0BGxbsk5wd
8Avy27G02vCtT/x6lxnxRU8B+4o0VrGI40yQzfXibI+DMs5siefElOK4nkDxJDa5+sEkL/oAnU6D
3LWLUgF+IHT8Jb0Mi8gUuFgAMv4UehlEF8SsvpBKsIdSpWBEIr5jGQi01Q5BbIHV11W4d1jBNvsw
Bn/dvcgGVEhfj1qFzRG3Hi+EaWmtQ8Bt9xSm0rU9C+C+VI2nINKAWx31pNw4dyo2TWDfEzCERWP2
JJrQTpMLNWy07FumMHFqj3AUdl1+W0M8ZmzzYWoc296JqW93rmOFVlpqRxP85P0HKyKIv18ezCt5
euKuLW5mC4KGJaDAXRhA93GkJ2deH2GDIfs63lyH8Iby5V+Fq5opR1D+ySFbjxE2lJVko4OEgjZF
O+HKnNR4yX8m/zyr4lXiKDOsv8cbPLUNbavGGhskil4rCMbH/KzawvyfOwciIS+5orJpwQLx2t1N
S86Oq3LmrrvwjH8YFZPF2EWtWLrBzum/Q10EGUZHjm6k59Fw6xtr/cg0ooluMKJrpmI4VJBFXJdr
mQLO8HzNFBchQesd8a5Udhvu/3ZiQOBticUvyFDZ0EUvTtKpIy7Yt04w4FPvrDKgLYvMVrYTttPp
J2ttR6EsCpGxvliG2TTaON4HE4c4A+5EEJWt3RFWOOonlmshPlok0Ve6azqrw4tD9kZsU4bY2HZ9
lmtx5cpwYp76YT2U+zeAO3rKc/s9JlJRKxBVR21w7wBOId9NibI8Mqhr7jNIybyWic7X1W+ur5pN
0SZCNtqnEjl+U7GFpX2/jpbeUydR739+K9NhmSeYLjrT665UK1YfhC/q0czzfZQkDGcG+xKp2ejL
KxmOt07xwTXwJtVG4ANSOnz/MO94WYZdQDjLZec7z9TuQntkwKobtAF4DAM7mFvMCfg7tnPdXhtL
Ai9bN56yAs+hO0UFBLzGYoCT3eIphqonj/x2Tzp8s4LOiB1Ql7zRbbdOm3NmVT8ODTW2ndv9h4rG
aI4kEhhZqgVLJ05+REDYcQWqOdoCSrjxO8+V11KV7/ch+KPDyOl970+bCtFCKQTxz9hb31lKForC
MDob37rPVeGvhtQqpSzfR3eVLxfimXUEEAMHyCn0FUL56N6qu0FCZl9JQVc3e4eZppdNjeYflfE6
pNuuWnNj4IIQPnN0bLNAyP54USnAhFpI63AdXv5cPMbtmrO1QSP50wd2xagZj0W+4glE7yFpVzbg
WUJn5ixszf2Hd+Bfyb5ggrH7ZwACpR8UbLV4GruPvUaXjzBd6dR6UQc+oXg/tAHPq07a7bEm4tCN
3PB9Q8Fboc5EF8/TW39E/+FxpIkqtiZvkxxlWck+w2B2GjtAjEjz3J7G0NJv226ggj38x49sk8MM
meD8y+pKEiV3+K4R3axlO/uTQdweVmWdVr45Pvf8fWrcvFov1VnfmNhxjU84n9l53yCPiwmuJJ8O
t5IEB0mjW5kYFMIprbIP8vqL0sdTCKs91T/nN6NU1iviz3fTtNID/Iw8HdP+V3ivxnH0bcRmcskq
nMpCjdChGyjqHTVNzhWVvrvlqNko/As5tyrNNhpz7Fu7c4+c2gkHjnK7S9vWep4T2Ij9lMBg0RJi
dOKYakH7Og8zT03JFAQf5xTsi7QRBnMJZeuc6xLpxQemkTo285RHZRYbkMnqDi3zA4E+bJROMhob
nMa5W2yuy1ZWAHxsAWcd3gpfFq3GF6PiAvxOln+EAYvnmLd59s/c3L1uVb1y2Ncwh2xplVrN/oUG
HV69rnDsSgDT3kPjGf4lRDCA0CUuGGd9jQBx4MC6ZSyB4RDAOk+4PxzD/8tUiKEHEeUqR1grl+J7
yOng2Dyc3QtoXwPSJWyXAA3Zl9uFmw3H2BljwVrW0Lv2re4PPKButOFcihnWyyZZRB9jLKAxfS5n
DFrPJTAWHM+/W26gFKr3MV6QTxQyqizsAmBESYOO3Ye8myk+/awWcabERnNGP02XHORKjsVqgPeg
UDAiV60JN9zmfxMmq3l1u0PmwwT2LNUsWwOJfQ8TTObTfQ4S+KNoF+ATZdO4AklV3QMPOROl9syN
DKhr/9N2Xz92GihLVDSRF+R4iysqfshPn+ccIRfCYUCnxLb7iVXR/I1kxH6Sjrp+wmvPXKyWYKTl
EtpwMQemtkwXSAHFwWzwo0LqezZcjDkJVBJ9a8gdOXNTEQTs7SowgoyNvMWVml/SkouBEKwhgmE/
V23TnQe0gUKMP6bRXORTCFS+pdYyptA/l4FeoKi5AfXO6JtW0XC5MQ5zZfjxyF+ah5BLDc6oDGMm
5+V7clNZSwe+aYdh9EXXyzsQBCDIfdFxbSwIU5cvlvY8wXcow9sE7feLWy73ljs6l1ikXLbFCOLU
FjbQHEZdw6r2LGzKJ6LwAGzH58McsSA62Y9RHiPSusDIIMpL5D+ZD2zqO1alh+opPDNR3/snKQfU
02oMzbQQ12liouLsYerTOImfBbXjR7fc0yH6ngzCUGg8fTf/PiH8bgVgyLxSaBRdYUFvW40OaQ58
RqnTq3SLjQ0jAphrC8gZuos+kXaKkorSJKlSRSkzJSjPz5EyypcxWjjYjjReA8QXDiUOIrxyWceI
tV79XsMLQmzU9A9gpwnMv/YS7BclJjGwp8qMRv83VdKKZp01bWBEnrC3U38Ij/QID+q+/mCeZmsS
vKMOVLeUqJTsXHsX9n32akSKrQWW6Ah0WwKgVFQxFcITPE0E9pOCglf9wN/exb9zySTJa28GqePy
YuqH9wEzq1v6jfiDX6tIXFzVT6mvvlCefyLjRNEMlEfPHxZBf56lfeZJSVbM7fW2MmcVflz3B0/B
p4jkxG4noH9DmPKMPCon/ElU4FsJQaP7P2PdevzZOx7NcpogVPxxTyngZEuExxXbe4bTJYaLEjR7
Pme6tgrCKRNv3imDXGRF4H0h5C8zS9M4quQE4lIaX+MYfJ4cyQciYTwpcYAR1tbKSdHqw+k9BNRd
XsDqmjCx5PON+83TJDLobpmtDGGA6q3tIzN7xgzdZsjSSrS1asOQGjJiT7/maBMmABPpaul4z1z3
3kuplX1pAX+JoTf8kuPVVu5D1woDpJLcmv9+kTvbBr2pAOBmXawBmPIDdrup1dGzuTAjy9gDep8W
GBZOPd+UhuGFxYv1RerIpCyqqSdNAnpTM8EhlARgYE0ZBy+p/bbJBIjVkpneq5UsRi9hJHwiTqEj
WbUVkbIMu5NJ3QVW1/UeFlGg1chvGDr0SvDI8H5PR6Jrsz4o+MJhsqnT7lAAN2GkdC6e7GD7q7qR
CorH/Idhg+1uJ9sqZSlro2p+MmzJNHCLukJTOGddmzGMSEKSHQB+dlhsWiM01XIWyN931HHwP6R4
U6SScaRhen9vuHOKnNWf1Rz3oVAQ8EeTvmwWVH91sITSY0s3R7gfNYbME26p0gu67hKpEiw+qFR7
goioFZt75vUj4/9fxzVYvkwA0KaXNeMYPSxTZG9bfrtj+rP8cpugwsZUiB2Pr70zJVm8xyDGocZl
BFytOYkdxUy8jkAeYNdaQNPjXTEc7ydjG5XJuQn/finox8C1SJYIt7UzqRq4zUyGiBmbB4KdM/3D
VkNFRg0d12eCeToArDRPZggZCClhufiQy2coriNJV/TstnKtgTES4zv7v4LuCA01HjRvPQTggeIC
Ay2Atjjdkn0ycazwXEcrK9/+HjawZXM7CKkwkUqFZ445wgsCCAKpm5k0GkUsrEA6tQeuEiukTvNJ
TNDxwraiM2w+7/jbLrXEOCY9IfAWAitKNPxFnIup/C2LjkYaWEFlZMosM3JV/yDzpFfHtLw/vny8
Ftxj9Rmumpk17lJ24IVVi2WKtDOfLciyoqs2Kk4m1XnZxkYC79dqLa1wBymieHn4dyB/+RI5lFXh
SPvuHzqXwGnpKsBzAqv2bKfbHs+BwCJTGlZsn7tz/bNiEy8qIS9luev2Ykg6R2ZyP8QJITYz0bCl
pOwYGcu2J2LE2lwtM9hQZ6L+g3DpkKEgjVP7BXgW2P9a/36R5tBJY6NurJgRY9VbcyPKBoKolPdi
iBSmlFfXzVMSMQJvo/XT+GtZ/c8g+dJYtDexOCC/jXDydVMxk8a++/R1hoiSmnbJhAPvPpPt5zdk
gVK2Efo806MM7/7+Cax6Br5t7vb9EIvtTwN/6zwd6iDStMPyyNgUSifJ9QledYqBMsMDhBPaX9Zy
XuQ+ypAAvc2FcJdarkgkUrpVrACVy8GqpQj/1j8fyl+dDKoYFojTtAlZLZuTTUSIGa2uzi180qx+
wVGfOlNWfE8E4ZjqVdL4tFLqGBgfgYSbUZ60UKsBE7xF8gN8BcU65dEyPrWViv4E55MlXXCNNME6
nZd0FQ+6ZxJLw+DWIz0xLZ4BW6e0b8yGg2lNZHp1eWZQ2QNwePzFm1Xw3NnujxpLBNBPFyaSznVW
Ku3ockLkT4tB1YqCoMw+p9o6m8E7+et9/TSHJ89hcJBJMWb6UOGZhPsLGD7w4FHYUS4DWdoYuGFU
+yOp1QIcMxSWWxZwIS7VsCyeQu7nxw/lncFCGv9HfQtAQN/hQ4PimLhB21BW6nOSfxvoVcf/Mipn
kONiEWP3mvGK/YXHDNt8sFcJ4fjYaW0RvtbkahGPQWyVGICbBOkTmlewbtMoscfMUtyH+wj3i02E
nMUd611q7xqOa5yCXN2qn4sVFWdCz4h3PAAHItyxgZ0o0xEslFmMiBPkeV8bqEXPiN/VfUHY2kGE
j5oNnW/GFKGAERiI1qLjNk9UQTBdoRHN0bYPnWHq15QkxMS1GQ3L4CFQMAEqwVM75rqxGf5LlEAZ
ATbonPkztYVte6CAb33pf8u+VEKFxWy0PoAFrZDUqILVyg7nfgEt83K7kmy0EJ2HhMWEYamJtxKZ
k9gkNSkv9OF1HatGvp+HYvG7MF7ZvolsGIopmk/k9lDkgHaYTUrp1VtbKTxnTW4IACt6Gc+qyqcS
2NPKm7CQ0WpoqLeziArlZ7hhmezoVLxsBusQk6mrs5DLKWs1lh28WIIXxC7Qs+YtUuB+JWdBMCIO
7A6IO6IgvY1OCHlH7vNEEBi/sPAAfNjrk4VtRRVR3oX4UeUYsHmaHsWoKYUI0nYi9bFkvgPl9xnl
F+r/70F9TCtLO4vFMLXA91eMawBCHc1EdIZVBuZUpj563iBdcjnZzcoIfsCbtFFn6QeShN0po9ZI
6qTOVAjhFBoD7+Y3BzwH+mIpH6/gHaAE7BGbIhJRhm1NaUD9CabIzmbnM02k+BNwej18Xeif3ZZ/
48ZTiD+gu7CVfn1VWyUfs/wu8bDdR6ElKyNMMypdiuSnU7cQ+D7Kon4+7fu0XHfw9nY0qT/ia1Hi
zEftvbHK7ApypDFePbdd1zNnsZdfR3MsFdwf/PN3y7F8O9r60krBvdMLDbjmERuygzJ3BH1tDfj9
OY7peLNkxCeRcy4E+Jck5VB8uJ/1eFjWFI+I+vTvaVgmkVMsPl/ztvp1nd8gowCRn/mwJpm/Cffw
vC4yErjAQl1lYTv2GORthDpyBPdN3Git7xsTvjEzKROmMggmcUNqYvrcWFwYJxHyGR0woYPlY9Vt
0ZHs5p6dhBOA1vrCKmB8/b9ejtylCENPShz2J+kuB4/fUnUYkOt7K9b6kpHJ/G1eL7Htn05xj482
TjjmEqlq51RjfjeOccXMpBjG0jZpH0pMAMA4WUrq+40MFBprawpUkHIlZJTaNgrG1Uk5ECn/KPme
J0o4ksXpFmm7Azw4emKXf5TaE1eMrTphn6N1G4VjYo8hQW4E5gyp3hHLuLSaa6HX/3+h+pj6lSPk
znnSnc4ew6uzxY48TDV9sD1d7cfLi4vwn0+S5dZ3RLsjSjIi99CWCWFsf2w7XLcDV6H+K9qEvzR3
Mh+zxqjltOu4w5l8ycqPh9Cs+/WzwNnZSKzaAHInLdzNWvT1+P5ncb9FwtUON/+k5blwouLrQDL7
0j0siaRVsy+vbKzd6sh1oUbdyZoJ2DJ/GLA6D6FwtEIbO3IsdCvZQGi+bRbQeSNNarclhO7ZmnpI
PdYpuUAZ3QsmnB//MJEuf2BYnuaRMkbrQ5lWG3pADMPZWsqOyas9xdwxzW3KOmHeHjvIcBpjc+2v
seLBnTsKI68xVR9Cj3JHX5fbnqz42vasOHc4fAkX+H3OuOvT7JyzihGGYtLf+njpGni35BkmLU/I
dHPm/+DFAHKLSh123cxxHVilfRWed63cDFq9OKXvDHSDG3e6HyLoZVs+PDf+zcoWel9YyT7QnyfF
4ZOK8mBt41/7pwW6PVOu+QhmYW1lPtBpKquJAXgxVG8NM4mps1K+08zBKnKEQ3wlMlrWak0HuGKv
SmWZI27m9gAzrXYnIDETYPhYEeYtX6y0KFHlwxhsP+OFcCVi/z4UKPA0IQZOXllW01ak359XQ/cP
xLfhKzzB3emg4AWAb8e4pPLBUx0XS0JBGXVPmr8dywI7Clw/aospnmIa+hOpgDz/e10ZJna1WIbC
f2wT3iwsMgYFx16PW6zuPLXnD9ZPy/+xYSNI5Oo60ccmSLFBTbOYIiG29bacuy13lMedNM63d7Zn
wjQVIkfCkAyQjrWv0RlbHGPueig/9Q4MWw5BsMDx0FMcw4pNvYTl5wZXfQVTXG63t/M1El79e6C2
DC9jJ3M+0f0uPTlqyYjcn2SJdK5p5Fk+XJuHp1wv+cuqhqvllH+sb1cqVoLnuvUwMOtF7rXYur7H
OL/tiaTmSIjl+ehm9Q7pSCTmgIGoyFf9rnBJ9WRAvmezq25UsW6TjnPQ2MZO/1rXj95FlvJDICP1
wDdNOJau5UWxmJhAkWjs6hRH6LKz3FJh0WNOevhIkLyyEFcr5ThCjznY2NTOD9VxZQy7MzbdFyut
pGZZA+WsWTcMfV+lud4Al/1oxhGkeXOu3sEcYz6jzkQfqCXhp4WVXfFoCx2I6gOxJdoeRauLpevK
z7jAmjQDzNR79Bf5ffhna+othGvq3LwmDlbBE8GCFieDv5mndSRItY+oVnp1/Yau14skpCz9LNNY
E9n5d1wkC8FsWzSzw7ta5IoqUalD2M1qvJVhHuhwrSeI1hsq/F7WYBWY9jsBvKV6u93dpXoXliPX
hfUjeFYLxYJdCjTp4yGFaXKJSRMoYDnpnU1j5U1gkWY9FaiMf1JzEcZtUW7x6VySHz9eAMfPJOT8
MAibgkBzNetKY8wkgisGqJTRL4sbRnIMgBK+Y9mYunb0xKaGk/IpyoW0+d5pXzmzLLhV+9fM4Pum
SJyl+fs29/x2ODghZgkIQKBnpItYNPlCDimOUXydsFN23uK8TnYgQ2fp9GXL0v74HeCALt/oa2Dj
AEFq9w110WQQ3CbiblCdgMkkEyGxoLyxMFoNpU4e+80anBErKPXnthrF9XMF2zUsqJrC08/SnH09
b8Vp7fn2bC3wyxf9dth0x0ZelsWORx9cAA2T4xCjyv0Ga5OY/tNdqkrZODnVH4tqHUjyJzOqmBlM
6ZucFnEGnIKZ0QSa4P8zphZebttL6d+3ySQcEGMDKyHBfcrL1FlSskgJKJtuwvusZlEevRpa0zbX
9II10P1KrPUTQoG+6pQuG9hOqIn1hnGyVPS79PE0KN/nOHI5Ki8ui42abP9R1A952fFUx6htgLlg
tUALtR2YTBHVnYeSaBHCIf9HD2NKdJHcPhKwSHgYLiij59YbtG4orj/EsSoVbq6JrcHtiwn+OP/H
Yri6ZRa/hj3aoSlK630K3GpKj160F7njVNMnp0j+Qql/fpImrCvU9ooUU1G+WpQo69w3m5Q2xrpw
cvymE+KEFsXdqDcxCknBUy8u4uusXOXytS24nJVAh73k8eiIrMhf0EikK/os0HcoDBGVJto9WoHP
9unXrDMK1kuRI40babfkioX9PTi2YDQSbzWfN9qorJ4/Gz84J7RcdOuxV1icrJ/NutVrCrTK3kQa
a1Q/w+VOEE98x2IvIsr6px4TsGwptSDoI6BSC+5jWk1xwNygwwa1/ohWIwyPM5T1ih92GYyGhxD8
ZcRHi1S1Mkz8DlydY7N1xf755SVXgmOL9tcanYbsu56X3Fput5Wh5OWXYpLsHNlhSQu5jznoHbya
0lgoNEzLP7Gh/rkI4/WMXDlH7KW9CMz2XY2WimgLR0b24EqQETjsPlHfrcSU7CQC8J5WGCxWwUP+
jAjaTFIdn4VIu+xC0UQUkArj8Q6rjvULyJ3uw+unnO0PzSDBCS4q3NhUVdkV6OOkgMMfIzabnWNj
ZadP5PujMUcceKk+vRBB+aDspps1fdLGJfEyp5wh4BdFw7/YdmDqV1s5+lKRzuUFcpejsCDSX2u/
BdXeDemFjTVuRY3yNlYTPFojWwCUhAJqMnNrdBLpPDk+SdLlWPqZxMcZL/cvIoLZyFbJaAosSPDq
MctsEpq2JIG3IhW91PQjrBTz90cZT/ExmPquk7WUsg/lM6mR6tBMYOVq/gDRYmI/nbnX2jML5B5d
KSWjW74AlcJt96vHxm+O17ajMTKZhGw76h6meGk67lUuM6q48OGg4ALRZQ7B6o/u2xupUdhnXcfU
yDVCfdagXRssDMiG/kHm9q3wwN5GsfLay56TQpHqyXThNGwJT3Zz7/sk0ywbqVW++iIkhkRyIH+3
w8k2JjEAP+tYHKh5AhpWIhLwxGOvc42nnk100GP3drkpCbIWEKz1HVrm0ZITNfkl25bXsf7TxciL
qNiTqj7TnPZJhVCeRn75FvecJt8TambTwr3sDQSMk4ScpommAixMCllSDApHhnZR4gmTDgO6vuyS
kDvOinH3p2SONmvFnGe4pzSa4bPlQLeN4T1nveNX63AJtu7djwxpWssNjG6e84Hnz40Y6LLBKOzZ
ko1izgJnxs+TAtbxqw1CtJWCiREKTLw/TSkb+Rs19i18QBeJXIun81hhhSCXytMLuRld2AF3Yyqj
bVpIq5SRlbhP/HyW2hXE7VnxlQudR9crhj96rPoYpNVcCPS3A5aqJxsr5f8L4Vg8TwKD4vC8Kv+i
khZbiXR4vt/HZkiqiaJIDUrZKYpkElUAp6TzmEFsw2a+mNXCJ3tckF/AV8hcrwo8zpNdqAv+ViYa
M1btRFL6kf9PzM93zaotZkuKz17NThA4ss33SX9ZqNW4bE+LewvQpWrA62wK4qSdau8ssf4c7rn4
FygLEDaWxw01i1lnS2QBPDaxKBnL6JAHjhYkLBFNfiPFKzza8VQsyRyHdeplXvcYpU4mvxiSuBAA
ddjH5KhHO/YgtOjkGf5ITYSahShwQdg2Frb6nIg2a9CloXiyeTj0NmIygmLY8IDfeRc15hY6zV6h
zghcEiMbHyqRswiMMmY7mGJ9eQbwZ1K3HdS3V7g9E/lsyBgNgZsXr9SrQO3VhqKmeDvaszkmalSB
YngIatSNc8PjjK+rQU65J7Bbf64VC9j4wGP9KVMyVRnFV0wKlX+dUxLyHcawFYXTjYgNVA/hrwKV
K1Pz02IwPCiJaA7ow09xl4l0vElRmOv+1nGKyyomVjhrj24tLbkPPZDY2kTVra7w2HkrtLDN9Vhs
hXf2TZ/qAzGHGIDOHQS25dMza/yB1CYSZieHPsZ6yq4gM5Y+h2RBqlD8pf07J2Z/tPSTHI8ekitx
IyDEPt7VNa+fc7lbgTSavSMBjwKpdoeCJIyLEdnUxW5Ha6mRfRKActvs+AbYycc208J9OjQ6F/4W
91hReLzaoYw90CWth7YpTJr0uJ34FleZ0sS+FI7TErZDv+tk1Gg5Mmu41bguy34l2iBfTOmL2n2F
psR/LnWXPo2l3Rz6jgaRd5PUTBHwz+6KYf8yB8HehlrwWrMlqNRl8kUX83QL+zG1L8lWxfGG8FbL
zckS4oiJMPDFbtTcFWl1+ASBeBAbZE/ISxaw+ScxwFsF6puviM1xjjZaN+BmlpzoUZ6AgX0tOurt
9QqmOoPp0hnD1Vu0YZZ2+jnXWDpis+rDl3sFnGz/b6E/ysU7AjyujMY8vjQVAgpXd1hBDpaH2ZOO
BoztQUb2GRinq1I7cNy0LM/49SLm3aTpuETknFgI08+47wGEvaGFh6Cnozg/4UvR2tTABHScWgRl
V/rk810HZqPGcHk7DooWV65zr7h8MWkR1opBBWIJzmT8/NUE0D8duQhoOAC0so8AbXoKpzCkOfFp
FPa+l6mCXNGOJDcJIqAGurIHELHm5X0dgVuS8tPGjOoO4V+WT37kBaIsLdEBZ+77+X5jviNOKmIi
BThzBps618BNJMzN2dF1jMWGVjlZQpxPRz9Wd6KG/pLlRPjZVszhpKz2Px8NRrfukrSz+KXKezyM
62kDnWPwwWFSFfZd5Sj4NpdNNr44VLaLVzxWK9eTwmdJifiWPZfZ99y1be2cEZ7tIV1Pife2bd8+
YL7gi5dMGk1O6JZx8+vYbIcLDCkX/P7YUObIrABJ4iaxU8UDERVdVtb/0DUC0hZ+oqLRTTWCFnZj
8f/IRvmjF/Ol+BNucJVloaK7yikVrZEFGzSjreLwqWil2AphYi1b5ia/ubfqtF1imkXs1zvHHlHa
5scxoHwgimsj0JgSlxn5vtep3VX0S+2DVTJTzYc98Gwk42eMtQm3r1HybECquzAkoG5pv6+L+9G8
TCB6as6PwdvPiCmEmDTNwzsVTv+pbF669GP/HCvFpZ7Vc1OevxVSa6mY5wsvjX7zC1dv/xGPrQfc
gTMLzhCulHmHPR/pJutWJEfvlTJYpSChra6LNLaDBs1I4a2ndTUaAnGgSQ14qFUY7TrUsJyxRBzX
b1qsW3gh1u/nRwRgzGGJ8xR4e5hhb2Fy/bDISTTjSwHt8r/Q36LIDvyHkQtm8YK5Pfsk0bvhqtq2
yrDaDHLpPYbN78GhdWgG0cS5QG5VoXDX0bqWyYwnL1V5GBWxvxDMdPLUw1yaXVnBhbXXNVwexei1
Qb7pCn8nIwQJXXyqjDonoTI55BsTDLOpnclxLR0k4jTZm3pUEFIISiVGdQ7Mn1qPbkewz9QydCPm
86lgkEbqqyOXoCRL9vBHYjCZ+28C3thNDsdkSOuU9MLKnZY7mpBMgDvAllUijVf16UXO/hMo4EXH
Re7Ne9tUP2227z9Xc8gMZQaUPpe75wkJrRj1T7JFYR7SaPHsO7IGh/b9kguiHikQ2ZEjFLscV+GW
2A/98fGlCrr0ZUj30WAU/u6NVruC77P53p4+u427TGyp/6gmyhoimC5e9qhUb6STSHQw+kQNbTY+
jnugFNFpBbhfXGsyxwlBfLzzokkiej7GDbAwwW0x5AWqk77RUSyDpfXhivoSIpmiw7+dNVZPdA60
V9Cbd9sVjzkWiMgjI+57Fq3YjlndspW9P9fPsEGpKlbcBDZcTwo5oJKVzMPWMQgmmNuDFvYhVcVD
zZ2lGYluRf5m4MhyBvKrwUOHbwbgJz2l4CtjoaINnRaL2R2TLpwExXdqWyMxUWo5rSUi1ZSPwyF1
Cpu2zBo6G9Cl67AJOs72GTxHgf/W9bZHcMmnpvBD6vWhjzjcYsSpSNMvL1t3EXuwNlkLD7u9dOFQ
b0KDU7TQy0B5yNp8duiP77eBSAfgiPt3QMpsqxMtIXB+xO71pbH/KVP+nXNkoUK1X99khqgKhJZN
BIexAoz4dXh8OQfkYZmBDx6VdVZnrXThLeUGctwdwajSze3kqQUcYXG2cABuFgQ9lBfb20w8xZ5W
/8x5JEtYKzVRmbrVEr9jygCJo140DTb+e+soThycLIKR/GFZdHPVhhvS2ww3CmBQFY5iCz8CZ915
arKvndb6Tgrre9hvJirRoATX8f23F4YaplaHfhAmJmVvDz2A+Iq5eo1j8Gm7/Rn0KAaqJ0LXIqjf
QfAhTqQ3qVztMpliZie1aeO9n9wdNT+Xyrw9oZFLA86ER46bz73pI4XnqMuZR8aC9PegHBQC6aS3
iFzitEGVRERbg6QxPxmETxDpndF32wemKymd4LBS9YzcBo99jRAfvQnkRWBEkaNUDxwadB7xf+a4
ITrHkZJvql+UBgArec3YUoe97g1aL6GnHezdIuO9U0liUB1nJLIYtfem8I1/T1jSgajrqHBh3TXl
4iFfTEIRCLpYdVTYlHFGmc2IVHO5vi6u3FPEhHZZTTqruGJjnyuqLLsr01dXt9JDEMgJtahPTWEl
6v0f5vj3B707j+rElBZCzae7TumbIF0BJ1NXNlDa/OL3EwLuLbiTECU7+fNxz6FASZb479wtfstA
TvcyW8q4tVSKMtwGRgk/FHFNFFi5hxTt8/SJ3EflmLc81xufr8maJXzk3jxsf9ZFiLg5XfnY8S3F
GmGF/oJiuKLweOvuULcTdXRW7zcm8mNJfRLR+mZsBQhKQOUT5z4uVT67MPJ6XsWk1qous1ym0PSm
hWQe5IFai2ODNqiy0v8tCR3I0LjRADstYSScqGWR3ObDqsstcWntoZ8IYniFADhvPVZURgBON1xY
ORJk18BGlwIPxPBspYS9xIwK9hI6MSRCxo8IhP910IDZ2XRb13pafZqQTdhKEyEYsJ01CbLiT3ES
Tf+/Q+kSxX1G1WuPKzDJhzRECnFhLYKQOEjfz4NMYaqhsPcnDttMFswL9Rwm055PZGMg3JK5ZeOB
T2C2ht2L0Cv9x2CHcM8Lzki/zJTu5/rMS+aJUiSkENvTvNbRnbWmmNXzAL9sjdiq1XI4cKJna69U
X1vNgdXewlfma34GsNP2VE1Ez8T6wg8hYtiGID1sroKqHACqEEpcdjxHj7aAQwar9qu+m3vwAv2H
92lTF40w44KPi+dV50KcjxIOoUaNR/l3Qk/Ro+kdgAoVU5WwvnTtY9TyM/7Yuab/r4okePkfknKe
7TIos3OYqbcm1lCJKSSse8gAWSqCphkJq+PB5l5GxA8kbs6LS4ckJkpGVH4AzE6GUF4Ik5vZa3pA
kLeL+nPc4WukQbMSwVBao6E5tRT+F0/WmEkPivAKHkCMv2h0pu52Oz2Ye77+8yaFgE2F3/1ikFK9
RInvj6ajMK3zKKNbsv+9GwV8FhJD6RqUpCPJdrSHkbMXJ8pZL2qtYBENeB3GJ9rzyv2UTft39GyF
SSidph6dlgCYi6rdY5kF7/BeefQKGnZBc+T6p7RNSf7CgGofpHy9SxYVlB+AvPSUvHdvjMyn9zAA
JKDauzLXB0fYRIGNO2TD/2vMgzQvK9eOpmqFqLuHEGcXXs6yGMI7owOcSV8NhuoTvkd5lbvi4Vze
NOM/GN5B+S3KUxFScl49lbFRdvqAk+sD6VLXiNzmWCW4Y5gS9Eh1utKJjh+NdehkVkGWSqjz2T5v
TLB0qNwDoy2OPhevgUnNQmbG0bCO9nDrkNWnb53lMUBdVkRMnHs8GRgWZ93EI/sQLSQg0cYQdBl9
V1uMMvSPjsHXvLSvUMRfZiWRSB0EkZLt/hWPUeD1SkjdIXqDdehHJPK4jOde0zigLScQAM755WNr
/JJfbGiDl84rgFiamdOJ2Qe+FwtiYRfkTx3z3OYt/TzrXKjBYERaBSKkvlV+N73gPdYZWsPHlwQ2
iyFRATJ7RpFlzrE0GwJ/tV6LsH3THvxRtaRI1ahfD+TAs11T+hflWC4gAijr+Y4h2Kk4Y5wAaLHS
0FC5c/MZFa0gxF1vVVtELZlfUEEuJQQnEuyyXEK4/wp7d3qTUB0pE72lDtzU/cIocR4AHAtAuYUx
8N1TuDUr7iXFdFKSgZzCiNNBEEnWhA8upVJohRuRVFOjNN/oZ90XM7ZoqyC1d4moykPlONLYVsgK
6G6wgctWsu2Jh60A6e8lY/qRwSwb0No/aUhPjhRZRPkBzI7h4cqzCgEZK0Z91VJL6vOo1duv61hy
vkOjFxxWOzVvJSatrEz46blQSeT7pv/S14gvWzTW7u3wgVWOVyqkEdpveqTfaQrZLG57PUpZKJb7
GYtdzTP4Q00mvn9IPBrmrDLNHGz+9pvxYAE4rr2FmUpmZMltuOSydQHPjd5dfhy/z+3HrZcBO7yS
g/50BPKiES6a4zggWsO4kRQS4IDhyJ2c1Ja6uZwxIzWRWJYc9IplvD0nLK6QnLCqNyrqTzWq2Nhk
un8NNC8NtqDefmkzUqmuPxfkxoFNRLYF5CXWpEUVPjgBDQfFbBF9uJ7dvSx8g8GVU8wKdt28/0E6
4DBnRbnb6H4kmdzlMydhMPnGlSW9+JKwZ7XvhfNWm2WRK9OK2fYV19TJ+B48JQGwQKHAqYpiiH+n
b4gry1bOmGNkt/nKc0jCzB/XW5A86k+HNXdziVnmFksAUVa6kL1Ke3wBTK7L3dRCW4bXZCJ5j0Z8
uqprOlOqNnwm2GUrsHi4PS8/bOP5pi4+jN6I9qO5YaATXe80d03SATP0QNvDf/+EYyjxwNCqR7K4
fGUMKNru5I/imPuV7dKjLbyPpSqPUb9U5ZeoPhM6MmPbwQTsiFMZBzwTuypwPFoH9yIz+a4R2gYH
3gfuNlK17ndtkn126pS+a0PxwrfmaMUaHoXoyZ5BM01I2ZX2k1FtmcDlhLCswjoqnngW3xVK3i7t
5WelLnVzihQPYcSQUkOqz4vRXvwN40AbUJisAnoTFdZUiiJNxc+YHEEdpR6v3YoJUvWM+7UY20Wm
s8qicTHQRPPSUdmJQMopnhSSyi83zhHPv4dZsXbys0bswvyQ/azenT2VZt1K5mkh/MKnAtoy3WNd
23/aZwZo+bTW5Av2CbSc1U3vSUglLcEBXkRSZmoYq8fYhcMT6DeRvFYdKNCA45m642mFKd1dWDCm
5WAJ9LUTpMoRoB+IJa1tFMlj5yx5dQCTH4Pv4RfahIwpVkSJe40VSmjnXBJxJVQRlJ5URsT1uBEd
33CCHxga0gMl6f1nBnBJU9dnaEFK44ma07/lKjw3+Yb5XLZq4t4hDT6F8xcPvEZiiLFP4oaZG6O8
Pe/tgE4A8zogI+r1mzjNQncJ69u7wJN/00VI3iH1xhBAOk7O1AS2VFce2pWoh2Ebxglyy5aAdtfO
Svh3bl9ufYmFwQss1Qh8aULdvg3X4nA2nWrdgrdYIc0izm09rsj1kBbGMHWjkbc7QWaGGc91fXUF
r95lwBSDV6wg58v0lB1OVg2iF0bmo7kiveEPfRZ0uAbp8k5CtSctRRN6cYBLhCS4GWqPHlpI1TGj
Y9kus2icnQsDjG40/rUR3ciQuV+jjzUIXuFPVblYidlTfeOlxKC7Eue0HX+Uj4jmvxM4Jyr9CWyK
Zqpf8iY0xFCMgElM8gMSBjm6mD9W2/UhqFLT6/kQk5gchZNY84e5QpRhgHlA0i5NKyWxQPnJmwdy
HcHrVw7aoK7BzfCEKz+C5EXRxeAVj9CDLqmieaDl47tg1K7BSYawt5lBOnrEGgCx5u8TTgQqW86k
0LNE4fbBp5QAkSZTZBnUMMuh9K0cmaXOug5ASuAsVASpCgq2jrCu1HuoWSwyXbNtIZwZqbI1pcTk
Jxrj6MeMYtJ/xnfZo4NEV0jDl42LCfhxzYpZF/QzsG7iyZISVKkMY9yqlnysU1xbYbEZUM9fEenG
84SSeKafLrBFqofASuDoCQxKssHjHJ/LvcijhK7D1zS11MNgqXpsoX2z3DlTsQcsLA0y1xaF3rDw
tthodnMlh9PcXAEsDWahEAxPPnMiuRddyXb3eQDzqFSVC3O859n6MUwsjpPehFKLcppnAt5CV1lF
wys4aPg9r/JdrgKZodval1JJQkfrHFU1A336FaP41WfgL6XL5JoOuJ50qNQjpvTVL610MjfZtqzz
2nM8ZGlDyFNTrskDTPpyipgIF/txS0zy1o5g1Gyb01qEzaKZXWtO+dIfAqnHtlKjrvKMNElen1Bu
LiKa9JcyJ5eTkwXk8afO4P/fY14h/7VpRube66mmcF4BVU+b/RLY7brBFw6ci+LyGRG0EKPddH0e
u2etWCQWKJhQCJrS7KAITm040sjHtFQJ208J0iTZOPtKFkpQXIb7Z8RM93BaF3iC42jhOpML5KFH
31BdS69iMiOpgl57sti2ons8tA8WnztZtZnbUtAxIMyj3TFqnwlobJs5IMJ0XdCBL85DJ7P4GoPx
eUINpT8xbEF5hvkFxfgwMO/dupUerWiFq1/ros6TLHrzhIUKUuzB1p5fNFo5OwwIrozHCdDKLhTe
UVSU7G19AMY3u4OgQhGeCTU7nmemjHrXH4nlPK5KZ3551ir5O5xXaCKVwMC2OUA4TwPfNwfhCInk
lE+pgJ0ajzidijhSwHIEgNF2+3QgpfiuBIiaXTNjKk4qL75+I8NZwvgW+ZetxOsmLQ56hes/98V1
AOr8SPeJ+oCjJhPcPP2g5jAnrVxH93YmUSSM6cAyXqmJ94RZE/qYmtlpz/RrwHGvtnDL8PPl+zBi
5i4woHr/DcLibrUbiJ8ijFsDlsJznybLT1J26Z0coTy82YM5m1h5daCOuVTDBv9oQ7Si3hwY4aPv
/df8yxzsdtbTloFHNu9QuX1mlEB8V2LQhvJ0ZqgJXSLNjeZQiAuj1BLWlmlbb9TvljScjJs/HKdc
+nkZyVuyT8PAF3YjLh8qW6kjYFTvYCysD/HQuAxAaORmCwwmsn2/114xGjnh3Fcmam6R4zPIQNFe
IdmARQY4vI6ASgzD72v7deTXxEqp82NOKtFjylCN4rcKzrBKuVJ3fl3VycCLeAZ0avRxuM85l9IV
/UVjQKsS7oiTY5E2JYx/rsluClOW7h2i9a79FTiTAekrJG70gKYp68VazqAFh1YFGd6tWrECg/hY
41ifu1ioX236FcEVhaRQuGezzvL5RgqQ19taMr9b2bVDQ9O8/iTEVo0uKz/rmqnjGVH4X/lc/7r0
96bNy9yog11AyXZXeaRni+NX9WYN0YuPs+6uptFsdcIYCgKijxMvpjS8cuE0HWCkzAbK4Rs4OdVY
d7UNg8mYAEtDh2tg2liwfJGTU+QAGebTBcc/W25+HFekddsPAGRHEGXaPfVE+D+4ibewLTcAv4w3
6RpFkd/vtaN1kwX1DUR5IjjxKCoX75Ef8zBc6C0FoBX1Ejt30SaBvhmsqiEy1hy2roHw7RqccmPT
bftcVvV3yJFPvjRPYwp0V9buW4KgoAjhmjmLvyE9EtX3Z8Nqr+KQMZgE7bKkqqJxIU5hb5sXzt4k
a+TZCb15B3C4W24n4JJRRQo7qyvNeJQJV8msqq0A66CFBngVh79mNe36ssE5JgyjLU1hZyTTflY/
nABNWQsaTN+5o04hGQ9BGDzXwROQYApYL1ohZkEGs6NbMwQtsVGtFe75BXVCUF1ZlU7q3vfFzD+S
Tbq8zgyuGUpUyeBgztY0LD0znFq+V01w9WiF1dvlne6l56+bgZBTsaPL3jegG8Q+upa+DhjqFxR9
2s/s5cHyUCDij4JXNHD85ZcFANVsE5NEaWcUw7rty0H51pRz9yNlVpQatTd5QR+N6bKJtiW9tIg3
NqHVgcgeDsm/zJH9ltxhBkfSjYsU7sf871IovkAMwreFET8gaR2DrMRkqOmJdhoXLbx25yWOMjeD
RSxhAdF0Da5N7coluLtOIkaQzpqlNKWdmxoAVhvQGz0F/dNkgQkzEkbFFePCjqmG0+tsZ6uM0BXM
1s54pag3klBp88sOXgld8RZvmosgxjYaF4odWZWpFcdLh9wBc6yk2PHAQCDcT0OVoMbxnIlhaMXC
TjEPM3khdOKK+//2NpYmT1ky1EDtdSTxVnQdoDN2fQ60rsWh2vULuuvD00Ompne3xu9ZE+/mMEWJ
nq3StkiFXz6vcahZj4PfWGjDfFB/niN1+YrnpgkRDdPvOnlmS1n51WYLLVuC5cgFXNIkIC86Uwqr
elcvFfA6Cjm3eWZvHZ9WFm79FxuaHgx1WDqWFFSoxY6UbRYt5A8a8MhCdbz3h+3rBS69YOWaskeI
tf09VNjXOMN/dMbsxQRlSQh8FpmZZJD3lwvwBTozEbG9zDLRuNNOIah4g/tlL6N2IaT0wmeQ1hA4
3gdHxLTP6D0qyQxkIMybC6rpTHfJF59gDSytfLPECtWsGn6miOrRyrKR/62VkWTth/wh9PS52aB9
GSOnWH/7+WlNzWiMJghYDMXLWs0kAUSpc0kWUuJwuvBE66vQsL/9wWfDItwJ/bIP5dpYW/4JYQyM
Hr3/XcO/qnATl6p68WiU79m4kC7Kvay2efwIubcHZzT0iBtP+EDhUs2+hVnCN3lGdzgrPvQtmDl0
en5TdCmJvsgdKoDy8h2JLkP8sa/tGJltrYUb2a6Hzmm5LjUFQliuZHA4wGUx6horMoJYSMsBioZU
3PMTwb6J9eF8tIp3v/8qDWnbANOjFSnoDrjn0tx/7TJIpe1yBPA+scVQJEkcLieLFCNwlYHdMlXQ
hZTLkFhIME82LNBGLaowlzjW2aR2T3YiQhQYCGyUOGISrY5wpVzzfRQMr7wKSwZpRIIOpyLnzQOW
P6XvqJhMZFEsR9e7fZzoJAeA6sAjC7U/2NPgYXuCmRWbDsU+JMyKkt6oGicnt/fNizl9ntFMQA++
FtlY+I+gGZfTjMbR0WpFfr5kNbUiMaiPh8lnqM00S+VcSY4bqPPyVI+eZyP2Xhm72Z4edInCkGgx
pRGgAZsMl/KB8OMEG/tutbwj0gXqHVJ4oOwlGDdTTqWuOJ4KnOnzdldFHqmcGGEBkCD8UC4tJEpV
Eie/1F7rKMSbCktsveLK/V2KTbLe0rZGJywe+hp58Odis/j5IeWKnA7Cx1wu8cwlONlrZxzzB60d
kzSPbkSmBunFLwpQJuWsZNivDibMOCE/z8NcmJmpwRImw3RUANezlPhDS38zRlxu6lRIJ3lR0Ndi
8hLxs/UaWDj+o/vmwmV63eEDcSH2mWMQVb8Y07EcTZ6lgoGuWSwkLugFstpwefuYkgyR/RmNfdxN
GeY3zcZ+w9zBLDBTHWQK0/4ZeAC4saeg12hjw/WS1LRz/6SqX8b74qMAhUt1njl9sBNRoEleGcEB
Xv3UJuE8xlNluh4dp4X9SBGw1bK5/xVortCsVd6m/PKg/tg09/KLc9e1A5EoAeP6zIWxKj4Q1Rer
F3BkPqPnEmsAW8oKnhfihbHuhXmcM4hVkVVWZ8+c6eGaZSX0WhscV5NNn8sNr1o0kSfR0lCzVGUn
5ycvPG3kT/8BkBa5Pdbvu97BXON347+fF+L85GtsDglsmXf6VDNiirD+h9jxRiEQlIveG9KqCXGl
nb9Ze5r+hhVJ5QDNY5PmQYZOLkGT3zl6vlEp3NaPFPWUa8Mnh9gJWGNNGwAD9bcujQCnhNAYkuKa
YgFWJp2QTzZLqZTm40Awx2HxbuvZ4doyXo6YBwWFbAMa9wq6w5DFVrHBq9frC6j7CQKO0hJIjq81
l40gGGOa9mKQu4+MMJNgHnw4H9qzcRJQwCEX8vBxHkiJ6mj+JMmAnW07DK0HW0u5TzX5SeDFEr99
pc80eXKsBECtkiLvnXYZupgpBgb0ZfWoYIAjVw47cALmb7H46LoZadRwGCkaFY0w+a7wZ9Nu7OVX
8tIxMulHCKzZABNbkH/BHvfu5rvwm+ZWhJj1L0z/Yl1aSsRvuY9iFOsYFxdDbpQqZy8ZhICQg0sc
G/e9uyXKs7J0Ftg84XF+waww95WLaXlSRFTVVrPnX5IpiVariRmJuWf+n5VCOFfAmi/3dd3MXAgq
w/BcxNUn20WOBJeX/PX6FPqsi+t6OkmHuTfFoa8hN/FFaL4f9xe5MBFxbM/bbKnjS1a1os4UXRTd
dQQ+NzZ64+v9+JMCgd2KwzthK/BB8GoIC4OOR3vrRYcuoQHG31f0XbTMyU5SeJlsnCU3tVcoCjUW
MOFgUB3bcUUdwmluN3JPffZ05v7Qfu3p+NQNwtW/otKgV/miRy22t36M+XCZS5YKJwp9XgaiQ5zr
zbcuhxw1OhbiiBw0DsQHmLnmeSaGWP2HWRxbVmxSphbtznfst4MUpq/wQyxS1QvRr0TYxoqOJR3Y
SN+UmlSA6Wjzb7EUO4pQ4lrX/DNXXVBpqKM+8hfqi3HjsiJVx4yxWSeaJofjxqwzoA6YiFuKZ3NO
m8W/9okWObXMPLr465qJMuoUXfgjPnLU7xZSZoysegbBEvzUJq5y6/IDhct+sGQUFABF5+KgTsI+
eiC41HP57reg5aVeeworFYEqniuyXp1lBMe7b3xFfhpnFdXjr8TrRncNZbKZGd2LiTPXI2AlRUOW
LIZlYbeBvaJboJQ1N85n3NEnqqcMbWSvFG/t9A7o7C02lHbUrnXfv0BSJ2h54Bba2ZxwL9a8KM2M
IX2x9ZMgp5Me2lZqO3AjRksR1scJCY7Gnf6khYxBLRiXnJeG2nZM3+SglRptSqvmaJCjQILwpNk0
vkMbQnnnTNlB8gALzEo4HDqMrMojUfnxMwuYABRRw8apOCgpzBAu9aroVgEgmD6ZPwlTFsTnf+QD
HnRo+yXnY63dVD+sx1rYaIa1J7doAG068rtNhCPQiCBS9buaZNmyPnEJmwR9Qk7CtNyj3Haphpye
ThgRYsVV5mFFdD++oNtvJwLtCp2MKLa3CjPTHTqHDblkWCXzrwNovahb8LZTeMSIWBoXlMkdmTrL
L6RR1zDfub5lnZBeLMv/WMDliOkSdRSccUJBzfD9ZcVKjSTPX5jk1q6fY815gyko3ke12oKuT1bL
3/zp+WVlj9Rhvq4Crcd7JfVWW4FMI+r7nf+mk/2AZmIqVl0srFmp1UbKmtv8p0ZxjSJJkuR05KCh
b6Ac0y2na5XTRqMgpVl4DVtEOTBUGz4MIjply04Ndz6mrKj+a7kUc0Jp710WE2zpKkXzu2H/xsYA
xRQadf56t5lIpMmZ+TgHlKXF8xfcbu+WnMSRK1dh8VFRVUHbhbJZxbf9VASR6aIuuk3JxulIbyWk
khkUM31vhjFgZzNZbdc7TnVCvvmK3XIxl2RbswBlH1mOmCA9FyAyNJaVmD5phubArXgLvzTPhJy7
tk8+x8bgDZRap7t249s8C6SNiRRipgZzcPcLjPwu2p5ybBnt1tpX2adwmFBC8qtLhZRZgX2yka7b
0ZAqtlM1dY85DOB/FScg+MHAaWeQHIUrqO5/6fwPyKtnAj2TIdvMhg0KD74+HE/sNqWtlfNtTp88
Mzvp0o4cizAWAtHIsvlingNWN+qW1Qqw4KU/s9CASx3ZN3YyqlP5sWxxUGaYhllwS+zZ2X4nNRbQ
diaAKMmKleN7Qkt954wr88iXx6imvZvw+HLM6GYRzc+kpgCYMDigzlhmkYS+uI/xYKX7eURzxFRw
iyBQ/vKIhm+nqwQuwfxOKOGySf978XQWup8oCDEQX3z07F/xRlq1BAnab/rtKgKsjwlgjr6kKikV
laOCYHYt7t6Ec37Asd0WI8TNvUsk3vHeD5QhxDXyuJ/J5zrZl7YXooOREeLRCUH6AhBVh07j4hZj
NDjyHvTzQaGQ8D/dOYevoTvKIERoP910KG5cdKKd5lJ8865+TEs/8WF9SdG3Iy4jt6KaeH4gYB35
TFtWj4wKoF3Rx8zck5/tFAMzdMx2QTJxhGoYS3t2aMfM+xN+7Ef8qYJYou91zrZ1BGLMkS0wrCey
fnUP93lGKD/wD0N9auBfwwAGW+kS75qnlFgQTTy48OysR4ioejInKYxoSfwa4h24iF4E2jvOiiey
7nFYxGQ/QWuT8q79UJbVpdp4nqw3Hsy1Szgju+w7oXUFbehDXe7N4xyDCNOEcWxIpL+eyAgbHIuW
SGQ6b7meQDahRraSBT+Zv7jk3X70sM58URRm44g3MAyOzmiORf8XnPxaXlzfqBZXL6jvHfkEUoVI
D2EClGlgafytWrgDOyzyTggf+z8Uu5X1EG166IKHi+TmLGnI/j3OnBQsdHR3yCtgcWJxPRol55Fu
kC6+8NEAlSZZvEE6a4XM7PdAWnB/ytIJjVGqSUktJQtKiwg+8Tlh/9XYjbFXUQxOXavyZVOZ/H9t
LaOEDuNeDX9wGivXlcFws/Pw60QJgO540VRX+tTsHPf8n0ZcpbMDXJ3P2M4t8cZf8kiS4HZZy2TL
piMayivXiKs2qAANPurHgl2fd2Bq9B41EHfql5wI+o43iyvc3cahFGupSw9MIEpZqoV/p0meFkZz
s5+JwntqL9d5kP5Xhs0+Qp+Kzu2NtFvS7G5xwzPP+azvJb6GWvePTrVqdoPUSRYY98R2eTy1548G
JrZwpgQ4yL3wlJ5vPdFQPNHvXXNwZOuIb0sIzF7wICiMCed/RD2Xgr7HBjvGS8JJcU5MGxLauem7
Szto24Qo+BVNbg95FPGhIgar9f8qMaS26GKlIfvXKNXjWk00vd2GqRxgjW3sNzwcled+qX/aoZKw
QM813jl1HUHqyvRUJ3Yah9MZwCVwaBePoVP99ZO1cdjNyXMZlf9/KoPYj0sFDE1FV7Z/MEEUG3aA
6MznvkiOjwG55+n7WXWN+Ey/L1c+4NZW5lW1GWT873eK0Jct42jxW18/E2qBorYtcKJHA7GfxCSB
NVZO/0U15xXUNFfvoaR+MBdzkIpZ40qNjRBUEPuat753dwRwLUzSdkk7pwSFnarYzJetOH5Mu+yX
VTz1fv3puA9TKFAvrzayJQAwRcx07g9oDIDyAkre38mtdpgpPCDRRyyfE8LDywXJv8eLiwn1tH4I
qxmtq7aveSMqBLmM274Y652lXzP6st5mTmkiztkhFLh1tKNQE1flnAI/eCzjY3z9/fFSIwPviiGi
CEJ/2hzAWJHqYFbTiWpJvO0uIFpNHaa8Etr6+Dxjg/OzY9zbgdk1QoXaC80RLyjim9r/PHkLwwtX
+QmTp9aOFp0NqsHp6sXqu8yJsq84atjTAAPhQHbns4vLC+iLhSXxFDVTKvPgiOmXtc8pl1IR3E4P
XIq9i5YW6CdIoMsua0vs+JgKcpCoffg30/cWLbeRWbefse3LHn8C0IL9qch5oYFHpY4lJJ5zLIbk
fyP1xT0ctIESPD5JKfdQN3V2tJChaoeZlLCm6lQ1sqLtKKU2JsbI2OzQi5mi/7JGgdy0gomtbtxy
Bym1snBl44wEKdpD6O/iuRvN7lKfet6NPiatm624qtr3Yc7cVf1r2I9dOWuaCxY7m/mCHJHGLVGr
Dwg7m9Fh8FkZVs0lc87ZT+3zYJNsBKyPEmDpzvkegO7kzt6PiPhSlyekBIq0jQ7LyJkJHAHJ/e+N
9tf4anO6xp3SOzmHAk+MW58N9847SrXjEZBjkPxeHVTZXUWdU2EEIaTvWUvHkBIVPjD0jQIbcPo7
aHu9gUiVXRCUuYQU6lOXOJG2+wbXcbmMb4Thi7ERzTYqR/QIdwKaYBaUFwQxlJKFASc+s6r1L4RF
OlcVy8nbofPb5nzoSFTQB68SpZW8n/AlaIlRHhicgrHH8tGU6FPwV/AZ3L4upod3FuTZBxa6XwM8
hnQx0eL0sdIv1pw0mImJj6x9bV+IxZX4rtlp44HBsENvKYOi9DOkuJqXjDk4SEVfRkNjshnANm8d
ijcc1HR1g4wIaYu4LY0JQSd8mgeMvtZCyPQPy+HFJmIziN8a3zz79wqytWlJdvahRowYMzfkLGmq
q8ugR6RFPYKMs2hSr7MGQdY8fj43O9GCuTjdqrNd4sx3XKUbTrB3Zj++Z0ob8gT1ayMGwVuWlfds
vVmV5mYumHuJ/SNHEYhKNmi0EyRk15ns5YobsTeK4EHSZbo8v1RfDuPCZX6+V29AbpBhIu5IDPZo
PgF3gnF2cz3AF7/f0eGVGeGWKqtRMUbVanh4WmrE4kcVhoR3V38LGh+mCUUhKoSGJ57SrHzS0dLc
2xhldj1SUBXCFh1bOrg6IDUzjxlUSwTcmnkEmBWO3/gS2Yg3BPazmbx8ZG+U+874KLJZfgOXcGH9
tJ+G1bEFbzgh7QO2I+SPKRMXkQrqtJ7pfxU5xQp1TdR9ZJBgNoMU38W6cCmOedRzckR8bGWH5bzz
wtp3aeYzSA399x6UEqcc1luOjS2F6Bpbw0IVwp1QWypfFW0L2rSKXxysaK2TjfMsUo43uI5wb18A
ErdRrI2A7/xIYhCuXSAPhei3xxBbF7hZVG7ea6sGnLGb3Gy9DmzNJNHDUdRi3olnZV+aEVryix7i
JpjD5a7eotgUQyO4ahceM0NcqHhPm8uqwRWqr2bZ2dsHD8fMwT6i4ttpKeYGcTMkN4kpT2z3XXHE
HZLriJGhpgHWWKIFqSNT728tjqAuTEs2VvHSWDeHYwSCY22xVAVTifEe78LjqhQxMzi7EIhzIIhU
aK7Nfms3m7yr0nTUifA9T2ejAkV4spTwTwUv2Z8nLFc22dm4aoWC6XPMwhGAO2X4zURyG6TnZTcH
bxcvDB0sLtdOmKNxO3afJAEBTVTR1WQHtY7hoiwwIbIMsk6KUnyTTS41oPnZqREbxGNME0HTLufd
a+/tn47wCd2Xbb+ZVmC71gYTJZ13qiPYleXJ9dBibwfKhdQEh6w+9gNY4UPx/y42+YSVZeS+7cMi
XUZnqDzLg1OYMWO6aVVa4xlrAfJXHHMzIzjFTqrnXnJm4b77YgorMuopTcqQMk0S6Y+SbCEzlF2z
sYBdwChsrrLw4t0DRk4MliLsmkYPGAdLO/0J9wIy1oYCsdDr4IuFFRB1deVHpX/SitLfPkm5NKN4
9+ekkbU3fBxajOnKYSVRGQwndziVZKu9kBARNdT9aloyvLq+uduySs9gGArzaiCkcwlQQfdLSdZC
EkB7Ygyvsk8pK6i+nSav223O4or9Opw9f3Q75/7lvsFnkirNvyqG+KI/49FVDvoph6Fnog4pmIQE
u0xsIg4K7lrdce/IZMUETPQ7Qnk+vP2rUo878xxPYEkKHKv8CI/yrvpIj2IkhFxvYt4nb2P5oAQ7
ajOoZ9CiSPem5SkwBraCYga1FBxaXHvkWxxxd4uS3FupPkmkrKOwY9l5bjECMQo+tpccXcGRYHrv
6mkG13qkKA5MLnro7ABX2PAhNoJxaUa1pGObNFGimSiZJgjFCaMXXNIR0hVOs+oPAsg+AxSYQpP9
HzDKtkpv3hY1kdP3NRTUXhBRy1FiwKv4Gs1fAgQEGpg7EUvcDQNzTq1lLDIPmyKV51XplBXnf7CN
MDjW3EYyx3GJ3baQwk7OuUZQ1EKYt9ziPF3Qhcy5AbNc2gyLZmq5LhPODRjnh7gV+d0iZvNHbf4g
mlW79JKqLIClHN/LWS0QENjJSB1eFGEnIKf1+/FB01Wb1mA9egyi44pcm3gJwNxJKbeShQYB4yzU
JYeyTvDoOg+FngP4xxzSUWwRTTiodZD+pr1HZltdurV/FcTqK62cktmav5d7eu8KQZwBFAqNApWP
ar0duykAt5uL97BOGP2Yr5soTmyFpyUamwJeLfjK8ciG62A1DjpFF5f33HwzGeH0qdFZSmsr0Zc1
ET7z7099PK0jS9t1zt0D2r7S++4w+kuHsjQA0qrfFj6hHZ4F77MIzyHloyDn/xnRF0WfJuk8Tq/w
UqPqbTTaaOV7Hnf9U0NCqqHQ7Mv7MNqDBzsuZN+vQhtiizfHM/hsqq3zQvBN5sshz6bR4GxSt7jf
zyj2cxz0mNWKi+TswRZrORvXhJl+h+057E5x1UmuIq4+GFPcEJdZCf5HgzQNDCbe/P9+ocNFIlwI
PYrN3D+7xWb7tnGpxExjx2zFtej1aP7g51d1S4aoroa/JZYhGkEZdiMVfiW8O5gf8bl7QWvYjfKm
GXSmDFc9WDlP72AQNMAoL5mdEKJE7LinpyRtspTSt1mxbUyDoth77WXd/OtTYDqajSFpVjoFttGi
YmlLc/xMPrNnJ/d+B8tHwnBrunQLPaGPCfbQY8uEnwcOlrP/4lQFab+yduS4VvYkON8uH4LkVbSV
4iH5YpxcWIesPn4tnrcTx2Z0l5lYDUiWAvDkejo/oP35u7DG5z1O6z5babi+XcUnDFMwrHu97px8
JlDPWjL0nmzu32BmUqEd3h/hFW2Zk0y5gPJkG8TInvdbBTZxhaojNIeUnyC/eoZmeHqzZ3D8+D1B
VF+k5Wgm664E3ywHGiYbxshxAjXVI8EisTlOY+GP2oU7Nxz5kKftY0Xvfb/6XvuXUkRj8Gn9tUrI
2F1PWfh7UMIbjqZfp4egZJ06dcecG7SO2WvGk3XyjHJab+tQyfPrtE7kj+5eESwGhRmg910VQ57q
HRKuIqymAITtX2wRbXvcBgfhcWJyoR5UH9vNghXuNsX4inK4a2YZw0OqPKxhTerQwiHtE6qi+hUN
uCi7fQq0nfHQJDcGmVFW5cvhr6fBoZfKac6c4UuEeuseJYGQAPmSAUsKEJienqfjSPd4iXIvM0wv
J/DuXHCnU+00OEgZ4d9Ucu5aMwKcKindZuNAG4JFL8QDFOmTr5Y0hdy7Ju9a7wnBe7Px+e8faid7
MrLySciJFS0EcaxsZIWgoZV6uoqDdy+JZTeeC1VttIeW6rSZkXYmZ/ZVfcqd2K3DAtDkLzJ2Mg0e
RHAsZCKx+2+wkergtfqmzs+4RrqY8de8gl4Qm3QKkxO28pNyWPnQEXS97IWdVIXP9Le+DLVOuvzL
JV2hWYZdMi5kn39Fdpchyv/x/zEpUkrRJh7qlNy6zfwekikus0cOlqOq+aoyj/6g54rgXHkIBFqh
NsF1DnkNKsqOdUzlVCKYR6rIQVQp/K6OS5upuJ/FJdm267lTVPIIs+u8PFpAAI/Uy0Tq30EG5eDx
K9p5YbB7NjpcnhE5B3wp+8y3nShrEB562vLox61CyVJAzij7zpmcArhEukkmvKUZ3ibI6Z8cVFhq
dqjYUNTMMSHOeXEFOVlcK0KGCqguhm4NVjEF+FFvcmnQooEDIVxgOQMco0DSKHY2rE5943roWb1W
ekpsBchGqNziOdFbvDzqS8nkmJEYgI0IEHtE4zsh6erY4O/8mHz7eYnJyJZyQo2uhVpGFzGiKDHk
7+fv5/6s18D93sU7Hcn6rXpQkZAngf8TH3YaKOMKPgkl8GAgKsqNptHRPi1PTqiMSW7zIETePqDa
l8M3NMW4Yh5l3wNCgESaRa7oJQjFn6CTSVxttdE3qVI5HYqi4PzllypKsqRP4bCqt6n59ZYh5uHt
/MVhWWXNsq6V1BKVo+61vQkMQFupXmP73VjAc4hApjzRLAPYJMNQotzjin4yg3a59ywvMP6ZtA+c
LAgdRxm5Ecwo0t2IhKhBdj/aa7MxAtvoDFqY7LUvrNC5yTu8EVNcM5k9d8bKV69Hpgi3IDekmCId
B3gcRjNo3zVdVItsDwLcuNKCVXQQ9bYwFrP8WYh7PSvwhNJOgI2te0ZFw13wDLr0rwIXI8lmcfTA
XeggQUzHWUYH5zsLRNXJyA/nxMzTIJ+ShVZC/ZhOSzLW9ijveaBfHIx9bOZVYZfPYo+EAhylyqZ7
AWp1B5ykDs4WwQZxbHYcyHIbI/OPUQ+kUvriET502FMbs1NVemB9D9312tlr0Bzo/w7UnjV2OSBU
WcV2k8GQsS17I0t+eWFBaZOfHhDKLXPaU83h9rp6AidI2lxj0YDJVzrsm9aiU37FDL9Z5QBFYzpl
arbB3EOGXvBdb1NCv+QtZGhcMFVske8pKuu57/rYrkVtV6XQ1wDx/h61FPE4ixg8L4EgSHLBwoaT
T2A1LpNJKSSZrGb/KL1OOZ69YKPKNgFXYy7186+IvYOkQPtb8+Yd5bLDjHmjnweBqorrZwkSBKuC
jFDU1an2yTW4NlzasYwZRAUP5XJmhNw/sPIkO/af2Yi+JjAAbZxxyCue6Em7c9Zg2WgUq6ru8Tps
g+RsyejqhctgA4+IMKOyZq5OqE3AJrFlFOEd/UW/zkCwyV38ykaXeYOKIpiGgvmaEBZOTR5ybJTq
cghJ4T0ctqvXFLvb6bLzP8G3x/LM5wEW6FnOkzX/wkN8zp9haihgha8AMEUxDPV5jqH8XAdhCiPx
3eGghivc8Z0Rwt0lDGXmmAj5KGPaHz3OIcvuMDsbefQOsza3P+AwJgKHwPeR11UTq+ifq7149uE9
IkaTQsl07nT1nTBsUoywItRZ0fUjTWxbkkiI1b10BJaoDpdU5Hl2T67klrKoTQlS67fsBVOO9eZu
U2u1Q0oJO7O8XOGDP9gZ+T/J86qANPA7kxmPVCA7Gv7qtRydIicsRBk80mYppzrGBytbSXSi7lg1
WpW0fuwGTyLZiVJFiqxHC6zVl2RnU4Aw7bnifSSfrw7uVAxyuwaEuGi54AnxhXcnIwiOZWqNfh83
NB9PCjBU9VGuIRa6WQr24CUJeqHnGO9ZAEudM3nG2+HfbqFLAlc5O+PkKRKnWcPXEKIRn7n5bBza
Rf1zoAC3j/LCQpyOWk9gThxPisxC5jmX5Abp8khwrHqcWwGyYVK3GFAyzlxJAE8o/YH0kr84A3Om
Btyds/wQMmcPnGRoP57xr40I4jmLZKVeSrqXkGxa4mdV9uiqZB9jvOmiU0q75UcUlhp5zO26GPRM
0mgXG3UKCbc2/tFnpQQ0x3rawacEp8yShudcmOs157uwp19sTYpS8RU2SbkO6lIIzYAst56Tor+L
qJUaOB0fX16xvAkZgDKEX0qb00SdqURvsow0fROwfkEM+wFHnxSDR9iNNTSFCM8TrAIaxRYB3paG
8ClHjz8a2KW8L7abvpJf8PzUjTRU2RcnmNGXHYMxQXv5Rjxtx4RN4aqy7ir6WbzY3wnScgjIummm
ENAJzsdKr67de0xo1cU/2aXpsTWEWM/aWL+l8HkL6o/g4f6vLXMeEVjal1bzQFPV4nCMSk1+gzRY
7mwTlOMboWO+KySGgtN8kAczE8pPxPK2E6sMXO9uuVqZcNXWSYU+5mzX7RboRJuaTmLXFm3Ymb2n
BMj3D4vgWNADYofRKQeo/HfBMEcvaFl4+5kD3W2ghuiNZyX9SKPCBmZdspGwBs1Hf5huCGdW3Ihr
tVlF2f5HO6qTow84edt5z+ZUlUICUP8LXtGEWmDM4Nnrl7j4YXAxMAzxQkHPcBjO2DshJ1Q8zvpW
l/UNFisBbENZDV9aPt/Xb2746EiF8OZGq1HNOt/JHV+K7CyiYdYpKV4pVNUCZ5JgZ+DsCvJIgbjm
6M74v0uErxj6UIcu0q4t28TsSBcolzZ5jCmFRGZx0l5dHRN4ZTpIKaRFQIBo/1eRFUN9r4kzzE4P
sWd03EOyDNuYu2mUxmByKyS5rWIh8STBFQAK4uDw83pzFW9DRkVlUyeO5K/amtdqahUBr3c9+sSr
VkmOd183Ttqwe1eKY3paF1jL1vqsIlB7ZsU/uix8rFRmP7+bg9UmofbNitF+ZDvfRxDMX/4F6XSD
OH9TcrcjC+eml9ng+aUZzkuJ4vU/6OtwlEL9SubY+9ZpZfADzLR0N6gr3oHxcFKg3ZIktuphkdKU
w70E4MPXc2NMOKIVjS0StkccFbFdYnS1C6t4OIoQj86moQ0nKpUiUzgJCq3AgnBQSATm3ehDQ//+
GRdlWpNuARWofehrdzkaC7kPL7Ez+RI+t+vFRi7gQEv1cKZwsGhNOls5H5GiqGBGeJ96nWF0aylk
LvTrpK3KlVrLmW1/VCPeImGMtMpvgCW4FgutSCFt/zhdXI1ofTk5Ik1GWqRR2sWMoJaXCcXDd/l3
h/LMvZpMwS0JbF7HEEtVG+RoaE+34o+K8iYEa3X3Shnu4A9l5/hAqqBWxtyOEYR0d/a2AZCDEjSU
qN9hjvEnsNfcqJkwalDV5kePLszGDpV1TTb6D4h9PU+ktyUd3/m+E4o8gsdnJlE9iTSMsWxJ0A0q
q3+Py0kIVxPyHOYygIduo3IZPIIcRFuLUviF1vfN7HfhV4+js4cZpEBpcQWxnctZxNSHWLufWKvW
ociDFKKleRyluEfbEVVcFh0O/HQulfbFjXShictkuIadYQrjcUaomMugri36HQ6G2Io7FaVznpRV
VP4g4qsZQS0lC0kDc0AV8swAD1vPhP7TeJwTZXXhry4ulJbZAfxEalqc4wOmC+FACDtjpN+8ObBd
kbxpthhNd5nV+Cfy4LZ20dOdXkl/Zw/j9mf5WOIKbF3qSDVteV2nLBZI8LiQxy1mYoVYe3NfiCHT
iVjc2/WuVh9QBuIodEvCR909WaIhJctFz/9clILSUpPq1c/ENNBKuqEIL85kGhmTdtFuzlDz+7b9
2wlAIadltV1+XdbzUB/DR7TFPdmst3LyZeS3IRCiZLXRwgu8H3PoRLg9r/+kkbZX4HiXdEr5W9DD
+hOhWTaJPySEpPBwGh4qmNHxPyZL8kvYIlEUQjTGkMDKOlbuvISrc1ITB/DVHm/yxv7P+3kDDjJi
VAKrq7VwZKwrwpEwlDGiiM+4bgTJiSXPVNGztVTVUwq1G6WuJDC9eBf2JUvdKNq1xIXoaX7CY3Zp
2rDjmGK3FenLTfJcXjBoMxgnr4FWgvxzJ4VbgX4hv5sDabCd7yxwNxiG85c72N9IhMXUlwrw4DeE
QBlzPzRDtvfiOG5/dy8HMaZceFfaaLxdYanVioqIB43VtSXZahAgdMqUfbtPvh1dbyidyy6UNjoL
755jXM2iFAxGCCE5bWHXbIfjsgMu1HKOv7FA/qJh/wc0dEp4g3jjVM6P4LjGc4OloCVdvlCgD337
mJMo36+cUrryeCHhLeFB4FeYJHkdxFAGMZRy627xDisqm+IJqcj51A6lPR88/Gfw2bQRS85nvcxM
rUK62kqbqeGg6d6DwyRG2TVpC5gJQo9marB/f7KV5Yxeih6Dp0rRmGPfmHmeEfPTSqgbduEFnOBG
U5ZIkP4Gfx7gqeTDdaap3A6mLoWzG1iGCNUOp9+BtR2vJoO1gH9TR+J31TEYtgoBsTx2RYpZwYLg
GQDTJIHJyU+YuSoT548QS7lHODZ3XQVS43K0HBGMyCU9q0vZJQ0bqwuhS81vRnnuXrTV7Xn+wLDO
Whoc4ZnrCF61NARdZslxuNVSpIuARcrjfFIUvLLm9j/fzS/rF5Vy/QfY4xsvTid/kxY8aciPj63x
EWCQHLQ5zelMHUVCmIKzegU5iZl98jIGOioyMluBmXvihAThCJsvhCT+P5RGuffRajyqAdrBf3wt
7iK/7KRp+GV/WhxCz6rCmvFNdAqls3feXskkbRfl72wwwVamYycyZWPVEzMNxfqD6jdypjqnmEYU
8oB+Z7m99I965LFuilg+q6+Z+bd9FbkckUtEtxrBTGdUwRbCbAbl9nIrGHhBzRapGAkI4DEHGwHq
c4fxzQ4YIFZcZwDFjRtzviheWSvFEmPgw8mNZwaVLbRIDZEYYGsDNJ4BevSs/oK2Uf9MfCDNi1hy
GhicUP1cJFNkgOhwG0DC3IU2jse2iNNlxf9UcBDwW/P9P2hC8FuWsgxMv2z8MWlkgKz3dkkkq7HG
hF6stRCu3DaK5OLZh31gFc/trw53swHrCbqzXeiIJaTP91ZhbeMFD5g7OaLONjIR44ccMcKM3AUn
8DyxdpC4Y5f2jQlWF8HwUwbSfYEdG4yOSIpeDD1BRQntTjacOihKkF+uwk4SlFNqDOHNiFUUkq8P
WGbALIY1RFKPQMTaU42Wg1OIDvnvpXBG6TGUZD1dV3lXi9FJQ/U/qZGnFJLsOAvSzpT8bJ400zIL
+EymVNbUGImawCkM/+UlMid+Ix4y7anXlWzIyRXj4UWZi0xZM7hhSzY9jb02BOhDdEgckx7yfXs4
lSdoKnuSF3XEu6QH5+O72zMNh4528wiPLaCdRtiYlF9HWhbojgIISjOb0gxh0cJsu/cReusORw0H
bEaQjUDhe5kOvHv6txo/7K/s5sqOZKOYJ6ygKV1oNgOiCtknDVtbOxgXtBwLb5Wel9U7OrtET5B5
1L4vHz4Yf9LlG1Ueqwpm3qg/aplrh6hCLMiKkJUIouewriPpL32TQDqbmfd7Ta6KNMHKjvQaJY++
dwOJaRdGmvbEaZDJM2yyQFL/XxuVe+EQgJCQVIkJe08WSEPKYQ1BalQCOzoLbRTYdYNVWyH1ocIY
grXR16mVU3VqDVzAsE3rnpXEz6lN32bgDJx7Cpdtoo760zFa+QN3SHQnvNHL8bAuCIJBd5TZJuZF
aNa6eMpCvwKUkjJWOELmazxN+JEIlsx1ITGjfqlisvfJPws/15ax2P9J1Z20ZwtGuAPF4bRXUj8/
6vdN43YeFQdVx9VwMsqFrIzo/flwBJex1vhmkHA129DYVwnY7GxUwWupYrNppZHS42Yc1qLC6ZeN
UgE7NCGiciA01woWv9kvn3hRLZ01iXmFHqz8OkxB2HNS8FQKVDwqUkkuxSOYrDboZztmLLTgn/B0
kzFfCMQxRlKlQeehT9IN/4e/Kt4K6Hq8xeo55ivgHAGQX8vA60Vs4Ld4XO7PEuNoTe6k+jJGTlfP
y0jvfZp0+qlDo+hCp7tDpTrMy8Bd27V/SABPiFT0r9FxWmaIVKM0o54vixVRg6Zgdl96V5PvHgG1
M6K9325f3b3KmBySmHmn08+gCpI4GpzLaQGfFDUC6tKO+MulpJMPiEnsHUWE1aZEP6jg+ufhuRTn
mBUwMBjaHEKS/BTYmri7NqwkJgyWxouu/jq+zw1+LRMIj8C5SMEq/JhZRREoiMg6e+qkDW1uaOqF
ZwUI8rHONZhk7xtn8tCfL80GR/99iespB0P3dyk1pGf/DP+IA7N8oaLh2QhtaPDW/4Qk1FtYSAfB
7tFK27CH1zpfays8wmZV7/6/Fxyz/Y6crJKnhwtWOPFoiqhNuxXTdocKnTNLmP04eLBmFAr+SJfi
1kErSiCj9Zs+MP+eCTtKGMUVyi4jPWQwYT/FGiVm4I7tnyZwe3wK8zPOBGzdeH+gFNWoOgMksAWc
Gp8fhq+BS0z5it5P87bkN/Z6kc/dPOF+hYPULj1QuxTvfCvcMDJIPo5aUq3RWMVUeu0ALtbho8+F
yxa+iY9gTt99JycrbicFUCe/H+98udXh5dGG5YtydtFFOGi1hBuCPlXwFOJuuD1UEQhxmoKjwpXw
SeHlOH75PIcMyOvBmv94lH4sOGcuJJRGxmKh5+gSXLJwNTPMkiMjqPEwLjgTQwtO9D7z13PBi4Nf
WAE+U3zYEqb0oMgIsH6Ga973vqzPAcND4Uv56AbveMlfRcUR+FvE3EVog+89Cj7toepj2z7irBsg
IhE6DLUZ/eR/Upw0NRgiMA8uiEAi9N96ka2bEXGEBwz5gKWMsPxkh19lJNvQmlVec34RzaRf+usm
S9oWq4jyaGhX9Lta2zWPoqhRMnmDqg4zvIp3qXU099lqk+L2HbRXB6A3xfdTKGzV4kQLcK5Hg3P0
6TxgKDqbOMYsjuZWG2EU/GKvsWZKSRqg64FOflKyK0WWf72cxhnRDdAlsgsFBIizxOX5Ml9AuQUQ
20aKAWx9eiOkvwP22LC4RjBxxjM/6lET6ZUdtfB9kbBilXOE5Xt6uoRnojAb9m2l5lrHFDRnVTZ9
M1MSLh69enucFk087CAl5+3sr4Sn5TkoSmasThdGEqz8aKEsj9vMXsN349wSuhYXhiYKNyyJSj2N
GbqR1EZYnF3AKKT/SeNy3vwrnrUhqAdIZ+g0rPVUnMVDfZMg8/EokK5+pvNuYjz+7M3mLYrCBYX1
0W5YPCBL6r+uHUbOzPM4ues9M3mkH1o7o8mY8h5EqySEjAjDHhp99LZM5Uyg0GTdBZJ/YvyCwo2G
eUgDgzr56DS5gl+WTzS4OFkZPK8pCYIOyrW1wV25JMlyEaXkKXzOP0TZinY0K/zQaJydOvjrfesy
SlAr87LGGcGiOYmLLe+EYjAknl8VKnok2h4Y/Kwp6UN5lDsiF4KZls2OOdeMC8dNF3QfVscqpRti
PlnsF11mfUO+fPGPbtYxx39FCaAie9v2Aw3a1sYge9Sgskb87DtS0uqnbFJ84d/BCAeFC4C/2Axt
iCMrGmC59avT/gW/0Vgyg+auCSoPlQS++D9n+wyq8nmw3iH7V1ffAh1RGHxxjkk1hp3ElEXubrSZ
TZFfFLOpkRuzfhol47bMtw2yHxk5Nvyn543BjRkkpprMJYFV2keKlxIwyO8k9HVBItJEZ/Q30dA3
T/iD6a4X2VqqxNtHipe037eFJdlbutRgy294HGVDlj8yHlFlauAxpULos57+ReUHc316MbDmCwsy
fGMEK2OsjJsdG4rMRee6TE2Q0k5gaZyoTp9GuFy818Niqo2fVHh42Wz+SxRRaiUvef0q5BwbQszf
Ip/Ck0oR+LRDsubNIfatzOQdUBItwhAJqs5/Qoo7seVI7P+c2P/oHwWRx4dcwI8ygqdqPE3HZ8lC
rA2rYd0G9oUNKUGhiVOZ5r9mzDgQrz3KlmO3JHVwgyMPCcQWsR6Dj0THDkc4Xqkd3DiwRMWJiJ0v
44S+tLEvC2ZvcnRPEdVLV/Dht7RpwXWizweTquzeEkXA2rXTEOhJ+X8spKhaC4v5EFYhN+hazEMt
0m/u4PGt+zhxEepKtYwuYmSdi0aBRVXCyrWoOvoYKqvVWPt5PSGVnKlhlbyBdsU9hE3669i7ycw8
z6IWsatZKpyrB7ah91QMn+K+7JWxFI2mDGsn4OLrYFM/wqAzeH9DYogamUK+0jzsdT08c3x8cugs
xPfij7NilRZkPzxtF5EEiVJBSTE/EhrlJD4wsMgbk2ZK1Xzb0HwgkTZO7Rcl+rIs0HAa0KbowKTD
dSe3r141m2DfWS6KrgmNjgM5iLpAvWN5Zu/NrcGPmXu/QOGsywcZ9HlhgA/0RxbkhmoL0d3hutMI
SXAO3C1hTp909HZ0yRCY7wztkyBklaP6XhYUw5dW3nz61wIw+dQuV1x2XdPTwqcZB2Eyr/UBGhQC
AAcs6ExNUTPJ1sXW1T6ssS3K2XCiOgQAbn8n1EvvxBU+guqlmFvV/CWAv8q0aVrqYbE0iZMSw8eN
VEwarfYT0aU+MauxQoToAl9QpjtUcepOFeo4dDarjzQrMKXWm+nupUpuFSfIadWyM2/CzoWuJjaW
MH4HiCJt/y9Jde7CfJgf2ASQBkhwH/PQ34bjuMbhbAITlLKwOn+qWT2ahmprrPjgFtdGHdpRdL0T
H7JImiZANwab53UBjNNIqIKL7GwyKJYNC14JRZFmTzeay80mTb3Z824lv/JegnMvwvjdX9Bakeum
8MdCezdRCzqVwdW/sxKr6gy2RcvXRD1tYyKUCbO+x6qNn0HPoLRm7nbo8xSAA7ab/qi6QcJV15z0
dD/XW7FY1fY/5jKWzqRhAuyoCoGslcmEHuG9+mZ+R5QJV9JWTQG8sieBWAGY1mrrhpeu0+4KYMX/
socuNXvh+cbfTDnpZaTJsZTzMtAw89N3XOulPXb4xtuXSJplN9cOrfCUdI7TEL9GRrAs9YxFRaKF
RiAHFOrArjGif1nGq+vK5e7MD5YoMiGqGJmP7nYFE6My0dqx1MrHsHusjpokWn/cCd34n9Jt4Ip4
girZd6L9Ip1U+iR3d3lYQuN0rJ4F48aB3oTYAd5CaMYgv0l0VhZS67Y9ZBloUeUVG4LpC74GpKdx
Dx0A4MASho6XHgi0MQoPlvGwrJijcuqAeY7/NrQnMVEcXKnKgVgOx9ZCQdAJ3XErSAmFm5Z3no67
Ev5auOmOxO/pMVcqHeipm0VvP+3gjaWg4GjDaYXVF1NSOneZUM+QkwEIUvToJKeoyuQSben1nXnq
XUfaUlvOkbnrV7gYMRgKisMf+/inr9KSvJuzB/sq3TNvQ0yUGk5WKyvGxOMIxC10eD3zj0e8DlV4
rSpzllH27dUCdoBy7ZZfYwYBVbqLIm//XIdFBWM5GA8C5rVjCFIrBShi2OJd4JXHg83aqmth2X7A
as5CnI2XHdCqRpCZVvXvraL/XSTLV0mDgLhs2LfpkyoRHTyvtuTWO5olnYy94xghhBJ1kwF+LRpT
KF83DHops7R3XcOwvRFfvi44wNggq4ytEJsAx80axc4cGKCOto4JQ6fhigSq+hAGIEpJoj42dg61
cx8g44gs2WYDxYCeEZ80FIHJBYPq50eiXC3Gmm8Vk8ce5orEe4/pLOKvPfzZZZb1QxcYd469ncmi
QBawz1hE6nrnIdGUNEO7Iq57EifZ0dMFvhzb9F2e/+mM56oTQYSg9z5JcwK+BfQb1ETzRZnx2q4M
ahXggCgqOCXTbRjWMeKwKOXnAjfmUh0fQyAEatNMqzyJNixtYmaXpZsRir6GLSD9JuWX8B/TSMQ+
H2+1mVMA3hPFqyPmWKKMHMIsaftSzRa9VVLBoZmNsbyRTNFhJ1CxnSz6//Z+SjZ49opUqQw1x47N
8Bly3aox9G0M23J0aVTctN9Ysh9YxuVoSZlvweE8TcQQOdA3GwapcXd17JG9sUBfnB65idR0Ni/S
O9qJvrv97+w5VHwDG/wh94aBr0D5wbXaW2hirIkJi9gunmpE1JZmWQludNCP7jMdqnD3bU/Yudoc
iJfClsXcYCr3b4vcZ1tfKsRitPSw9JbdD8XCVr++4HaIc66xyJxHQ1zBFjMnk86DTyhnnveynwQq
gPpZGmpK5agYwyQ9wLwOm1ktKcBhZGjDIZ8Nl6NmLBjXE3GvaNFGSpJulKCzCN2tfkrggogvbGMr
mzSaupl6zlClxqQM4Q+iD+u6qpURJdIyZRrKQZ3vhHLPFD40XHiIOnvAUPv8G7GCxZAwETAXI+JW
Z7v85jw50iAxKn6DVqjeog4aU33zwzdRqlv4AuLsg/EeoHS3G4+yUwYVhMpnAPhrmZU9dpkG4PZj
PuH3ndIQRsxdLXCfKnhpS7b4wixQU8rLHMhV8Xn5rRsAwG+rktsH+Nm0U3i4vQGZy7HzaxFhxVM3
Y0XwM9cN6EAWYgk5oumjXQDpcja1Tj9h7H3Xpp4+lETbRb7mKqnCzUwUqdxN8+hTqIJx7Chx+pK5
2hon62aZN4odWTXTODY/KzGWbIyuNTBRXlgp2TzEl/pL29URmCR8yx3xPwQ6rBbxzS0lxsSztzqB
A1BVu0+NuIVrvfbEljcRwlHrR+TQiSVkucGmEJEKGnX6XhbdzYepgSkcTsdNxgqWCmoixpqYRvB/
h/tFCszqk1c1kippzbPOVx8NkYNuiaaxRFk3DIWnQZpWHPoMWTUiDS5AxLPv61SFV2jjDVO9+34q
H80yBWYEc7xp7LlpkPKt60SZsxZsfy+K4DYAxVDWpc1pp8PRqrPjrMsuKc5x+M/Ob7ub+NpUE7Ki
tysXe/k6GEoaZo5PcZWdxeoy5y7vELvi5tGyQFdqYDQo+MIfWOxgSdeBKvCauxVZtJDHBrm6fp54
3oId1OE3MgJDE1+8wCglPQqtHZs64W5oCqxmGzWxfIWYNhxYr0/qzOV/wEbZgHrS1VIqOCMTyjT2
UKBlvOSwvKP/mCuxuRKfLzLOqaGSD2n4M7JB4OPWNT9Jz7qjyQRawzP9YPMV2UgtfVtMP1KIny1v
tVbzV+q2+ZF7UXZa3GlmHT55LS7mpvJZO+l1wIjUyCBuXhlnkqggbzFvZkRr8Mrtd4YWLHO/ibPv
e+T+FZlOQcugkBtj9NqFlOoXuw2d3M7SZVpjbpybLwkl2Gg5DCvbw8kX2ad/fIrvxStQDtsla/SU
FB3/o3vLEwkM2wsYVb9sAybNjWdvaf8uZelkv9NksED74D3eEW/wNOeRfb0ifayrU22jtpnW7uWZ
oyQpcKfUIJbQwQgaRhAxaSk3UkwVzpH1WxfskbI4t5FUAiHTWdrZLDDm2lDvuVsozM9XBleTUkVp
GUmFb1wOmsec8YpZCV0gXHAcgvLPw55WjMV6eIbj1GqnQfsNQhOW/PghSa8YdiNJXd4hW0asu4uT
we4n8ymVYppf8nhdof/QAj6pY/4tGbsJoNegof9jYlcL38g9J1FjHJs5pvndJqbLfMhDpiUwReYR
oxI0BJ/5g7KnW5H3mhPQlm8EqpKOrhTBwcum+ZPVeXqvWompnuDhpZzJ1n91+wL6no9truZsdphW
jYbZ0m4tK5I9IBOnXtFr9l+9Z5EYFK/Uph5fRmdNZCrxC+WNssSz0AeSmgBV/riFa48FH/gf09QU
W+WqIa9VGJFvsQMTlCjttN/LHY40KkTMqGa8T2QF/IWnLBw2XTLABSs9i4NyQkPNty3aRKib+Ncu
vIP0pC2nBr8GHcktlcgg7EkDKpKgvMwglDVOLzoIIjpJHO/RHCcrnAOpOvpFIejWMb7+LxVaxuOM
RwU+YVd0HYy9hUzRYdhI2WxbD8yAW/7UIpzQ16ITdwHQpZQI/IihpBBQr9qnB23YMEFvzmSmw/Ln
s7ICDDXCpnneNxeknaNrlOcr7SqPqqavDYeXiDh+TgYcXQoTYAUhNJI18l90u5jkwejhdEolsd10
BjgDA3F/V0xf/oY7sw0sP3IRAvLLxeTMOpNfPW9aT1rn6ikG0GTJgxXESoyhqgBkQwE8fnw7mm9N
2I7yoHi5ID9vaDXTA4O97MHJt9uYA6x0wAoRTNefQ6a5cfvkRv5khGW5yo3qUHtIRu1Z5wBACtrO
XupMOmDk/9kTstYm6D7KvyGeRUN/zTh/SmvMTLDlF1LqWv/0PanV6OS8q8EiELn3F+PbWODgkZhv
r1Hm1xqxR7dppfPA0av/4FT9KsOIXs2xaj1RzccOBlO81cQwRhb09HoAHjsHOo/dvb35/zZs7q3S
tfMx1kRNTLpFlNZlsjg373Bh36ajyjXIwzdXHGgqiZeGkax08h2brtlXfP8Q9VBhfIC1PKGTxzv5
9ngpDsFhPv9En2hsAluKlOQUJKCmCGpulmTDEni59pKJhD35BKTeHJ/HMNevjBfb2rZiHSkb3do0
3oJMOISrdeVxdpUA8DbkasR1YXM0YCBD++Yq0Hjz6YR5Nzfjo5q9qRdjR5ypba8+3ZhyR3lrABpF
j3nBCkwmVrY4Oh9Ceh5iUjFv8unm4j8dsxEsle40ziwA5+rQI6XnQVFbVDhYzJ1wxjPqFb56v0/e
QyUWIelmVy4RjEt+Tec0hiz1btkqrTtlgkRtIiIlbONwoMMJD6mWIjsUhPUQXiMxIzOXDQXJlI+s
uhXQq3ZVQ1AhPdvit/7dH/DHyjTZ9UO4YlxRHyEOVipA0CrlTYPPle5GhtcAbkxQVC1KDw1jJiHQ
narNarW59RSGGom9VkG8joREM3ectdz2VFf9xqltN/MX+KkxTvW2q9L4UcrzZ0zMR4aPYKJrR2Wa
fR/lpLvyRMpWpuRtZpBH7Qp7wFrgD9N3TP9zyEhMAaMhw9S4M/va61IUdy4cN6rQg7oHCPYpn/60
VVRHMEyHajasxJfOMitrPblT4D1iYoDgU0ajdqX5b8ifvOqm1k8iyQJ/ks1d3rnNQbddKwjzz2ym
BMMTej7ELwut7736jf85sE4/6mqd8Km5/T1kWGMwEhywxpMBkJKIajaj+1wplmUxe8RW0kjNvg1Z
sa2kwBANou71juaBW/6jrqiJKoItAJHU7xsYX0mxwgZSQCeW+BEUDe+1a/paR5tN4fiFlIvyowQh
t59MpjBF3ArnAnybpSvGufS5PCcpIYxHMgnnFWeUB7KsBhpM3r2+T1ZpM/J/6DA2CPfHGNcE4byo
ai/iEpYSgvyhON/ulEJbAB+fxmI1lJSfEIi2CsIqQsXMNzix6tmgFDHX0kEpVkCQikhPLy5dWtKY
IdjgZkc2bdSvpN3AgUyPeHlm07drbNEi66NCabhSOV6JSRKsivuXnmHV2D/5HmAJT6xEyr/wQ65R
GuGMgTVmx2UkPdE9+rPUNk4JZkIZEmOrTquIGPo14aa2GkqTnFdbXdEZNbZdva4mDwG6rY0igsFm
j3IDGB7curMD67keKJYca+31lwMGYv5jvxXUhnKvdFQG2+BggiiRqBJSLygJ8GDyFz5xEnLdMXBR
beVbyf/U8p6ooHwKJw9Da7xR54DDhQyZOsKnWkld0lSwiskO7AAJNdDd6a1tJcN61+iYiQbVCI3c
RYir0oLIEAdSP+2s2RW6GngHtxIezpWeXXky/IoLGBdLa0zG6oSXdUf12xdx9dNe0yAlwtYWl2CN
bkFyGFPAzdvin41+Zq63zKV2LADuxeZFYFFUntmnA3bhpCFM182vfPOo7eDW3nbIuUb/WFqS6E+l
IZODHEGvIsLQxlAWNe1Jbeh1n7ChFmSpokUiQGx8feyU9uii/zl8MpIpUvKXbAm4emFi3rW/9jmY
2J+aCdtVXDTFrHvP9f4LSDpTjsjm7J6VBexeGT5Xw/hXVf13veOMLQ+I2EoLWwVv/UpubEiaX0HN
Cpbcs+c7ebFSq4k3io1/uoj31frzmcfR3UDviUxL3XDhWhTwWQB/6HqUfWvfGZnOGzMgxqddGEQP
cUqGlOQt55AxZZZ+0d3GN0Zh662DUsHnp6GNQpQUsPsd35IB6/msaMRu3MxeeYFhTysKkroS5xUJ
T5JLIY2kfBCxKRroi6DVk3kV6R62wbe58KW7pOrzhl8pP1ZoT3wBtnsVrNfEh8l8Sqb+4YxbPM1C
jcnEwzB+krsAXwgTy+T41hGFPUzXi8RcozcKH9k7OSbT3+9vEqrdgUjyLSJMai2W86zDCb/07t9n
5HxfxBnk3bNFrMETMwTMZNb5V+kHt5uPWb7m9d2OQTvAmF5pmTcYFyY/FaOe10ohrBJSksPz258A
9V0uESGYQjaprsaGVB4RA53u+kTREA4R/sumfAmDTOO27HDyXCzp3b+5HKdeFTmSmOdhznNz5mmZ
ACt/KNqqVnVA+HmvpwUqrR8vKDY4ojOmZksE5WWYHPJXBt2E45E7WZ+9As9eK132WNVusapQkfQa
KGqZ98+h5gvXGjIDHOQanR6rsPtGqTsJhpfiEnlQM5k7J77RYfHeA0cRGIFzfWPGss/JEImUex2D
a63WBlDUn6FWIOLm1kUFCnRzxowU3tnITp3J9OrKl3cOzEdKPYJJPvn59Lw0Z2VnZef9wMLgqT7V
phSjVdEXkM+6A60/D4H2XsjDVvJbYCAfWmmPJhQY5PBjFgsIxN5t46MLQwe1EesNY14qj8BrLQKm
0R30DPI40uK3RgFEIbboeG9LwH0vBtBYeE5BF5OIcCu//2SmNjXVwZxWjN5hESLwQVaS2f231t0z
UVYnUXlLiPZA4DXZK4ABvy3uEgYQbjGR2V/6WXsJk9yjDc7Cn0/W14WgAvVlYDjWktev55ogkkTh
jKCTwFhLLdI9edp8n5jTT+khG9BI+J16Og1Tdw6s+C9j9SJKd0r0qR2PFqF71h8ORCKGD7cJTkRN
HuX5wsliCyToGoO04e0WxQyBp1Ji8Y+LT5hmRwe4GeABxLGSaoLEY1a0VghCTZhjz7lSkMW6FEFu
uWcEGQQ5ocKckRIsJ6e2St2QCpoIDXXmA8xBANmMMHxmktQlb0piCYKDSVkZkd5cZHda3vBg2bh8
PyovwiIxUSe2rsTcvKmHElQ6+bqIII3OXZr1x/fvycRHpwjj45jjI+tcSwf56h83zpi4kRTaYXCc
tFBoUhTAOeqee9IOTOB8qq3dTqNd5Xvz1bd8VdNpkDxa0KQCxQ+dtEfrhRAchExRP3QFg2RGqoBp
27Ssxxk8HkmuYk80fziwtAVBM6MaW/E5OknQBgsMKe3PLMwXalb/i8GGdGdijFNs3LPDc7tfU8Y7
UxaRetZ+npyTZ3Qpo+GyhZdG6i23un9xX7HCZ/Qd9BYVeGMCMEeE2qwF9ClTk9I2xk8zxdXCh7Qv
GWKpCatSj4gTTQ78WXlU+loJtOz5ZTmRNRdb5eGX6wm2uZ4UQJ3yOUhaPxMDtHXPMxwa2F9DjCE5
oE8HQPfE03VQcRBILZGODm7TNkZtIiAltx8DYHIUOPbf7qELbhllIPFH9GoiN19QCVJCVxDXxxPp
1J+6pP6LzHLsVE/rNv1fXdr0E9gFkPygiVRizgu+XfzCkrsA4zOj991Q49sMYweNGeexDA7vu+Fp
FtPIKSx5r+2kUfabiiDp5oiejrtc+SiC7/gaFrX9fwE19r7+tRjZ5Jufe1zSyjRCqAxH8x/+mACf
PGOV6m7uLn4AZ+7CGfMdXtXwbhEVwNF/BMLqaDzuyOJM+ufpaF98IBjp8dzW8enN/lUUmZ2iOo/G
z+BUhS3yXnLtBhmWH4sLQP3dcf48mXLAEUEWyVgxAQ9kKsif1pX88J624RU4lYVWlPzaLK0MepEQ
egq77hL6zd+anfbSQAqZxTaOQ5fmNlTkQXZZFP7i7vN0Mg5wCP8Oor6FLtQNkz7z3uCgeaVt0QJS
ZjWsAbLqcX4u2p2FD7y4uQo9+FrB+YpZl/fN8xWdO7UPUIKgCD8eefC54tIVAwy1aZVwgD5wXpAo
2FzgwseSnpUn9WhfQ9lhlVtvwEDZwYCPi4V090HDNA1r26MQBeJonXuaca6aGwySgmH8GLz21uaQ
vzEVGEYUned4OPbnknuuYQINk8LumVW2MvalHC/KFfzwJqYbDHfUJDQMibuOI09m/tfTA/Nj9Yad
jR+9QuemVAo5QVClrr6O+tJRhG/s9aOOpq6fW8p/cmXlTozULutnMvfIa+P/R0KWW8KAfhwwGbfb
7Xrhy7x2weztumYS5YTJ/6+kaHZwC+oDVYS3ZGmb4QeIBRDhnx3JqZDhuLMpYsJoRSI3fR+lBzqx
tN8JQD5v1QCuA6rT9VQEcu80FSYcV9oeyOtEKweHw9bNk7WECUHQMioUwXHTue+JcSMX/ZjH6rsb
WOZkylatpqLqjUcFZkBDzAxPekg6ZJZW2ycRdZHKjq9wdu5f0VjB5L5aBWanJBeCsJGb+Fdg+J6J
l4PwDOkbpZsEynsDP1kIHKkGFpLIIvl38I2VZieHULx4Rt85+jx4pepHgTYfPR/QBCbD06ncqP3p
Q1wASCIG7a2im+Sh1wdcO/efe5o7O31xJtPcRhqz3kOrVZ2mqbcr5dXMXGa7/M7KhZUigBpnVJno
oxFhhweA/x7acS2jvpxLE9OlKLlMQZ5wK2pRRTch15YAJswxKIN8W1Nw0X7Lt5aGXeViTkGFy7IS
uEyVjjAIlllmi7qc85oLmuSUMMTDaAsBLomD8yt7q8koSdXH8OwbffVN04c2IHL18l9CzFCxE+Fu
5euOTlISgooLOdICJy4iO7XnbraDiB1N2HZ/32iY5nAIp9M/vfIcdMnjYa2iKkxJh6BA/9IKn3lM
3vo2XdEQGWwWLhT4GTjUFwen/GOaGZeSvyxl1Ohc5u9RtyNQcpVnPt3mj4c+O/6W8f8gqcdEb/fT
TcAImiLK/UzB0qCnfT8BCg/xEh6V0Pq+ucJnuqe/yhlH4xDwz8W3UI++4ZwUpiOkFfR966hu0h60
W8AGgnL6D3xboKBuySzh0W+ENDAyGi+7H/GSzRxpoQ6EtGFw+pP3tgSuHvU9tP5iNOsiULgRgt3s
KMTMp2HTBE0aeX0c+u9ANOE6MvxfDL3Cwkzs7DWWkebcwnCru9lQe5QfqCK5lpZYy604xA/suorS
Lmll+m+tcIZW4Vk/XTmXb34iMkSgkMJWSI5Wpz0we2Z6h6+9AaUN/kMyRGkOjIpbBDpqCYP3gioO
02QgT93m45lSLIHZ3QUXvIVsJKOJAxrb/FvGx1b12bg7ubwZTZ0BM9+txEwzsMy8U5xL01u8YtCy
wHySksKlB+tVGAnw2UEyqMXBEWOTM9jX52z4xrpc9Tz1HlPmMezP5ma+PEEY2oeVKsXsAVex/eRo
fDZ9CHgna5TIIIiSK/vu6eIKPdxWhMOERqmE5gDvbrP9u6/wymrcNgIzjR2wt7f7xiXFZmy6qxSP
EMJFI/SaN+qusK0BUamh7gHAS3R9F9qbB01khMuUNn9xK56zAPPDJaDT6Sya0GyE0kp3gt93NQJm
Vn1es48RYHIb1KM2VF/oxsUEtTtEwbur9ySj4I9ZB1HYZIzO+NcV2u9dytV+ppWRvt9vsk3dnwx6
v4VbvnCOIeXL6ezOr7FxWaEq9/8abXTDhiw9pgx43U/5GnslZMMwJVm1tUdMO8GsIRKWBpITBBSd
IMnPUDklw0RZ2hGo3bfZ5J1WNbOGT7wNkdS9BtUAxx1BxcG3E/gZbzAJ0bKt5evEwBEpxtn8m2vz
FvLMaqNZRuVk0BpYeaYiz84kONKtG1rPy+lAL0/YPdknNOcxkPbKDhL84PkpGGYgWTSQxmJ7I2ZB
GQX+9pa9p/N1bn5fjsduupu9+vDVFlr4CllsROzV9obf9uRktO/9YLkHFgONy7Pfqi9HerrQBcPC
E+5cLdc0ivMn/aMwybvqu+ilgonPvohwZiBbKVMeiM6tJ77x9BckwoFD5+Ey5St8y8bM99HvwCeQ
mAhybqNe1I1bNFDBomcZRca1lsdbpXoO3o5sduSm0E1wbdesduXfgNAdeg5DJCNVDLbVoh8SQDmT
UFHom4AyZnpSkOFr3UsKcZ6okR/P3p2zdjzf7IkkAO5D+otdKXlOpcGTav6gGcY3Cm3jGVtQjzAR
51oIn3VTeuXY/nqKwK0WtBpemK+upiFQvKBEt03PIXhYH409lwD3eK+mlHD6lUNCw5DeUkMlNie5
fLWXouvZgK9r1jZfB5/YXh9Oca0JbOif4WeEAPENXfKUnkCeU4cCwqJabjudIQubHQCqc3YnLjiM
2/5CPd8Uf8v+ZJdJ3+47CpYuu4e7hL193xjQbHZSjGYopEpT6iv7TlZ2VxemYP9C2rLWsOPN1hDp
yc/t0OJJw/HhplZSK9ijc2oCuihXL2iGH1NLmawWm8fkyM1uekipmtDmqGB/017+x0TS8rXXrvSB
blIuh0JKxK6OOEiqdx/idX13o2UDTPorxDYOOEZ49pTXhbRP8JfByZExe1RJAMl2fX+Xx1N3k7g2
xSJPGJpqz9nRBPetAAqrnus3FA4Rt4JI/CC+juKbRkLrC2cgbGADf1MYuFxwevWHkK1G6jVg/ZhK
UPcEkhSiLqfeYptjHvIIGMvNw0czK5/iNVpKvAzNFm8seLxQl/ibw5yBLXGvFlUDG5TIScnunFMN
EXpvBAcSBnUfSGABJbrzqvTXFBK9qWtOHT98ghxXQ4EXcUVewD/7xhkZy1TlCPDm9/Mqfclhy3/3
nnZqHaEuh/u9hV+8ke+IBX/FC7yJisUTCxTlOfsRWvrLFQL30mDqVYV0tJ6mfl8nv8Y0nRdAD1Q7
vAU5Le6ae52YITpD9OU/opaWXUKbYePPZ8OSHRcXuQ3PqXn6LCQu87tXbug8fO7tymYV6Yun2EBK
UJg6nycSJ/6PfmtEIfX7WLrTpfxNnLkQQ4fsry2hHD5ZBXAiWwtfHn2eIcmJcZmtAf9FhyQCeUiv
MOji3RNdiEA+KvY6JuPgc/jl5h/TguIjsm1BoXni6wmbF4yBYOZCzK63F1sFTpRRnzoNOR5gD9RT
tWZtMpuO1ap8kU+QAnb/rh7tuo8b4dmzGXMPAfx4z8wHSLuewwKkBf1f6hvCz+PTzscs/rPnEbVC
Bq4Nza6cjlzZ/e1Uh8HVbtliVa0LfOeQCVNhTZS1ZyBJN4vBnQSNPqgPHGZfZYelqAbK8bvCf8ME
XNfDq1hQ4PHYmFjqc97iUqk0CH7+TTFWs9vS0Up8c0TyvzVRiNHSNuS0p9pxqYb4MGW1/3DlK3Gb
kaSKhIc8eCLi7T0HBmMof1LJ1fEE1u7WcqBr2TANzQNTylVzRPl61lkmnbQVL7uqBwuDxP57Bxil
poOAPaYoZjbrVGXgbH4k42dfwyQmIu/ferHpvZFfXgYSbFjjCs9ObGupKClV8LL+bQDdUmB7sqNz
du5a18ZwnePD5KEm53tu8xZoR7TPwA6BBqVT7Wd7MVxtyrx8V6I4KQYdTTDqtpaA84RVEVqsQmkk
dwEdY9/fFQrKvZXXEP+BljDu0GGHsxLCBoajNtau+jVnic2TDHsERSysMEwTUIbrbnYD6Mlmm/xc
KiaWKN5Q8LWYr0SU0vHNFZztdjyVaIhlDpG0eUD+osSqfC+t1TVrFUr2khmNcSWVOvMGXOJpWMqN
ppa54XyeSgZcoKNm8DFDxfgMHwYaEQyuI4J32IyBKR8V7cub/rL/D0OJQyi6CXxD4kgg9hXdoyXX
XNJrIbdJUpvI85czFe1TUgXV4gXOVFPX+ppuVmGwpDZAjxyLDz1Z3CCKaZBAlVVPFSA1onQnWxwC
d7ECcVY4uqL8JHwR6Kn0ap5axLdsw4IHSn0cOv0vg5nbKgRfd46S5vuUZorGtSXdWnCAUkaX+fps
TH5OQFOzD7Q9/UXITILCc1HUwqI2v78rng7YP9Bn5SLm2UNMHA7bAtPkZ+lnZW58w2m60qEQGJUf
IdZ+/uL61Lx6HAiZoBMILkNTj7uoTTk15ccEDagxDmltiMDpkNgq7frJJgWdEyQ50XTkWHj9ntoy
0MNOuseCfd2nKaiXXdFTMRTb+xol8Jx41SPathyaSeFsb42+NkCBp0FZzHZ4d8U9649jptzdDHmw
qJ/P0pg1JaW0N7wO9vS/XfBQtfRkE5NbZxMWEKhHnJRioBEMah5oApJKRQJUXIBp6uN02la/sLc6
xYy8UYKzY5VImADn7bCxk42CBNy3X4nnZQC0bEuIeAmNHyvHCCOmHCOTi7NgleHYEg9kT7tDopyy
fVVTSF3vFPwj6uPoAvI+e2P4C7xwtu0aM7oSeKJ7MEH5RrdHDxxMuJ9e5s9IYhWRsCzfAdj6M8bP
i7HMI1L7sXwIUWq8lJ9IFqN0uF+eqGEr+lGn954YLacUW5Dh0Drz4Ym2vJa9TR+xJEu13wv+1/lG
rGtOxAUdoYr9xK5ckG8eAJUh3cB0NS2YCGjdaD544/6F5PA2zH7qxtU6DQi/+LGRH7gF9W0Pw0qP
/XFdkdZyHGPPv+DLa0gaLhldTyZDVboHi9z9e9xWccbb00vGi1OglRteooK9ZQ65fEoroUVoNZto
CiCDobve2VzpegPNnhIBHVS4qtgEsHKTVSnnpwSFK+8PXQ8y75vCHlHY/IFzF/pMZEVDiLc4buxD
mviEBkrS7CEn1grq4to+MWme7bf15J4koBtH2oQA34TizPSn542DJnQkfOXB4tf2j4f2xJWVW4tT
OkIqRleg8FUrqRlg2ZEzZamlyokxY+JGme+tTTeHT50n2g/aYrwAuQ2jgQbD86Um/jTomLoxWAhf
stXG6IMHRyYNehwpHDWmE/Xe22xswcu6/X0JjekTUqJBiYcXhjC5tawPbuwJdP9x5t5OiaPcYRM2
KeIQ6956DoxCBk41mdtfkuNJ2UesQ5TUBJZZgOQ0iTzqn3hm/0m+RoWRqmLDfW5vFQC+H/MSNwaG
DJh+4RTs6DxB9YcoKWNjmB+r6Pg7nSc88P/NDXVwUfmLGvVCa1IcCyEL8YLtn86K3uorFxMAMXjt
EuLkehFqKOcPgH27H1Zp0pA9iyv8M5SQEmSb8LvJBVZYppTFs/j5saMgx0MV0FFGpCoxM3QlI0P3
swS2cDNAA1pdzLq6G3XxQO9IjlNHGC9+sYFrhdDeWHOzWkt4O1HRK0NeSPOErB2xyxQhwTnK6r3Q
dgDiNZ7yhYgw9G45JRiACz9uMjkIqkAa1TUydFhCuuZfMXiyb5O/xX3/ujgji5LpRrRgQbvutX+9
IvxD1TeL9fdPs4l36/9eq4K+QcB/8jTu5BsqRFlolr26zpYjZb9eLb7UaZCYE0IO+NCGKxTpxDyx
K+wZo6W4+EtIIMe8W1pmfpFIomV89zRxiOm/CFlVbYfu3NjWxd3aa3CQ97ID+B7J0vnzGjy3AGVd
zwOa8MqcFszIg/8MtilkZI6wrtmbfC3+QHSdFFCOZotvpkvWzKdYzfEcN6su9Zs4F6Xm6v3oSOqQ
A//89ESWLenky9KNFPsliH2W0D5rQIXa/yts2U9mcU+5J74bc+oz/gBMYN5yCwLZfT0vXp30hU4T
FBiqV62wk+P1dvYRKXBL+FDxrGPPROGwIj0AMltm0woXENmPcOYyuNUpbboZpxcWMZgmTLEqp/80
oiZSRHYyWelFee8aUuzqkkz+9AIxWQ49FyBOG9TajowmInxaDy196lfSbTx+kM22Kue3mWupJy4/
Id8MeW+mOvGIk4ma7tufOsZSv2/87RUy0HEVCuMfx8ajn6RsCwzBwG69guiZBOIur6qjP5+iWXjz
gckAvq3q6IX+Yo133cdhwYfQG44y294rnrkJuDTKWVwC1z9pQTq4dg3OlS9BCDPgAjZQB3PeELjv
nwFCGE1UI1yW1YrYNXKfxqtfzqdzMLrY5qlskMLsMuzxwVKzVk/mNwcz39jZ3WBPC9zUc8swKMjv
uqYDMqjYqagwAMI1E+rglKlSG3/tGnS+h5oR9YmRhATno+hbTkYF6JcDSrW4+PP0fUucLU2ru8rN
k3NOxAyK337hXK60pd+zwucOFJQjn/Bd/hFAzrYra2vpIC9+AAL4rQfdyNHEFVQ4C27DrBB5Aa7g
HS5W2sIIXkPGgJ4ObGU2OTTwnfuTbOWoQH8rf10G6uXOZ41eM0C3nCkrLSnS0ZTeY78cxJlCvOJX
viePIGbAmYUx5kIcr2pNIsKLl9Xs+4oZywA8iCD2x6IYiRQHMVI3WzXJrTWO/W9Cke6In7ZJNodt
EeRfqQydmlTS8ZadJ1MYRi12vcLXCU+3z0JDwxJOZoPgkvmsQXttJqrtZAqhF1D3AK6hmf3xGQLX
9h2FmjXhRiVoyyuGDiV5z6LFS14rDuNvgNhNAT2dYTcnj4JPrvGQlnU+yyfUFoCAC1m5ZaddshWk
TrToqeitWJrnTy7e5RPUx6ZCFr5soyrPpUeBKft0TI1m62n9DfoTEuLsIJfXQULI0+UacnfwLXRw
zCeVS2BKC1JVfLegYoiS0VwRd8Yr3CF71UVnMpIOLH5GAYfx+dIVe1Bqr+kVRvDRFBkvGwY4OWxz
GjxGrw2VlTDpEQfEDQP+3nzXGZP+zGklSzG0sKI1PJ2cjaKPW8gHYgUGi1vIHew+BFXmiQEegutl
kt31v982lwMAqTji+w4cSamkIJgtDm1Ji5PRK82NOkJNR+b2pQsd2G9ILH45d1b1RBjmSZnmkPiL
HMKoccfKYqCeiw6aGsy4STsDSF3jxR+OTPAVsfVz9ttg+VYaIyJEQ3A6l+u//pO3k1mWzNolqqRo
fvn6SngBHCpNV+WgbY3h/SoDuP/gXuj5Z7tgviAyhFwUsCooEmzEZ5gbB4SeiNk3mFMP1EAD10fI
F5/h9cKy/iW8dPYiqXdctf8id5vXewtbuWylSgQqcmUNAmwMtodbo8SIWbCeWj6saO5VPYql09Mc
LAlCGQUSfZrDuHjC1/B7sXSkhjMld2M7mWwzy3QNlj+EOY3jZEG0bmmaAtkHKJ4ADB1DD4mXjieM
YD/i+WsQRcI86LHg7pWS+HNcsNohcP8LXOjLnYU07x/HFhA1lFtARr0D1R+P4tK7MOK7lkkEey/B
LKAvJft+Ea0yzZw2pbBuSdN+r+XnudobTTlde+J1eJahokYZsQ0EzXYSQfsmaYqhJG6xV0GnIPbl
UMSKQsHLBGwZOjf4f17eppPqgQ2wdGiFH0JZSW4+sw+vRVUO0ma9U7Afnga3FzqNy1XAyMhYz1iA
ymNCWK+rsC6HFaajdfj5WMimBdBdLMRV+7tlw3iSaAu9o1BJEDPONz63HwCHBYngBhrY6nYp2FVA
yvMwt2Iy6sYDsdQEfxgve+w3xcBjmzBUYVFv77NP9BuE8MtI2IGWIJ8td/gUiMy3NCkbQIX8a0WQ
jND5QAp0rla0SDv1PlvjF7zHtgKz+MmoehbFep9VIMm4l3MsmOoHECLZACgswNmBuMnqfKLO2lYX
ah3021Tg74OfBLHjVx3sS2FGPZk7E4WxcHqQPPNANIs8ia3DDsA2zxNTqe95+snT7vcyrI8+8+4J
jtS5BBEOeIQ2OM8p85RP7upFJx0yHeZXy8hzuNBXt93Asot3E8KstHcM5iq1EWgJJKt2VP9/iH3Y
3T4aLdq60ZJfTvDvNxhO4/2iCqrdp85y0r5dtj1zv58r1NNKgyt3ht/OA0nC/41tz7rwEpciM/Yd
gmumgOtlA6LFEk1LhhfSUxad6gSspO3m/hAlq//Xph4oufVJfTndbNWjjlYyNFrOVUDu3W3RdBdx
1gPFaNd0m60HePBQfnF0J/6RCIcY6BoAgpq4uE8sdLtmC8Kr1+7GLHkNFOBbQgwBwdxEsAdi92ES
xKqWpIWHYR1xk5EmMPFk6mQiu+8ruFufR8b+EQlI8uQAH2Xu7MP0LMR5XgkP/g80I1W31TnQkT2O
lB97hThtsbecvidUUiq9KJmGLTNAVmeGqc/r6Zg4UN//1md1gAcGTynQ7kJb+JhsXb2XenxkMyg/
R+YzV8L8aYlDV5ZYbx1jDO4KdA8vD6xfXy+pSjbXi+VJ8umjU1q5WRCrH0+h+mhPVKESKNAGbOiL
g0Zc0EVgNmNqwu4suRDTSEnt2OtObi2F8wu80qxECbbztLlAG7jRwbqHSbTjVfPbfMOehdSr7oc7
u5xqQvLTHymd5Vg8wMpGjLhQjB04XzZ0nMEKm8HvfBf8AhGZRAn5ejPkczTERtIFfJxUy8G8pUsx
VZtzpNuHcHV8a0U/VJcRdUu2O19YIRHK4PqeJdnfUH78LRq0Y+SCNYsIaIDASCP/Iw2JMnEBF+Dx
U7g/IPPHSLdYrY/chFksJYNZ4/GTJDomXSiAjP3EGcPveoT4YvrzBaIiKH14jr/ThyyrEBts0ccf
ivJ7lgt/7J31QTMF/MfyO13lW0PWGIPM1DuJx9QtxPW434L6xgNdKh+gmEoIK0sc4Bv+fc5+F9UG
kktEZf1qCrnR76FwyagvUnBN47swJ5SgxCOIdZ97YakOVI1eQ/FjC6lCYEAbOZN06lxumHDn1foW
TDzuV0G1pZqwgpvl1AOGmVE9ne16PTQSOwLF2aUHennyLD3RbqqPEkX6znhgeY+K6Py/Zb9m7Dtx
AYtytgUWQF8sEgZoWDw9E1OIbcxDDwZTsZx/9jUPmx4h5xaXb8bCQ9kNjG9AN7dhyvY+ekjF/fVV
quc2LNJN58SuBLy4qYJbdEP9zgTgg9cl08SFQoKN7bVzKN4eA5/WeDNpI/e/VJK1xct36TJmy2wH
1taTDyEvro5InzFL5fH91gQ38AsQIVi0czGCeERQN0WsWmQd7IZTfIWNLAlSuNIdTtbQi7eEGl/W
x261OPEqZbKA8g2L0Draid40s6zZgNV0cD/diSsFXYhJVNZRq6Operp1uS9NYOTx5RkR62kG+AS/
OG+GD3/uOebX4kfwByTHqlL4yYZzlBifcyH+5xa862lyy9iKsGrJAPlcBLXLJ3c+q1MfVOFBrV4x
JifjvzzMmMD+rnWHcKF6Q3UiFfkzaclxYyzjlfOftz6wO5EfOenFnlaFjCg3OrJmXwyq82PkbOEP
c18JQl1Wib7IF3DjX8sf4EXQtP+98TFj6ZaudBr232eqdDvu9yiIFh/hMULm/vhpo6hyLaxeRPZB
2SLJqpdZI6IfByISOrSsfGwO45qRloxjtsumIDV/aFOhIiaQ2zJ6T1R8xoD1qpn4FWN2zWF1mYzJ
AAcUOCTm6R7Pc1pbOLv2XvaO2unCMYh/o5Xa+0GMiNHAyxF63vhaLAG8VXUAnrn7B8sldQYECsut
zPBQGrdK5fZ/pq3MyXuPkIODn7A30z46aeS1KVRgpu13UImCOzqCkCV9t1CeyO9goBuNfzV0Sgyk
r0J0OwpKF1JpnyXPblYODu32HEvfxTk8iUvAJMUsY9ae1nfGxd7apQcARtQ3KUVYkdJUw2XXO27k
yrv2BtejvJsVE4JS4m3tdpH5p5i4ITWbHsm02cApFy2bP6ACLllKS9DMBBcYsi2N3rr2HIDJLRTQ
jN2a3z6tCYE+93IUSjPzHX6liCllo6GEwo61LEfZEh9ernxng5+U9zg8/1r0B5qkWd3Muge2DSyx
sMGyF8Gs0US9yuImDB2c2iMzSZqhdnaEiGGSRNlgjxeXoZQTyJyXQXlod2x9JScLQ9+MV+BOaBhA
hMv+m245Gg4wxZjxAc0axx0T5Zqok3c6eOc9bs6n0808ASBnthLtraAFq57BkeIR7gpRdXycM7vi
aVNbHOJDkxstwY8zqs68Gj5OSYZB6e3Fx6ZGw82EahFL0oIC+gLk5MsAGXuTuy1ljrtSEy47FAjl
Ae8y9wvODL4kjR6K7JDitbYCoDPzIGySNh8CWBoWQPxqvp1VMSk0h+THw/+GRQIoJnZvXBfmJuVA
zg4epyw4DW+L/0TorSuW64jzYntQsNi7d6lrZS/A58drXy8wmFprN/1pa7ECIwzUbKqUdPI4jrZE
6QU3L1Gc75WP4MNC5+8bDZKdC8M943Gfv6npv4t3zmqPt2FlZylVLA3LFTMM/0npk7yEihS+u119
sKrNnZk8rFFHu5Uq8cWexgkYpV2W+YNyICeahJwJlpCheZz59WwiC6ivsFfdy22P0NrWCdwnC7sa
jNs9k4GLquaQ0o/LPb/JW98B4rxTpBGsD2Rwa48s97v57oIYmqi6wFIazSzX2h7trRP5qGp290fh
lL7M60c3SbO/n5dhVRCark0/l0amRxxEjD926wnhp+4RyXf9QFNZwPhLROqoDfrf9Sd0GhD5KJH3
coX1G9Zmysctl37uOg1GNTwJUI6YJai904XDgjwOiYQh9w5Lhf7DqrU3EPG2aoEqcGe68kr7gUO7
n6kOzBBHjdbxUFXEZixH2eAyUhncrXpZvIosgg58wstYA0Ntmvmd0d5mOmYCNnkQFPkh/lkY6tJg
MeYooURezDly7pKNJsxr9NC36G/6fMae4QcNBoeuIh9M1NK19GAP9k8VikAGRO4sZQE5Dsh3FecM
dmbDMvv9EFqRzAXSzJQ9rXdmsnW1gWtIjnKHUfk8zwL/XQTyrV3cHW3YAUZz2LzDhYPjPDEkU60i
16+CbUpErrPc+i0xODLPjcTdz1cbY5aWdE3mPX+ZLc4z4UOjv5JN3NAb6g37q/aQncH1XKrw+yma
6D49GApvN+P07KrjYRIOi+rAT4JmAsT8G/CdnMHlSEqEkZ8NlHRsRayuHBqtFuT6zKZ1iAKIXpsv
60NErfbhJ0EnEE/+MPrcEId9aXMBzyrDL1b2K+jDb1kzHOOYhmYoFx1KyyN9l3kEoDjtqlpjCX1V
uma0r3vmsdjxlgFODerDZ7GePWz8eGedEdtCSoVS5MiVk3Nky1yTWoyp+TBvmz7X1CSJBpYEmz+3
/rY1V4cP5ymaVU9ic+P/zA9nFh0N9tQl1bq/6KkcDPJ6fUaLHIP3gpV5N2hpT67Pc+//gJdgVG8a
S3buGgUYTbcyuhzX+YsSv/XhbIGXK1j+6163oUAgqQ8L6HbJsnV4DGUn5d26XKA2RDz76SXYVaH3
bEwoXqPupAGYJsnu2XlOvYsVE2U4snNeiIjPAtKXmrqpHokRR+PJRPk4YFdl5uiqZTJs1MVMcli1
CsaBTo/VuOKh2PKdccizV0SplfIxV1lhJaA/8nU/7Gb3PWtSpG6fYg1+QCNC98WsZHO8isI8ZTZq
bGE+zdm2Bz2hkXN8uT/ca3MlvaBrFxCnceXVfFGcK2yaPlZcZqWjg3cwxA4LdfHDUocIKEkTISpF
jFe+8+D+kdkhVU77fqOHCP6+Nd20r8uB9T4hZ/2Azs/Ja0/EDfllnucnUnrwBWEnTc6C5s8Resx3
Db7b9H/UYods6QH0FX32MkyHUlLX157YqAjvXfaVW4ZzZdsnERQgbocsRBGpU2DE5/hHpBkW+u+m
S+i18s5WNfh2PNjHG1LQSCpXcrFLqEevvsldHGt1uf9giVjOU5u111nN5r0MeM6xRDDyxqjaW42Z
zBCgPDIoltSl46YtsXHgLSueO4Y7lNhs1J26vdEFrCPcxNl50jUfvV/vADfAUtwZ6v637F9/nQWM
/eHPpq1+HxAlWLJL6+Uq2H0J1+/CF6UKpJv+513MWUwwdaD/jOOk2bbDOmtijzLyypnbcsXc3W2A
YzoxW2P1R4TiRCnlaCIP8bqoXhhFE54PCuOt5Qj/KYvCKS7Gk3DMvuzfHgAG4Our8yiHEKHJnYgo
lmq8W8UXZDFZuTVbb//JmjXSSfO7kHa6dwmoDg08IKTO5OjLoTY2Mm8agYMD/Qh4Roo8zNwcogd9
6Hk9TqQ1BoyvVSxhxu01zsfOngZ4schAzMqAbVfkko1igv2C+N3fYXcDNbQunJZ2oXMh9hBBaogD
HHz5g8SOmkvkYLiKhcJcupGBTCBW+JXYEt4UVTV0Wg+Jssj1cPpFwOgutyWeSWONAVg2Ma2LJE51
9tUqWxUktkdBLJpSg+fNWpKQ9A5F+LVGZJQq55B1n5kGzWbCeAbt6Af9hX5/ZNhiM0N87R/vEjuv
SNZKJlWdSMs0ZHl6gofA6e024H7wxkhDow4kFEfcahqA4bjCqZly3+rTIVq/5ItQt/aYj33vF1Qd
o9WB6hhPu3iTpXJobqmxJnunMD4M7CpZbHLosHaVvWLMeX20JnDpgxJI9qzymcVlORdxcApQyLU3
s8rpLXnZ+W3ETXVaz8BRSXc5LtRU7/MRfTwUj6niJy90vzIolIdUIkK1W4N567RGQv3yyeyyVK6U
8eiQVkPJjSgs1dT26P/K0fXZCN+3Fr8U1jF+4Zs7jrByCSqx1xW0b8HFIfY+NlmQ3bBCBg5mSDag
HOMjBQwkDTGzU/wyUZQ1BTi6rDlBHVwcZyWTwLzQOiTaUSbnSxAFxLbCgzPdXD2r+sne6AGfxPdW
K56xPSywpHZ3xUVyl7K4eksIGym67Ys4O6BQNEqTfXmEtHySSDeM/XNBAPfmlxd4WZ3maeJ992Zd
KAGIvXhBZ4r+SxayPcE7ifr3o0PWyA3t64ttsT59UGrGVlXC8DdgDPa/4BZVEUzD6GshzTPut8pw
JAcfRC2sm9KiJMZt1a63pi5U1aEuxWumoZ9Hs4bIuf7IM5wdYXmorjRkr0YscbgZmpm8lf1+0rm5
hYmLssST6DXJegR/iUBpuGMEfXwlkVQXAq0uz2XV0TOzWvwFgcptRdDQjolX8aWhT9DFanjDSfBp
olqCFbmLxa1Ak2smmYq7mLcIHlSJ1g7bUdwBLkNbL7t2SjDPCBFWwf2ZCCkuw6XNC2Q7rcZJ2RVD
87ty04UUKZ01tw2cKY+KnCXk2oz3c0vte1/cbs93RI/AAPnthMhl4S5pk01OJJV52+4DZBJ6BifW
B5tv+UlAHxT3pBwVxdNbSYxNssTP8XiR/AaR9CVIf0Z6DX5OP6rT8PhUI02jufN1XgsXmuN30DCi
MpvyHYNSeVYr99iFR6KFRmH1yFKoQvbtiQmNnV59uYJr0Qn7b4qZhs/WWJbexC+3wUTXeH1RXC62
2dd4UmgxdWyxubjulDIBSeWz0CybWI7Z2s1M9imA3pPLBu6e9W0M8xzYxwtPtT5S79noShUNiTOY
ouXGwI2MNGvIVmMVXFh5mVPev7dywKlYJxwFfch2J/8E+KfO2Y3e6FhfyLzKV0F2dsmsw9LdILdr
9GFK+x79EcX0OwAp1SgxoaPrIcz2AuYPRhWIRh3eVp9VWBFLQmWfbERbXuiO6qt4xtnzoO7Tof2K
m4BHmoa3TS9K+Q2njBwWjwyPPl5XLotQJTtLi33ySD9v6yW/E+T9oiYVUlautDVU1DoOENfL2uQL
sa/doP7G9+aS4U7wlJBPCGS0sEnn7jr8rnvxueS3VczADZxWnA18SxlZHccMQmCwhR90FivCtbXJ
08/HdlepdAd9WbNUsl28+hQ0pv5vQGtH0Bhf2IIGXJJG6G7gMaKS9JoyGbaPBeAWTlm+A3SSQD83
c41w6Q9mWfBGCNFooqZMxvGXueuqIw+YXm41+/9kog/QXL47F21oQWdZJLLu+KMF87NLoU060aVw
cn2bEn1HsR31uCGmhKMb/FihZcaffArqCjItNcDPwxHHTYpJCevRUvPWhn0EOVLDmUURiJ2o58Fr
FQgNkiRVgcWSUg/07vki++6OOK96Q5OPx50pP31QgAmeUY9qv5gBa+/vfzWSs+a4NsFps+jJ9prQ
GuS85nYm21J48c2jhKO6zWGAS/EqZja+zjzGnG4snu5UiJ6AlvMiDvNG2rNnBaAYTrHOQThp0Aks
h5yJ/5lPYgsHNYGvV4jQYIVAcX1A8gIT+oH9rnW/PT0aCVZrfh6FzIOvxhbmWlFUMucwJG5kcfQ4
gGiBUyLrSNpeGjXw1JPZB3/2gXZTgH5rRrKnt6yNdar58B/orlGeq76DcxGQzkdPA3ubJGUWDk+X
dpmLe0QYTr+i/C8PBsznj3ias+R50vnGURFkuZTsG+Vn/80sATu3LundUP7KEdi0YH3OWewKrGMI
1Cs0pFLK5IeewD+OsHVJH1I7UxR3KfQ8jL9h9RMaSfJeh45y7rZ4WpFnpEQO2GWdphxoA/y/aMwx
J96yYa8VW0n4pauQ1vCNNIu1d+OXWnM9VYj6z04lFgZjDAE38ehvVrZK3mmQ8dIGMzugAdRgxPrh
JDiDhO6TOOhLeoivxRnJ06xaEeKJc21lzsp8N8ArKgHb2ARQDbBxJ3hudmKmILaogVzJQZFg6vfa
XiofM6LweOlYGASx8PnnfRNFmdX45wYkCf9WHJotnjgQszAeaVKAdGvzkMHA+up9Mw9fSLLI/TES
MKZ8VMGPb4lTOzUjqwX/h/VJVPz9Nc+yye9G2Jm6xkMdQNbBigsbH5yxKPPvfLsgydG4qxWm6oWI
7+xpiT/lpprFQtcUn69ywd1rEGiUbgZuKB6b84f+qDsIOsEfZhCVQiHQa7Mcn7ok6zVcRe+jVyn4
lf4eWPuEUHgq/U6JmqXuzWln0pRd+ExnNBIjnbTG67l2yr2J7jHsH7AbHGYJjLnvhsh6EkEAi35u
A7Np2bP/9Dr1l9cLVRPxTQuzJ8rO1xpP0CV+O+pA/HTt1jn0oxgZ/VVORoIpJm8K0ZpZTa3eenM0
zVspc8Hr4kek+HnGmZk5ir5JMaMJlGg3jJlKS3U0nyV8bQ1DxPukifnjpvlcSlZHbiAX6Tj6dQgm
ixygFEZNWB4Piyd6ZSxhwDgqxgjkIhYvP1HKmLUn6ZLRWU/hLnv3T4hbMICI9e0Ityrdeqs967my
m/LRqG/htZzajph4aiUcHVYM1auc9yFUWEWS3mp72jBJEgTh4Wd4tummm4zl0q/VulUjv9MFjc0Y
Zt9x7xAyCxKeKM4g5G9ZKGM/e0B0zQPfGqX8gi4qKg4Z1GHFnD5wJeCRCM+IyNmlnC0/RDYxYYsC
kbzI7lNnHDw3oNYB4c2BWJXPJs7wsXyqPordCCaMlfCLJzDlXyuMnx9B47iw18BqL7OWQVRWhu/h
8us1pnmx43eXFTqU0wRHdl4HaRHdTCVhgH/Qp6t50uwkuuooMJTSR86w9xeGAJ8V6DmMYjkp4ueQ
sg5ehPKg0IZ/t5O8OP7PZiSy/qcPlXE//xJmAhLxDwRvxD6ndJhEEq4x1S2OB17IvPgWZ9HoabuH
W3RW3mIgZsKXMEBSTiMfZjm4lC68uY65B9VHxXWclGZd4J3WiaqhFtCBZNiAU/oNEuJL1XCq4h7O
255OByGXW4eZNi2eL0aE49pgFkrXvccDcSwdxdyBpzSZefTzKTkjGL+g8Fnm8BvH/p91WgQAj3ky
saGPfcdoYPbpP0cQ/PnmuIgUKSajgwhxKkgrmOrc2N798TCQz5Z32ThmQCFMWZuoce6B1aMhfSTw
qSAAk52f/351ZG2XFgTv368phMDlXS5+++H9qPbJCFTXOyEY1FMwxSs+jWHc61JDNvz/2hXixRx+
s6qApbkypaQVji5ndz0SPsnrksZ8VTWDSrlG8zOdR5EaasfOREWEgYieZHWjWTuHDJu2EGQHRn99
rzM/JfxSPUV6f6BroY/RktfkEL72XICwrPBSKq/fulChi57SQByUVLAnhaqsOWarKc2ZMc8Zk3Z1
7MhTqFISE449ixVyimKXk40Sa5bP3wu3pkFHdSdvUj+tYbUB1ZnnrSi/x38nspsQp29km4irlQMl
soatmKrbbp3cF/Dq2ISRTEla1v6vutwtp86MjJyrt6C3TWDkQ2+2vCkN0wAHnOhgjz8ZZRo/5EW9
5Hkw9AcZ1Tz+hqWJWTQYhbImaC0s1xiT910I0LMeZ7OnELQnbzJHxXPltoolDUDB/6lF8HTfeUTp
D6y2xifWsz+OoPdNDdRQunFn+Fs/UUlytcksF+bSBQLbHjmfvVVetwQrYszhcmx1nvIxMtcQspGU
uftLt4iFKa9n+CFD0yHE/2h3u3jMVGbGgA0whgFgI6pyZ7/ijvWCE1DxEYv/CWfa5zm80J9Jay8J
+kx8E3Q3TEcIt6dpbsRdphzhgmpZ1f6/hiD6bXTGXcCWupDZ/y0IYQRHKsGkxQq1SQv4Xf6uxsd9
ab/auuKcfn/REOnI2NvHgrnUa6+7fhi1kDecqWUkKVXd01jd63WK0z6lx7XEvC+JUSfnrtmWX/te
zI0EHWOxO5iB9BmfSUse/Pa41gguZifbYmCANPs1zhVtDMaoTO3upBubwVv7L4KVhKXO/ruNhHrL
yaZDPcINT/8el0iMpOHuSXmuVxfwIQDRjSwkNMelTSw1O1PRnmCkKjA+o5qJrdSOuMoYJ5imFzj1
qDMO0nWje9YX9KkSNLLEkRKwvORUEzsZycp8eoEW738MWGThoA1O/kEw+ff9Boqr4nYML20RTE+G
2yTCfwwuPLAnH7N7uk3rGGCpiDw55iwbELHRzNnmAjjiJPdCn50qzCoQAibnMkLYxpMYGy5z7aNf
XefRynl+v5HFfPysDoV15jg7xPHeJAj+1A3uRroys+YKcxqYl1n4esV1r2PuhE2my9MBfn5QcQrx
muAXGQc+e9+uSXvi4xorgUwSY9wQXSq+nLZrC4slIJy9xBANXj5RmlJ4x4Hbqs2nsLhNwcCy9Gkb
nyRKIA3HoUes6gFID19WfNEs6rfvwA38vs8GPyOgK8fpuZF61zoA8RBiSb3UAZdTiGMXmNikpWxw
U2zDcMyk7D2Faz/bcdfa0vZU2CmWcdJDfsiejHBwM7VRUrFWOOtvFFa1VJ5eUb4FNBiYGlrflkm0
SamLkm8YwWop6L5zv/sj205bRzsLy9kyMZtTAuVzNE3w0voC7WM9/I6sT7w4Cl19vWdFG8Nvdv4p
xuJIo5gWt0DWi04SjReHEvAd+RA44usPIqYW6ZkpF/Hr3Hpv0e+GnNHHjOvaF5Jo2bGOClGzGzHU
ZOo65ksJHa3qe2B57wYgiEjI1i7GL18kLWil9pIRfkxE/seDUs3w00oYEo0s8SwxLATEuK1gGuo/
YFpKNVgqDtADaHDNWSjVnrpmmWxu/AYqPqe/JovO6VhVsoADuLvzhzj7y3RaErwwIvh++Qc4SQOx
zxvdweY9x3DuvhVI36lfOak/3mrVzc798qzqhPOMDOnVtg+7bOQJxO3II3dwHCxNYE7msExn5zsv
p0294uflXYYiL3ChBkocUtxDsOomDwpb27ijVSkC8kQ2oUofwCfe4R7rLo4XMHTfdeQ2cvWotxXS
iykrkOZxbL4o/sVyagDF3JvzscurMrspAo1RtJgpoZ5bNRzUxPfa/uG7oL/sFcohtkHUd3eR97Mj
oaFFFXVUZROl4aXX0nsfrlNy+WaqGGUpn0AA5P1imRnfCn70+1dtych4M7pIgb66VPs2N9L86a2m
/kLDHcik4jJVMpNH7ASVSCqmyClOybkRL/9dBAvcPMnlr35XYD9pcwciY1tIp0zWLy1qEPEd9ufr
XK/vtb4V5XWcma09ilTMx4CXwakr3OxhAko5iHZQj2VRFHObgPRGXJQl78t4QP2aPaSMUGqUJqu4
a6A8jO+Y7GJkDJVvq59QzbkIUlLPFAkABKmxi/7tzEZnTcYc6WHbqorbSCDreuggHn+5uL/KE/oH
SYkT1MY4t8NbpMDL8yp5VSMZqSnYfVtS8HWVH2r3X7b913R/gee7pG9SJ4u86BAi4n0Bgyp4G1ug
JicnSu5dH49SZbbi4uExqYV9aUuQHC8bai9UfsOvc3+dIFi15S19pRmxKpO1Kj7W3GMZhqXJvRUF
Fsbpm1vg54P4kHGj0snD4HVuDa1XDTaHGEsyc/tz2I1HWN7X04uN6pNXg276P5KtHt/GgDDaQrjo
jQ6Hzup08g5wkwFeN3pJ4n9tHkkVkaMUgTBhgrCivsrY3T0G4VoqOdKYHF2uJ0Lu1Zjyw1VTM28n
NWfFWMZ+fG15BS6XS4eaj0vzeBbyz2XoK42xNXrTLB9KmwQ73FnkmFQ9FqETFWAcGPtnrY0jPJsj
sfILI/IyUnwdfKxJf+ce+4VyOBb/zmcKf89Eo2lS3zV43ZgpHXvMPD3xOhEn1CRjCuZSZjiQ664z
EzO+wfTUhDG8iBeZ9jhmkzjyr4JSDCa3xm0tsut7L0+4QSvm6zAXBHK6+LVCCVCNb6E11TTJ1rZq
FVSnihKY726QvrmXh2JeUNssEIsCJmajsQCgzNqC7Qtkgsg3HKWY99p1TtK6oJa1rBYmrJFZOvlH
q6mXVxl6NThdXocVYzXQ9YHj2WTedQoeejlM2uZ0D02glSFBBTPL/K36Ljj+fCHqQG9r0odmcJ1e
7i1AXsC5aa6CAG3riYy5Ze1XScK0HKZqeFlBA/OtDrP2ohQMQYPMrET8Q76wDZ5FUdIKmQogFem6
FyDcJFHV7Lj5OCFELVai91CJhGcxNF3wKcpTDYj9yqw+xjbIxAWVVXkEfL0Miw8fqDMdVSaPkeG3
u670s96ctbLQuP3dc1DmgEUiVyOn/Vy5ELEx6GMh/hkUQ8SMxWNreQYtOiRMGCnXCAFMldbOU0Hp
B2pbhDDmdesLIRklkaITgVha2sIJipQIgYlieKz4hEMyULobCeZZJrp15PZQEwhNFaPeewOeX/Wy
4qyyljZBK0XSQXROOmM4J7x651LVx5zN5Fd7/L5Zlm8sj8gDJBJIFNo6GCHTlHvo5IAMybN7ftyy
C/vHzyoKfZ7g8h6nHqT0lkOd0DWUDCObefE/bAGmxj2r2RJc0AhWOB9VUHtDyjFC6Q16wXVHrg6/
mQ3vO8beWj8zLhlNpYIj996dciqbuoyu83eP7oS0ntHzUcU/MFfyUqfvG8e/jKDAuHkDeh7UxDxd
k20ettXDlkW6NOZY4XxYQvfGVX2zvMh+MOGyqyjT6TC+ZGwpEb4bd/k5euNbszEFGvVp9q9d2JDv
LuhDS3f5c52yNsT1sCQnZq1VYKHSArOKy50YlzrUXOz5ZvilFklBV8aP+byhKSKm99nDM7//BOuq
fWPOw/LZg9ct41/MMddwxfsewtDrxTO4vzjrcOPHlSmEJERbENubai4QGDi4bFKmT9PpKcq5zL9X
OjYL42rPVviIzmP1dXd/At63wojlyrz23V6+tbt4SojDvC3hkCG6AcJRVQAQw5iA3SOwxutt2a+P
E/Bzu6QYbC6t8GOXgrSNMAkXepQzPgSqax9p3DFvLlX1QaM8uEkfD28iLujz//0mTlnSFPeEW75k
mygyTiLyMEckkt36bj9L5gV5j4J//G2SwOLcYAbtPchoICSuQDh5LQB/tVtK+JWlY8JEnOybo2tE
igdeTPTWVTjXNqvXn2NzioaeKP2Q8VVrhlxuV6UojYR/iOCvSa+5ERNPSjWSwbjPFpqNnoyeUXl7
ogSTYDw89Wv++7SkAJKVoR11393Hrd9UhMk5/ZXz1oijZB7A2s6yTekhfrHGQHvJCJPU/tjE99Md
oVM349KEJeNBfNUCUb3VvQntL5H94372HMLc36Hteg1WkMm2c+ddAjopqS05f7MZW9ZwJa78OVl0
EyLLt+PZZmC88PNlqZSt6hEDBwFz/BqFvdbQ1aXxz1sy0hW574rEh3vGhmMaMvC+DYp9S/Jc5XZB
BHRO5Y5y2MiUQzdEdaP+i8t4VxcMCrkYeK9rGmfr4lMUN1xVgMe/Sz40WuYKlnf6gr7dof1ePw0W
joEq5xOmyLdyWXZAsGm0PGsPPVkxTuguR1Bi7bz03pE6/5T0vnGHVJqMoGc9NqJxkop3vSV6keG0
qfItrYtHypP8makVr2Iy+7/OMQGUTDqewl8OKKxVWK21afAa18lML+dNsdfgVI+w+XqVSkPv1FxF
4KdNYdT75LOlCTTj5MrYmj+lms1IiUds32n/jKt/waQtwHDhZ2pGXPeOif8uZ8JTtVCr9GpAm3t/
wKD/jjTzGonOfN4+fgfeWvpMj2yK08xCyZSQAsQ+U9WzyZwOBRlvpRqV9f1vCJ1KTuSnZNI3kdB1
jz3q9o6O+k9oFoSa5zrf44+bIZ0KJMppRjyfnixaQ3GOMuwS3Mkj+RpAhivJQNjOs6cH5FSJil99
FU/LqaiXnH2mtaZj51pN4Dai/iS2vuSEyexttxR7wWPHkxsR9sPSlGnBDkSElyxc9IP5G1v+D7hm
PMTbtMoH6osM4vL9LWymg9Asn0FF0HQqB+3J/Q9JOLlICKCCdL+n957Ax/O9dMpac/rfGjL/g+dm
E2X+GVZTPnGTbCA8JWKTTaYeIKOC8dqKwrqsyKOfxTwKbsbD8rGDmFHaq4V0gnPlYzv8aCuHQQcG
ctwl2xDZb7DX4NnK/RRop1TVLbL4++E1orqo1D6j2uyYjZ3LqAsgrdwh004YeU6U2IMfdRqM1m97
WbdvHmfD3Ag8/aNVKmIT068vkOS9mh6Nb4iPJu0LvU9T9HW4778KTofj/Gn89UuFvkZaKZf3QZ93
qA7Xs7n4d2uii4QgmFpnIZDxqKxnwqaTUYhsCrbnys1xIIb3cCfHf6zHblOFnRnn7qrvIa9lBp7E
VSZqSfZbzr5ynL0cr2IpNyFOPtFu+7895HXEJnTqtaofL5+gkgRshsf+HMbGKf6fSjTdVJ5fM0mr
tHpg5Cv8tBOR3GKrT+JE68GdP0b5QjRJ4lJ68Gaq2j7c059KCj6BMqwERyytF6hE5MBE7sTrDNkx
coLW8nTwNAY8YIF8G1wH+9S8/xHucNYcbnwtLdGQzKal+6DJrJBz1hhKfL0k1ZW3nht/jTPnPabE
CXsb6Ah5QETIBNVtgayzbX88WCV2ymET0AmW8pMUll7n3f0Wml4MeINrNwqgzcz5dfZkssA5NCXu
mY+FOU4MYkz4ruPwI6S2zzMwxj71GfaJc5fh/UCOhC5sE2kAD9TMFtAcpaZR08P3TmIyO0gYHtWq
mCyhaJNam5VM9cjOZSHkRb0WhRMuOMY8RcOJ7bm+XrCogJa0fSM2WE/LFmWF8fifsJL/w8+yBqQe
e6I8/c+4iXWbCCOy/9kzWS/++bFZ0+bsiB49NH0oDTdhLO4xzl7bsvziS5ZAhDcC1xIdLAvmea4X
M7Jwgvm3r5u+zVwlyfeW3ZA/ByZXndVmyXAuEvBxPq3EJ2kYwAKUMabGE5CI5/5BGAbmcgryqoYg
28dKucYljjVmonzNEqQ0Fz+UDf2kwq42XYuaBUCXLzCNebygTI8UPOz2aDwarvnfkDZD3+onIj3e
jdgfE6v8Bj/gebTrAbQK2EUJJ4jd7f+E53tFkbbys6BsRWHBx5+JRLNeoTvUpkT2WYwQEQeNeoqB
Djqao2azJF8CWzXhya1AzE/RTuCvnnFoKSJLn4wjMNwI6qHH26Vamjm24IC8rQqcDvFK8PgFMxyd
EzFi6YnuhC+w5vcVbE9bXSKlWDicSiE45+0kMmDeXbfq5wcyRo4z8/O7LDjerkHXIfU+UqZi3Naw
ZeL3uwYKoUZJ0J4T16bwwtPUOd+iNOhMGfY/neaAqsJBtmFFW0C+96oFHrFYRPUAm1k8PYiNSqVz
M2E8RupyNXa+g8GI4/Xayvf3KoEYx2n6S9gCzR2j/y2V7M6SyeSO2ybhdWSiACyIUxPME0GgTE6P
+P3Fe+hHAAVEQPiCJCTpqqGsWQf0CTyeKRQUW6tNrDB5pGQawpvDTFrEj2GE8OV6oRkN73c7kKwN
I6fzgSILj4mc8VyBvCVjGH0a7cwqnrYmzAZYUumSvMkluYMAKDRxODgRIZLStyv62KFHopa22YUF
vBQ46K3voeoR9V2K4/8jqWYCuBF2EylAKzBi43IIzzn4XvsmU4s9Rl4xJxR7Y7UFs6Z+blvoUmi+
8QzS3m02WnljJ79gY9S8Rmar41H2P44cQiR1Tl5yuwvgcqyL7ICd5FIVCyUlCG2LWp5yn1TPfvqy
O13q/Ub81MEln6BsSXQhDiNHE+oCX/ZiUWMdVBMiQCv9aEtcQH4QIlIi6yF52V6JlHD17Lbuh5Sl
hUvAXZBGdqzP8R5S9rAAWC+RDZURqie/i5etBs3uTI1B49aLlXH5nYuhg0Iwf3JJZyUxkhjvOwiT
H6iKed4miOjlx1Guzd9aMxxiCJyzS/3Jd6Y4vkNgGsCJGkU6bOj7LaD8eAw/GqpWkbW0G5zgNicq
pPd13+sPj/scJWtjNdoSSTWmT5poza5g/iudFggeDpGCfvcnThos0a+t9GZwHiTzJsRmxi+Cljtz
XE2pCLzHx0j26uRxT/IkCy8wQOlLW9DN5oDmK7fYjuxP5L+ZTQQgs8k8F3WN5r44DdLt0zs9HYFu
yp4J04c/R77BVQXE87eS6j2ukn6Gt2TM8ALXTTsgPe3F70V9qleumZNBihWteQUqtcVcCUDKrbOu
/LIN5IIRBJ2H126kGVOIUMWEcWpPpTVyfevnf2f9M8o3tfVFjz4FRSQ3y08Jc1kc43GS/5+7B11F
3STD4J8QOm2lIhbQVCnJOn2eWoV4kwjmvAQt7qm8YaqiQ/DVEzyQ69lsLnT8yYrzSyY6XCaqECQu
9a9v4t71Bx2AFr3WR9TYcHWep3pZ+CWLB8mgkjgHnqCmLx9nlOy3hHduVLDssYXLTTqrSdSCnn6o
PyI3oAeokShIcmVdZwC1omTAtGzjBYJ6GkGnojdK2VNuypE+GiPy8AKTs/U8NFksYC4dR8MSI3os
Y4C3o2gDEU6j/cVMiUeqlyN6zsHp7JHOQZrbeQeDgfnoN/Z6vBA5cpkLWgbxFQRtHuIAzkcP5ANs
FS6w2Ps7Xp/rNM5iPkNgMKqv+IGMXGzeGq72XRn/uPt6FHKFLF59KGgRPQWuYf6T+Do00pISp+Bw
lyC7H8z/wEjk+AmOmGbrD1RSs2RxLvv7189HGGpHT6tYEO4xebSU0ECgx8FZf7KFMq7hsWd92Mn4
A+7w5aIEJIwZ0Q096HEP7RyWoej1RnM9z80NXfpdg0KhZK9ZBP9vxC/VtY/kIlPpYwMpdUGxdZoT
FSp55878Ph0gdHaoe72iV37Z6iUFipMqMlAgfjf9d1syqKimz3gzC3hSUoCFkzn0I4s4AyKkv2pw
XRjuRJtrDrKKhNFc+BGoU8cbOCOsh2Pp05fP3WFFN9AKYXd1AlLrPt0W8Lztz1v5J+rMTb88709h
RrKkq8j8Ewf+naUTkIgzJco/7MSanZLrQPMq5pzINHSCX4NsVIWzUb+GMFRMt/WJsDjXzbsLGmdX
Ne2nB651nXtOFDaY/nBo/qVe3S0Ykuqi8r+fLNzTvWy1GsaQPzBVmzMNlcXgiyzm1E8JJvYvlde2
hsZ840QhnPwTZNBlMRHCSnJXCY79654xkpG9wWedhUaJHhH7MVmkGbZv2yeOggmjb4zH4gwcfz1O
9TigxGMG5cSJoV3YAroQi+j95udRlythBeGKIbfxieL6E5JhC2zYrSd8Ug3RlkF2fAxMI+RkPgrp
q79eeQ+kYr0b5wcyy98l1MVZtMC+SOcuIKEIy1yhoPEDxa6ILGeMkFWhYJsSPEY4Adz+7/tmnouT
MLrr00Js6LsIK3WJqFVUvtFd/UaT7+oHK0NevtjGC4PwXEImrHEO+aIARZEdA594ogKwc3o9tFYQ
pzhq3qXj/p/PkrXVHoggRJI8upINriLmzAl5qpL21K2NZTb74yETdMCvLbA2U7XNfWdTaLmyUYUx
pUFzF9jDMsxx89fP1nnnrBf/QEtKWXzRcsrGUuKLC47ctYlPtxU8o09Ky0riGovbppaDdyoT0HeH
WklTBnA6Y9vknrGw+lgC1L+AzOJUGa6afmIdyzRVxM+rz/t28u66afPx2Yj3SUzeaFoX3KhpCF2Z
YrC9IlzgH7TMYhBo+rWHwXPnn4e8IPBQfZrXGTlEcjDeQRVm0BNWGf540TbC1QyDKr3qSfb390cP
MQneFaBEuTmulEMenEacwljbq2sPGPc5ZIxiKjQUE9zOARluO0BlnK7sKpPOKaVwhmS4BDE4Z/bi
nRYlMHbACW9j+LnT0ONtPxGDleykCVwWlSmQRP0gT+pP7Qo9W9fYz2jxMUBa7EewFmcihd5ckSOk
TpNeqaixK3tlVb4kFYmwE0zcg1DRbiC5uFJ2gGzsTAFHJXCQSOBsfLsOQJ6c+ZhRAUb+9VnhEEsC
JmYgnVT4w9pitPmBTNX+u81ccNBmUfEJkNjPsjjkenB2Ak+QnzAJJHkEiCdYh6JNG8pptZjwmsSt
I4IvihSTpmDcB3IOtR++WUyYq/5MBGo2g3fpNOSTYS3uX1PqkCt8/tRzo+ikyFnW6XRl/o8ZLrJm
smUo8qyVaYJyHBp4c4KrTL2S0kDuHy4ZvdUKQRnwMmTIAoJcHVZMhM95gIK4ce5k8uKNNhTp7nQ2
438xjETE9fqrczmTvayEEoi8G+Tc7j3Tfb9B49Q7GOiDOrVaa1/vHhx7H6wYIQVJYPopEXf6ZnvZ
ALZb4cbgcto1wxdNdXwxEC2IhM/Od9n5JR1Y1zR2mWdPvp3LvmF8RugUG9fGh79ebC22Kbg3iX2l
twB/XOkHKspRtXajwfHQkXIf0Wmu2eG8D3jFq4P77K1i36ai9GfGAd3Mw1oG66TXECf0TWPeO62F
09UFTGy96kAzWR8dUfkVqIjn7oWFzqGWGtPY3Ifiu4ypOXriXpFVHFs+AuxzSPEbpq7zE3bHSRiP
G4bPWQtCXa1bS6GHnQsFvQPXM8FgdiIysRbXp2Mz/e+FQ8amkJuD86WiPXiBi2kwKXf+2mKIsybZ
gZZgrLNCqQ2jO6P8qyWTEGgT7QyLso6SRuexkdvSmxR7x8zwWGG7e+P2MAvRj50aPKUCTDjni9JB
6qghK6y53R4NrSpKMZORehpsLf7OFJFZVBE8KvCvQ3IjW9WodmrawmVmWFmedsCVwJdinzwWWpEe
zihSx/93SFRyesLQ1+n07cOa5Ljr3ckUViNwKRQdpAuz0O2RuGFfbE1Fv97KH1o8TgBbaHDTZWi0
pYhg0cU+1WcbyTesQ5yRA1BGrM3apdcKmNvRRtrnuqCnhuWcu1yoCjEjvrNInQZV4ocuVGWsEgzX
+dmy2TufDFSHFcDd1+T0cQExznCjMqEfPqAZQBYz8bZgmiz9xTNAekGlAIcL8mWR59c2uV9BBaWB
/rxNInEKuJqrnWDIYliwPMnPiiFQSIV1rZP1qCoA7GjkdIEXj1mgoF4jVc1+GSxSQhSLwUMPFMfn
sCmxFBgrsqys93Gi3YMbPyW83q2V8lg5RzHa60RpwQ/+wJfI8iJagpG59MSm5K8zXlFCacVS9KF/
jMV7f68v4j8snUVWMbXwkELOYAA4eYWhu8/MMdynvPqZQdNYcvjyUqSEJmbT2VUIGZOSAlQocohZ
ZVPrLJyJMUOfuY1PtzvgpcUOIsTRwng2miUh1JMzi6AI/5KWYO836acMGtpMP4xXwYfemkAy9xfS
XUgOVwe3DrqMyUDELQOfthZUpWHFDkzfVuWowMcdQFWB/LDI6oNPEPsIX2MB4eYdin1HzW9T87c7
xFi1845Ttawxu+NcoBl13ngWQcUVFnqetfjRhHJEubFBV9CxBLM2ks7eMbSD3CUmRvSSwI2EA2Md
a/4S2E69AjYoG3JYGdYI79CNZk4YtGzEubDTvMClPs0JQdNnTaVWVJBBIBYxK3HmTbnNKaHQmYz6
/jB6huHbkcs+uNExqBAKK1rPbGYSTs8+kXo1i9YJGbrWhWLd6SCagq23KjYfpPJXCYfNCzbsMJat
lnTESvWSqe0T8/GmSe12cIVrrSY2JuhlAxdzBG9TFRAF38xx/e/10zbiW6bQ3FC0sC5dBv9nrN90
k1GZx4XPOuHZjupdhiT6hXLu7z4FT5ej885VnfpTtsCRXy58Jj9EmwHagCir5BSMI9vDZYmr+H4v
wYp/sNI7hvfjCwfA2BBt8ACsom38OYxmLteDRjUqlMdTUNqs+79Fnh+4tycIStRRWWL2reGK1XqY
rr4Kyr7a79TiEdTpLMBYFJXse50oW9wBhmqbyJZj55Suo+qN3PPStaynj9xekgH8/DV5z5I9zuoT
cCoHNE9Ibzp1wYQimgw130iQXu16KQ3xz10Y8ZI4n0JZsMLE7mL8C5vTSAvJbj+CnZikcweCYoT4
fgcaIwT2wad2BpotzLnbfdF0zHv79lisj1SfUkKbGSAouE9Lv107ShB/d8ew72KtDfOkpaWpI9Zv
sQn9bX0PeJK3vhS8v/kms0jX/MqtSDNA8aRiL4q2rTCIqQJEZXYMM+ztyTysvbHMlnq+aTIF9MY9
VErV6EfHRCNLynw7aXA4FQ436Fa1l1aKV9gC7d1mvQUNKIH3zkK5EDAIHbquaR1bxGdYwBSI4oxX
6OVSarhVSEGaS5lUroN3JxIsXaXZhJEXoClJDZOwqaO0aAe9mPlod3mS4b/p/CJGTqclpYCx6Sa4
XKSy88xs+OuWq853fQv7WTGOSignxLSzj/xc40qAwNw1vGmY83NJJ2+fqostwGPZS98fIRSuXzo0
USv9nO5/ymdq28N1sl0IiNaKi9GFQYleM3SJR1pDD3tncoGd2B6XjV9GAyAbpS9Jb06kvTIyYFVt
gppjQ1E9JCYqrpn5ZsJD1+j+yEMc38iVGqRnoO2JADw/fvxQf6MVomPhC/1jNpyP3Il7eLs0Gk5C
n6wdC6gzmCvE3xZVhCVkrVNG06O0enyYM5oJeOd7eK8LDNC13jYCFfrQh7eVqxgUh5SpdhQ4B7kF
GO4G5p/k4GckmQw0hL99co0XIj5JFWWPB77yPZK6LEEKSnLpiUguKhO2yMY58ApkBKKXXBzUoHPC
Swa0Ggo+vZHJQDyjUmCd0ya7EIhO64ZqI03BxrjnmccCth8qInU973GAlkVWDavhS1SPBhWB9kus
QfWkmq9eKpnVy/RwT0SIdMPrafOWzZr9qhm/YIRs9rWeHq4AU4KedKTwanbo26XBMiSQoDalSIzh
xEvNDZZJFR61hRUO3w3nlQa/5RdlEw0c54WNjpY7/nYDA37qaKDCZxPpVKAheLvtvxwIKe0xOIJA
XVxVgQ7Kb5qITtSwjOmQrTRkUVtiS+SMuy9vHCAa7BqYP/6QLbv/1RuiEvW05K8ZZqLxWBhZ4PVZ
rGoZEcsMdBih/KGhyxmCjJxhvT1IKlzkk7L7iWXRW2VznUFqF6A1cSHAVstqhJ/2rKo+jlIFevVc
c+2RgZs88ZrJ8rWWr4Qz/+pNlJlG0qs6ImAADERDDMFFClx5CEL3kw0hczzm/naEbYlddLgYpblY
CV4UyBBLXfjwXIFC3tWzSsxlLNwC74JQuKie9tv+kNfNA2IENR+YBMvi2XHCOIhB++7Q7Bip3jDU
r8+doQ1BpMkwG/qFhRqDyOEleJMyCMnr9r89fm35nVHq4iCl4DN4DZm4l2MbP3S4cFbNpgglI/3W
YgsEFCZRJ8K3H/wVv0WC4hF1Jexd8W85+NxJX4qTj40J6dZ781A1GxpoMKofqLLqDONseC1XKGdP
iO+N/+t8SlJlrGq8BPFCy1ok+zvOIQFnUoYTamDT0EzbLOjhiOGHzKSq8c1iQC+/E7T/a3JL4OWO
mLJ4BuRDyF3+p79c13HyqfsnPHLhChJhn5YMesaGPuEKUBkywO5UgMnxqgsXny9IMYXDO5lZGAwX
zaG6A9u9C7aArWgrEVqtWSvU39LexmpFhXfDj7sCu101P0w9jkvbSY6x+IZ/9EOMSX9alH7ztxTe
vAHZ5Ody7Aicz2zF0AOEhvwe+rvasd+q4CwtAl8lQb1oVFaFf4oBTjXmn0IwfD+CnAeZveTUSJAd
0KS+gJBqIjZ0N6vABWyCgYAgH2+0jejR0/Sod8eQ/wPxWlBMI2bz66BBbh7zQVWC5G4z0IHmAnIK
WRxOQexGtoHsR24V5WdmnrhNHDKIYZVydzEDJhmUkrVVFNRtzDUa6enbw8x56otQWvMzC8099BIb
orh8SfbTIrXQsERMW8nxkRNffpCKH+pcHIRH6LmWpjAZocggRDTkiTH3zhy+S+8WET1RO/rfM4Gu
bDx4Irz2MujhIlbdvJ+WGT+Lll62ELIoAWu/k+SiKHkMW+F86nSOcvd/25BRy3RA6JkHI48cuGmF
01gTvsO3LSnAUSC21aq8SnOklwAqVH13r9KJsxquRgUM8OcJXfEF4zo4IXtrCRbeiUr8w/dkBIKy
2klhVHLcUxakF2m54uvotVuZlVZYKwlNC6UIEjJsHXteg2nQCpi2LlHwr0uy6oQobQ/UC8O3euK1
Z8rc/PUmSIqiD0VYSuWAdX5Z0fH7olV4gjB4xFtuEORKTEzBRFPtJ2Gqr1C/piz4o2MHzjvx8bjb
Tk+mh6Td59c8MOShvZrKvVGysKZc06n/VWf+9+MfxJ23KRwTe/cOXvafNDn/QnsGgmH0MkRATGOr
IkXnfBlujBiuajYhxxGGD3jxOpV0bcZ7lsuw0KxQOor1kkpP4PZrRdHHdVF5swhFz7jiDDY+Y76e
FvR/h++Boyxf/ASYERM+o72xDt65fEOnWyzzlTNtekgucxcCP94m285bxmCFXFic96h12GBULdsP
z8TDwypkbMkY1KU4PImteCCoPLB+NbGDAmI2bBCJe3RBqVsW0B62Zfo941On0+qq7P5MnKn90mIX
VmE/+d1EibV9RXZsVj6GuTS7XtiJdhW2XN2raq5o6k3F8s/HBMOdNKmCI0YcCYvZRyEqLn2BhaBP
Fz5A3I+1WsFJg8oyaYr78jfRI+iZYHuL8UOcPA0iaVYLEDqSl03oo30K9PLqjkrBYtOpECjbSTes
ZUyFzFMFOAyejWYJh544KpN1scGN3Eyo09h0O82vOJNhPExj2U7cNwSg7jH7wjSms1tOGk0mkWv3
RcqppQhh64QGyV5DtkBZT8YRz0wVfPYrfOgtIxgpnoKtW1sWpBI6FS2bes2k4R7NmWmzJVFZLy+X
aw9D+NA3EDCMmwAjabV7JSimLnpHoj6fcNXCoXur2bmaxmYlYe03M4IyjIYSaiSem7Xld6HpZIRu
dyp4XTnVMe7vL5ic3ujbdGaYSt/1e6O04NgraVY5Ho2g0zNFdsJN9shaMvfpiay49gDVpC/yqoxG
mRmL9dL2yAOjI4lyNFYwrCVcDt41Zfep+mMOkc+JicoZNBJg/weBjogDxxJtP4e+hlE4OuIKXqap
2M/I0Q+WtHfoGO7xM84kNz1czb7A6R9EC2rlxJcHaAkWzy/5yicrIAqlgiiq4SaLig2m7NYw059c
TTzGnZhdl8LURc9MOR6bHFXUswkL8yB5RIgv/Il3LTmgA5hIr56QgzRYYVcLHW7JQROlVfdWa16d
xNnCHv+OPoe/Ptr+RnX4tVL3BHhFyL4YRg8piIoWS+vn3ok02W4DzggbJSqKwo5t4kqMAbdn27uT
0FuVQ4nN89LHnOC4F8l8f1NWKabDG4ZYJLAdiwJ4WCrutD3I1TSKb/3LJDWwEGx2qk5y8XVgs5uF
cSa8E3qrwbMsRoxaPok1R0xbMngspatueYo10mgpWWOm5l/xX2xexLkkRd7g7US+wMZWxyBTv80X
awcDwDqhKMVoc4cHVBJAfzQd6q4/SmhGF0pKVqp10F4lOA+uvcOQV+Ra1nbMPknFXeQFYmBRD5fU
+C66hpvWqZ3qClTBjVfxtFSyus9wWLLeALJFlGF8wHbCuHeOG1IItY+Uya9LAzKfn8vB6Qp/nC8x
fd4EyTFunsIkUlw0KC9IJ34HbCMZkhSQbqX9rJvgSdWWd51JwnDRg3A03bAYVIoOiqTiigcqoUsU
ECcA0Yn4FWjmPm1YEpj+J2oW37RCWAbnHBZejWG9kxcHLRcxdSqptKnDgMigB6kyvWKW+NaQiVOt
OnwozIXVhyzRcbKAfAVfYkvlV2juTTfhnneURuHwC8UF3t2DNH85LSPI6wn5sWplw2o8A0OgYmGN
cCizM7K01Ja0VTwVJf3vVxIFPYGq8sTcPd/ykuvh8zhpBdMr+5xjTTAYFnMx5riIQ8iZxUBrJXez
q56gLsuBcKYERNqu9RU/AdaJvCCAzf99m6Wmk/VOB6+NZKrSh9/lekEgekuFWkmokpzwQrNF+vva
SsdJDeKv5/OaOhfUg25nNJ2f10wKjhf1xP5P2zzLj6Pnf49seiz4bJlcr7dOnfvLGQvSwRFX1YgA
0CzSFTIkNesfraFB7RXNbDRV912y7+SLhGi1tZTDqKKD1cxP4MlG2Cfzu6LimyZpGfW6+0MgsCfA
joyHMkUtEIdFg9vs2x/ro9ZnMAfrLUNToWmEqoia2wCU0lP4Yd1osqz0cj/HOpgUiglNvz86wl1e
Dc/sD/wQXjs55dF01dpA9DTLKlCCNAPUtbPy5uaVPQExcSbAnRraAylLZwhWbewtl044kBCimfuW
umtI5noGZm9vwn7DJJgy2VaNbUYGtb7oKpqQOzciDcfY6gD9dmvJ8G7JLQEB4XrM/MTunpexWOFs
Vtd6cGF9IstQGY3HF1ysM5lxiqtH2iWtkixLtvnKOHDwwSnChqxxS7IsXeTkWDFEy6UUYQu0OKtW
tETL6X03B+hmwTGM+YZ1oIDWfw5ye5xFCvBiztQo432AOibIYKqIy6eB80mxcMWIhNC56h5IFRg4
EEZkI+43CzsiczRWVTWZAhI7QF9CkzT3yC4pmWj1FLQJmdWqrLh6+CQUELOGQjaMIUivpFAeoQQL
0sUDpzOFjL5CH/EqUZ1OsbC/bMze+WqS+N+qj5cHOy8uwsj8MVRp7iLpgxeGPmh0aZGR1+DqfN+G
UR1s4OswNmWASqRuxaKQuB7i1UfaSiftCNcSsLNQS5UiaNXYeomspSY7DSe4OC9n9AqkivRWJrY6
QK5wBPN1o/oiC+86nFCuSl6g3hi+fhPjfxuYzCi4b+syST+c5WV7SJ1rc2YHvDkG4Wjp9DJ5XWGK
wSlucfaC6RWD9sS0MvX885pGjtDKO4CM/gM9th+6w/WGpIJwl4P9njyUe0ovp6kZPQt1nygryk+3
op5/dNW68IGc+gHmKucA6O7vDr1U5hx6BZFZbOvB5Wh31k1/cc1AMG2etsGnOa4xjcJ8C+XO8l/w
viQJC++COo30E7Ft65jsJztf6V2C8BDlj8Q2QlJRDVVTHbuEV2WnNuk4JiyW3YIYDOdQO0/I0pDz
qR/qfSIGahwTYfihlaMLdsY7d7ic/bR6ACQ7e+b5HqNE1WqQq2mnzk3BcRJXhP8VGWBkPFe2RPrM
dyltXtlV12iaqvnyQ13l2QINyq31FbRJueieCMf8Hrzc2JgBqkMoRhRyvH+7iWvZcN46ctxBQ1Yi
qPkZAGmIOu8VyPpe6YT7RpD2GcW4jFC0C1Ip7q/G6uy9HTet9hH1SI2yIdzMMqbYRHgRvnr9fUhh
QLx8LrYmsc1uIee3HKnl+s+xJvV6c+6sSOOc9MhtxXEUe0KmBKO+Ect0siUZD6ZvLUBCFWZgVuBS
TM6+owKPfhwgz8uwRN2LxOiagqZpAlXYXgjpA2gqARuHd+jdYzpLWIj2hCnb2zOV70Cq7oXvmkDc
RxSWkksENRkmbP58XR1+z4KGCpDTiPfJlzEJts5fa0WX6YFRe2R/LIq/nrX+SwXICw2cgVJ5e00I
kyqcPJ+0W2jAFwOXD3rPBZgZsMKZxN69fyxLhU3BM7X3ARAtdr8yxFmvYJauNR3cjocW3iACYmcD
c6yViiM3mztVwpm7h9SH4N9cDd+2FOabuCDv1cckNr7NqW3huMk1VIBOaoV2RFNc2C89oTP8Sev2
PTZ8yWRDPvc/RB9+ZZpcmUUgD1jhCyNPBYZ5HNODI4AvLpHS3WV6/c2uHAiHx2o1foxcExJrvHo7
soZeFyUf3ZCb0gHUaB+93Pb3xr9OV5Za5RxzIMsYyjBlzKqw8hs2lsFAN6Mbm5iJXj2WDN/Vk0Uy
aZZ3mqHtETx4Tzm0jLu/OocZYVCu5jyBUoV1dpy0HEIWlfdy+jJGt+Fv96Jg6quNxvAAdec9JjVX
+Lxaeo2x7Yqvg2oojgL9GFwktjBy1V2Hrc1cx2JIwXUdNfDqg3zjadsB7NtwkIZSg98RXK1rCRQD
MfLZNoaydRkScgUIwbGR4NAXNS7SwJ4qBGaLFGTL6sovLnn8JBzp6wixX492o41zt6AwggegqIcc
HbiwzqvJdXeTVFtFe9z0X/pIX5xJGxBarIj3gV+J+nHA+EKBvZqgML6NYnkrbYzt5Sj3k/WpFRCu
maIlV8OogMN8CSeIzz6zVIDwBDwR92Eqz0Fn0CO6sXbZYHHwQxjEY+bzLDJaWVsBx08cKxFRUrFe
MAEzY92UhETZ5CAg9ixv4AMxxgDBj1WRaR4zjjQuDhH6bTh97A86N6JcU/Q5sDTg1eGukvCOgUVm
2UMUs+Jwy8VM6k0tM3UA+RJUyT5J1eGvuNSrOJxkmyyrC8s+VQpffhLtJ6VrtJqUgGJNjvWq4BNT
cJCqYO8BrPK9ttBCENTSAbZkKbGX9dh8I5wTzEc29sfjj2jOQQH+KoWGiVg49/Yk1/EB95p/s+Aj
J9tV8ZSgAdoIEoCdtClADlD6OHsc5N92hcLKHyUGKgr92bcrPhVIl8uh0v4ZxXHEUi42iHh82b/l
uWjbKW9YBkZpmwLN8nLWBp266QkqGdGCLie2D8Sbm8esnGG6TgbBL5x5ZV5zUfMLF9KPdNcQC1CI
vkUKr/SvsFOq6wX3xrlohixdQ+A9gopoP4Clu1ZsCi5zQ5YWXfG5bGUJ9n2iBrFt4dcodK2i0b5W
V97e4HqdjmwUdNH4jYpnQxTyPs/0ySkM3Qn46+EcdnmGRgBjuUckq9ZLTqxYDJcoMnB6M+KyPpKy
2MpkEMXu+7nvc5D9fzx4I7PF/o3dbR8sfy+8CY30G/adBzZnQ3Ok8JH5yExEZDRSuPyS0fSEtGzs
LCxbJR1gkyY1DsqcvnnbT1MrRgFCBo0BJFDzYvV/7czVB3WTxDtlHwJlpMidTJtxfRcNiTMggcoT
kCIiAFbb8FS5Mfh67Q+2GONDTGNp1dTzW5XlQ9Yg/104A5qtLyvQ4zgeZ8pjp5x8ZhfxMtMuYwJW
q1zcBx45pq0/rx47qy+iE+wDnYj7mWHNieRlEBw2jwelWVYypGY7YLtueNw5MU+848grHwwuLCvk
vg5lnU8nGTswemttbhwgVQsYbFupGQOyR4/1vjj1PLcWHBCG8/zs57IKtVsTSPemCICJIxHJj2W3
8z0Pc5z+sogDzlNWXe5EfR3LnrIfWZHyw8ccJYZSvopY2k7hxVmxGCNdqUZ1Wt7Rhorcigww3A7A
nathkc9L2DcDGb6CbOIYgOY4fDVnL90tVzqWHH88l6FC8oRi1031omIgI2FVh8mHCQT0AAxtzH8w
2PwhGCwhtqyEcIiCX6NCSlnSwdlZChzA2vmeXM0Qeiti5TCWFBmeQHBahlLPwGDqZ+LkUss4XaWi
OFg1BavuFf9rpqnYZUupMVBRFLbx+QOl400xDRM+Bw0wGmBxh+IlZ6CqW6dY7GgKf8lB0+XiKuJ9
D37C9njiR1dq2GN4UjxTegnPvvCfIg/9uLwd23ZhIyLT8zKBRe59r8MH177PEO5rncQARIfQnT/n
/zqMpCkTrJ2apWc+l83+p8Rw8ts1QLedRIM+CUgUMrKDckVG9ipYnnW1Uq1A8c+uCLp85YBzJ3wC
oC9yGKOVwqAyRkD4Ik7+1GABTobK0PioddLS5yTWgHZz8dWnLufn8G/jMUbShYLCNbGHLP+NId4F
sXUT/Vsb6/DXTSHOOQNwzLMrhS5HmSFLW60uRYk63HmeqcvRSFN9D/u5amj88ZqkGbRBj7Q+EN4f
D/IW1OHqFY36zLKJyDdHuSbFTHT/e9B3fPA7BaIju0HAvkkLGNfuiztrukSlUNsm69R1i8p5jSIx
G0tS/x+4Dl/ClY2ej6SiykTwxaOe4I8fNBdT/HT5KDklDt4c0JSTOnBs/fu2Vq6v5ReJPkD2zVj9
1F7w2Z39nCtvdRpQQgm1Up57DI3OJ6cB6H2NuWkwXHS64N9TSVmE0PDVJ3PYaGH3ybXEfgoQqGUn
vKhnFXL6GPehgNUoGUqlR8JVRUm308jOxfatQH8LqFkt26nvbG2nq5ExXaHVlOitenJzzpfN6D/s
UZKYL7UCXGCsW3bjEFz9baHNpqlyisuoG6QXExjGaWF1l5yUigyPwz6NGkUywNUHE8vMq+jx7mQS
JaDW+xvRkZykh1moz7tBemqxGDaDLTmwykemF1f5fUrjOl5JPPT5GOrN44GxSD+D+l88S7ujTo3+
9IX4yqSKIBENplZpKL9zy3j7N64kSxq9lfxFWKE5KBIzjllxthcxJrHsRO+L201+iGcGeHT4K0e7
xRpMCP+laOLg1M987TBpp1RIfSUf1ecaprFBOb3A/gBykINShq0I7aK5WXKIHuUGS9iYXK58e7DF
IOt67PNc01Ao8oYSKCpmtWUq7/gX6PbeQhjOGvEqBkimdyCutllf+Whty0EnP/dnTc0QS0xmntfd
LjkCTr6sPaKkzhJib5ru01WEi2pE5hHQG+Yl+FL50xRggJdG+NCGW2n/aJH/NLh23R2hH2ZcOS9Q
a4nxlKKK8vaprZGgXcaepczDYQzmXZqYoRH3FxBAGb6zjo3IXBjXkMTB4rk9bRxCSvCoGP1hofx2
lQyW6r77O9ewj+m/dSGfkae8ox94wI9gCvSzRuyxUKQDdox0WsiwKCh9vx/Yfvn7H//EjT6p4aAp
0VliZff3X+AUjJX8rRuENRHXmt6iRo9vAN+gfcofxq3wQx3nK9m034daa0WCmOZkov8khKaJpSgF
VJpdYG1VTdXBB1e0ElJnUrQBVxjYCOHHDRuANmSW3qTCFhqZEEX5H4WzqxVfv8+wWQnD8hrPO4O/
BgXLL8uy4XQAYKgYtkQd5WBHUrMXk+8wZKVAhgl+Ofvxp5NkCi3ALqOXnVIJzOIX/QgZdOpUTYi0
Po+x0TI7MCAzTvJndmUtXUfm+7fRzJKZQBV4h1+OTg9y6XjTfnrLMsKE7maMOKtB/bNt2OOWNiBs
J5Mr00fni+0oRXEC/e55OI6pLe6eFqH7cyeTykLh95bwcEqpFLBMlx6U31FVsx5s3PFdMNtquIcp
3DPZViQNWNR9dE4wBlTVybAXa5eN6m8jxNIO/0eIUN1F3HtghU5AJ91+msOvkgdrn2zYyTWq8QHO
LWOPefDS89no3jkXM+WhCwzwZQ5FBT2ZbZq9BgyeBHkGdoE2L0j5CTexfLWoXc4jRt2NupQqnMPG
Leh2cCm87hes52uE3Mp2wDBmwUJb1db+s6rxvaaQ2JtM/KpR/EqNIB9pBryvuiROZgkzCWldzCbO
gIjapLd4fSVHyjXe/OeOOQhlWhFdbYJbPzho/NXKiN20W4XkGVu/CiHZR65O00mrDycpNIejGr10
ovAF3zSR336TvK3cDflbpxzwU8Cdt+orCO9aQz2Z0Ess/1NZUtzLRGoTSBuO42RQoPE/uZ4yLCc1
3XxoOvE6+XDSUqNsZOowbadowp1C/eH4ZlRap0Qd45uHJ7o7bMA46pnjmoa7S+Qc+4f6PZjQ02vr
noev5+GarEEJvKCu39LfbA1KD03oGnRYGoUXNFs4yhCtYXSNkK7NO7faUcqQnzm3fBF7TrZ+A7g+
FFrDjoEuvuIvjzspghk3n70KihMFIrxIf4z6qIPD1CYqDeJd3+48BfZOnYRGvFOVqnbk/DHIbTAQ
nw2EpV0sxEYo23PN/Cq4jzjpKArqykjd17gi70hCkJgBe4l4nQH/Ae/BohMU7fSClQZQfC3+CghN
QCuqxz3OKEG8kdmBCC45Ahq2cUIT40lCgCiVtnbakc8YZHLFA+jMq+rMukYuYWp1jG344pCzbu28
zYcp35LwC+vI8o9F7ZRaZCx5AqVuyCMvmc2w+o5LXOrUQgFxQ6HVvttuP4Yrov9vpTAxGTmQp1iX
GZ5QKlN3EaLROxSqKkKZ3bQlc/c7CfFlB2lkbhpq6F5RSzTzbiD+KBoQM55X4TxobiILXRcGWLPQ
z5E07bwyVjREdLNa9Gqumy9W2AvDBg9FaM77sv1xkY79WpdRsTlGNznhV5em43mzilVWG7pVim/Q
qm894tdJl/DhHuW9ShyT8J6vFC4iEAUKrHeEkqG+lBDVXlMcV33rLCMd9fwmzXcHBUxG2lhCWds2
/A//sKodUfp56Tj1RHxW77JYpb9kSkJpinww0daG0QGjpoxc9ZRKgC3h5+8Oi9kzndraJ+uWXG44
qOv1RaWejLvOSOZqnHf55zXQQMAHs/UvsqSpvpkKNS5SaMcN3rZ8fWPUwKkYH/5qGCJmx/DAGUGG
Y4XtNi9CZn40yutk8Feiv1OO/Pcvd/FB+N03wjW97PizOTtSbBTklUOCxoeR1fVQcRZK9wHz2fYF
K9BgE26LuQbmZshWLWaYPVVRHJPxvij+pZHnP3V9lRIyxYKwHA85vZmcRHkhe0XlFnv4RPMFd+sO
fnydL3XUcOO6J+7ouPTr7ty8T1OxN/8wjrsDwOncZNBCuAmuwmjKnrK6nOkW6OEFmDKAeVF2MK4r
4HExuhlm9FA9NkV274AedIHL86NKoXeBI7PFReu5safg9BUjs17H8nB+pMHWfJIISJsvGMkY6Em4
K3sGwjz/5U+YCgOsAjYPxY6JFRMj6p8TS6m1O34edPJ3rpi0OGpo1bfxErMVduX+X8hN3N80nejQ
1r7nlv8mInv2iw/kk466M+f5hYNhyibSok3Sg3H4gBwrnHH9Nfu7dQNQ8iNsZne6hGwHHxyAKtOb
V0aioX8fFgcOJuJuhj7weh1FDF1h2ew5Ggh8Rk2qtUKNVQK7VjT2rppaqf4ZlVfA5zi6evijX7er
U26HfV+8nlHT5CeK4Cjl7IXswuXySq8tbABRjA54R3jp28DDWGtbwBwmFodUkHTYAOAOR7TVLZ+p
zIyOcX0rtR1rMAHqnZfyTz3HnbwQwjM2m7GF7xDaQgyefAwet0wHJGxLk8zsSJyT+sP0hveigCRk
WOH7DdhYvuzEGyMneWWmT1MK0NMmMr45ixw7giQHufB1GSjtvI9rk6AeizWMHgCtBKRLXLGAHzUW
jTK9zUZgFya9OWrn6CJ6Avc8lzYm6CBoTEeAjjkGQh9RE7iG56gBfSCZ7P0G10ScpEyF/HAeqdRR
VUvsYiovWpHyEhkCt0m+rXZA5hdHoqSnVNzp8rxbd5/jIQ+OaywMP4EKdqXPEW3Wu9o45InZoqkd
RvvlWWrIkTm6HgwTnznoCNN45JJU+fZZ0ATK3DE8NavyNWwBrJP0NczOd2B1AwRvXcxNPmFfeND2
HNhHcVN5HB/X2xfhII3n56EosolR8qXX+x9mNMFZXwzadZprxF3qpa9kx6Mrc3HwW/Db51K3BTy2
J3YEHU38nX5ySjnE0Rs5JWwTS4d3ZLa3SdZ9OhBtWBGbASiO/82rcveSH3ii5h97a/lBvOFaUW/v
fiy6iKrXzg6p6vc2bgVjgF9aE15aQYt6Ht7c7YX5g2MAAPDViUb3W95SNBm4FRl8TKbiA9rowoUt
taGjNQHJL/BnCImN8C9YMWgLqn9gin9mGKLsCvYvWphZx4h1p7+/3qt45AXaz/gAyw8YrHDOjkml
PDz/qE7WNgQGesd2YJMrkzXEvZgUPh9x4uyVsBpIAMWfesNYxe2ooc9KeFITt1AfqkwP7odP2OJx
sJnQM+BWpXLDAtsDF2x+e8sEFn+Ahb3gdfKFpBOSBWXEBTRo2OP5L9nRSnLM2+rrPnOgxdYFd5fn
HddHufIsmnUuGbRz/CHhe5eR6E2NWDUB5htF1F/xTEmLWY1clDEZ7fHIGUyW3gGoEYg8R5zF2ptn
qGhqm3k6CpoPan618FZ0NjjKDn1ptb8ympVczuUQZcL5bgr59J8QfJFowk1sRrx80rjqby6sMZUw
wlycmL2hoV07KNVgDWTRzDZKUHBTIOfDRz9oZu1Npa5Y+J7U7dV9NsV6FAbIlK5nbro7CvhzX6mk
ItHCRrnl9uoREVvUuiEAvopI06gY/8qQI9YbLOXQDNj1Qb+tukpHQ3punZ+q6MEGXlbwUtON3O8R
fI/d7OUD5J1go2FsulYQtHDsXChsG8/AMWwEysJ3zCr8y39kXl0i9Lm4An8IoOxZnaXVnuJRRViV
IBhd4aBGstwnXqls7UVXOfXGPo5x8oQv2OZzl6LhVjEdL3M1gdKv2Nx3hjIxebX7LU9sBCwjAchs
fJ/yJXMpu+r7cn6/bg2qjOjuENzLDwvU2+y4LOi+kEfu0B0MzK8Q9McIr+1qy0CleX6Pcqe6k21/
yjubdkKAWbg7Bplcfsdvo1Mlbo0Er6aDVXW37GaQJp7w+NeAnen4aUJQ0Ine1mFOt+VkuOtUD4aI
OI72zqu/yK4bPGCyFUUamBaHyRpcS1iwY5rHdn1lxFcTRWrVzBb9K3RxPhHajdxLINulAd2gMLX+
TljFosf+XJVp8g5/dygoMUq93ho5wGSbtq+1h1y6d0y50D4B6FYJOjnCbFCC3i2O0RvE/awuluAL
5mvNs2R+0PFvtrftLmNH4sAV5eD+7vP+V3qUfUUv3eavlxHrseZF/3JOBjJXO02kPxeEWGHU4P53
HhtZY63assbXs0O3Iva0z8msJl1ZyaT/VccP6u4okw9WErb1n7CBApCcINMyaz5KMXBjaOxBDA88
rJvF6sRiLuT93J+rO1Zhnn+KH9yopfDrH10fofpiFgvEtjRWaww0tKY/zcJPvYD4OrNuY/kBYliO
dnlG8hlrA2HpzV8I28M4FoOBlJALAFim8q8oEf33UcZsXdocJnugS/EAwuDBvg9NTiiA+bWIXF1C
kIBtOS2BqPraaBjPChoGxrRgAWM9UmZqatD9JAOBdfbbaavsq+itZAh8VE2c4F1Tp1ycEoXOjxYg
IIqFkQjunYBD3AV4sEw1Lbioc55vVq5TEADFUm0E8meJtOieeYB1OZ3y6C5oLK/Kx/EKjw4AvQrF
PpyqGKw7sev7XTb3cdEY40Ypo3RYcNyfXlAF+G1Hqz++p7FdVOiQ91xE78eH1/ju0IY2vYndzpko
ULe3MiVfLIuLaCHzDlC+E2yqIvayd0cBxRzfL3a/yadRuBVYoGCYIygeJowEAAk3TlRui3JaFtWA
ZTbiViaqSfdbjBIEC5EGEw81P3/UrP90+cG/1seouKw9/O9Eqzd0e9KgSIUbrGZh1kBtJqdxOxqW
gP9mBeXsUrMoqPZaJGjNbK01ZJyzZWsq6MiFIulG/2MU8rRJPH6TTutdXcM0PevI6IwgFDGUsUjr
yvQybzNlemwJd9saCsXApUSzZJeprRJb/E2nRIa0Dui6UytN01yKcgCeFmyNpPrKJ0GaF5rR4f4n
1n8ipPRjdux6BzyKHkEqRd94sZvJMK6jEoT8s6ZtgyUgXuLb4UcsEZjdHBiKUQQw5TPeAHjYHS/C
+/dl7EVRhoHDWtvBt9q211XY+qtk5viuHXCC+U5k0J6ynMhuWrWP30iF13MeIm3GuEMS2z4+BvYQ
a0rKqz/Q0mN0LmHc1HvIbZu61GsKQ7iEhjSPqBQyD8XK9IpzTYqEiGS3loKW+HJeRWoSQHLwi3mb
imPzshXlN3HDy6MCifgaSM8GPUvsgun0C6zvLg7S09ZLYhFyHP/tOKiTSHeZ6wddPtwUrZQ//+Ak
KY8LY1XueYK3Uh8lTUh9bP7Sd+oU6/0HebDaONiVooyeMmrJaEK/YpN+1oitP7hNAdadbyxgZ+ye
z2tiQgN0cDk9Kq8JisYj6+6k39h2/RZIhA9sPDmJW8eLB2hQARGe/cMagBwSi3V6EBmnbkIV5RUJ
pGrnxYTXnMu/lsyrdzJMD1PszIGUVMjV3pMV6aepQ1fbP4hxRepTq3Vak2vNeBaeamqOnofUQ+aq
nzRGrHuWedzv2B7nuzURAvY6/pT8HoZlOQWYdFUgfnauw2/LII0OOwgvCy/UIKOg1pATd6SfyZUX
SoFNUVP1MCwSGWVuOluZUBY8s20DgiUtZPVsBxUwvi0LnEw1cZXb/WhKqk2nXP2TXs2qCmFy6LdX
LpkKhv7ZJlLblbQhBwIQXIvvkkd8L2QXTwQ1sCXNUL3gAXICLzLHkzF1S8YyNj1WSy9aYzgXqx0W
PifW3SQJqZf6G8OSzhAdo3NPB/s9Va3TXMudblESuGwfc+jtLDsddkdGdc0w9Ehvx+EQvCcsj9X0
bz2e64dvvZdbZViJ9Omr5SM0y1CHPo5pMhoi6K4q/WeQYVcwfyUI71sA3oojRf4N/5/NXlbnkpEc
YPI644BCSe2JGdsSBcZwM8bzhWoZG73XsHvXrKm6B/Ttt2Mti+szM7QwdOfPkpAYCQnsekVI3jD2
qDbJlRx1dPNkuErGP0lAFvFraOSqjtRfl0/15JvyJFfa5qgABBtwFoHs6csRBCgo1GQf+YoG/36j
B+G7DXLiUlXNXN4ytjYI35KU61J+q66iIbCavKQin147mdQ7VBwQRfNh6l09OVHJOAky0gMDM4l2
Y1rlpH8r2M+VYQ1wHwuxsUxO3SmBMi4rTjDKQu1uoum+sajHW+Yl3I72CphnBPelgfmg/IpovkaE
PTb5/gNxqluIB5AS2Zkjoy225L4heYQWJZb2feb7y7Auwv2N6znYo3ARVYazh3WKcRzsU0sjf/bE
LuPaqipv/582xSSw5OS0DIXu4uFWbL96k7wsH8NQswzvTaXaz1jSO+L+Rvayt1hq4M3MaI39brMt
qek8NxK44+5hF6sya5J/tfZ5EGtDVBpIPuAuAeBx9OrNG+pBfOkUa2wnQcezB43hWwEwnLzzKFco
A3YOo5q2cyLDLqqPjT5Zsr3S1eqrNjGyT/B8fyQhUUTCOoluuCS3bbGj9feb44ZVqyTjlTfZrfJP
pdbyk0qOTJyb/Ga78amL81OsF+no+OaNanAYdB6HyFUoVI0F7nggrYeBuizlTOehn5Nc3TW+cACD
YPTFsFMotSaV2R4IthA2REqz+Ul2f4rs2Bu9QRQIBvZfXef0qkBEcP1tJm0Su6mjKXyDWxIQdw6/
HOHoydXONiskVoHJNZVar2RCa5zZtAPgyXNlYX6yhN8JDPApLhdon4Her8WBTgwGw8N8eKP5sLjz
38/4Dy26aotaPrSOjqyiMPtXZUUm1rRXq/bOXYBof86sLf+u9FqmqnaPETmF9VLhF/VeUuDg0TY5
+V81iv0qVrW7X71R5ZASddmPrSn9cOfR2ZyXhWwTStcLX+/dQtofyLzhLTTSWc2qZWfYmqwB89/P
cS4madIMfsYyalNzmCxIJIpRhYqcJYL8f1ndqef7neEsFsrOrLO/6+COrOoXVCWhBj+dG04KPBJW
LhqXpjIpG6ZxMabig/Ai4Zcw+HX+EDhfl1ff9UNGLJC9Urp/s3YENHPa/fQfMbLbr+KAH07qf5Sh
9/NynJpeQ5vTfws64UT5XWoipgkY4ATrK+6AioYCZm4jPBw2W/KG769tdhSbXzYrAVJ/veMyvsOD
Xv37J3ItD7jPbDfXx/WcZngM7b/ukU7DQjoXxnFIK5Pdvc1qFC8IIFZOk7MxPQxpgfdQJQIF/WsO
ezPnqR5bVSr42bVXOU0gdXKORaiE1hNjdM+FSLGkK6oYMNJpVS0+jYbbRmfWG+F7IhCz7L4DQc5C
ENHRk5rpk7wPETZUsNHvkONBlPBjETOlWIisNZOCYWq2j5YWunpitKoOPSaqGyWdTdZOD4mVvuvm
48bkGbM+70Bt4xLBKGavQvYxeR8MTHh2Y5W2KreVYfWH24t6QXWYOD0PsVcd0JrNEpWyngb3Q/PU
luTk5EQQGvFwE3TCwamkIPcCT7vu5y0iYi6cLD9e+HiMuEA1ouktoeONr9VJLcrUiNJUwQJ5/rJf
x9e9pBEuzg/U4N/rjFP6HjnHFAFshuRuC9IQPlV20Cd4TtTWDrqheoyJRU291CfLN7rnn/MuDNR/
W3dehOh4f1CTpuoDMns1i1kuLGOtF/BtvnyyB1/pM+VxaO0xZQpTluO6WQ6eqQu7EXiCYIF2cr/i
OHU93W1gjz6gC4N74zNbAJI8a66pkMM44x17v9xRNNFYhPInPXXEpDeBEu2fJFz6N/E7HGGstam4
1FVVGqUfhE/4wQeiODeblwCuWyLhSdW3cdOR0kGFcbAvszwhEOaNBJft3Bjd3zxMEuVxBODIuWtP
tBYlb3CttOXIML/Jq+CVm5BGFe03k3AsXWo4cFQKK9Lwe+0uzsp32qDZodknIc3aFFDSuG+1SqRN
dMPQfHm0DlZbU3Id37l1w/VwiYNUnV+AEASskgAO2rhTuUriomCt/fpr90SP1A1Y4XhPnc8IZ8WY
eBB8/FPnDcb9UXftwIjrE4xZiocqvNKKNFhSKcZ7R5hFjXJXCQSmze9f4Bt/Bvhb/PWP5YcYmOLU
15jr4YGw3LggXrdxIC9DONK2ym7Wfh4QOouOhnf9OibeYxNAQm3/zWy9mIthPtI/82FUebXrXTf/
AN+cQyps8duAeON+p2SIUh0UfzxIKDCZTEBrK7mwvEHMwjlVUAT7SSAN+jI0P5L+mofe3Hsof9wW
oQPYSqrLyDC2GzyyXgMR/AGxJjyNsOuFhQ/fDxPKStQ/YoJHw0Iuv0Tes0XG8Otb1jWNfVkMMOTm
mJK6J2xd1NDioiW3ugdrPm6pE+g03Ry0lzJ4JK87MYOjPsimBFTtnyxEdaxz6oYD8i59mdzhPEmg
IDybPLKdc1qoMnLZdGqgtsqONMwnLpFhVx3lJN/+kMkxZ/z7ohQgcO8WZ8SnqBSkJ0X2JpoXPkeE
LeHBV7jXKWh4f1tjTGD2Kj42+tEpO0JWZ5vtJfMGJr/92AzTwMf1m5eXAgTVFPryBUexZcGTEgTu
3siE9jYZ9vAczlfr1VXT0oBsLA30U7T26WEMBQfOuezFlEQxOFanMfli7l2DjsT2wtI6ndSiT7zB
DsUg/1fTCqDgI0V58oklUc5yEEKf6MZsYc43NSAksW8KEMvhYiDtGi/YFDnmZDzxfUzPsJzdGPsr
vs66+yVLy802OgT4ghZAPeKBzoQ8ZmLrGFhwqtSIbhw0Rjei/6OLj693pu20k97rn5Axn08P37ja
LIgRR3+5CDzgrP4zZvq+XcT07TGj2LoWiAF+2xJDwTKskDduh9mWCkoLOU50K13DuxZ0yv3tKQkk
5DfJWnLf1vX1/bWRDDbK50OW18fWaLg2tYVTcG5cer2yWOI7O6Wsj2w98S15hf0HJaeuZMx6zPYm
S8TtV7xuifgVWlIw/GolohjlhLf4RfE/Mcd9kJJvedczSQ98lekh9/wGEIHVUZJXkZBHboOldHny
qGllR3pZGtiYYqkIw+QvuGBAryL3aDdo+aJtxwYhIEZDmxMvHfSTaNyP1uTCCS30EVpucliBuBG2
uhpmnlb/rvKEqpdj1CVSIFP4ePclmv57aQOVy67Q3JRbarXyb3vjDo0fXuJPuij/81CIVkGbvBhG
BdDrHN7RQPReQZEetQ1qNauMd/E5VfUCS9iC8Nho9x8KAs4sCLTubEv1oSa8+8TT9mbujXI+MuEJ
txqGcnZc1aLVDzys9G6ri2gwrhZ+L9R6ZtnCg94+MKj6F+XLmlZSGrL4jy12EAmeOcaJ41PlaWuN
FYwNvpzrmtDZ79BTWUAtSceezDrMwOl6JABUKdYKawnlJpLpCdp2i+TBjv7DbmZcrMtlY3rASIDY
E6d05fOxyLmnY6JkQPBa/jukL+jkDQPMmVE5MqnR2wBNhMFEwxCjFpnSxI7EWFEBsGyMh2ypK3SP
+ScZKUANbLxc9KAbdCffmIk2GmQkjQPTXY2bvz9I1Djk3YW+fgdndh9X/6rpVA/B5LHu0uTjeVCf
CA5XJzHal4QHAIva0BB2kSodQqxPOWdLcvQr8z1asJdsErzwi+ROuMCYxDjaUjBbkLD4jgSgLpMo
urKTXiFMbW+yYy0SSj5aZn7dNEwNvJMJPeRVIL4BwlK8WT7QqGbXvN8fccqJ+2luKF8xtR45cELy
IH8SPFq3uncghTPntVaUDknilR17MqItcpenPCWvMSSoJ3prurUwf9Q3YtCocU6FcoTUCvCgfFnf
R3rU397Gj4QUOsz1QtRA64fCKyz3CQ1i95Bsi0lu2uR0VJIqujO/Lyze2tYZXbQUPKcWUd+bJUxj
qhlyb4XMVOwwj4elBnl+jkSQJj2w9eeDfQjh4dKB1V3j21Wvx9u6SenyHRzlKHvEd9BHk+Me5tmw
jnSN1UkmsaMIRyqsbSe0TEkc6D/kv691VgV/HOQJIuHkJvW+ix5Ud09gbKHAdI/9Rf/I6lZx0W+y
dHQTK3MycREBJxEjoOTzR6e6N4x0ah/M9HJ0xJcPrAJcgF7gNiI2Ahp9F1WxHjIlEH3jwl3fcabX
r5E753I5SJdXy2w+9Pd9xNYZ0VbgCFHRYgAexHTqRklCz5Meeha9H/jg9gOvKxAAbrClHklX/Lb9
zoplavAou6HIGy2bE/dKo0a/TpiB+51mInpvFE7QR1u43VollCspCm3vzU8hXCWR6yDVq65sSE+g
+t2/KZ81mHd7MDvJRL3k0hs6rN+S4MtRs52Jv4FZlGyRA7U7QC/lS9gDTknXqR8dlAu7p6CuFu5Z
jpu2xtm4MfyFvqEAviVSSEK31Y7pcF5tAk+VJ85b30ybrYbCCEbwY53jakV86vU0pWVu2yGIHvXj
hNbPm+JGFiw+twQheMACk2HzsgIB2LJJsKMw40m/JH9+jh48uhLqdaBANAv/c9160jzMfruGZL0R
ps5XOnG+M2fQYfO50QNwRRxJ7qzl5ege89JAASDAGehzHwAeGXf087xhgO9CTQvV2pe8vSRK1L3d
k1aO7l98piVXIQVWezauycgbbcXnsAHfTWian9cSwYIfb7OXRXZKUNDOZEe7xjHNL/mjw2+CqyWD
f7aYyw3EUEIOVXKj4T/SBCKsFXsqrrxUiwAgGCSwPt9FHs3XBIjYrvC4BWlnrL9q0ksILj7/xSUk
c4z+ZPxusYV+GNUB5S+yNoyVPSyEWMOdEwQWl6TkY+uXQ+bZMUqdk7DrhlzsiEdE30YRI1iWm9pp
LKzRdFlLI6D+SEm5VUkUgdTNqo07KkbvEYz+w2HlA4aVGsYmml7eEIRotb8kK58PSvG+5qu5mKCd
/UBHKexye3955FQ6F3elVr86MsyLkJ6nVbvBH4fjaP//9irW1esdh0EbswxUGPtv3xhe/C/KqLCg
ZLGwaO39/RpIMn3In1C/qcy1JUSyFTJhZ39Wara/sleHNkx3nh46e8tr96DXI9/0o/BiCMyr03Xh
1M7e/ewXtzNKqA8ZwEAIUZADUK1DgDygfpSFncOCydMhM5DaJK3k5dsUbbM7kZonFUepGH/btJQ9
RX/ddKDVsGm5y8QlARzzHgYwxd4iWI137ZA/RWZ00BjNIJ4mR/DhCueTG9ccJpxXzjbiXoJAZOVf
NPKacLqCEVXV/ioDaMsbRUzgA/V8c3M1lhpJBWtyq3JsM3tF6qgA/+vPyYTAxzC/0O7qOjxlhdB3
cyaLLL4K1se9Rt0xut30+WwxDNNgcXhuhJzKZxTQiPaGQee8Th72No6A6uaPUoP5cBOO/rA6Nrob
E15bCCtTTUjq5mVOzhwD07NWL7gE6rSrtn4KXPtxzHFyRtZULCHyVcRiH838GiOShVkfsE96kiZL
Kb3WQJRvvLrDL1erqAqNjLCZrSNXf2jcjgozZPdH18w7g+B0sPf96E/ZUmCYZ2vsQcSRA3+6qRvv
xzHjB/C21+Hag2NXVjpq9bIwSvqT2fnqSoOZ20eYqUA60Pkfs5UQN2IxU41vwY7bWVhTzt8xaBSO
sMTpDUgn5P3yWFZ5ZzZI04fSKOprrAXMg0ktaLHkavueEK9V4sgLJZyN9xXEQVGKcmQQ+KPBqpwh
96tEBA6hLxUJgm42TNEgnrGuA3Q604IvEuzBH9g8k3WkJ+RX2vF6gVszM031HmzmoyfbB7OaE7LY
HwQZ7v0PS8+agppJCCMIRc6FSEpLGzmbitfeSmep1UtfexA4Rpn66v3Tp1ntIGkyhdGPLbs4L7md
Pp9iymKCFOBChnDMultteKaei8p0sX/Ki4u2RWlzjLRELkI5j19TTQkhioaAJ/BlAc8HiviUOf9i
Vo8xryafVsSbKDnscx0ay1uTrXRZy7TqcnaKEV7Wo1Pv+w5mtyUq/0oeDPXIbNakPJWQOz3C/PbV
ZSo/Uy9xSw2lsFWSIL4B9dcfiGlk7uxE8hjgDTpv/fjeDkk8oAYnZRilMEqvnHB4vaiB7Xmu4B3A
xQrHtES+5lajEKmSQJuTh5bv8DO0bjFb/IfJOk/6j/qxwpuZcUY/efRTHZAfjcj1B+lRbq5WKc6q
IVyc3KzzOuHmpqthah66ssmzl+T2qs9qlXA6FHk1Qpb3pNi9SVGESVi/Wn10iqeby/52u2vU7/Y6
ReH4VbdNp0l+TUFysOSkHD6nnfIvio+O8czmfy2SvtYwtQqxYu6bSLS87mR6yj5AUHCK/nFXkkFe
fMwSmfIYM5CyQ3nXm7NiJldYIvThq1ElNW7LstBuEmevQnne4XwXu0zFsh7YZsF6H7i7xRNP19RW
PUp3pGy6qjvyPs3qDbsZZRPzarB/qVWEOZ5+KxJqSS3uiROF8PBc7eHaHJqnA1DJE42k3D++G/N4
ZtNlqZAKeVKo82w1HZcbeIPkuief6F3BfncYhDEx0LVx20CfZ4ms+V5b/jrNatWYKDsYVLEN1A9m
/hgScxPZlP2ShLKW8WQPjLo5ZaCuRXOKTGLbfFBzXkMQi7TEJOZDgMuJ6KhC6Vh/LKFpFEq8JEnf
mb8i1iBP6mD2ZL7cPCwsWbEIq5TpKdXowTxHPftj8flAlkOux5TQo0QotPEC1vjKsLZ2xIxC76R9
kKnwYx6VicB7Y+n8ePy7zXfxLtZaZ+rEjmRfQRD7kHNRQ4Av9drzspVbVsB2Y3MUOGWM/DVLrLJu
Jux1yFF9YTOcBnbX8RfiyDdLMmo944AtLns2hf5nvF0fKwhzsmcb34j4bSRN14buEYLgB9+9HYLU
k+OQcVdRIMp0yFL+yZpgF3HIBS3S871EPpLnw99sPB6MpNsU6yzFm6VCDPRKCEMTsUbC8L9LmWLB
/6gjipn/RnFezQI7A3Gw9bWpqx5+kBTu9ztVGZd5P9kAugjF0lCEestsLCIEhTfQpTBWYWhZPbVq
5vg/hCyihPk3iKKBKk+ZuOYyQ6wVLXQVmbqty18e33s4VG9uBIjkoXhiG0quzLXtM0E8xMdf/o0d
CmkwWOlj4LB3h6fpxthl6nGr9Mt5mMHoW6MeyTK5O732QgJRvvJEP/zOBfL6Ak2Ae6kb1whnRMN3
+hvT3yBUCjN9lITpYy7h38GqjkgCY2Y53aLrgvFslL/c74OuByQeaVaymW7hX4gqEobX6hDCBNjx
AdH2K17NvMgLc63O810R+F738iQvawIQKhrZbyMySdiUMuYfxs/953MSDy7a7ru9FONRKuYvKcQk
KaRnSz6jcm5Y5xYl5r+gF3EQmBHW22xYPMQEHmaNsyMGnPiYa+/oL4W83GGkDqbOd3uSZV20Tv+G
jlRHsherNwbuYPvtbfB+hNW56hjb6JjXnUde1ybRvL2C9jfd6/1Hj2BaucqQkLkviQFwy0NVsRCt
CpOZf+XBpG398LUkKZz9VABzy9D/hvJmCykCwkLdmVdDOsliMhOTTcZyni262mjtMGXzKAa6v+/r
kj8h+Qhvx5dzDZFC9SGb5RVgqqDGgV91s+Ae5ppgNLk0VBzvDZolKk7aCrC7SHQOQWWsKhmL3sfS
mzcL2lM0edHKPdxoFvnV9xN4BBlLuDla7HOwG4e2h8t9t/aB/jIGqWVa0qV8GSn4ujahfsmb/idt
11BcrTOP4GW7NPmILHS3wnbJa5/IIehzBNL85d8A7Q84xFpGqGwHrAAUiz2p6e7p4b4i1C2P5tr3
1XcRVcM61ipcq0GwygQFHODO6ImHzEStV6DI7sz04rOK9Eu3MtHOEAXY+Jcgk7Ix+N+gkqX/G5xN
PLESKUyYfVpre/aNUOF2WI3GPhlb2QzX3SdtIlAcgxKZHzQiiJMNYZ47rvWRjXkFoZ6OFlEo7vLb
B3OF56QWXWJ0/pop0Xy0YJ3VxVBuJwfZZy8TU8UMVUHCtnOkfI6FUtIzDzOzBbl2fsvDS2rP/YBV
kraUn9A5oW8EoDL2oS2U/fsPdMgdPFfMZVdP/LZ4zeUoFTHsipHqQmWBDE5mjVkm5NVdpLlDcbEN
RnBT5gPJsFbHbre7oE/RRlh345VTE4mjFZ6bbzL//vzTx9Pkh1CyMVmIqJirDWfMayH7vyFPHOTm
5T5zVVWPYVhIftT4CtkZSc+yC23UzyMzVv52PdOA6+cF1Oy7ZFdA1K/7vVkrRKClxtgsJlyACx99
jYlhsR7SKnKxBGfndWpydlsvgatW3y9lBUFqYnwx85HmjxMkog6wd1nADPxinhJ/wUyv6lfoBtHO
o3ple4RS9nqnzzaFZNrBfLFpoOtUlGFxjfVParAtZZBUHnAWBsDAYKwleOgoEw4AN40937qiJWfH
HaNPCl7rLT+cxVQ+YbBgWUWBa6/a1XwHyh4h2Uo812ZDJ9Aq1BtjoAjDlG/tvQlSP4kbHynGGawU
l/QhFzHHAz0seGcO+pLq5p/ylY+G4I2NfE9bjp0oFDEieF9sg5wZXssktOuqSa/ZrKUZc9y+igM5
T3KfFbR/ex6zWp3PVJWEDAe2+FRAiKGVq6Su33xwv7HgbQ1n73DLggn+krNSR8fl30Y1N5S9iCRr
wDTdxfUIkRi9uvGapiBBBu00mAZcdX0MtaxTG18ZHyBFXUHj5SMtCDqqwg4vpW4ESM50C3IN1Myi
frtmrGjAOb5hryu0T571WDIkpY3ffda7zGrLypwSBc4p8A9hWnVJF3pNVhv4UqFIp6SXKzl7UtdU
l3Vvg9V3TmVLbrAIlbb9xxYHAeM7gy7+PvqMj5zbvM47i6ddNtsUYYpCckgnSq2AJ3nCsY1wgXpc
5TpzF38v2yzgGOEnLvkYfWcsp+vdjXGPOBvg/h4Tl40xsGr4YpFknf4SdU+y7MMYlSxwLQfEeKDt
+Oa6UhPcFYPpsVNoYvl+ywqQONs83/G8K+UT6yw+yO9RyHzaA2JGvWqGxEK+LYqbxiBByVufRRE1
yLElnp4b4rHfvCdz8zD3WagQLki+fKdjS1IQSmcqR734pOtdLqW2FNWabHd445GpuVDMmxgWjI04
bd5NOMoesgFD1dneTUi9rwHfBjUTLfliLAQ5oAYzqs5Iu5Wj5mA6NAHhtA6GhlICZ8aTgmQiPRI5
loRNpNsjssYifnTwzHTi5D9W1p8nR2JIRQ1N3oPlZcSrcRi48L/1ErxrUpxqxqdHVd+fmvg4o2mX
jLuxeS5s/hrslWHi176F+3xow1zXjppKqByicHNW43w8ag7bptoqinGkOQv0bFpdYr5bRtQUlr3d
7sEoe5q3UUZOEKSmzX87aX7W4z8wHHTclIx3EG3lnUHN5Zo2hWlxzpNt83Hxf5keelIMWqjPMEh0
+At2qdOmcyB+ndhe1UwjqaCy5PQcfLaXhCeb+++T8+ihPxXbfBvSaW4qYSFqQXRqtLoJlH5LdsIY
hcxjzuOI5uUKPIa2WMdG3gTuKwPudNbn+wto6Hi1qzBiCxjB7aHra2Gf5qH6wUiOyoq+g0GZLGxv
p47eh00eb0PhevAmdgH0+gWFXbZNi/MOeyRwPsxnWfr8xX44Bnh9j3bZlmd2AlqvrESQgsEP3RTM
yIok6jPXBrbHuiqM+O5a0nuI3evnXqsEFIPFQ4W6CuQdbbCLpM7Zyt7mw78y7zY/cjv80OJYcUQs
tVIj7JLvcOoPNj7d/yBsWNqG1ek/i70ucRfwLAo5xcNhr5CGCvO8P9sRJlLvjoCIq47TUVGG14YL
7ubORcOra9gYPhygeUrFImxJKaWDRQm1WJR/ODz6q3DSXWfSqDE4Nl5WY88VyJpSkVKMoqJDVbi7
s8FiUCAcQpSciqo+W0hTUWetx84TETbr6skjI09ah2mdMQmLufm06WHOxhzpEzfiAT1S6Em2aOOM
dSD47kuGir2ztR6hTnEyVWmG7/JwiczZYcdFbmmvaCn3k1qwH1gFWTdIqLI7lr5ZgKlRBmnRsIZn
pSYUQx1WelfHWXesP2no0LbxBQtRfyxD5bMXnC9mxKRO0eabeChRo70QFi3jwZFvMbbSViGZZ+2a
JylrJVsAgxZUO7P+Su0YCNojrulFO8j7CPm6C7kddY4hhibo2c0IdbTv5P7LzsN4jzyCFPQLxASc
STqIv5PD3ySZjNArnahdCgmMEPaV+6yhR729j60G0nuXimQeEzQNiWLiFbsq+ryJ/qoe1Gw64ElJ
0d0rTJa7+MS2VaRV1/PgIZZdbBgOmnABhPymgLcyv9SZN9aVDR39/31ta13+wP769i46kuuRPPiM
+GF29QpaO5WEhrkPDJZfMVBaiE+OSfBczgJzWtBCuAHmFMT8Rm+NOUJPEO+JHsWFt4+3gB0MZECF
UrztNZ6hGglpj7dhlEuGVwZXfnB1jJSgerv6dg5rLrTHL/Fpwn1fng3u5whhlvfSKX3lglGSvfBz
+yLuoAQibgM2WdivJ6iQe5aCvMVW0qBKbWhC0ma5U2C4FGPpcrufWo40Zh+2BG0qS36nlvsfIaz1
yt+7uHrAdDWeniXX34LI2hbMtoS+qF30nXuTXJEsagCXjYJw6AH/YYzDAtC0GWg7yne30K2NC/IF
L6LuqC32SZVlIG8ytVlGOjbQ1u+MgUUJMKrlPpnJ6hcwZ1jhiVTB565j68vqmvUGsYiI2OOM51Zl
JYD8W0RNoD2YkkWTcYvoKkoAFQ2XcBjZPhOotSxaayRKTeb8IFrv1uLmkKx9aga+ICST1pOQ6T8M
0Du2hk9ks/9xkQ7shqSdkBhOiE+xsb0rbKot09oz7mqULkoT04kmlcMozeOYTQBmlC27EkiPTGT7
zUKlJ+/941JENryIQQ0EdvcQMTgFL9F+LzwcL1tyRy9fJSAGBd4ioQXEN/yQcs7TkniMM63Ah8bn
7meOHxwbUkxH3CzJs4cnJgttJhnJR82h97vlkBLgrFnVx1B09tOULBLgMu/FacQ0pNSnOAo2cKsB
LpBSv7wZRBvcjjetKovRr6hQ/Y4ZmqsEXxNg0WuzJusQ1o/jly7hWnWuvIamnKqtddzJsdBvLEx7
tkzfJRfQiAvHCbUkZpVTs97OFvNi4oJSw1DwJnECzzT3lv3t5TNPQ836LywuD8qsZILXoh492Y9d
4c+YBY1oljx/uXqkESLTdK0BxOCcPU93TB9A/9DJT7tU4y54c+h1h3VLp6L8Fy8oXsEohLUfgrGk
YSxHbBO2lVC3bFq5ZreG0QxB3/apyAMWaTxehrbZnbgiRmeiqguXvivKexE422CmOGDWhKw/trY0
VmSACH8dYB/0OmARWICymsPW0ih7zxofBRYnb3jKPeScbCHGcxxWm/OQhD+9Ci+NVQpstM8fh/kp
yxbteGfV0q/htqZ566sqDKGr+Rtjibjei9yV3WRk934/8xWif9Ne7GKHGmJLGJxKlTx4dMNFQ+OR
5oLnank7eddyiAkj5WFBAHfLZkrJ/8mF4J3CisP2AnmyIjQMZTMduMy64GMroD/2eAtUV+v2W88U
NvdOqzJ6eTMzQN09TQivbAlvMysZMKbwXfx4NEJAWh6reVn9oeYOzlUFumf8A2YUGfAXTEislfdI
fYFei5aWaXvxxP5XCEXKV2rZuMlRVwnDI58oztl2/Vd9q7Rbo+YUorWwqe3+D3t/I6R5bod5lEsT
VFKU/4JqaUBfPYkGF9CWYGpZ0YJ2zxN9f0JcKvllDK0wkJ5VptOfnBeTSzrw3lO+vN4N61Lu/0s3
Wntry9acoli6luh9gOHYxixobw+jnMz3R1B93rw0ermb7CFDVynVgscl4cpNPDXLtcldw9ir2oAh
UwNolOPArUqkQB03zciq4tAtdI2HpFhFxCWkgY+wMw0O1NWk911jlkftKEBcgm/2HdegcmCOxzti
IzgMeU64nasgeN0baQ7o3uod7U2OsPJcNmq6AgROgGDM4SCVEckq3dQrT300ja32k5QMKwH3zJAX
OGUj8oOrcUPxioHj9vWFaJ32Ph8JN0qN+eqczMyGOuwdPGqzRqcvI5TpILVRSo/XfRsT1kCRpEiM
8FdDB+U/iChEI9fCRxQou6gWjcWFAjpeKyfhami0il/K44uIjMZdciqOA+tD6TjgpCDPtc7Hvn5u
DC1BeLBLfOlclwt38qjDBtrZJX1GrUDUqewRWcCZFzf4mRd4gEM76TSymutVHoE+tldaCzsmxlN8
2Aq9rnv5jBnJBVqzMcNBSoSdet3RTWW0TV6IKVW5LFQ1jrQm80CQ3KvDxmCBAOiyXVxEpKIJm8Ij
/qNT39fSrzGSUkrP1mDz3fB/7enDnIigeU2BFEuwLOrMZYMUfZL6dxU6c7m+r4WF19ocy8T/6SPS
YAequ/ojo0VvGpygsFw8/oj5awpba9fXVoHQVpX4UNxyEfcYF+MXXX0Mm+UFQVTjLzHG66YJUaOT
4iniMAQMkoz93IVsvDw/M2Di8gnSUcI1aVVROQJVqWQX4qVA9Lo3IMoL5TPpT6hwNZcWwoh7PPYV
2TbcmHVhDGf5JaSXb9TcmE2gSHmToWJ26lOZdiqix5mshcnC6yQifyJY08FS0O3tF+kSwsWpApwY
9Tm+1URMIpMUzYY4VrjNxXr7DO6RoefjcHy9cJVEB0uqsLL90UoWBJFb73WZhGt25SlhSdAwKv/i
27TOkRQoCxkn3dSctMlg84TL06/ubjJ1upYhrlwCsKF6fUcsx7EVAF5QzseM3XQItTi8RLb5Pv5+
dgBRQx+PaQnQansf0f3gjlVlIUN4VmMcxGb8RDhKDLs3zlT/KwxwqwMi7ojIOxhoUG/mNSRM36/W
ztoUX8GpoTY4C+stSRY9kPkMae4WLSsUQLYgGX43ARExU6B7xHPn1912sq904QO6kFY/9V2p/eb4
4MoEE5V1JmL4ZUh9oIVzsElcY2UiHyUBHy0CwXY7kvTbvW+q3+xqaEU+t7aWGrVLZoR/iJq3hoY9
cYsXmizuL/NFRm565u/E/I6ZUL77Dfi5q6hQbBPib5xPJKjnN/fDrImHGbvUjCfyg5Jd+GA3wn8W
1JYhbbpxsPfEPGVnztmSbJP15ZZf/Qe0HPBhDKT8/rPzzW6PTbDTAVRONmYjuHyKERO8kgwuBhc3
BeVlwKrDyyPzYPek+B6ea2TaAqdr3V13Zb+//bNuD8U5s4OairVHMp6HOsE10ixwzbxjqO3RwJJM
67HT38CpR0RfyBC+xf+EST5EZBkBcdV6yDsuNyn0A0cr8UuY2LDf4sGAnEn9bgDz84HO6Uz6fByu
xoHX99+dGe14V4mxXI84UBnI/PSvlHPD6OcuJ+k/4+0CCVvA0/z+4SdpaF6O6JGvlmBqQtfXClZS
zuUlJAprOCvhSPnlyLcS0sYO6TuL4r0XvizA+KIUHU7PeFX959XJO+hpgeqAbR+EDLB89dIH/2if
jWW/N5aJlYToKTcsh1zvWi5+pItN72Hbvd8mPcNNc9klprYC2UT4USb9B+E2hAODsxMtVLfGG50C
cvs83pEVU1CBmFOVF6uVmgLJ2bhwYljR4QBty5bSaqyNczccyPM+0ednMjUOCeYbZBcbXDVie4kK
K3/LBflzNUk9oxKSV4qNqG5NgbzHqARaxCtyKwf07UtAaN7jTK5PcU6TOhlGSpurFOH8aGhL2vvR
NOziPsshf5UKITZ+fFU8LR2bWaBhsQ11vBorV3Fsbzp/7f5ZDxbx/uOCIz6cQ3L2ICAGlE/GM9jm
wOeRYvtWH5QzhHjo1Oce6zdbzeRIKLOcy+0PFq0N3m0lzW61rYRrNwHDPZ1RFKWcBjmKi8/dgGH5
mRobqHTNB7xea7WFR7shkJOI3mNHY8soi6PhQP/TEn8YIOa6Q50lu1pdOPeumM8Hf0G0yOcvgW/n
Hy5OQbTJ8QxlqvR6ctsRZc6GtyqNGMpRQSPtDSmQ6Gzx3BirV81OK9aTygGJbMdf/LY8mgMmHJza
3q4O2/NPZL8un3511dSKGo4f5bZj4uf9NpxwRC/1FRAMuhpPLSxV+yF/mJURkD4nhdZZRkjwwEGK
8qAH9MWLZ6sDAoSEnhwTDi5xAukReiQ6JyVZRS8H5GzHjfkOFTNk3CefB0n33/bKAOzESAKUWfVJ
BOvHWhSRGH7f8DCsPUUQ+2GcX++tVzFvg+BlQ2cQWr43cDLbuMXWLw0vCmwPA4Zr7MUGWGdy2zc/
gtcal2+mU44YndirQGxz/cA7J28Axa31qkmnfTCQCb0Uoj0elI+9d7fnkKHqdgCBbFxKPbkix71B
LIQIe35gVy7AVPtSfZzrxUZFjbTUTAuxkoFrcC6Xo8pOqe3LRMlpmImJ4NQICI5WPtBnI4SVOSjF
eTJbPpu2BZMlrB7Jd3q4u5+hT9VpoOnLW21UN56UdSoPplcoN7qn5KHkRWNdY2pqB6Hj74S8Z1ZW
Wpi+OiIOwoFUpHb5z/7GbGPcHQW/8axylcd4n+UcUFS7dJCXCGO+Ge46qZxNhwmSP+0tNSrDwAFp
BtdOOJGp2hSkXRgsY5euNerTwRst2QgxlVhI1jVxPRUNMIsDft3qW1zQGGyG0UtJ5aWIGwchLFZK
1tHvg/eV7wN6ZSCzbtI+BKD7/g8mXvGiSssQxY/15LEYMRFMPUJmQgtke4QeKqNK+MIxuHIUHOH1
8qdOlQpMCMUdVxfdQbKaiJ+FZsQb/W/mQxmIo+EXgxPevTFVj4pK2RSAQX7CGpCAOEiI7IcbKtbC
BvkyM3CKNUFZI+b35bERRuSzy2exUJewiQ0GfCWy7Q8xTGEvZJP1vp5ZyKYLJ7jU3K9vxHhqVX8c
mYBuVjaUU+WNk/3/V8ryF6VeWmW8hXOduWubzjWlW8iPBOP+fhnDZErYnzOz10NWK2BIdN4QJ2CD
90CLs8qjV04Lah+OWGKhNgrKB4WUAvHRfwto8jJkYs1Etff9cJwfYS2gBlY4k2dxth7xKx6JZcV9
E6VplSlS10vu/+yu9nck0GtfJy3kXomzD/UplpBy+x0yiPO8IbyfHI3oqrjsV7M4kLD8c0wrRChf
qLGRlMBX3c5G2Kn7UVE7RiA3lpzcxT0xE6UcTmSqRdMyPMIO2rNCOgWZgU6b89SVVC05h18E0koc
aMkEpJjZdYZrjcVljBrgAfVDcYMRC2CtvGOs1hzlVwNi3kzIYnc/O+k6r7vt2ZYCD0an6sHOGKyr
5uZUIOdo2JM/C1r9Q+umY0SBTCO7bKfraCCLEkCb+hKb1IqlKzBbHWZtaQHanD1fQ8bJr+AaAB0L
k0xf7WABtzn44M+XI/AbrIsAv1chqBr5M6gC9LL4wNC1/pU2+/V1weMQH2tqtc/31eCy7kSkvuUV
QUjyvkMT4OpzZnLEebQkzzxs61qT/ji4WhILZXWeGu9/dVhzPhU9sbh1aG8Taz64rxopVEuZpobS
J01Fi2Nlk30nLiEfBFBDkQjgmpAHP/dnsO3xkLhzpJe43P/UwNrsTsdn+dNLTJhFYj+9FBHyZTVa
yOtUZLPYSBcq9t0U9fmzFyr0IqeJn7xjdB+65bNxr0yxnLt13dUOlIRzCJ8piWl2E4pnAqcniOER
OH77S7rcLRAiFJ6bI2jKsvHmxZoU/PTZs0wAYt5tfl1VxmrXcHkJi/Ndi7rBwmAKKBvr2z8/ulnW
iGtMLZHnww+TR8j93TVcdPObE+hZP47pof5m3GRmPRugjiIgI9tZcDgO2ujD/nb7uKPAyb1XY2Bq
AK94Q6uAM+EYiTagqzHGDFeXC0YpcKnsBdS65PUP8336nfSBv55yUoHblSrPwK6mdlppAwD+uFvJ
v8nMa8MxDZ9CT9UFXTICqZtQ1hPWGozdr6qLmCrMHT7RiK8Nx89PpUwXeiJZtZGJ4s0VV0Y9RU91
wpObiKziJUzItpEmvD3ih8SBLjUPTDSJ9KbCDVt/U2406GsXaquJt1pRda99K0OiaHOcTk0JEqau
rBs6t2/RiCwR9cG314LBu3jxDzHUxIeNCCAL5ywZbE6kz4P6qZGjjhr5+QN0AyydfB/s5CQIpvl/
tHbTfpeAD+VaYTPox0CNY7VTVKSecShzouwQ2HfRCmzbxl8PT0aZaVLzdzCYHstzH7QqRX1lp2oa
FlUQ24ybCtcOK7RTKdF9ry1rfrdpFgSttmqSynvikzORZmnPrS0xuoKffUZ0d+dU38qKw4wB9VPn
bTrN+BLxO4d0+fZrO8vfz4yDIPPobdqsbQB/xrPpTaDCZjnFUFKB3gfgzEmKaI0GyDSXt8lZgUaQ
3Ip/Zu5fBELeiZnscCEyy0hh50mbvz6BJaUoSmNw4gSOpG7dlLD90RiBDppQ2hHHB0oVn/+saxf8
Z9p6Ioqs1g3tA80gdGVCaGucIKZc7/3CNQP//YVIZCXWKzioZp4XzY3wxDZnN+Kp7/JCVQqXwy1S
lKkKtejvu3pzfFUh2ELXqGvRgyVxRJoFpEP4oVvoxXzbm3xh5VdMXqCdBxeluj5MmcJBUVmrazY6
98q8sdb9ds2XbcgoUUYoWHN1sntk8+qpdaqTKo7Dx1oR5LlTVLJSxMqntrfy2QrZXX2ZZQLXfQgk
We18Cu2OgcP+SEXjVJKjQlnVByH8/sCi0Cq5SnMYhryRH7Ev/aZF0HsX+xhAfuzOGbhf+xoVo14h
YftnyMaihgjPxVtDYwTv88SMoLs5+l9s0NIyFqbOvgHuOj2nolazq/SnayBHJz31L6olY7T905tq
jYWui4pM9kb2uJxTIYcZ9HCLc0y6pdOzqV4lfEvSxhhYDQJjKgo5pQNiPG42JFXuou8toL/FCwSl
XnRvsYcqn0iyT9C9CDzdo2ariUwK+P6a4qCriwwGdSpjZlEJ9i1/dqILGiJHbJnwcQ6Z3dSvenDa
VnyL5y6OmE8DuhaAtunoz+0mFSxK8kotQdf3hH53gnzHSUf2E/VUBfRqSqS0uAJETuzEdYetVI0q
rpngkp+7D3kU5/Qv3Df4RY+zeVEABxbYZULnkBzcMdFx1iRHXvS2i6PlHKWJ3mQGRqm8/CT7p+gD
kSOZFPkNqkOaZzYWhz5ONob/QPHYG1jXNIUN8CMU7FZTnai/OHjZZ+fgYLELqQodSIvDWnQehHIM
JNUK64xme/QaMyjFLzpDeIjJj5nwB9F8DEU1GOQjeei/96c15SEgP+Ms8UQKWa2wXpiM+eHnKc1+
4ViEtlg9/o0pmj6eqDxI6XigYRDFyIrINVv+kYbNz0l+Hsr8K5UYAmjlJNv7uovFSTZgtFc5pDdl
P0wk/eSyoRFJDxkgQ5qe2H6JiyugCrk2LjVY5KLqCwXrLyYAT69dzQd0JOwOzAoTZdwz5Wx/B5zE
AJgAWqujfIx4BfTHGwLfRqXstL5lAI1u967ECUPWE9/GW2JTl2KHlW/HJ94X+FaowJf0d8OdITSL
YVyDDk1OEYtRlpeEZWvsSJ4iOYSjODbpwH3OhGxu155eRZXmD6gfElGk65oDJyys6Y6fkbwYdczb
myxNFrdNCQ2i5WjS9664wwF6OI32fWdo7nE4arqeVIIFAm3JO6si8K1LGf4l37ppB9K3B4Y3aE6X
4RBg7uB9/vXXFM4NfW+spG9JkcG568QcNZ74/Jg1bv1LjpdOu4ttNObuA5r90dSfLa4nE/Nktl0k
eQpilsR8VdfgJRCc+9zXLJUuTiywoLFEKu3lmztFCFgIcdD+sZ4S/otRGAGEZvC557MXA3PiFcpF
rLcihD9wve6WTRttg4ar2qbWjTyCt0shdXunw5GLRoEB1wv4/yW/iKSkV3yVVeyF+u4nrcbMjnCH
VOnOvneav6a+bUh0WzXrc7N8N+nV3p9w+jlGTlIiOhboV5CWRZx8HchCsjc08j5vZsnYwB9I2bHx
6t1S65SD/w20GKE0bN4s3FCzDaoane6GsTBoqSe4g9FLB8/jlCjZovpNfXxq15UiIrW+q6TCjN8+
u+EbW1NAbD0SkeUugCtX7NAKXT0SkCNKL4J6oZSCU8wBA2IVrvbYfyOB1rV7Y0+t2evcqpOxyYJi
YRiMvAZzLtbP7avjwgeIlhX7BYFLvvluGFraxbqVEWcaZ5mIAYb9ZgL7DV4cVI/5oX9KTzpl5fLO
q97IluFWbI0ubz/WTuibUVx37l5RDFw4Obi7GA4XqTsn9wke7B4mFWQCfP+H7BNNErzxNvsxUkqW
ndReXM/geF3RvHiCSpe48bayWSBr9jjhkAuIcw7UD5P0kdTu2Mou4YrpjFwbHBZgF2XQuv6EZCiy
XvNcaLl5BF6xuguEqABwxdZ07u07obuFkRIKjttF+beFx8VJedXKCwCcvs5vUiyNjd4vKbQ870rc
XLIHq9PbKJR/uaR0zjXPMmNMWBl1rj36hcb9x/EgGnpT9B/X/9SJCeYKwTXadSOOmLxHcIEe8vnj
pvRPp0euA7RAgcr15kbycBWUJeI/mt/HPHzHXKH/Dr5ZEEcXjw8l0BuDf3v/xVxh21On5Zmuzrsb
uvo+u3y2og6a+PDtuMYMzGc8Wq+N/stM/4wOJK23UZEDm2EKHgjLMZVHwVJMkb9hH196/jKgFB1/
DBibM0vt53HBpWBdJey6i/Qq8RubWH7j1o5+zFVxA1I168wFqo8Ak4mU0mkVenSOA06pBqx/R96M
bpd0djhXHMPJJ5RAsV6Or6wbEsB7xJdnQa/FPK4DV5jt/pPMv+dVsZIQFgyF/gL7exycuxLlpPt7
8n5IlOi+HhtGQqfaVwvkQqds2oOYVI8YteH/XlZhCXtGBdzkD+rGbHwFRPXulYZ2zAUVlAnrk5PL
d56t9QhOi7QMQTdgLYOjHY1e1w02HyYBpqN/NAwcqgj3bidTiq2L1XT0UJ7iF9fVvoTKI6HJSlCx
cvLFuNn7uVVJIAY5CbZgQtAa+G1dND4io17WtgXk2ZCp1MYRdYEex5SPQN6R+rtbct3myzsVdIT8
Uz75u1tTfELNIHcMBcvrMhYNTZdEZOPi+Vfr3wBP7rB2Xdb+kveuPjo5771zbZ5CmLMKO8z4bWzV
+YswWeMctX9k3/ZOBtCX/G4Q8L2oE+HVouEPMmlt6u7oUG4stByGB71OzS5GPyE0nMePIWDCYeEu
ztUORZ90CJsd5ZSd5SpMZMHeTxz9LESaboOxJpLzm6X/8rAkTq78v06To3VpRYEgqeqzGM0MsX7d
6SglE7trcZLLxvpBSW722bWoUn6V+8V0osYluJ1tmV4YhnAW5F3OMeW3bHHFhD63NZYEa3ImBtRu
Ap5G9VJuMDimMVGvkBxLnvzu3WE2htDEb3b3z9TCU9YXyKJAtqrVU5Sgznq+49v6t9IqhbHDjYB1
oTYaZnLVKMmzrCWQZs5oh7fZ/2Cz8aFciwQdBDhSBpTVI2Q+Fxn5SQJlTP9zgKgl258yoj9/HDl6
swqvY605b3+Obi80mRxKuGdjuQEX81Xxgm0DT+5uWwP1nazbsDn3Uh15zJGH34fJrX3G8QvnXeHx
SEk48f4qmCPoZ6yofvxdQeJsrpyWPAtHk2PURlah7WIdd5Q2IZ+hEhkZoD1rSbiInjxItLJel7SI
XM8n5iV9IJDvpu+TEDsZG53B8qibRBEF02NoQGO/o07YxHYH/7+p0gAQiDd0eLxqNwuhW/zRWbbp
9akg87j3hAUZ9m7ssZ61ZglhaT9S5KCxU1gVvrU1GJIyiS6XgZ7mW5gHShVSF2UrQyOXc5/VJHem
n6PRRU4nWFYj6tXXKR+0qomiUHqrQ+FNLbhw+6WKs5LNFsCRNm/S7xdLa7gHz7pej+C5gxZ5zpg7
KZeOGUkaDAt3wKiXpejgToA8hWZABDG7nQojQ/7AWn5PBqfZIUEI7Ywh0LxLODiAB09CXBrKxpXY
PzpH4XzaSmmQZ9CEpU4WC/7qpSgRhPf567G6q8N+Dm5pegNG43UG9nZieJA1sj2QbOfGPOXf8En/
0C5C63r8izyjjgdEMCMNw/dPy6Tt1A7ApYtJxpqWPDv5w9X+KicDTNvmRihtX/A4ftAqItzUnjEM
4KqYo1DA89MznrMVSCe+0etacNb0msWKGryCcEWJ/2NFAsqCK8Fhn0l0oouXOrEdW4y6TFKHTdYq
oKZEPfHx5tR8FnOrZvGYMz5PwVm+n++KjFDMtUHPWtzX6VbaufUswZHUq8eMkCGImXS/eVQEBuFM
0PUPB0sD5UXeVcdE7rsw1EvSB82/Xs1HRexdReVd9POf+zbDisKPdUXzZiz/bcUg0Kj0dY2WmEak
zrhxp8/kHfEITRs7ioHGsHQyXfoP/JS5kp+q0xUMFli4bqLl/qPhDVXcyb0XRmVXs/zEnTmVg/GG
GP1IzUYQo7iCm6DYAtOtoKSlcsV4TpZLYi5aRqIRD/7qwss+GG6wuaMMhd4DafE2ZrVWpAuPu1af
xf35WoFmE4nq1fldM+Yak+CfddwlliKqG2WQopjjYL5QogMi8fEbFQZwXYjc4OuG+tZrqXyhHl48
1uwjDVhxYAqfbEXEfkEkKl50Wi17abndy5U/3h74SG0x5byEVZQlADXkbftiOTkV4nvmA7D4Ql4n
3658uooWeIPS8OtGAvkTaHXmYsZcdDYTBz6PKBWzMXie5gi4yNiBjNYeyhVOXxnTv16Jvh9Z1xQA
UMjH6GDjcNoMaJiYOLVS5oUvkA/+Xo94e+7wNYxSWVgywe0gVVpGgcbjqVHm8YHxTCfRr2dcPnfc
aIO1BSOlkZ993dFOVVy2b7qkn5Q+LOy27czzNXdQeOZcXfwD4SgFqutXoVI/wzhj+NqFnsRFuEuy
Fybe+/nxXLSuCrxzqk/ODle2pj7JUwSzR/Z1s2C0cIIZCjQqvvhnxTPU8OAiZY0AsVIqJ4Q7TOUi
H6+uDtyET5u3qt9F9KRB4Ez7ziERdxl3Izr7w4zazdWvxlG0xbY58pOCzpbfHf+4KVjP0K+oJgni
97hwUhLgNTOlUi7bfg9CVLa3CrRdNDTJ3T4ryFLCSCqMNyMQpalDtXSJV6yC5EbMLVcMn4LMpB8g
BPlXSdC1ZVP0p/zk1C4MmGZP4zTYena1i1rJcrjNO4hu5jBaXjJrplrnoDqw1JQfSX3ddcwHNx18
m+iAtsjmKkhkw8XoH/wxrF1TW9KohWs6COiYDLnjTOQz4+n5I1TPpqHM5ITJmFqU7a32J22W+wsX
mHlgkQc/B4PNjE/uB+XR9rJWLJk96GOMCfBKlphCNx1juUFuTQBODSFWkBm4xU8fDOo36KPhA7DZ
FaZYYUJXzr0MQqAk7OPAbXQNMNtXJ8SlDOhwFNMNv2Bn90p3fMeYgzS23z7h/RHEn3L52wpu8/Oa
cJVJ1NlPZxkJbE9lezJrsZEEwUt85FiUlB4TjYM/A+iCyT7Kk6dHEfLjTCriT/Gs1eWlaQvG4E1z
/kiPEsMmksvvUveIYVYcoXimksk+nf6V31840BPLIhFb9CD4GNimosSMssfxQH2ckguimMvrMTDw
9tDFeTTS2wuhtY9ST0W9+1wM0DaQfbcqKnK8wxFepvyHf4JvZrc3M+EGlR3bCuF2X4glQ1dpIbx4
tmXQungManDlRX+Gf6N0He6q8kIM/6x1srhnX5+O3ep98O1HSQmMX2TPMUoqWSOiBxkUsoYbzG5M
2ked82ErClgyrZdM4xGhZqCachzbjaHebciLWSTJBLhdRuhKxfZ9sHpH6HDs36+9vEcY5pcLu+3R
sznmNCEkVVJVOIb5tayYHs27oUdyGqeT9Mz+DANFaJ/MOBGpPlo6pA83LIz/CG5DR0vK161VuE2C
/bXiO6g7Bz4vHf8+J6ATCZWH0oTzPe9udYhqUzjUiVSRo7IojQiQgalrrUrr2qTgVF1qlYEtVsIM
jJn7FbundTOCEl+7wXf6cpa04ADmSm0daa96IUZb8Mie96PsHtmSLtejiaozQsRu+d8U6+sf6njB
3rd5vqlGG0gXxDmC6ugJm5+gjdACJh33zW4lFDD21elZkQvTAAM1l6fTwcLzxYfw/cmXpfwiWY9I
Lgg6VLEl9Y2GxqOUHMQfnmwUz0uIWdhnQGSPp6dr9I8PHLLTBBof2Oub+KWUnnLyKxQtUdQibOJB
ERsYR9NuaUzUL7Ai9CYQG3BHiwWd1FRdUZO1vNOTum+cyhqf7HyiL34NVBvuGF3TcpaejwjRtI/s
mR4Y0J3U/POqfpMnXFadC4i2bvVt7clgxNQQ+nInOlYc0P/JFPwpWJKjRC/8ZZEEbAjB5N1PN9NX
I3O0vSq8MWm6ShbEtzN6euFVzTpXjyP5ofiws3boC+q86c181JN35G0JA7yaxnXMH3zpSA699YjT
dj2Nw12FXOJ3F3uLvayGtbf53tccuZhHQCXZ5+4zhQptZAihLbT2uj+XrbPFwwwRvp41QHTDQoup
IJjnjcYJ+zbhp/DlDpbGIjYdCkhcW4sIyg463X9uE/uwIk+3gb1b1HzsSVLkRMLvluRhjXASNE/C
nfvASl1RJjDbPImJL0h4Er3zkqiQLMSCKBldHLEKR+9aZe/D2t4QCCTkRQq1boIJBA7VHkWJqqRa
IgvtxpUpRkf76jpZKSJaHU7xUwdqIiJTxC4xubYs1PYOytrE0gz7FDPFpsO68v0W63V+Ppysa/Tr
7SMkwUisAEOzvmyLae42vzR09dlYImnfTYvSnKshEdb5FlRIb35j6gRY6jm3HuHvsJNO0YoT9+ji
Wmphnn7bOxHhY4vzpWIvnuxOoj/q3rD5iKDQtyP/j98DwHvsunTRJBr0AfWGJLVXonWvX6IuPeuR
XnpxvNECZu0kgeA3QsPK5kR91QKM1GVUl0JRVWeXKfLzmrtgQ8t5b9kaam37+tTGb1uW/Af2JZ+h
759HXrbR84xL7j7ykP0Tf7ugK3OFLos+hrtmsFdO41bUjkEbweLip+l3ffV+jfcNCJ5TkJ8ZWBAs
SqhWzzgsCBUTvHvbfTnEhWzHeK5vh6Khm+a3pasrQ76bomWEZlpKa6yC6FzcGMjPM1Q73SlO40tJ
O8ftrT2IAv3hubogaxtJTa6orDD+DSMmBxihgGoq72Kc/THTk2hrvfB1nB0l8KcR449S2CGad0Pt
qe7Oy1tdPJYmCwFCs/aG502lQE4w0E7G1lvAHbBM+MtXOHmTPurFta7LVhSYFVBlp3f1gaaYidmv
Tq81KH7x0ScnWD+l6XsAOdOX0vdS0Vy8ZidRgSDpp/tdYux6E9eFdsC9iSjgCeGdJmrvxdmhXlAm
wMuguYrxPNidIbMZKJnmKKmPBDrzON1Bgn239qRQkO4+RD4mL5rsQPNDSzs7lXGJkPX/iLD4lW/o
IF2w9yr7sQH6/qGdQ3jv8k0wMJ0YlPFOZtIR8vzA/fXdbJ5kRDL+PsrbYvkskAybFWxLe3PHurny
mPqLW2MNPypeceFbMpSx0W9qsZtyLObetmh7piqqnSPdLzuhjHG1zMmM42jD9cgm/9eI9k9h/aVB
kBpaWU6HYv0ceifb4huQBdW+3Kmjmp8svLCnJlt6OaIxBNjQqSJ/86STzGa29VNSeoEy7aKCZ3vE
rcJ6dUcbbWIqV4Z1RnlciT3AZlNTijJbdtp+OUioLibRwV5fM0g+3XCSst/8DLo7jz90Y0zZJ1rj
r2RiO65VHr5FTH66vEqlv8jSPtFMkmW/gzrrVfYN7oq/m27oAOw/r/30Yu1CSYCV0u536pFRlONw
3H4vRDSuKJ+qOEkeF5yLWJmcBG8ihPTcko93TwmbDmW3eiO2N8/dAyUR0boOxllrRaAfZzyL4Org
NAo9L7Byxkz5a+JShU9HJlASsVKuHP6UZ3MUyuhsW3A/CwtUVKYtyXQ9e6Z6QbPxhUFWF0nLiZKs
nLQCTJvd190kScVYkd8L24AVUQGWwXgQS293Pcm/oebzsiRfdjRVPfnfHG1Ok8KgvB4JH7E2oxBw
Khhp7aR+K2iQuyIZfkhwDk31RMtojroInb4WflvrX2JqFhOY2wuvFmvY8+nUzQHujojOee3gGJ1b
mGFU/QeBFyzr8sM1dwxbtS9TEW8Km9ZxCZDiFm6ZQRGGI+OitjomLyAOhiBKeC8maJQB7j0lGbAP
+uaF0X4BE5Vtn33s5FFLR+RYhnc7XBsbT//g0hpsJGLUiRF86q0x1vxXNV0RyWPf++3NSdM9FVP2
t+Mx24oeZikFB84Cm/kSRH+hE0Af5ymrK+cDmVIWKJpXjBcLuMtvwh4sNYNfpkiOvSFwo6JefUsC
+Lvx3QDprNcUloMfYCvdjI/RJzrwgzK+4ijz4acVPcabjWZB4Tnh7f39traySUKba6U7YrJPwwBv
3jxbKamg228W/Z8QogPBBEn9bvrLpcLOKiAYwTnDV6HhnzM4XErMjBi14UK21S4+UvY3rsadilwv
GUyU8a9ltd1lzdi0hU5mKnrdaDUdtDpvxfrtlR71va8Ro57PuikirAt4nN+6aBbBto39Pq8qEab2
Bf1PodXWybJARWsiAswWZ0vXHOJ5+eRhc9jdwC/aqm6g2+yaAA9czZQMlOyC0FUHZWD4zWJkqhry
xVb/VCFkIph7B68VsKJhIRazqKf9Rbjd7w5Wf/DddoYp43mKNtl7s/0qG4+BFkfqwaZwRMjS1GH0
Q2B+hCwQKShJni5e2t+s7P8hFFplHblu9t1blnyEXjWzPMUCaRPB4GVXtScLc/RTPG15+EuxMFMB
T/6cQMaOX0RFT+IXjf/DcTJACBYxYa0zHT2FMt5r1/zGTQU2Q1kjTa9qINXRru2ldVKpMBDacRzV
8STDfQ8vDwNiouS3g4UGnDkEBwu0emhboNbEVHSCPj38z/0OCp/zmLA1qK5x8d1vw7y0kRC9bcIv
qoyZl2OEtTeNsrGRonzcaaG+3veawyjhX+lcrClHfr4GnBp4Zz272ByUQSc8iYjy7mkRUZkKrWN5
Js3vnzO5OfzCz1vQ3ydNuAiwi2IYGvt9bcD6ao0+TCwhXxvA60deAQr+bRGp5jUpigO9EheRMVZB
6qALr7PyRFaAE0pjG4ZQjcK0epR46gR60dlIKTLbzztNRnwu5cixoQIZmbKuV/L7CwIEt079LGGr
MYNDVreVi4KjLZrQaRzVEa6Sm/kEz7T1ScfbGJplOwzLPMjo6tnPD9bQPfrPC2oE91XtuJGyg7br
Q0ZAY24mkm5LvFOuheZObKkOWq3P3f8EBIelz166LE8TcEGUcK/uX0fPBTkxYw7SNCILv8TxRu15
gN3/l2cY4w7oRIbyRhNRNebRhnu/EK9l+esmJWKY3LcJ1qs6+wBHYuozsg+26r9ingQfA5Rr98rM
WRDlosHcTwAPLmYuGFjAX6TgBvwEpLrB4e0cqNKaJSaQEy5yd9YVHpQY2MSZzKLUwQukdkavROSP
pJVOungl4kL09+a+ZKdbyGJRx31BRiIh3CNfAn9qTjpMAHiOu/jxp8pWwNf8Xbn+iK1j3OfRk6Po
4o1uYMJv7mTYheSjWt7Yzej9R5Zp4YEGmFFuY/fuQPGCDrQfxAb33M1Bad4dCUMgh56eBaiAp+pF
xrM8iQSPtqGdimjO5YhJkLu6DNQjruRwUtb48cL1C850ld2Wxy8HuO42dvDWoGZP26GUFLBEmI23
PbPsiTzZgRbxoF3AdpIp0kflQYCSpuNQEJKuCOeSUkjbCoZf4q+z2Y2fZv9pBDH5AJl/awpiKYyt
tzZOvjA5V+zCFhOGo13HO5RnKJkAJOYt2WCUJTiIvIAehsnJGsZ6hWhlfchlRRDO3HXPag5T2VVq
1hV23OHft1/d0aYNZBvagX9wE02XrIzf65kDf6Qefdem5RAEm+ZLRWHvpAlISHPKazKt4GyQNxT9
rrsU26mrhKtz37OySC00RDMnObt0xrZQebem0fdPeKu2q1YZ7qjD3CZwunlwZqT7Doa29DkZR/Pv
M8euF9ZAG3Co5Rndfv1kS+V2gOqNhh12QeIke9ZVuNMkJ4Gv/rYAp/BCp1/XqMr5PHOLT7zhCFXy
YIs5rT1rBJd7m5AohYNB++KWipae7JvzOxup4LF/9MA4MYXDXqFxcvwvLRms/ygfQ5Sk0H5O8DJO
stnbfSXdTIDS1Uzl8DL5vY4KUiyD0ZAVqfh5onQ16EYrGfQNLEcSc5GbAuTI6o7Dw8vQWoso/P9f
MNkyP8VbDwlIBiqu5GHp9ApqEBGuI4Yv/qFd0Iwy8Whl0IUr2j97eRfcPXPYDOc3sCHk1EguseVl
CpwIsQ1ytd8aR39kQn+ZGae26SDP1p9MiiixGwD4CqieJ5cBuq8j9sRhE5ft81kUFfUmBxm9ikXc
Fi22fXpisi/FTl8cN6Lu/C4mecGA0MTnoe2UtWeH2vbbr8XXhnc0uZtbJAy1acnXZqW6h0I2OQY0
lyjWFPkut/b58wlLFcAs6teindfVB6NO/jiwuc58ykjOog/D4s0iA4j1cKpkARXCf/xwyEVf0B3N
Dgx+VCxy7cjJlXhQqpHu+gf3Qa2jTbFhwSPHRYdizAb5Ui2vsKyeeSd67dCJWBjSBiytYKZ4T0z7
nbg1scGhoGMAFFf3+UVhHjqFESv8+/UGMjqRiRNewh/BWy/W5mPmLQsSErkeEvKdLR+OBoqrSNLf
LSmGPW0hfTLsmxO1mjLwEuSB2tcnslY06eQInf7wXkMj3xiAO2Y4CvKlpdkPu0i2cIRV4eMRdirb
6nBs+Cbd9/vOQRDzeLO5wT14KQ9yIA3aZLrQHvq+1Qbv0rnA7/rOAbXyde8s63NBywWt999sm2wd
o/argpTWtV5nvcsnAXvwCaBnBK9Y7ZXb7vLrAUJJDFiXcWaYSiWVsldHCi2AIGdr2a3Cok3h8+X6
L1To69Bfd4LgxKzY7MMzOxaBvQNbmbFyMy0lLB+2nhkrHS6pXhh3pTGK3z2wuXEmRk44PJkS7T/R
WQQiVWOARDgaTDsNfLgE5AGR43ZyHQ6oyxu4/cA0H1WSylXfKR2eY1xm6qExyfueycub5gmuv7Eo
eNQ50M9JaVmZRvsBiLgKddLways85ooAN795gCLWNvQ+hpJ1J21c2Np0MLs3Rhat2/a80R7D+98X
rcZ7cPXM0DhtiGIE+fUtEwyyCFxE2MHWarX8Z7nlhAHKhKigsUZL0Z0cRHkC8tkCJi3LdzoWvxnp
L1F5lWDc3lVTWuk7ReB0Owd4jjgz7tODQYGw6fw6dt1UwQSl6kBmn82px9mr8pbxGVNZRjJ/de3d
jbxwQ1W+YqiHDzrNZNHeYNSRiTTE1ypoA2Z4ub/1UcDyogNVXEyUZTTX+xi5m+P3DVUL+isHeiaX
u4NNzW8MPVU/7CnnZNjI8GlzbVDGvXPateZCIJOfUrm5+gr68c/PoMDq4dYaKS6YZBycjfBPWYnw
vHME8REY/ppVDorrCnGiXOT08E/jcWmhrD+zOOA++SsTDjZTwrtujd2AER6qrpj7M9aX733fd3q6
RUmHH5uDlAmQd146NbxsbAY0aMhRZd9qNiEfC/2I9oiWQdV3vkdPTBbzq54oImjrqAOiiPDNP4hc
JX5N+xHtv+VqH0lsr9RKXqzwVfUlsyA4eKMy3BYCt+A07lzW1n+sYcmw3wDo5Bvk69zgFZ3lBXVI
/TrE/a5Fi9B5GSoggqdy1L0MAmfFdwBAZUSoyOPYVadEaRazenYTPKtOkq8Ome7OTDyl8ZDAF9CI
OXCg084Fo/mswuDSiXrrXa4to+UWu48B8HOFZyvRN36AM43gysVC8MhjICHNpsNA8Oe5OQHdeOyX
yP67v4k2X+lyE4pcRBiffBNUpuSqZHCap2RgdYCh+GeYyMkgEBF488KG+bSFgx6HEuUm/JDj5L7t
r90DU9ok131IvZBIYl5hyJdVg31vwWd5V1gdnLqJFZiMvYmC9zMVo+xgjdNwR4qobFmhnVVPEgrh
08YBzxrs7Q89PFvoALMFtkW7apaeu+Y3xLMufVC8Pm0LwuAENojSsgKrLmhL76ezlviSEebF1dUn
iXPrupVZRGKnQlG/H1GFpwhEDOdy1Cwpd/XTc43m443uDH8SZrQdC9OuQrrh3qp+d/J4ZD2yer94
DT35yxvf9hzC91SbEklrfJRxfkNlkI3ZuQ/r/z4jzaaSZnT2DM+MJ/QCQkHsY1p/153QSUoNOIgH
IqOqj6n+NOGsNwH/U1E+nRBfvvs9tGT70Ml2tsPv4oqMeO7OeYRIjRAs+RCwm2+EbvykQDv9curs
mc4ynFPnaQCvciFKZ7hyGJd9WWajoR7YqH2wmmDQz2qeVHNanWgFiuHtEULYmwrEQBZIjWw9NydS
pWAHGxYSOSVPhP0FjODzvz7jaJ5/ycc61Vye4QFQhZlTOoXmTFeAKfSTrZeC0WPV8sdUso2R0tGP
Q1hn7ID71YiAkJr9rjM6WZrWiKcecyeHt0C5nemOguTO0m++7fIsJUCavIiF2yCsSBjA2/McmhbW
Oc3KyaKmsGIkCcNJJuspwOLSNppBLILfUQaPzWPA4qESrPiZxA7oXPSJxz+D/t33jsY/AgqCoQt0
XuHobvLU7FueDvZqwuG5mupMyq9ZgO/+rxlYAbLUPTVoDzGoAEQg8ax9NRAaXOL9Vt3RHLv6sMbL
2ncbUNLl45XQzpr0F16X/OLfhQsaq+iHIOGa9tRrvF336qvc+J92j+vEAIame1mcUoAuA8b+akJS
IkroA7us/vuWPmO/OrWCkIi6Vk1hOkpf9lorLNqUYBkEE57exDMsfRCER+O0DCd+cd3U+FPETThx
KdQebCaLtsDRIYC1cYZWjlDIgMjShdaxuJlazpJUtxecCVmEsuP3BkDchEtvhtUDrYjqf92qn5it
PqEWTdHufgOEhSvH+MomvckNQqUtx8ZBblbtWx+YL7ynTFXH+RXQrUIvVkGLCdNh64o9MiSdmgPr
o62IotGK2UUAfZmha9hIUoTfUePIFnLKkmlNA3V7mPZR+EoTeH1vUJzMR51OayvXQYZtkDNlTlDj
6PVVfbt81FHT5Lz+RIcsWRiogxN0P9lroypU7cdYBDcHBiXslQJZeoWhjIDyf/6sFlbl/0xd+usM
+ipXWlsEacBf3TcPrZd7ogFQ4ayF5FsKiYs+QhQJaWs4KcDMcSlx/uxDKn4GSEEG2rSikXHc6J2S
SLevXzJX00xx50hk+FGv/fdsqhLlrz0x0/VkL4LsIfljZKAK41yRCttgLG5YijiXoyMZ4aKH+b4j
myzWr5qHph0w6igCtWsECoJxnIHewTOIYJNheED6QR/sT54bxgJ/+s9Hr9VaE8CCwSN55+dgpuvj
GwLnmsGswaJHLWZqP3z37y1EBj1Xo8dqp5acoFWumjmCAtmSHyTcE8mUsj18tySNkcH1ZO/R2w53
qWxjzfz1UhqtS/lxl5yqLe8N3aza8v65QhulYl4/37ufoVGVJqE7705cA79/sCuh4z/Q7M19hL79
TkobbYz1VpTH247CYO0nY8osvXg2/zs2Qutw/crgJINHL6MFXnt9WHM/Pa5ENCk8p3NVy1FuGyyg
qhsxB39qCgQ+kN63QrnOzh4vR+/yxAwnut48Q5MjEPz1IHFhCa90+EWZc5qYJ/2GX3YgSPzTOZRq
ZBYKo9ErvY5ZbhZ0CenrMul2K+SUHLivWBPRPVfq/Ttakd/S7U5UvMFihbSO4bYni+2kr1rDnIaL
g4/imyuVnlAcrnMQhKaexCsnVqpNr/1/C/bIMBOjs4qj6S174+PocIO5eU+IwUX9XVtbyVM61FBU
cNegwU2Cx0LjUQxHRYjhImYtwhMYvouI45tn4Tpaa+lTt3+staQv/qzJi2txGvKKj3rX4sGWLlYf
VP65nPDQm2ml3LtDbnfzzrZOxRjyAnScI+dUK44oHzB3ucXV1fBMN9cU5WAzGqcMIdf1czgyfZtm
znTFu/pfJRY+U34d+qOnO/1BdDsj+Z3Rye/zXxs7CK4dR2oGJANtKwVG/Tp7ivMv/eWNn2x82kf7
Idn1bjVGYVyKOUHiX6hqqmBJoMSd6zbBc2PPMfFKOvQ9wmi+z/FcM3styrgv8oGDbqzhpW9S74we
Kp8jmU3jnU4Kpl2TXshHgMFxD7HQviICuaypIgvhx8/KD+rppOxC6QA3mzIE16jhmXfjq/8pZkWZ
e9lmzLfsBWU8kiP1bo9mr8lVHMcyPq2YN6hWNDYeuShp8f6zK8xETBwiMAW158yjpRVUB6h7tqwe
45z+jV9JsIRAip1W15wZLn21CSMaVnxhutM2LXn25RHQwmp213XWQmxj7A9NJiHELXrQ6jSRuXFY
wy1Jzfz9V80bVNcZIYRRzKn9NpbnTZ5w4UZKKE4M88lTbJzSNKlOm5xRS+miRQRfXSfAv1gMDFWx
jk6QMDJcDIr6ZzmbymTVQVUoDS0bnk/aJR7hZ2bc4flptqVTc5ozn8qih4m4qPKkv8T7PgKnqVlQ
//eMJf4NnLQ60kG4FTQ6lxh5CrG1KIKctjuZ3BImzofvhmhrlnp29bp8elwJLeVOSQnbGWjzAyF1
d5Dthg21Z81esA9t+AbRt3VPJr1YS0HswDfJeiWuNMEOWdPflMq32AjaGXg2MoXZN5PJSV72ydzP
Y9UKBjggV0+UUGCVjHjsqu/AnFqfHQGrflXcytzvmn12WnHG8pAYCfND0kMK1fy7eoXkxRk7yBJp
BWejYagdltYuTEMlGjq3vbscEe3GEKQv2RJerj7xOm3qcbQEi9NJ2fbyUgbj0BzVkQJDXGYti4RL
c+eeQ3RG2brb2IdCfAUZqNzx5MVI6zpVclWwVZlaRvUvaDuAEV2YW9EXIEX0f6zj23j3ljFq9Ea+
vW9DfSdJHD3PANYaSq2VX0A1kWVy9kkG1EtTn1XNlPh4IAJlFCuNv35cGQyzMo4etILDatfpVZ33
EzyCW+jPLjSXDoUwRUEc4E/axU/K9coZKR/b3gmFZ227ZprHdHTovViSMD/B9CMNI4zAEmx+Hr1e
qZEuBU1WVdvhaTKhGB1U+nrX/w6zE8IQmsPTHXEPEVfsDdjKUIbHI3NQTC68oI4x4LrcBajVs0oA
mxuNbatAOZRYN5HJWc+PlNqtfHYiZY2qnou8YpTENxoR8qZ3gBk0jk3DcTRbtjG+piklig7XDT9K
NR2VyNCsM4uWg4XhlvMfKaZCsxnLhfX18haFo8c+FM7N8Apb4dm5TsffMguDgTd5Z147fygS75Oy
GJd0Od7rlSpWL0LjUSblHpdDzTaCDhHWU1EJ/YRQUgxUbqJO4gY7dQwL+FVt0u19dwxkOZc0lXal
8CMSg7RLxtSMfPf05VtgGmmO7CEGGKQ288MmmcfVQIcnLabnqdUJoDilwfiVb2z4gc6QyjAaIEHG
wG0Y6J2afPP0GBlNjGU9dvngJM8q823dxTm0Zm9q3kLtlNsQkRhQeEi94RkEEB+4K0A/1/xsUkME
aNKd9HpAHrz+6FwWDw37CkAKyiubO3dpXbW5Pgq/6Op3C9P9F2e7GcggRPIu8+qc8aV7EbYv7Yn1
jvlNFFBxZoirWF/wMGM1/qqGgJV6P7h289vk9CxYGPiO6cxmNC3+uhEbBqmmzysia8gEP4GGoQrM
1b+Kh01CW0JdxkiCEytMueqSnfazlbXoJqmt2QGzqCNRHrgPgFkdM67SPXb/P4edCeEevLwEDAtq
Cvin4DBU6IxH3Pk2VOhPb6bNNct/sbPsdX3xe14FbbIkySXRO6Ff6Wkk+76bPWhqbMNwU0WfmGmb
blLSGoCL4F+RpoJtqtm+C3BNDTPHPd945EWY9YOO5o8lnfPTG9nRvttN28pCEFRLkl7nv9go3zKZ
S97knwrzq7uthTwcJI0huxnX9B/9EE1DAzMzMAn2oKGEDyLti1l5vV77PGCBzj7qX1F7y6WM/ZGv
tnUB8qLbkA6YdTAkgNkqkNzoyTPE0nWej0RK9VqDCiwF/RJhqHY+S+gw6YSvQaPxUgftRNx9XrM0
uO0BGBZ+dLsZoaIXSSrwKZGK0iqb1jzW5JKIBV8vdXvip56V/LjyDFxSw1dvb2f0POpcHLgZAY+i
4F3SxNKIRn9wnOIO4jEZo7Y8Rs5IUPSQMqHsS4/6L0xd6HcE8P4GD09Pi0Xa83/VZ31mUt30H9jA
a/KcANE0BMH+S7/ERMGTH+s0XL4twwKOSg7jXPpkR0R0qyXWFej695xYEXeu940cCsZVx+KA8otL
e4y5DZLG/walgmIzDRzavq8jvss+fW5iEkP1GcWGrqkNImuWfbDPk47ExUNe/AIDu8dwvGSlgWQ0
bu6isvnkwH4P4md06yxXhdyalzZbLQWEHY6LqCMbOVOek1fsZXi1HCDnwMJsb64uqX9VzplM+T8J
CXdMkmigqH48SX/ni+l+A9Ms/hgCAGceRZeXLzO5vimeVp2aOzU9xQ5619EEVcXceZe/E5gVBK5t
RwQ5VoCPnPM+eh54rjSVzGJH2/1ZWt73X9Vg4ahQU5HqfKH5GniGebv1I/oSwnWDn0WZGJx/EXTR
v1XUgs28hkj08a6cpV+ubqbGOjpbAmX5Oq5+dx+SObyrSEFwWrnhICjVCBsarVFH0wUALK1Uqluv
SpiLhuXbpkDRBkPXVBNI8nBcr26/ZyL7lG33r/EtHwcjbmN95fVaWS5rfbLNh/4eD0W6pdLiJzL6
N2kd6q8HRm+xBMsRsRWV1nqIa1EnNc34Zrz+wSqj76k+9wnpVhTsRFlGmAF+2oyiodBRxo6rvqaH
L2uRZRDr0H4pzAp8YD9/DCUAs86MQKyf6ZpXVYG0e8H16exLh+mmzz8YW17JFJR40ZVXVMPoRqed
HOEuEJd/xuxY6wbK1R+cl0paQkEMXA83JkycTDcsEQR7uR5Qx//5cmTU6m6YYCwIaFrrK2mzdjhg
BPnMxJf49XwPmCxdwCWp188q+jDqDnIxPTD7+3WmUTE70kASxfU/SDeyJhnPPn8M0XGWFWxmv4T1
hZA1PEl1IyQbmHKVU5rhuX9cSOEW5iZBaxrW7z/Yp23tbwOE8SuirxOkwpRlSl4E4O+zpvaokv6V
B0ahMfoTuD3r6OjF2KIdC72e4ojDpSmFRfli+oPGDep1ZlZPF/g9FYg1xRf+jzjocB/0gFPhMiqV
iz7LjzkYBRxBRJN7C9e8JaMycuqDUtwHSDKFqrKi1thUsiSAquuTT4Bn5uy91pi1OBo50AGgeUyn
YaKqHLtI8oalymFRs+KyErmF571y+JlgGGWRGg5M/QrxELDdo1N9ihA0PhnKf6nV18CZiJ8PXRY5
q00gVWC8VQYUwBKc5oiRS3FiFTxtu3e4oWAm3I2pC3U0boI91PDKa0UsCK7khcAlJyvQbG4NSZWj
dfDDruuuenIiBTqOujFteQ7yy2xsCophbcNCoLet/WP5rnIg6iEnNmhVANv7kHDcr2RXHOFHzPrT
IqxBPRRxaRdlEQ06hbSkIuk1UEON3ywYePsDJGE7puHJLppI4diqtTbEnaUyUwBG/FM+jS3NA5jS
ioqwueP30TeV4BE/wA5tW1oPBxYuIi1P6VU5qCCuDht2TJQZFQU1cdFtCwESDPmeWim7RPkqFcc5
fmO5vLqrOvX/tfPvghm8dAVChpZKKqJPo/Rre6sYAUJLmGVLrDwJvfaNR7rRjj6cwJdFURCZhq1E
iC0i2BChVX5aveWwzTbKr8sEUrWYKaeg/DClwEHpX/frEis8G+NhPzIFmEYJCD1rUxhSH2ASkMRm
o+LDN+A8MggXG5K1gLnhCFiOZQ5sgLpkmG6jfcNA5L4Tsunj4UgDgQFXZ0I9jJEpdp0120jJIMmS
+x7DCQMEVsJGh4YAIx/pyxPHBuKkFUZ3YrevmBcPN9veqR9916gkByL0/Ujdm21jZj+mQDsWb1/B
YNqDgYY7OEBaz5pv0/7PkfuLu/Y968XxbgHUwmBSkDZDFCAtdImXg4kMASrGii3BKTo+bL0wecNm
5JI63tp+AZyD3gQow8662TmlEDfRSBAj5lm92teKeNlnpTZ4ZZeXn/fByk2mcMbeno8acZQIyJs0
a8rond8xcYuGEpVEkrc0TEYKsrvz5WFP6TEpCXkT9NXt3DhcHtT4ntW9diosPk6Ya8CJIJjGYMgE
zOaNZqrWBCR+CE6HZzk4Hn1Gnj1vU17nyJKOD2j7jZPrYIOxgqG158dZFG2aiy+nppApIdeUed3l
8voz91LpAL4SSoMQzQygql7KuB4x9Z2U1rjQ+gj8m92CKkE30ZHb+T8AbJdxnPo8Lgc784Sc+3yv
XOqbieC/HLKgjvCmsUJP/D8/sZhh5rUVlMV6DgONQeRtyb+PY5ggSQDSxQX3RiYCebX2YUiGAo9O
yRr1/YINlPn8OjhPymbm1aF+mqTKnWrbHQ4UsF6mNkffHYVf46FXFWlPAreif3AtbXtrXPAvPL/x
vyMGd8Zcjfm+bBK3GI2OsGbsJ0zWtfJz1Zac1Lrx0n8GJROcMh9HOClX64U4lhLAGEhoaPB7dKFP
/AXgLy+GN8SG2Ab8Yw4y2VvOI4CKsDwh6ndQOvUidZEfcwgAS1Jpxvi/tAwMiMF08sUgsfELMtj6
45yc5os4b2D2f1Oa7f7eSfvu+1r8XvCPmJGJBLa/gvY4MfJklC+h0rtCVgW3bNni1G2AdG93ISkL
gizoAtPPI+A3Wx4MdEiaXcf9HOnNhtEhDfQ8mz+L/ChmEFGzWTQZCODCw+wPlPRjQBjb6ioWodpI
LSNlmMjNJPDOlXoK9MH0caP8a+pVRtsp1/gq0VPFcDeleJqbnD3Q2cmxuoH84lCBPLCiSs0211WA
mitiQyRxlBZolxl1naN+u4c21Dktcd3Uk43AjulMa73GFBuYaHhSuw0rRpPeLaQRtXgXqJ+42phf
rh+gWTEbCp8uo5mGroLO6O3iROcxUo6XsDIBWfEEutZP7artJZeZsV4zt9+OhsdanzuGxWeW3yHa
a3Sen9B0hQ3XQZ5+01w8zcUh5jEG41Um9bAeGF3xwrM/qTVMJzlMz8KYGH/ZfqyfAAQYp4mraqUs
ttbX0T+0GBYzDdrlEFqCgCcrifT0bG5KYDGtTJkdi2ZihWYJtFfswMaHhpajaOxvZ0ofdkqBjKUi
szWmbmSxjVSIU4pfm5vt+i/32viNkEmdJUM2p+MA7Q8ju+RN8dcuP03RoIZplHdYV9tQo7uBkWbf
4AyAVkLHW8uf4OhpzcWEEwGrc5CbhpaOLmT3x69U+zmC2K9VWpqYGtoeQEYmfG91ZzQuD1twXe7l
a6NDHoXmgSmubMtZy+ps+8a64v56HSk/oLb/VxpruL4xMDYnbKn7vI00r4a1Lk7GsXlXFzFZ5lw9
DxeV82JLIdjzvziAZAR8Nmw7H3id5F2Efk0uhqN3i8nYUb1M1SUTcl7BG6KCXXqjUcnnyvN6rJXP
/7+Mc2f3QBqxYdO7AsBoOAs2mQi62tls49NuBrhxIaxhsb/RMcTjj6M+2evFfriD9kEl/+PaQ6yr
Oc8uumBG9TpxgF+Jm1C2FPpJIPtAd4JQfzK9C3gmT4DxbWxsZ/ISpLiQ2G8cF/+WC5NcgC4C1d71
DZ+N5DmSUeINrB118vXqpjRCHzcwRIwlRnPGqtCV0GFJdFf/UubwHfyyGHJ6kzqWVYLdbcETEh9p
4LH+26uxjvOKRDfhI6Gdi9RDCF/5zqfx+sJV7ufGZUZ3fmY8B+Vtm+2lWC5clQbkA9HvBoXjrGT/
mP3JDN7VlRa7Ufxa+uKCMczKR/LawAYCtTAioUbcpI0aFhkFCvdRqJTA+6Kp0rwWMex28lAOsrQJ
Yiqc63yOPySPs46WSnxdzMJVARF8Nx2nkGIZLUyrrC3e86xZpgd+40X4h3k0sSBqYgGz6JiwTCH6
j6s383NFK2+02NRg7yU5ffYi1fml3l1CaD7Iy7VqKfT1ZuPXXh1ak/5mUUXHWTgqs5Jn2Cepn6n+
9FtOXmQT8J0vjgUqaPzFWq6ldT+wV5KS7QfwAS74hmxSKiA4Y5gREXmwwxaXxXS3M8xJaq36DQQU
zRwKvQ2jzSNWh2L4Vuz98cyYfzoB83uh0+206+ZCxoNG5DcmpPK/VBmToBw9+HQRVBluqVXCV/fk
v8polhRTwiSiMxDdTzSja9wy9HH7Ej+Ra/7EO0JKehR9kt3Bc4zJ5pJOZWVRSiT2CbDS7ecM2hfr
v3QkbtA1jkSep6PKERlDjh3FggzHRcNOk/YGV8Rnt+cb4FA1YUAghEBRjqGXGfd2hBQrHaM0pRzR
r9omJTJoaSdSY9Y1qogvP2uDgDnOci/isC9SujlhNy56zonEvXn0lWXW7FVdCoI6gnJwi4EeCAIw
UW7tWU7Q1+4e2HXO3f5szahq27afbV3h7XnAXMpWrtYJhNhYeT4KBAD2AJ9Nlr+Q7Qful8FCDY7u
MWfg/61HRf6ZM/mo+1FHFG3qEkjejcg4Cd0zIwKvfBISRHpXJGDTpIfGk/BEc7sncuFLzEgRGwWf
p5uZaqc7rhA2y71U7Lw6enNlYIJ1cy6PGXigRwmag4GCe265OW1UkbGzjj36S4YR2GwJ0J+XdVjm
UDI+7xxgirPyaB3tFxqEXUCbfBc+84RavYqPCwYW+PBLQ3jIM3e69w6UqWn76IklM7imGw+me8px
CyDotyQMn7tZG/JK+3It1gUPJHm5LDodAnz8BGoUFdmTCgjLdk8naX39bMhzyvBX5zd/L0uE6jlM
EnQK9ilNk0zOSipX+w/gW9WpjdiSIaFKtTR1xPktNJgslGRbuznal5BV/FPb1ZsZpJ5BN39hUNVt
yj6QF3o8pRNYviobeFMYkGy+RLYW6oL9wz4s5Lg94j52NCcIl6vI6LBVkjtDTeS4iZyxwnSQwQ4k
JVC4hPHfh1KymWqh44Co0qvEVDRQVbBecPByFoAeRyRzNl7IZntfoWYF84vwC+0inrtI4CLRLa58
mBGg+mGPuV3ry03ezw0B7/MDOGjjs+L+CzHmBt11/FASzFkDZTQKXmctD8ZNrqSKjjf9ksZa/G37
KfUpYTuLxhVwYkezwvZIPycxj8FmJaGPZvCkPhSB+TRDCTldGv+r4ezjKaGizVMo7TNnjyZNWfZY
6EJW76T6p6v9DIISBOsLjpIy0bgPpDBZoBYg948SZIgpCti61EmCas3x+snzeA5jat5Wxf62NAEp
EUzkm7Zp1nlT9KTY9RqSUSld8GU30+vIJVAOaQIWnY4OAkRHra5jiPbCp0Is4fiEj4N7U2idrbhw
cHyro1VxQwPoZ3vdiuO6WgmZVYKX/bNn9YKwrg1tNh5iiYnTIXL/fHPppSmQmdg2uriBzHehhsu6
rfcoRN6DyFJzRb/9YZ+SRfSWEI85nOJ8TFVZVLVWvMjHud0Ge+4T+5bbZrrLRis3ElHRh5GkSoj9
r1VtsFAwqG85JMexMlJGKMuxxtwJ+HhctkIitsQEX5hcm21lMZd5svFZW7EyDmr8z0mSvZ5dn3zV
0AltzzCJJWbidui1/aAplWSzjt/GRgVhZeiov3NIw9k6qEg3dJrBJAefAEmRvhyFMyMfLM8lNdTb
mVljtZTKk04StWNa0nbPpDgfLzulFX2Eyh5B7UdQT803tkI29LsFZiC2Zh3kvMh9B5g+x0hFuC/O
QwzNJBPEN4Ky02Zp94TgGf5rTuuHnT/41RqiYzzMrAgcn57S6Akah3C14PEs31I4zm/sxURYB55t
nD5CnpQ8Z3qLGqhnFw+jJeYKBLkro5/HiUHYGXOQPlgA+2WvH6VCkM9YWI9q0xC1t6FAVDXMwsCe
Ck04GgVPV0p41E5j85cxrbsgfAw/Z/8hMAZk7DcR14KtiS4XUTxcXVONU8Ojy/snMzbOWzir8g6q
ztkQf7elZ7KVUpMYvWpmr478S0a1Mq6Z+QSgpmjS4yX5G904vJdDW789yWNpimwrrrvEhh9QVLID
oumFaH6uYl6Y3r7t4h45KFTUC8VhmN2fg5pTG/XW9Now/ZaTTh01KOWgD7t05lew+jW8/OkReuRE
wYESu9ZwE3d2L71l67ysR6YfIEpQErAutvZWGrimAs2m8+vVHRVgyOiL5qz4maJSMDpunJl/6PG8
NKfUvD29Pz0SPVWYYfiga19jCk7LW+1+6EjkpZFzOx/FyzUOSUKqd33ddubd+6ugOEraOdA7ooHj
v9PG3UxO5i3DJFF6DsPd53Q3LlvEl1lGF9xyDtqhoefjsZ+/RuwDngeoa/6ksw6MfWi/FojZsdVW
NNtOGfQshy2k0dBqGG1te6hah9LaUQpFscHVgtX6rBz6aPZwWctXWPcti6XAiglkZEdI/2P6lCk+
sreyT9M8rdwfiaAcBFFJy0d9rXeoG6D0dfaZYBlz1XoQKzNEAjK2wutueVeox+ONJNbeXK6o95i8
Ie4glVQuNc9eTaw1otTBDtbu8j0puLocepDMwVQX+smTs5hOfqCz9xrNhCp5zXs9wEEPRqz6hOhx
mntvxua0iEdJjTgXKac0Gd/dmRKqmhyWdeEqnKA+1icYKepI4cCantzcIux+t/JJ7qdkXYNTWPfp
UW2SoDCCiut6Ph+UE2HbzAm73z3ExtMEy2TWE1y6FLtfNEe4xQvY1fnoB1Io0YHNBFoIdRy4MVuy
e/CwLdBwgJY6JycFlsfUMldunzztVigKBBHfpk4jIKzQsOrsAf6fZJD/2nQuPPB5A5LiQIx2R/XP
srlUCzsg1rCdghr/zZSODJguKdNzy0Q0OKMjCvj8ufbBNWVQa44CtaF6l+E1TkW2J1FrOr/5LDWg
9roRDBz3ZxcPoCXJ4itFCPir+gKqvqjVfJDz0IqHC96CWD9thIo510B6p5PahZkrCavUjusSVbeV
cYwaRRKnr9uZhtQYAJimHrm/jNbco7RHXIRqQr7YIPaedUgtqoooJC+26kL7QYwolQrTk1Cd303B
qnH41Dy0QQdIZnsZ89/4d2/lBbmnaR++9ewso+kC5RNpNJNe1w9FNVrrk1CyITB89mHSYeyoLSQ9
O5QqSmtlxTmSy95QB7geXIi0A75sGg2W/tr+Am83H5664ulVVV7WGkPRs41A6IsG7PZrKP2tIMD5
SqPtcNcnhgRw0u9JOCLlHsvEMdzIAvmynWIue5giBcNzLAnfs+BBnJDAa+g9v4LzK9ubzP0sh1z8
Ei4oIi8r5kBfXQUihSO2GNzJzkLlVCXWT9oExUev2WQvQnBYiZeKIct6yru1BkJyGg5GBoYeZThY
LBJIgfmfG6cEIQDZ05H0ajCPBVx9sNQ2CSyt/XVPo9RxKDILiLSiV1/JJ0xM1ezRA8/4ECH/1mqW
2OwdL25AJNSdBsFd5yS09rR4qWZThhiYnhob7H5FSGIkNghrhfywBAUsfOYYAoHemm2DJv+bFXrM
T/booI90wiFiC3yVdzakipxcrCFJAjYGfRMOARJZvwHjcLFZNs8j7xDThsVsAflBPfKXuo6AhfYh
j8AQmZ2i2aGuomMMFjdLQnFmHRJADc9O++2ZTJnfgxdo6EmJGMvFd2owaJGAdIZQ7Z6ZtAPZjRDz
V2j0pd8hxViVL0DQJfTd+z2g04/+SesG5ewY2ATv773Z9ubcJkLo1gyCWOEWLCUIDHmsTGywWo2E
A2WYHOzPscLhODl+HpkK/KgI3qb9neVyKv1kOA7UqCx79Rifjw10THuEcc2LdfzedlcP/lHKlVYr
45Umsw+eH32sLHdh8RxvGXeVq3Pkv4vCp08qw9wdS0KL664P97+rSRbtfsqCBeyGWYhI5jd2hM0j
PdB7j5DFtyw6It0odTejFGreQVdYA2/zQIs6Cx4ohv9X22VHZaFfaxpwx219DePgUYr6t6pbMn+O
kby8aF5sSYornCdsOY9SnpfCWb39XkWtxY/dsYvbTgtmSDFkB/f+w4/2u38EzcyjQQHBUn24zH/c
bnsaQkhQy2Pa2kXsjd99GCUY4hvEUMM7DIUfmbln6UAGobMt42U1cvTd3gyg/uRWs+1U/RnX9tGE
oaUjEeEUduNkV6xHiNVl3XuVBtvlySnCJmJ2/Ni8T6VHUFeU/zf932U63l+wTC1+JPVsO5mfniAR
kW9wKYytfA9iWB7Fphd8qwwIskzj3HW0o1Q3vZbOcUqTetbbWZFSuSoEoLFizeP0Nr2sJ5lChaKD
dRuj7F7GPPdBaABfqhnB9FdbxPjcYAXP+rBaEGj2d7x5xofNt0Cb2SnoMzBCcE6OwgNTCohhiZM8
NZyDXtlsYcipbYkEM5UpFTqA1nxSZK7AhXNCK5Zmxeb8Jw4FICX8invt64a1cZJDbJnucwag/1cR
ZLga6uBuHSSv2ZwcTiTgfi4BXh69kBZ9W0rcSyHNH1fzLf6mN6yEkpOx2eBl2EZRg6fIjnkR9OY7
fMOq1OXq/cFrzcGm8QSBRAslxXnTJXQliZ1hi8gPvTRH5M2ftaLEQz2tzDVlHRVIHkJw+cL8SArS
veZdBLsY5lKoFfyFQuTmjO+nc1iQbZ4hawYaooaa9tzAUJUAdO0bqLTgqgnjS7R0IFGj7w7f3wx1
Jv0j2cjCV68ZzYXPRXGhy2PTObihIu2oLDvctlyXjxpPkWg91fwc3rL/CRDcjY+89jdZsdguhEG2
dsDDp6F3P0ePZbupCxCyYqWOrvZKZAMYNVzV8/yf7PfSqtjp76cCp4lQEFfwq4F1WJVKBs73oZ3U
csmX++kSDW8E0sc1V5+K2xbLcp9c6Ls6qLJp5t2jyY4q3ni3jmdmR9DppPfx+VgcsJXfKGmC7m+L
YXdovJI7Hn3/De3i6kXOXcfaQFK5IlHQvHw3PApvTJ5zzeqMWCAKp1/NgHzp2h2R3w0SjptfYZR5
r+4HNxvEwYT73yurM0WZ9gPBAP3c+2NHGz4WfUShwVutsEwJDAP35UgvlpFDpWnKBThBLSMDiqB+
U/1ezpegWUksZc5RtBHKKGyxyphJbVCWMjJKKw/UNil+kBgN00a7osd4XiNxZ2Bwk88bK71HabZq
yjIejFEL6kv9Hvd/jZMBD/5gz6SOxaCuMyTqmVllv/XIYLPozLfj98C22zzBgaIGzq8Yu5o/71TQ
5KdtAWLbUY7+PHvYsyb2haM0XoZgrvGZFx1Tnw5u8pBuu0985AwMchy/SjfY985jkNMTm6BUx87L
EBmZcmF/9vilBeCADPd9SuElaeII8tmWZ54FGGgAn7iM7ByA/LSnRYPLhyM2fuSPRvn+BPMj/bsd
Ltq1kdCKsQA5m1PsfYU8eA64Jx/rsxLXyOuoxHyK2vd42OqMwxDzIH36g+As2Ci/39g3nkjYjDuh
wP0nqsDlZXJNoB97wEgZTM85H/0q9wiwfeSODNsY/4rxm2yfi3M14Pt/Vb1EU4rMvelZmeuyV1AP
0y0isI3skjrgXYlJ8hflkyAabsOnf7d2xLEZnX5P8va0DArI7xjYrWgXQ+sVtdensRNeR+tWh46l
A2neuWt1+z3ZL8Usd/Ffr+L5EMUZhtEfnf/rGILZ2QsQP3HxbZ1alD5Mb6VScsSSE7u/4CLVKhFS
Ndq2iXd1lmKlpZQg8E0qDR7ukZkO1Ka9B/L9WOUCtQ9svxfS6kDzJTkr3UZaRqQsjN1tobCsCRt4
RBJlgznzAe8SCoXKW+uWUQVqKQnWdEV//Wv+zLVRH2M1ua9yYV80dgGV2Krcehyv1bLMB0S7Z5db
TgTz1tgu1d1uXcu6KthPR7QZ80q2oQcd6sv/VzZVl9CRvpmVyyJDbfFHHWFwn9ulssI9H8ujz1S/
G4JKRAVsvIVPz9rgi8E2SGGnCEtvjXFLSrwohJFUD2+B3FFQ3vzCNCQBSLNPi8eMkb8h/8y/KOPp
U+gbUzDc30f2y6imLV8uORnLA/+IVgN5C40hJ3Ed8qyD747v5ljXhDEnjPq+x5jPIj1xk6zviHsy
Io8Kl0Y+vi4x7v6K49nJiFAnUCRvRFGBVCvDrmBW83AdPDTUc9wXGxoC05BqDp7ABwH1ii06GCrc
RpQmLwAyP+6iihmDvd3gmFVsq1hB96We7YAqFcOni6OexiYOkzBhU1AyDAbkpSXUaIvvlNl/HStE
G9f49ZlUVCFVjPDMUudZKi7ZaubSVDN2dWH6OJAR29z6vBGCT4FiFxfLaTVL4Ith7SE22zXFy+2F
xQA9niZK9wEwaYZgAFa2AJgsQ1ceUJa0ltRsYOPdiLb4kS4bHwBdAfPSa0GX7bWhK8Soc95r6OLS
3/YWUVGIMP2Vr0U/S2Jjnb6OBSEGUF4tNi+nmAB/cIlFEakx3ynNfSZ8up/mKbHsjRAEr3XN2dWW
oibeS4xfSwZ3Dnpx1xAr6WA17scNvEiUhA+EkuvEUTRzBDgfd0Yjsz81W5rfZ/ofjScVi7ofNRgX
kzSYzS6+TfpLUvRaZXtY9CBYeW8CUE2rj+klmI65oT+fcARdspr0Weg8D2IxjE501XNst/SE2yIz
3R6ntJB5PcYFUv9UB+R8ySb/pYYtWEUv9c8hyL2vmt4CfcO8zDBeHVtKsP6HaNnU07ybQn70y6Ql
6zP6bxr49EACi/lEuj6qQVnU//LwUrXgzaMCh8q4Ilys1saUVGwvNmxp/5U0LFSnUo0UY21s9SF4
R/Fh2VSdAyE4BUNyLU2RrsIuSvCL4YRvB7t8H/ufEfV81RpR/m4kaUt30E1hmkutpywehEnKIGqK
mrbcEy+uOp3FJQEq+EorfeUaYcD02ho6ubXNMwRc8/D7uw0Q49pnBHdOwTXuOLfCupiTRNRGv1EP
LHuBNJKXDG+obIwySDNqHuUjB3hqesfOSC0RpAVE06f/Izof0cV2Ys4jWZPJpRrNOdZC8cMCN5tr
2S/rlcG+zLiOKlmpsW6IeUSc/EBYdXbn0SrgC8UBb3jtFiJBXgNInvMI0+7icytigTYN/Wp4y0IS
fxaLCSuOqijOjTTNpcFuvJzYBzPbB6J1ErX5dYTyujy1q4rDJ1I6i7VVRp7fNp9gix93+OCI2C2O
TCIrSZ64DZTHp8CGZYEAgMF9qQ8fOZM5rZSUhhY/zJimp+5kh7DIZKknq1lMvA3Gi1jnSxmhQY10
9+HufFwrueIn+rG54WVwlHGOPhMLgAuf6vaovXGhRWLvE4VOQQb3e/abUB/ZHBAbfJEXbi6tPcXa
sclh944/uWtIcSK10hWilqt7FOGJ1xFhbmniv4N1RNpTHtKKClingx/l/XUezaz9oEVcRTvztf8A
gs1yX7NHFpNt8fMfRekf8cb+IC5YE336aWchbQdl1jIcduY6noZwsi9ZASsj8NKarK70m9TXg8Pr
qm5gsxPqjtBXu19BQzqmwwen/zdBNFCeJAuwlIVgewjSAiFiNsz4BisxndekLjXcwtGtpSyHbEc8
skoTT3F7seMSlHMtVQKv6ztPE295F4588jv4WD697LTuMV7e0Ue3n/R3Q4son2sdFstX7HojLw1F
U12jLihqTUA09+urbI90LZx5C9W9E+Ie2DW82MCc9ao/CeNp2RD6HSiR+thppWXVo2AtaA5hXDZM
L6lra/RhaoxaXKDw2KR0Mzi3XKNCHwXeP3gJ7Z5yscJCXmPxbx7cZOPzx250jOx2o1gXu/ajAwMc
1REHPKraL02AC3Qzr5dpoBrqCj8KZpckYfiArqfOGgHhYrVpLRadUI0wqCb7WFWu9Onu3xdDZsn4
rYWtzTzwIGgFZFDYXZGNp/C7ReTxWLT1DUX77UtcKSfr1NE5+V4m7lrWbROhlmCarmwcoDkAZaks
GDKWYdnU5nmOLmlHUWiHcMpMH9BpjBioAVBnHTCu21K9Ohs67krxf+s3g8kNr3kz5PBkCMumEFI/
JOYa4g+QpzKjXFZMMUAbA2+yjbN+yANGsEA8P5jk7KqZzw9ud9cq6PLaH5V+S6F/KKvSldwxV9tG
peZGj2uroaxK1wlJZ3IM1NKxQvtoTEjb+NYT+/CyPSlpNr31x1n5A0LG+GaKr+T7CanTyjZ1GkHu
QgUIr27IqFTGzMNNiLL94w/J03SeETIrZQF/C0BjYeuw2Yu5+35GoyToNlHJguJTTTnUP02SSFyd
+jsP+0jq8MRBQGQm5Y7Aa6Oqiip1QvmwbnnwV1AjXeh0OQNi5fxcQ/dpLYbTPonPHkUa3BGlPLFo
81GTo2/U9asiYToCIVykoq3C+VbfTG75p9KOoCCKpRucAwrjHgzMUjMzdoNBJts4oS0zHT12AhIa
QQL8DRWaOF8qIDKqWzcDkLzcDBuc4PDqjV14DNaOCMeH25LWc8mDMrEazQskrlqul3UlQ4lpz355
2iOVt7vZZFIOOKEJqJZPHWqF7r3PLJcxhGp7aPGA4KZ3pgRpqElJRDZ/mcokyE5WDxDAJQ8Eg/kG
uHdTWdqGOXK35yGiWSdYh8W3OcSbma8EOrGsFBMC3q47Mu79pupHcmxawXtbdD+COMod1LosgilM
z9ptVkUsO+rnHLl4jHXRvxHYBmjCSOjb9EibAwH58hWj1O6dbS3q5aYLAH8ncEMIGib8eLowswXH
6qNj4Iva4ga43mSrJYj7yVAuu0wdc2G32aGFGRDBsRrIFp9pnQbGutqBGB8FDN6hCPEH4ICASPKb
UdrwSUFtPx+T35zWTTyfr8z9rxo9M4tyTtcIt67IVs/ry7ErFGwW9nj/qCgWTOe5Rr5szcOoaQl6
6dqSD1E7dz9TvJKLDzsrgNQmSnKlWV8jnYOFasPjzy3srP+Tso/6vFb6ED2cMdrRh5ARLD2wVGSE
1uO9kuHesOZcljiaSfsyYYBJ6kvVz4ly1/1pIoKSJV64ILFHx+auGSbFDe6DNKdQHU81r+bDM3wF
gnkW44Jz/sYik80sZQ1au8EJ18sGZW86H1wBB8xSmdec+WsOuziOsnAcPZYJPfGWxqvUaF/oafhr
NtO2freWb9OQYoEPxy6CA9PHubAZk/B4qb48fON8H5Ltl+ods5eti30A9VoI89DsSWSfnxfDCBJA
FbxNN5RPw0DEmAgzLhOWqFKhYi4RtlRxNM/USxYB00BBq/8K8jsKUHL/8Tuk7apOs9e6uRSBF8nt
Q2BsZnqyOnQh6VcssGhb+X5GWLjvb9SYJQL7zNraQ6Y1PlSqC4y7wCsnX5o7srfJlYAPQaC1+z4r
xcgEhvL0HDLa9Sb8XPetCYFa/G+jX/2XfD3ikX7GbEqIHFAf4vi7j7d0e2fualE7Z32V7yn3f7X6
ZwnyC1cD2iNpPfR9so8C+Tp73i0HYU7ZtO10VElhZnY3LStLfm8Kx4pmQL4jjWgxNLGUvNFvsxmG
r0oup604IE1TRLK7xfJLG/7fi6Kr0x/Nn+vojj0y4QaCCyvNhYhur3W4TTclbQDpPoa3/NT9jDRp
8GcfNWa9Q1eMi+DAYwo0tb9bZk9EvSXLCNUn6pg1BcFDt7T85BXRydns1iKs9LLdYMaNoPV/CnOw
mEN1hFmN1fg3dYSpk3ZW8so2NchlDb/6/Rv0563H0nCjD0JIuGyhxLJn654fn4BO2QWoVuKhdq+a
TMnSZztih5Xjd9smsiVa/4VmO0UWsOGxmr3g4BGvoMdwPr75i1SYXSXuxW2IXA+wIwhW9aIHS+rv
N/QPgfCSZjBO/RaXzi5TDvrDm0q0sf4QGLvu2s/DSCg/th820Fmo2RtJ4E/GKjHAn6vD/DZjuRli
3HLPywSOpp3nwQgBqTZU8g/W8j4DFRkiwWhrujFEXj8ceu/af5LQWTt/5beAyqxFQ0wGlxBU+aob
qEJjFSD+yVZVvVYLLArCTkw52FxstdDyfsk66ANlqQIqm1g9cyD1WFTMSA0PoMd3La87T8gcg0QQ
vD881UsSfBkP9oSSKD6lK50PRi053G12eTKZ8viKfebxbDMsjJIyZlwrXb61oD+XRMh1HVMEUv+p
vo+bsqXBwHp4qt3Eghe4BJbTaRPXVJvdqbY4EzaKwD5fFOvP5i7hP2QGDftz3CoTPbG9AbgoR7Xq
UBAnE/naCUH4X3gMPLA7kkVeAYt6j72ijm547U4CYz0wQbBvYb62m6LRztrM1FuLi79Jp5hc24zh
sGD5m7Vf8IAPKd9QX3z0Y4TVV1EiWM/5SMj5B3S2V+InV0T2k9vvTEPBNy/gDQPwKcCp9B1JXGku
70sRz3ZCNAijQgobKEqRKpPpu8lWISjGFdDCen4aLyLS+btwwrVyk4sfwZYX+4KvjZGtIDFYL1lz
3C5z9yBLm6TS2B5oIjSpHWxzdRhSAcab6lr9rlWGc5kNQ7GGRyRZxG9p+LM3OT9vGlKrcbbndXt6
W7yR6hH8HL+kd/u7wle41exEnWPNaR7hYJZEd9YVKPbyjMMi07mrzku+EfHczyFiqzT05laXBsrD
jxILjagPMAAGO3q+I/5H32gXf9XnQ+TlafAK7wOr4l+r0jcIoemt1hOY7Fv7GfZ11AfQVFwTPnb9
tFPti0mZ1A6uDrks7jEcgO4PCkRJsVqoUokA4f43JFS6RQc55G6iYwZ2Thf7SpSP9TT7u5KNPh0Y
kOQmb0+cPKDxutBXZC/EXjqC+Wj1JatGAJysIB4j8sLpm9rqh+r1ToZABhicFqmSefNBuBpADGWJ
C+m6e6DiH+HxG2aIdHWiNDWcaVLIaiTmCy6mpeZuvSnETiHoKLppn98rvhizcXhllAAVP+3OoiMO
Lky0TpKXpBPzbBwmiHyAMJV++wLzRkFH5r/V7ZyVwdEjIuAUnG0cyzqGmAOjaMyKNuA8CMg0DyOP
UVJB9DzThCJ2jD4PcCFBI2SKFC5Bib3r2ls8d7WMW0IZCAyDeKyAXFLXoh13ZZdqM8Pse8ByFPIn
4d+hOGq/MxwBsAp1J/u8bj3T4J34M6B+5Itmah/72PnIhsyGI5n91PtTGbj7aWPD7LgCwI71Y/vv
vak1jbvfJm3Pozm9YqdA/5wePfGSvoGluhT58l7ZkI5fLAmxvKdaONtfiQClavG/kLMK+c4fcX3l
MsAJsr+gEjUQKxd7RYI7ibIockRntFo+c2mbX+aW6+ZzYgjJuX/pkpECqmKA172tIyblXuXPCrQ9
DqwkvwBuYO8PKiKxs2pbrXQNo+yT4brnyJum4QhEBLXiZH/7oGpmdYDm2mZZknYFQ09egdaQ2WAK
6PzARWrQB9j7mYgYno2H+PMuGo7Cb2MjjxalRp8FYcV4wvgPSvQKGiiLkrIKk4K4S7PlzJ+N33VG
jgMjK9J9eXtxQCbHB3Kskx98nk4hoaH7m7oeXJRwORdQQh9HWuN1IGnpBfIPdWomyfKgWqdFswVD
WO+24cOv6Jvv4YtmsKhX12/ACQTsfZWbe/V0jkQVACwUNwUoPQmYeIEDsE/OLBT9jKMKXy3qK9vV
JwzV1JHs22hD6nscP1JYuLUDoA9ABUVzix3wqKfw5kERIQzq8cQlmCT/XEmC7rgnBDNTRgRx7Ml8
Tm6aSv52IqvHNB8uZMdF9WsLsVI/W22QmBecivM7yZFYAHL5qDqqOcI1IkejijwcLnZcv1eLKUjL
JWw7PkunvKuyy5BKh7kqLb4tPhQg8C7Y0dONT83/R/P95YQliMPptNZbkVVTSOx965P7DKgME01Y
nPx9JAIimhJz49NP8hoMEwQj7k2nSOesW4lQFbxmD7lMFOg8R+10HUqtSeufPoX6DraQsCEb8H/S
N5d3+GhuWwHZJWHFQWp9g/1NRF31f0/nGrWtIn93fTwSxFF2ddOyo0kcyWJ+N0sRjJEbQzihC5NP
+4Q03KgI9bVAl9c2YHrSBXc7TS48/BXU9jbYM2gkjgRGzaKo5+yYo4TdRZzlMJ/ONZ8F4kvthem/
NoPmuOj4At2BQ+YZx0IMPMYUbAnQF/DEhEOIyRy8NU1OAZ2CUVbZiQB/frdHV10oxRYXMyUvA7HO
0UQNt6MrSWCVXBpHc97D5vL/fROXCegtXc0Q70LuVs+a2aw0EkUq9jT2UpL+hChh1FE9TywrpKLo
9/kZ8cypi1I9klGQwyUVTuB4mO216VCPLbMLRYbSaHiBuFPAgOl0g5QR3oLAejWI3GgcjddkqSKS
GZp4T4pB2Be03ZfLe5Pk0n5DOF6QMl5Qc23LPC8CfR/YjhiWpkv3Z6f1KId5N9/wRZ+iDgHH3wqd
7LHkkmeDTLVsMXJV05phRFhFVQfHUiILrm5FZWSwYAM5QdssLW56PYDGRqj35tPyt3T7hyiloPz/
dLq1A7UXvTJg9VtH66Kj6PC5E3/3W5zi6KJSr3ElwqwET4Z1UZNpP1IWSjHeusPWxf75LF9AbByq
pTkNPlq17kiEojq5MPH1g+AS5T8LCp3KvVEiDzjHViL8AdHXNJ2gEUaMNZjUQNYRGhTcL0e9g/Kl
90zA7jfZK1p5r391R9MWC13yyV8t3x6sJm+bSXYxbNX8U8dCWMN7dthL4dn/RFNWM745MXIcaXNS
cACdgeTOLkpOC5OZ6+L2RyFuXDvgtYIk3HJz2QjRCxHmHl4EAWUrAwCyxGCLCAcF8KLfYqy/+Mki
X9xI5pzXlatTs2betGteV9mDwzJ3PuB2EH6G/mWeUeNcOr+/PutwWl0wme4X5V6dyqSQx6+IwzB3
2qx4DpkIK6/vNFR73l3eapZE57TJiRBpAXhTqMnEfkqH4ETOYdLray3lDl5MIXc6o15E7hYaJsgj
SXyzcwhbtN8Znl/0dCuMK59va/7medEIrSlDd2L95NfoVKIGzHEpMvzWH9Shuvq4xsB5TxdFF3eJ
D7rxlSvTTCZYcg7F7dihffe/tamh5+SB4uyTFISTS32GNkYTCtbLKcDiXiowSzdi/hIKvTtoYFqj
4Xq/jqbvpNdvNjFaZd/tDmnafDmiOAkb9qgZRqyP+D+eeP85hIhYWTc/gaZt/bpyaMIjS4zlhDhR
+Rx9Jpfc3NSd1QwQEfyxMWGyQjFW4NU4n97qW9tMoGWCu8oFFCLc2c61WuHtUKRNQiiAUDI69sL/
90pa2/THqu3hFBO0VSYqv/sxNFFLv4VU1wmmfAJBJQN3R5VsetCdnqHgC8kvFdKsFo4sD+XmGwbB
gZvgZ7acCa02SL4z/oK8KOs1kKbtEE60CQpt5psuTT2l9wVIZ2IDXrg2l8qT5vSKCmXR3DZP5wDM
TR3PYgwI8Fz2uqqe2ttGy5MMvUNnQc+AM6g6+VVcJ7xa5lUpeNFAbIam2QDLX2DfmFDhSbA0pD3u
6g/VnQn0VqKRsGjQLaC+xupavpo2tFPjnp/6bArIpZPLWsTyWZlPwI3vWWKeI6zWo7k3jfzWY2dB
tEY4DIHVzKGOKK+2GnbioBQbggnLgZo5/vQTxP6Bl3suA8hxB5jdk1QwwpQv1q+wumoY4EzWijdg
iTDlNPwxPfqJDHp5oMKZdThlQUIfX7O8cFbf3t7SYG+Be43RAf16fzdkeU2SOxz5AN8PwCNPlosC
itz46xd/J1Bu5/nbYNURHEK0eRVkOo+m2nPjH/kMOnfuyvc1hNDltgrGT4PfL058f8F6b2UpmRFu
RRBHLXVYGkG2SL0aPJMHxYPsUXb9QIlM93iSZwUpzIbAJfsroEO4oXBozkR7jJfZaJw0PkFLIEqO
e5Yn4IihdAICBq2sldtNMGxFimFPmzfYDCqat5QUsDxnnMOzwxOmn/XnCybfT6iErVCA71wlTFR8
NB1uG4WgK+mXuvA/nszPaamnAtiJ/UIK6voAyve4o4PVm5tt9amQnvzlrRztl4NJLKJI+DsL9K55
BnD1yGeS+5Mw3t2RK1cHbKki4RBw2GimRW1EtF4IlgXUmaLp/iY5ABrVGWJS+jcAMa1uO5YgLVLd
fg0moNjPvanrAHRnFz43SeLAvdWvUktK6j0nQjKElPzsnWAjY4X0MmwHNDGmikxzwIF7fQ8JkwHh
8S+7Zhc3d10Hznl3U1C3wJyudNiSwg966+W6hyWcXpqi+7SfvveubBZbjlo1ry+EHCEjQRtdk+Y+
gyjgB95RHfI4oAMaxStyAGwP7kZ6eupSIzpjgdAO4NJ21rpEi2iME28TBrBs3hjtV4IilVo606PP
mzEBy0pij2PcpxWticPz/onEsfgGx+3+6aX1Nulz4kK6eM6ozAB6V4rTuZ79PFBtxd4ACFLSHVok
cj1yYtJo1iciWFf9CImAWhkjsZkoknayQ69njjHhWvBnomaQPwv2WNgPlG75wwzj4KuzTi9WlAl8
BbYRfoVZqt8c3RrdtramgpCz7uxsGhthrmoHNkYvW5b2I66tBnRUDWJ1RKMYQHvT2G/l16M4bpRI
ogh//PKet9bf8y+f+GknQRrFXZ8ZlfxEmFtnof9AWY+TunhWp1zD+IDBIZHsMr2Za0HlvB+bKB53
j3qMVITnnsC2+kpHxISL7JW9G6HcWPG/1HGbMIW3PLyrAMbmfeUeVlz1v47/SA8q0JimhaDvHSBh
ovrVGL5Apc7AczN/uoQJFUm7OllapsR/9LGucd8qr8TtDtqlmBIRrJAEBEv+aDaFFfnWYza2yIMy
brrPrJKZ3sP1P0ZkfTdjS55IpC0067lvNs6aHitblN3PS5pl57mkG+3MKf+kr91cKryEaAWwrBs0
gL83jzQ5myXsh3R5+b/vKe6yXujn4F6k8zS4h0FqIRi1gZoybRdDf1MZ6GJYXtt7GA54HX8aANPz
iEOgOy5FXhHSDMiatBQNHU03LeWrfYa+BPlMSwewQGF6Hj5Nq8eBQm5FNkMIbPZrtwyiafb+tDbc
f8RGQQjrIW1SGtUZEv7uEgxG35LMmbRG6UXVvCXH5Y25yu8iqA/+cVnpnZ5Ylu4ZnOndq7H1R19G
mSqVu5qC2rxXJyPuCO1SydeHQp27rHhE4OLKeuqGFiSafi/dHM21gYqQ8XahtGzvaTZkgE0263rY
uyJSVFm2pyTJwDMHvU9ZPLINy1jeTBkfybz2DP4pdk/cFXXmXyGY26nTRVH3omtHYRTssyB0YeZ2
RRp2xi2/w7dq02tKK4sQO9vgVvSn0wiHP9qGtxJuUgmUGzyMvDvGT1W7LQ3w6tmZDmMejpWLV4uJ
cppwuWc3OpJHSFL62Ewc+1dao6T+upY3Imocz+XD9F4sjWlKLLZXIyEbNzdVe/P8chbyET42SfFs
P6HpfpFxvThsdi3naw1EjyMP94ky2hLdDR8+zzSDO1XhyPC9dNmAen7xwSAEzLIJjUC4S85og581
sUAnmRBblib17KObCdUKQ8ZNISpgzfmXKru2iJ5Q26upfqw6oD0TnO/05Y2R/t/+krsZgzGjhXjm
Rn+vEIDwqaqjmiL11EVsKUzjS5zlAV5wwIF13Y9u9KZPagaFfFk7gLLETAfUZLXMl5xY5kuHz/Ds
0a52Td8rkxrXWFSXLvEz/XzfPGLAnrOflNJVhoKRCl2F663f3xwmVOCQJjgCW8YQfiqn6jPM40rc
2RMr2J3iUE36/gIq9WrKZj1aor5XxkD+tOuQrFnHaiN2RYoV4uAHPxfiHGxlbBkWd2ud7xwRHlZu
mIw25J+mVOANLSuiXZ2rLdVGqSOmvRK3gy5RhGAo8mn9Qhs6VsBCVkFIpK/c3/FbEksHm+FZ9xyi
/rvVMna4dYnr73XBSOhm3xZPMcNNJm62x4R7scmIZD5yqKORYgDk7XAqk5hW6IK/enn1S/1buDgp
q1bAc7Yj97EQ/Foax6c+BfGvm5Kpq+DiRpKmltCPDvOJeKKau17blKz8NzTt54JbXjQOqdUSa/T8
84TzIt9S6r60+VON5kqt6MJdYq3PEMwYqkc/XyU+nP2m9i7x1oV0PAfWlWOHxohC8Fd1NS6eXjlB
Vvh2sbjUUh5XChvOQ9hohTbaFHj4fit8gOmMCJbB1dLCSJuKl3q+4WQHPBFdmoKJHEpJ270bmz35
3wDdpUUlw5uRyLqGm5+4jQV34i61ReAnAGOPCLzMCzThWVjzoeIyz2iTl2JA3pKctRVni4Q/Poe7
R16XI9r2GZxVqMFRBhCB6e8G93tH5vEagK3uDfAh0gdbx15L7pKkXwgOzWoa/70Vpg+xvHsJu76l
ktDf4t7FP76ydiAp7EtDpzyxIu0J7VF2MEjWAF9ShfDbYJXxOV/9SF5thXSQK7w9eJ+orKeDHnNB
mtsu+EQIEZBGT7OcxdeoXHJeyzK+MQDqbzV1fyFSfLCi/Xr93nLd4EBi2i/Ynh8t1bjwfShMCmXz
M1VgjBLRDmBHGdALl8uRm8VzjY5m3jpT1Ull30f/WFxqVU7hY5T/bUHsSBoRsx9HqaWBlJykmOmc
gv9yUOUFpYifJIEO6Y3IJafGwgN4ZqmHMXgjXLrJl47Mbcq9+0m3ZjiNsLycxogK1s5O4B9yyT5p
KcGikDVNw1CstSmzPII9euv+VsGPEyEtgHZjjgCKgN1TSnlQnu7t/GDejm3KYt99GS4pxYEJRexy
qbA9Tb5iUgKwqsQa9e/oLHEBFAmGMSyL8WfId+okU5nYlTM8LVdKyGcvMpwHQCmb5bEZa4zC6vGc
OZmP1FIdp3RQo9lTvC8hSCVeEKBUAInlXhvIhwXGUeeNYNgi6mwsyAy8St243+qbNrqI5vPBGkpT
fyo1XZTBUC4gtlysaFzw4kV7Rn56j2hCG/pazREhxKF/B3JX63WMRIjWt/LQyPJfBqr3Bbd3UL22
3XA859Hzkl4V5jSyR1o76fphEFeYYB+rClFwdCSfgomn5FHERI9V2SdL+G8xW6etckhLkJNwfIqh
JSeA8j3a5+gykPdn6PQWc1olG17X24Li52stB2m+nKytVPVP/2JAfiB5QRirQ4slwLZQt2fWH5az
FifNw8qggBIZEH9fBeglyKtir0KP1jCijMggZA3XZ3AFCs7tcxh+GMOsZ6+ULoPxqZEn6DPgYWRx
XEigEvZmYigLSs10Vyj9djf1/Qm3SMBJa8xgASekBGVcJcPkt0P5T7wjQ5KGxqy0jzCxV8eLimyS
yMFAvUron9qvuV6mlBf1HbqCw500OpPAnt3cnroW09JPevsa0LnZLu6cABMGpBusiF5DlzKdSg09
kyKk8Euw41FUWjGuoAGmdy/ibWJwyXpfSrm5UTDzGiBA2DSOVw4XPD4WTyjgfqbf9cnxV3RiyvTM
DduHhzxY+X12CihFpEgaioKAnYdc9ETLwym4qzvw29T+SP6/Ct7SUQyAoMHGC4U8dFfa/fXnqcSy
zz3Zd0Atj6l0Gr3eih1yF6AGOwqOtELTM4p5LfeOsJzFCGwzbofLWgm+q6u++mi0nB4pJDeVE77i
XIlh7RsAQZsL1XqOduACpLk0y5w9AR1XXeYyRsnLpIDLS5w70Op5sinBsodB8Tt8N5ga8aWBrLeb
bsg0VFYJbXQQZmm957B1t5UbdPivQqzSQV4uwwlwWrYwoZ9GUarvnuEE5oLHuda/yFAvgdUkL/o9
Do9EwFIOFUVTmNzrKCd7PZqxCNRJvmLVv6Z6EhTOFghh02hnP0A7fmg9ubdiHeNssYiejzUf9Hxg
9idmWOBqnJ9RWp58DsuriAfWR3pPHswRgvYvbVS7Tugl7nYnG7xKUS19XfxJrmVLEFifc5Y8qnTx
IzrwpscQrRCeuaLmH+cWt5DGTz51pJVqptFuVPU/St3s3uuf+Jkaz7xMciTPuJ6dmQZl0YYAywBs
bF8l+kczt2mmQs0CA+vDBtJFTChouQGxDosz+ZgX8PnEhb0BL3tctWlIqiJ691JBHCbb68BBoGiH
cc2lpVxCisbN1yR31vM291IaG5uO44R0XWuXHgAhJr5E6rYZ3Yc3AulpHMa7bx+JrVOctrH5DYFb
9Lj+p2q9hVmIqvqJVIEN5UkczTx4H2lj7T9i1JliudzzZq6TGa+zUo+oB2OpUve6doXGF/F77i8x
7B+790OLaJU2gWBCd9kQL2pqkXAJ/MYYwCJNJy75Z1Wooz5NAxTiz31M5iyyuhPgcBz0VCwUa78o
5W9Q+9CDfQsio8SLerHyIU/GnDfVEKDbkm5dKiGd1XUYoiIkZShydHe3hieXFJYixddxTgbE1DH9
O/syP4EhyKw+WyNZLZLZByobfrV3ucJejYVfrbK0oSW9anNMsq5BuM6eNDFzQhq/lQZh4WfZEUCK
ym0d7GKOTyJDo9w1/85oIk6Im9yGKAD4qzKo1aLP5X4hr194geZJqRXOLvK20o5qsivEWTgkfV2I
H0JthTJqbhQBUIc+SXAC4Io41gEApmQN8KQBWwRPNlhkxVz1k6cafIFd1mWbazA163KeGqu7wMb/
M2Zu2+nvPbHBg7y5KOvxZKoM1d99dAgQsyc8NfQDNUVpJlw0S4LZ/4AHsTdMJScSSoSmW8sUYcK0
HO4XM4jiipuna8j99H0jow8m8625vPP6lCb7T0tc1o1TQbBJRWYuMh92XbutOxtqqUNsjF7yv//g
vTSn9QXdGl8DpYHhGsr46pZvFKu2fyB05DyGcsfV9XmFzfLyMBeZ5mIqqq3CsQvSB55Hw/MS3Nkw
hsciY5eMEX/K/48LpMKpERuy+lZEtBCXZ4c403LtchKjLF50Y81uStDM6e85+n8j1mYOs+rTVAjw
fb/PclPFBWybxsZ4yIe1HvbaF1HdjNVaQknNd7pgFbqHOjT9xTtK6xsjIr++5eKPdwfbrg1yag5z
L7LDEnSP/M3PnZlipUl0E1m/HKp4ImL3kQ0cvtABz2uf1ZwbRDWru1VD1C0i6bEcEKkXOE3idiK4
5ff2gw0C9TCwPzRVlQxYQcBeeYvbtJLKj16Rj39EkmIuC9LNvk2xjJhIXpEoeeTsAIuiaK4T4pKa
gDgQL/lKVeWsrCmWUuj9lJojczt4SAGqSKUZ/1GvIQJKeZZu0WdbrUmQ29jLJn9UT+wR6EYGKlG1
DtVWIjXAFvGk3diisg3NITCkc4lt60xeOipIDUIKk3bXdY2/+/EY3oAmtJ4/FkHejneMyjC1CXzy
ENn+78LZXtJ0U0IJzV1uILAlc2vSsU/kQdcAU2c5ahNNx6FKEEn3exkqLzxd/TNFR+bHuuMvI4AG
gKrbMq5O4K2Tt+58MmrpidV1TKKJvm22cMBZAJojHVIbLY8LmUmuZSjKbWXrhkFqp6NA27RsvfM1
nL1iVwsB32mHqFWQlstbV1IBJ4OH3tcaBFiLqTc71Bp72p9TRpYFGSei/1/PS9YVbXKCYGXnRrsg
aawAJASvwohmV43qYaWueQNwlwn9mrAGSCmNtp7Al4kdUzRiZl7DJ+/9QJAi3DXV75Upfqcg0QEG
kEw99W+QYNtZ+/XiP4sXcSzvZDOOg+SNfhTM+tr/bNSfJIwSz1gjYouX7dZt5oLQoEdB/eiQtd5u
zYq2VMRxD8IOYuN31ufLYk/LVGr4ltprOoewamBJaJG+sG/+KL6J2YsBLplrMN7VeQJKyn4A0r49
l0bpGbSYOAFjRTJRJXzG2nLSmD6bRUBIHH7HrR9F1qfdiIDqFTquAmUrtl5ipeOqBgWbTjivZg8k
uj2XBltkXs83tRQ/N6Sn3+EO3Jov93IxIO0YQJnznLkX8fgQ5aCg8NtFbnbIY8gy/OXvKl8s2qr7
yXkr2ZiU8F8PCQ9yV37YDyAaxVQ1YYzP2mr3hjtdX1Vni0Ah9mbZ+SE55llA89RdfSEvY3nu3DRZ
aVbXb4iK5O6GL6N8QzqyjDnw7t+PgK+xCBXfNWffcVnp5YrTy1O9jwAXUVCo8oMVG7omuumlkPCK
euMlTZT+pYAEzz9Hg7mL+KY8aRV3nYBW+npzXVgnbICh2p7ikZVpVDfTrRJEC8xWsMMAJWgMUKG1
rjO79AZD99/QE1A2IBajdz6OHBO0tiwRF+x9slEzlukKS/fxGaYs8ggxY3F5F3XolRtkKfyBN19Y
8yNZZRD8oP9qQIjqyISnx280qIVNU/9+ZpFILVsabjf2rKlY+GlL0yZaPiuvzIZd6Ptyng7M+sPh
A5aFe8L6VOoX84u1pxb84yXrE39kee/iBwWD+adplELg6kkGaUVmGG7ITsxxYATrAWteKXsO9THc
zskEAqK7VyxkkqzYmjzhyQJ/rNKN49BjvOY/0AABZR+8y/VzcElxr54XRK/rb2j3Gc3d/SgO9pf5
z+c6A6NfNdqRszMNvUOyli5N2YbWgyKk4bwnw7riwtuP4qYjhQeA8ey++Orx+6HVOfgZtqHiPtTh
TDrSWI4ybxvlemW8DqAYAcEfZLBoQWfV7gJas38YQ6GYa3FB/e+2d8q9kCpjKgT7KJk7EZ2SYH0K
WNq/ZKSHg4RIb+9QnQNoIW2/f8MFotNpNP+UxnX7s/L+wa3puHuIZWv1DZucm0bHScFLsr1Jg37a
IeWxG/m8307HUR9vwpfW+4vWSgjg+euwAlXM7wwahAe8otbfHauVBQl+Z/5x5HemqKPcMdY/GMeC
nMEwgfygejiKShH53jihOZ+178YbExaT1PuwFE6pEwqnbFRtcljaWDEQhT9dmaDcVYh6iY5eS5UL
2Ldbayg3c254YSjWh3JGQk0A5MU8N5TApamZtANH6cpVwSMxz8SpZazymshWw9qiEGYj0gJdFMLx
ug4Mb8N4XsmGMfvPu6F7h0rMYydQeazxxBpjsjSr18AJCMhQmwobUqKOJOBnRhqUFamOexhpbMdk
fNQjK/DFnskD+DKLjWXPJNL93z9kBxtVSrg3wIRNY3cBESICGvdc4kLYnLNL5H981idR0BEI/t04
OxGOSdI6Rw5yYYrRR3s/+0nIeF3ac4kCcnVZrpCMoVL+8jUslWZbhkTUGyRPdL0fb/95HRJC3Bg0
fv5tcPrM/MF7K3iEO/VdqqykWqzLdUFnrjrNPC267wyavMZ4dTAgsPUPNPgQp8QbqlcmFJ28m6ga
2kCdj7Mro/nPUsXmtrmuowW1Yn86PxOmaAB6DzT+3aUdPdO+CTd/plHH4rGphuHHxaNIcyu2Sa7/
00mYGmDGVl3J872NBR24F16ulKolMb2jbHJXV0GDhfw01NogtHXkXxIe4NJzMN2aAXZKk9k288QB
ZuJKU7wiBxpFtjxG3IFKsaPm/J71NCVTL8uG6K9EKDoEDKaizBQxynmGukQVEl9kuREd/yvJq9yE
U8p095XxxJYI9pdQJFKOk/lo6h1UUORWCzKPPWEiiPqjR9D9uCkADwK9q2J5bqVwHILioE6inj+A
d3VOTJ4ZUVTf/2jCsr3kI1Rsq2Ghh1daWGvSrjVTIac68fWQ8KGQ+sCRvPV9gPOaYyy9aWvW+g/F
aV0027u5Og2a8KcyakFm8aGV1+qbA75xKpf8DJ1v9S+cZP+OzygJBiqeZcpROuac0WmhdeI5ofBU
j4gC/JzOpU+gr/mxvBuHxnNVj3IVr3U5jQFxgdkN99kFPoLPV1AHBJQa0KCYNJphL4IHQreRFhah
JEQouRfumGJCVQ1j3tgse1RnT8Wr5WawkAByXk+5AopWbfyKr9qtlq2+UTa4kuc9685ig/jWhrfi
x5gHt4K1LTdNCK53SnNi4eAV9hGFN4vOLzepWKwdJuOg+mD+VwGecAiieW9SHle7Sj3NZnq3su0a
Wbbi/OUtbx/xzAJff0MYTyOA8SxpBqPo03kqzX6yde65oA0obsg9r62BonBWyje8jlp9Ih+jcoRX
3Jd7RW8c8sRMWnW7PLVFtSLqjn2MdgmjuP0w37hY7ihFEA3wJfptAoG9ABrs3lq2AedoXv0GTE21
chIGc5C9H+DwkP8t8Er7/H5UJbwyjejuAoGwjRSGRyFLi9rCNyGmEHPVpeYMxWQk0pGg+54K6KgI
tQGDzz2O79zCbdAWL18YjmsW/BYQhPV1hIU29mFS9d0zUO0eLh1WissBuW5FVZCC5P1JQjOnoEjS
mDX2oL+B6MHj+UJkpLRyhDQj2mnad2XnAKPlzHagmpuNH/2S6OsVw+BRbvRbCo9SkDRIbBQMZtr/
tVzU8woF+S+e2i97QRtxvycLmqHCYCGCIFDL6jAzQ+WBd2+1wuYg+if9v5yktcZczlwXFLVdk5GG
mJ8/rbLRZe9BZwtz3SYYo+wIGC15OJh9PZtQblOqAvVyB/9SDQls08oEL4IQ9GzF8tb5qaYvrpgc
HToNoWWdqiRSTCJgTPzpy+kJuZcrbHiHlvtImgr5CKVik0jY8HZftNtNPsrijRD/SNZ0Jv02tB3E
iBQIv5rFjy5FTPIpYLrWb1ZTWRhBcjgCxwBnLssNIICzH7T616BrXDWeu1fBSihgr87NdlX/FCvG
vWFgxJVpcn45b+JcaxwcZ+IVJq3GM3m0yJhqtrU+EP/9J5Z5mIDYfYHhRwAojLwIZeUR8dovqhds
DXj5Y4sPrJn1Dhq4awej5jWz27/+hAm5h68cxoK7tbyWoy34PFrWW9HIdWKKea/6KRnBpj6LUB6o
W2y9seDC7baYfgEeCx5PhYHbVZ58S4bq7HXRhVCgtlnBhZ6U6VxgId1ws2A059bQNbpUEYr6tcjq
DsurZbhEwdEKJ9AupF9zpSO1sqFvpCj7SAMK+RERrN/WiaTzgOhr2ZcN8GMDeS72uV2df15NvxMC
ZNitv8uQt/bdcuZD2roiJfFtqHQIO6msPDlZcMVtsSaNOpRtKCgYhZ+x6+uh23H/5wOH2Iv0T3Gk
SpGuk6tnhggJRrE7ablDWqwK9jQihcOW8tEzI7kRXjDaM2luL4xfDh/XqFoWkXFEENNUxtEdoi/P
M8+AT8bBKQK2+TLwn5QVpvTTHI5fBGVYq89wRRUesFg1rUMhFdysPnKMiSe5qK4RgMInnZfJ8icC
bI5ESfdukfR/DxWTZTqCnFHG57ZpZ3ThlS231litxbe6Vap1m0qL1E+Sav6y7cVP2U24hyfy1E77
02UqiM4+6sLhm14nqAH5RpvkMgKNk0ahkyc5oMkUzzmAOxj1LMre/btaCb7sk0jUwc9x19OyonUZ
1ar9Ld/Ty0IdAtgy1mCZqdx1KGCEOgQS1iUpKwe+cOjOUUYmtTzqX7Vu34nSrcJKPxhrJYo30NmR
CpjKv6kH3iXFcMydHENBbjqwYvXNU2cdcf2JZX49pw/2EkwI8Q5Sh2tu5VKpJbu27woe2vSmpEil
AOl9T8qm27uAePjxi+N9lPRhH9832Pd+7/tp43e8IxU3rpwkFn+eUXqJM6Z+Fd0cvJs09tihDHpG
8Bn+bfGiHIRH8+mCOFm3/gZVQKfElHlS7qWg8AhdOAU+fGElZYij0i7uqLImZA45pVu0cW8b4wY8
Zt44lgyESLmxT6SO3zwrOYtyWuNQ/aJyLySZuvrYjCQU7Rb4XJBwK/qoLmP6WaL6144PHbu2VqZm
q7irbUArz7XwojGRiGfCctVbgHOBHB21Dml//F3sedhC6bHpkL9/W1E5+ctI+EAnp4czY3WKpU47
PVdqSisyUNjN2HmHgcIsxHGMU7Ssic012+6WyuYpGXUHkSVjxGVPn8clBu5Vb6sVeq/JSWcbYg54
PXwyCMpcn1yxrciRhmezh9QNdH+MIVlYel5p5u9sgJUVraFtxLPTnBuowEzCh40VMed038WNquyC
ZrdL5jI6g9jOpaVkoiyWfaYBNW6P/PAVGmWj3QdLCIrQF1+n8/b03wNhIN2lGtBDoJGb5oQlUoEs
nJfPXy1Lr2OHoVyDFfCsgGvRSiLZTVHpEK7V/9dYG7bW0NwM1qUHJZeNhgxuXdhyyaOkj8msgChF
wbkkF2Zmf4QEM7G5yRAt2Wrk7U3lBjxXaVeFsIEUDsf7LuVELZCIFxAhXsx4UjXBOXbYINszONx6
pH4GJNcKvd9fvbpIVZ4RLS6+skf8dvFJ/96eMYq498P6xpv1iUNgQaJgtj9p5pi2uDsLcLmtZzsF
FSsR4cAfmmizyXVPgzmDwAltfiDr3ktcZnTX7q8Mn18X8R0hPnLd/d0xyTqagEZK5F7ngZJI7fq7
oQu0XpJ4ZU7DlpzdBk+kC9v/29D3YOHnsZqJVRyt1MTSIzjZgYlbejk0A7bruaS19ZFeaNGzfWLz
dB02vf3QXo3sojQ8RlHsIyyTSnn2uiZZPYtmQhF2ozUo/I40tBfuAiBgDAbaFrDLl3ZjE8//tj2s
t1owmTTciPbMh+7eJUXZgmfOqiHul8yaL1sUc325PX1Skn5CeY7dVgBurYUz0nxWN79Ezgym6dgb
9NaeKVW6YKtWtI5cZhx8ko7f7L2O61K28N85YBFj3SGUb78woR2+c3adUANRMWk0HxxQ+4Xb0YF7
xAj6M2kGklIyP4cor1+sGBsLF8fP6iJCFwA+/e56WS5ZSNWKf2nqM3s/UkAAQK0fumpDLZFzcAfo
iiHKBYB0jaumWs26KKzjc8Qim+WVKW2NH6HHQvXhE1HPYZLbuaq/r8Cx6bWOUZ/6HnEEfeM4pqq8
bEHGBzK7uByZy2ksyd1UTnEmf13I/BWoP25xkHO9Ei0jjGOkn2USzpbBR11v7HwQQs6cxSxVijfy
AQgCf1H+LIPbx/jvmN/WvZqZ+CP/3YXK0td+IWqF0Noj4UfXHSslGoSLSKl402dkUnoQCJu6KqGR
xO+VXHBL1pXmgDOCzR6QXQW312ov29iQvjrrTdURCLR1xM1WlEqZLFFGIadeXB6246xeEoS0bZsJ
ACJ0ramzLCHqPs96K/tAAyz1k/pAhveAuVucSyItDE3Cg/wrHHS0McHZA+SwklqGHuu1MQLtn6Ao
i2uPnbdtVApOxOTyVa3/YyzY/6cxf/an4XD68l49IvWLPta95CXZNMPnbLg1hoZic0FDvQIywsSX
2gM0fVx1Ay48mmmvdpx7i8uABefRdEXHuruNlGbOodQZK7CIWZZUftW743nBvUgq6GB2gpgjk0ze
Qavmxn9kahuhUEVNMBftOASX3iMmepw0mtRF7H58SvncOqqMu4Z3QcIDJ0OlbjXhDTgPqvV+dwEs
r4UYAyUxuovgfY7lb8QkSdOsA8yeAAfV6z2uowt1J8zhYV/3p/JB0C2u7kOVypPZkyST5Crk+4u3
wNdvqmyaZ9kX6ExbjoQRRgxVQwg2ek1jj0mgaEl5JDWyR0Slv6iQMAVAHhqKqmv/nQejQvjMg4Wb
7wVl3avbES/y4U9y3bc1x4Pv56HVr6ca0GIhgV+h1wXSrGfe2P3x3BLpScDcMnyXOaJWHnV7CzaG
qK6yCJ3lyYkbq66nwehevHRwVuEmb8i9jtjvyUzxsMQdsJb28CsSuHzPBE99qnDE9FHFDvgkwhIL
gSNZVHneAs9sHylgnuTSYgBTieW6IgpHdhYPcdmz6/DFtPb991fzhPj9RDJHurv0lD1A37527QgZ
TGuQnWMpuqszXgWYQLDLEOfhnM4whUmbYjEVoVAC4zXLbx77N98EesEznV0EW8NLhscB9Gp6xZ2X
Q3/vIlrILl2eR8XmUaq+TtFlY5sFsvEydd0mHmBMEz6cYLl40+UuLwUELOfvwrRUGozTrvD7JHEJ
YR39+iD1iqIYewjg9yZy8zpAkogau4YxT8Gw/O/ESnD9JcMz6OPzf4nVS7uRyrnOFKfj+J42/ood
ZFajYL4SxIwuVF2e93Dt613A+J943QsWbf5hhki9FKkrIfDLRwSwNIw19AyFfcv7uSnC0vgARVFG
AilM8q47CoSzKZzarLxc1ZOxEBkmEVHaAIewtFzEMc4Nbk0vG8MAZThjh3/nZWiM/TCYtZyHWC/u
0kBpIBIjsJWVaiT6QhQPlXmuYppEgataVhYPza5vjHJS8+BBIT3jMwgsshAjrvJOzm11R92yYJQk
2bnozkxR+s+QNnQWx+++mLs1KZVSnoEmzcB74Ny5VqMtXKn7PSTX9W7zR9BlG9XuyO+azypxQrFZ
XbdFApygZ/ZJ9eiLr4eMtajZvCjaGz1MoQP/kDi4RS49/wxcp+L7p7399q77zirBNmyZcySOovWO
CzIXZFGUhiaIQa6U2Qn4HyHAfodNKh44YXRz0IRHYNSGL0qmxs5ik1F9eqU7pQ0qcc7vJYpM0ruM
tG3VbqmkXnuxr9JR4kgUtudslLvU4t3cZyvYmczQfCrMwN3uJUsFvXatuzIjN7JpQUciIg1Cm/3h
itsjmmFHdGoJppj70FTIzb3wOx9iXnE7ZaV0OWYJ2E5ZRfxAgSkZk0O1VSN5bHLWUbuxOL33vayf
Js5woLguxNnNN/j0Gj4irb4DOzIp5tShF7P/EOS84YiBWmtVSyXioYoVJIIy+pvUxwVXD/QTGRpd
vgtj5Tws9jnSC+XJjk2rguiblPq9+H7D6Qi6pah7oPvvF/sUEt2Zw15JhvBaJKK1nnTMm4fkSiw3
UyMI4pg8voAjgXL1hyR8IS9vady/mEiqEElHNg/BTDHqmJa64lb4Rmw4epAwxErtJJs6YVLH7V5p
YGtFqv3TeQcV6YyBP8aV2bB4UJxj2vdkyP0NTmh+azCVKmgnnfpyZFwif76KFzrwWYKDzccOzFF8
nrAspBoYQwZjs4grb2V5OcVwsxGGUItj/UG9n0hnZtY3eAU6wekgmYXHnbxY4YQL5QFRAx0obWVf
/SEvCJjuRq8J8w/zKGSPc3j7hn3P0GGwNNxRuo/Tn1RSgWlxffH8S1ADxgCBDbkMLlQL6Kmb8kee
8PACor4YqTdatD+lFVBhsGNv8u6vAsAtjXp9bBF1l3rmwccfwR3W8q7k0KD7GIA+1HPYUat5VVzs
pticNhH980sVO+UEbM/laLmvjCF1IJazfKZixWyVcRIdlWZs8yQk7rcCOCgVQ2QfSh0jCgJInToo
fm/V89VanYLa8rkYr4jT1/YnlobEZzZDaQXZ+/lMb03HTLFExkt1Ed+EMNOelRfeqZ3xExeOJeuJ
jr5iTPGNwJEfh0s2mVwRlJ0claZ1bXQVsUjX9JrA+heKpL8DlScDUz+eRqzWlCjVQDYEHSdWzZDb
HdktCXajC9azsjkY2grywWqCOM9NKGhHU81RrSlQzpoSPd0X8IQfLDtuhYI2K5NM4h8lTkd0UqPO
aFt0FcNxEo/CP2hPCLLMVEMfZebSd5j4caMJisIkoeF101+zwQrMcB5ri8/tBp1xDfbVGPQ0z8y3
xsRpKHljk9sCupkLjDlOdn2e8plnVTOwIke/KJe15OZTN2/AJncA7MvzO5lxZA61a6QnJ768PoK/
QC9j6JjII8nAIcfz9ovO+3HQbfHTnS7UjIw8UrSpFxM/ZuR/FK9HhAvVgmp87jEW0d5iCmm5xVKa
W4c3lPGAhJcBPlMe0Nz8oWzgtp4aaQ2y7JdakVFgWM03CYEeWJEOoqfMrNuOWjVSsY1DpBIUz5vS
N7Fo2BoaajDWm9U0Wd59sk/HVSHevDWB7FuNvThzu70TJW8c8scqLGMlIW7oPtnqOYzWgUyIsmDw
a6ntqodmxcVzTZaApWLNXjRL6ShUPQ2rJw0SFKFBbg7vMhNUzhyoUI65hRVw3nClMChFNrSPnxKD
Hu/ohgcIRHfM8vMrcrfPzQQKOzHBLB+C8y35evnMysBcNkpPa3+++aLVfzu8ZSCYccBh0QuanF19
0XbrRK3+2hZQ0+4yrVdy7eA6EtfkBs4p/QIVxpFWAQ9awlh17adupEI6Vc60FfUey88N0BoVrd3s
1JonnWyxa5e7RrDkMb+uLC3ZBvSc2v3XzJRmEYRXqh4aFFpwMj7vG4YIBI6XywkYopLwpbuXDPVu
YoUi4U6LkETHGqlZ1/M/2i0az8lzLOpFeLh2SbtQyfV3ShRGJQZreIzM8nVRBkeAIA5sKw5Z/DwE
DDePvCoZw5l3G4ZS2iAdmhm21ymj1ZokWatWrCXRH0Q89Btr7QXXHKInOfpINugNvRwnPpdXmSI+
dsWtojl24vBNiWYcSzwgbsnLUykjPaQVR79tf/gaATw4VTzF+j5ytXRYsk5lah8oGzMLwbX7bKDI
gRKATV/9x0WaCeUm87SBEDayYHD77NuEDZB41Ea3hMi2qn4NXN5PPBha76Jg/3vYym8BU7TuCm07
YmZJN5LrH/j0M3I5XrJfgPSQM89uw/2f2EtDnbDnZJFHhHwFxkbHeqfD5idamxjUsX7dU+Ionr0n
WK+LzbaS9T2jEZX4oXA8dUHC6FO0IAve5OtnCb8HqsYfYySuCXfJW2BPJKFxEJakJOV/dQSWmujW
il3w2GzA0MGuZZzmfw3moEYRBXzKfwx3fQxUqIvPDMqGzLNqT/w+DQ+atg+Fqg2vjKeTMk+1YpS4
2GWe+RWk4mV8DVY/h+w2eHm8D5VaEik+fE+V7QGZe/ApBGlKEQkH4MV+ZyOyjSXR7x15zK74a8tI
3SznuDR9JnQf3VX+TNtHU/DXAJ95RhchIEEyjOxNn3e0Le39E7mzGKR99dDllCq83Gie/8EfXUlu
8itFlY5tnFhTrLQe9fsGV+0JNddJfN5GYdzYeQ8nZf8Dg7Abk8jD9Ot355WAwG9hKiaDGr1WmzpT
bMQd4uqndqBqV2Q5IExVE6A+IMuh9p+TV6ERj4p6o2YOXV7KTjmZ60JKhUHz5Vi+qDWCZTMZAEK+
8fvAc3NlL/gw1WSFpDwJBFZxSFwoyTMTeyJV49M3Qek7CUGJ+acsoczAt002eg88hgm5B/Z9Rp9g
5SZ7NZmHt/MYgDI8IVTkSHmAeHScvJI3yjLOlLMaXByN8jhTBv+yfQvwHzaKalxElvsn0Xdu7lu5
Zvmyp5c289ld65/o1+JrpeNjkAJQuTKziwXMnSgH4U7TVcHH5bwFkgCwSekYuBDWghbyX3TysEKZ
Rq2jHcPzZeqCRHwO6lKM7aLiq1FGEekO4g4Sqfck4tZU2yA5zklfAgluJsokdNpGsVUGOSpG+5U9
99l1M5p1wz43XGhrf73X5LC2CKbCti5l/dJs0qKsY+Ez21e+l3PAwoZcpgsa61zjS9Oq8OVvrIMa
ZLrKkh/Mlb5AD9PvsTpFi+k+tQXskWSRmbATgbNzBStcNFVm3qIs7/OOnrkrGt6Hijg7lk2o+Q0L
Ygszq3q+E2S/PR3lSehkRx6UqQZPuCwkn80uxWMYpXplhh3MAD1iwtrVDfNUUAlaAWctXDxuxFFz
UEwFc2CfROHGV8Ad/W7iEET02+i7RZ/D9RS7qC8FPAE7uGfNc93CdCfA8yd2ALenuHyh0fvhQgkt
Bh2dfripWJG3NTv2zPNPKm6WylS/+5+LuxnfWKFMpMk57dvksWv5g/Wd0AupgmqkFDBcXOExWSp9
10SJyFDT0H2N/obZA0Gn5CqeuNQLj1+vkUXPa7MANlaG1uupYR/CflNC5cBPWyDAFYTFR8n20yji
Ga+a7ZnYlEcotjkUpwAsEH6Kw+VzWdEA9VOG8OEbT85CGynXvreNpOZqYT+4nQxUiPyr8kXW80Ni
wL9HoCsLn9uPwuVPfgwM6lcQA5dStuCE/7YJOxH/urAw4I81Q62MCjL0jXX5OePp7pP0Z3b0uIMj
hE706t+3d21MocVUP0FmUx36oUdmOKdLV5XYuMUqiVAbiAEZFy0w1UxwFpPidLJ+hReshbh8DByo
/vanpO22FNDEAXHSHUU7W6+hDfaSS3AFobs9b6wu6EZRhcbRbJ8oyilW/YZWCm/wlNm2M21c2H6i
OuX+UcUbTkv8ckoobDuwfXriC0pU1XLB3QbUQ+sh/Z/y8JhhP8wSxTVA61SCZHfOMGuoO41Rg5mm
odgpYo6lOnHW7pPkJnl0KlxsvNP0k1t/wwFSOyLfQZimxLt7L0Ra9C+GoB2C1T1ACwR26wWOTTVV
QAZ1fTcCfrmKfHo/4UMRTZH+H73jIno/Rscr4/Jxfrls/hwNxG/HfEZ0jZGJr1pfz2YiBjDQG2ox
X3+xTYHAIohL6OR51cw+cFxMZGRL8AbiLdDwR7hK/OqNiwNUdxk8169TkZy5G208vFvMGqI794V+
GUNpRlDol88fUXqI+AbjpMtiTg5jmE3Hr2sXQwxYuwjIh/mC7H4H7CIWLA6LwB9bbZUr8uIsBezJ
A6UtUZcqn5Y3ZeyP9HH4/v0k6eBof94jvzWRe40ZWYIY7nUa/smOKDIninpgJ7BnGgtdYrd/Ivog
mc6l2QiZ7PwhkzMMOW+E+OidqJFNBl+nC9qbAKqxoOX1G9xyiq2io8HJMqGFg6vIlQvtzOAavaGQ
bji6n2GTkjR418YaWy5+Ukav1Xe8GINJyTxPe0LnDXLNMLhOqPbNKkb3mVETycSbfgfyTzmMY5Lu
n3/7VRmOzZOtBssLEHQ6Isq0aORGlmdACdXwQk2vT0QB2j0j3UBWXom+Q70Mb7XElTpVmPu3aKAF
HnGxJMpAxxUPS+fHXLArqnzIW4LB07Qrol9jK4MVWxn5KNWEurxaKwQ8UCYyt8qpm5iQGINOh5oK
8HwUuuQPRKPhdX0AAQ07jqNjT/2qFuvTF4dgthLJn/t3Ac8yl8NCtDbKh3kCUo/2fmJlVFWyw78M
pNI42d4ODXAO7+IAtE7SIRn2oeJum2Pv3I2ERjjcLd7/ysuL0V49Yb3MjBMKDv3IWYIQyoCwZgkG
+4C2olvIYCZpmPdAJaOe6RwsQEjXNWUusmF3W2FBy6cdUlaoKBRWvITQ8WvdXZbWNfJOt9fGOQXU
T/yKpBvdUeNru6wEIcR6vME8CyLxunuG/WTu/Xxc0bYo2JcJLMVDJvSgQ8p7mjCxhWleM1lgS3XK
ukIfHs8s9BXlNm75HqRnHzWJmxY3SVzANg7eNqeO8J3Yqvw+Ap+ruvO6KBhTRMgGAK0gEIUh1iCw
WDI55Mq9CMY84++IBqYUDFMTkSJiE+juLIx1mL/UaCqvALQ8lw5scziFIc3VfXH05j+OfvjFX8rg
u3Lednv4TnJaldWArbm9cIx/f9h4D3WzIlkANhrsh3gVUgg/BBcamRAF3R4SOWB84QNJCvz9YQhk
Xr/I5V3E3nDbhiXADtRtFCjbE/IsLb/XtXlCpM/Iuue31rMUUX3td9Ys589iE43NFPPPHddJ6m7q
2erdVeB0IRQuRUdRfnzQBZW6mDUvW5DO0l6Y51nQdnfId4rA9zby8UbPTXZ5ybZj1vFaNKLQJwHE
0HyDq63dBEMBaRffiiMzCbOO6aPVJPO12dzIZfQEIkYb/S9NnLoXbC3l3nJdmfcN8wTo8Gf5rnht
SxdQxI/riAQAjWzezLcRJHskKzXgiNcodp0Pt5a1xi7DnAqO8cMO7IEfsJjczIZZI5h6d9U9R74O
HIpTks0D/vDOoOdh/btu3AGNKujJjK75iiUVtxLdITmxg0dkhsCc79n5YbSYyDAnrlJRCpyO6fFY
zGy97hs3wGUJTUMPqv48HqbrYQHzMpmEYznPek+avkPB4bzR8soyDfBw1SyaIKOWR0lK+Ns8y8i5
oMBrZkua3+zKGRy+RMRe0qBeYCbZ5ZTBEax+LXuvrfJKuPIGcQWldsoavJ1TXyl/XrtxHBD7z6OT
gKG12EpupYiScfztSnYWQgCsxd85/KIP9QjQZl3vw3BT/ki/oLZO46WgIpMLnxR6P70TrG+pZ5Vf
81K9Mf3LxCYmN3B8iV5+tDXG83ip35GS8Ia/R/rIKElmdfywg3pfnJKVN45EhOAVE4Eu2FAqWTcL
ge4Re5UBen/F2F54NWmhHSkcC2lb5KHIGyEr+5QdxinKaBTXNiSYPgkUBkz9bprgOKhCOoOWxNje
Pu4r4xnH10eKy4MJsusv9p8r17DrC2+tejW02HIS2eYM8tyCQL34tc4SNV+BIFoJRQoI5KmUATHR
YDb7ceuJlC7CmvRYfrKIh/Mw7And9i/0EXW+Df/j9hToMnwxBcBT52EKAI4DRulrIGKwxYqBcosO
4TyjQedPX96OMwjtFUGkHoQsBZyujwZzPVr8sKRYfM6Z9jnOtULYgpX6BssEL9OrOP0lgfhGeaxK
KJ3HhSuTK4D+uLV9N3n0l7XKRV/U9LJy77liA+u0VbxoiLVbkDwGMfDcfZYG+uBAW85rgWm6UrYp
vCpjm477uscsL+z2L4xnafrAIcBdO2oYWXKsvXub8BzAjp/gteqF8neM6IjnszW6wecmpxKwV4WH
GpekoqmYzrt+n0tnQCuFlMgwysdkES4Qft5tVtHqQG8E24tPDBf1hCC9H6glHkgCmxlpquDzgQku
PDH1oWSw/zB7N8/zWHgdES3/lhEvInHouZ8cQFdmaoKHf+h2cVtSPkjyqErhjiZ+rE52BCy83yJB
KfGTnq6r/gOh0R7cn21ig27gpJWwkYol9D18jaIdpa/pRfekbHclFRxyj5r2YxVuvhh2BqeRajVF
QPEZ8/s5YeVNnXbfAkB8Y3ZOCDUCuK1NA6t3EjIgZapqFiarkohPeugZ/XuOTCyZ2xkmX8wvtLhp
CKgblW+jlOBQDSu9eSThdDf4AOG9APf44AU7CLKHRBtsL+Tb3jAMzlvQuGKJw0Npm0cThZKQCxOv
AIXzcsUNwzgRaeyCNzeqZFdpi9J/VQo3oa7S85Mj3P1zt1K3+5WkAGDaiCuVKK8po3otUjyn4GJb
7YNnby1NxjxZkqHjYVecrk+Vrs5JY7vCPNOPkZyah+YzncKeL2qLe9Vnlj9r0Zg3Pu88RoQ8unu5
Dh3HJCFAnfhVEnqVup3inQnV4AXQj9/Fht0VGbO4sM+iaclrqqJQZpCy2doaxqbYXhU2QC8ziwCx
ErInmLbq9psmU4Gk9VkarU8FGBXr45x7aZEvQxO3k1ntfjeL8QOuZrA0GiFLCjVJN6GaXQ4duwOT
mqAQ5eMcVYpuk92q9W62Oqe1T6DuyAREt4s/eM0VOZuEOtV/3GqV4+9JShfKK7GVo2l+2com7Prg
0QDvFcilvo90mJrmzIjjIpbQIBxXyYMFBo4C0QH525f3oHdrEugqPxgGuyCT0kWz3eB68Iv5Mlrx
tMk4ZenbjDNaPr0KKz/oSQeiBsgQ7u6knhV8N0VNfEeVYmQyCzTQvZ1J5d09ZdfCOOG8ZKBqdJxW
UkAJQIi8mi89n2cSvh2myCEBqPUMjKBOcCd0j4h0roLzTnXKWTgo9WDlinDv/VmoxqSK5cPoDY2W
/MypWMfbx0vdulUCBv/hFRB4vv6gVKecNaIR+ybOB4No9/ngpoO/sSrlPIkNTbMD3cIdyAvAf1r1
3trMhJTKRDQdC6TThAKn81yHr+Qgp8cuXObd3uJYw+cJDuoSEMBCjl1ib5B2x/g0/nMkDzCjGHdU
k5AqRbmoz1LZGfjj6LOihXIbuPgjNgLW0xc4aJEH2R2F6vcTEOWFob7L7EYyJBrrlCXyO81UMjFN
Fip+VgoQAnwMzbrY36I1+BZqFnyq+OhUaFoGeKTO4HhoiUgjjoRSlncKYMmX8l5HD5xBVqTWv9gl
3R3WgWa3Xi1KgOEfBd+xYbWt7uoKU5vj73e25r+8SVcQmZmm49c5i8/y47jkq6cJ3RyLWDhNWQN+
Q196xdRwxTMbBwP5N0nQ7I9I7Xi/auoTmJNXFrZQlVaop2hojIZyfQ6m28fLSn31j2c5OufPWPAM
J8ByVuYwDwyCxmEKvwniwqDJTwVVD+BBXHuQFVMZAzrT3pKAvWtc29Y4mN0+03oQfUifoMIkK3ct
v47P30xlYbn1jKPHC9v6PI8S5ct33zmb1q574/9+uILsg+6qcodIpx5EriwQKbe4/FYmQ8MHyi0U
/D+55IiITC08rWIauo4UybE0K+XCvqfFOkNBz/6rLloqTFXWIYUaIm0IkhoCiwlhCoeawsWMjbnY
zskc8HPRAmQ7Elohag6BlbQOhTpMwB5bNXSlxXpvo5MZ6sQSB7GYUosxiXGr679jShGUZAmwuWAp
Sbr4sfio5mc2phOOKlEYVxAsSIIB7ctgQAoMyepVCjhkUiJP9f3MslN7YLXcBTB+pEEe7K2pUOgh
Kjb5MkSff30vgaWyPkYu46Z5DQdnEYoD/BykpmMeN0TOmKZQ+1Ba7+f0eV8QjZ1NmDoTLTimUA0L
kEiVT1nhvR2PBPNLFEcE1h/u95EcxNR+8A+roLOA2s1Zji6qhD/7NKc1NBhMXVFYOgNz15NPHyQx
hg4QMM6OjY+WdIfJCl5YQZg8bZgVPOpjadt8l6+P89Ob2JXS6Y7HjF8o84vdSsxvV+rHk/c+xogQ
+NKSSma1qBrBWIA2nVrd/APWzOn7Hx/VovaIvoa+BSJGKL7kzPRvX5WGKY+alICAEID+wGAuCMyE
IbCsQM6DXOIpXJp6vv3dzvGXujFUKvMfgRugK5lHOvNi5hP9pv4bnsExNYiWbxoFbKF1qH1QNuN3
DoxYRs+vedvPQefINvvdIz2C3aJ0kjvZs9ABx+eU0OlLLQmwup9JPW2mPGPnfhyg4taTI3saNLZ6
ITcoj3NOqZJLdoF1KHkM7DyRP0wlG8m3qL8pueCDTbZ2tfn0nXLd4qlJtSE+L7isxScNfi5Bdo5j
jXD51Ge8hYnezTUUPoa+R5nWgICl5ffBB7yf/yuiV77du4tKWBXHdMhU/GKpNdqWeFb1B+QKERdB
hcXcQi3VHd8MWxR2JECroi+Kb4bKV25LyFHb8LFeuAh0+cEkva/lGR6IEJPKu4EfE3HdgdAeCpdL
adZiRC6KVI/K4US4VJIookUZU7joiLRVl8SdnnobXT3gmO22YAzQ+X+PQ6o8ysniUrEhC1semH/T
VVCscuJ5Jfs4X9CkVd8lcwsCQQ731qw4AA+qkrL0bDkOEhzgnQ0hwYWO+S7uOkahdx4P5t8pSqhh
L/9mH73Ru97WB0t+uZg/LrsylnHQIeVNHTKKI97h+g++VxXkcNZ0dVPyS1nwiO1CqR6bBKdZGyNc
KP/8Dp/qzuu0ysJ6XELjKlrGdscoLHvip8qONv3j0mCeFjwpSXWlOy7HDOHlOmuRCc/7D1hzndKS
22HakcmNjXKjU2nlmaAHetmuHaxHxlwUxu2Xif612XEbqv3nbLmkTmz+RgEfyFw+Pt7gBncr1ZGD
zAX02KxSZCEM3jIHnRE/SPxRgZqjVgS44LLpHyztahE7aMBvTmjPSbh8+74fmONHNewoxJK27T+M
GoWNJ4yvSLsqNmaaN7KdHFMKmzT9Cdwr9AejlDyMAwoZSZUQq2AyZGYsKEdurk/lLjkcvhD+mB8a
Y/dKKbSdKOOYvXnrK+rInZVj6G+k4rmHHzUi34JLHAwfcUX4uEnzolds6DzMatP4uDQmkIHZhb0t
yHdPgUC7bqBf6ffyMw7KvmslIr9g/dg0Aus6mzY8pBdncTRvwEOm0/Yk3rDEa+XlFrvdFq0+nYoM
it8C3LhpyQgNmlAMrrdDwIf80HTsHLrWNO7TZrKeJ3tdmQAvHMFlbYLgnGKeDfuQUk8fx8wqI8nw
fnWuHehLjo2WxhtcSGsI3xFgdntX+W05KbXlJ+qalzCasj99G0L8bVqvs8+B78qFNDv7QbLJzei6
E+f1xO+JfTR84ac2mSZ1wjiBDbwbk8Yn/sx/eulTpgL+IkMF7Sv3JkPZABDcZhOvGADWfOm8sYgm
lBuDhp57w/dM9s5BMUuf7+kEnNdoZfTbxXJ4iBuIRwzhdOMROIOaR6VKgIMBfu+UWbtOWAxrnz5E
lUhWzXLNyxVXoZxI7AU01hMhwZBk7bJGeaArvkZF3fuMRWi2h9INzw5j2fo6yFjrHQAjnJ7pNHva
4VM+VcuofWdIsAWDqSOk5gMDr3bV/g5cOBC089hDv/52M5/gmCiFBavS4eqI8lbnKZdB+JoAwFTY
SW/ZJU7wFesWrHalKD3ZoWXxxAW0htLec208dlZpykA2G6thhhVWqjDbLRkS4jDiMk7ceTIsTdn4
0W+blfuvMhkGQwU0QIMA1olV6pauuEOpjAVeEE0aa/DPUDkUg8dho6tTMko8GzCCxF1zM/pdo339
lX/Zmd6voct74taDeozRKESHnqOF4GucQQbqhxprRtGZdRPpD36SvH6NFjvWslIwdEvsHytk35Na
KslxNZP6RogRvEAefOiWox76W98yc0rmOQvn8IWTScRQajV267+0nzbaKjBTvprm/HnY7GO1pHEs
f67Swmh/SPe5FzkEUDVVEjlQIpXK0V4tW7tEDGLxEARDWseDdCvtEE0lpwW5qTTgeU7cOuUz/SIu
fWtbA5sUbnBsWoO9ZpkdEhzVoHEiYz+nLerzFHhJ4ZFoRjNorS27SFA9/53Y1aCDhZTFUHUydGGq
XYFf3RFIP1MhCv5lxhj00tKp4P7u6YFHW5+gQualIHHmIYA4JDQ+nWrA+zrxfHi0jj90f9/mQMGk
OWDSljRsf1hgbclXf8Z0NrsvL7ORwdYYRmeyq7edqu/bewm86YHKn9ivDcqqSE/l7j+pS6j8ZPEj
36E9zIxNCYX2umQs9MhDoTI7mH1GY1saK5kp55M3shSgS7Ao08susJ531aaDFyq5B2mxKczwcX9e
pAZZ3O5aqjKQd2H7EuuqbhAuutwojOypK8mPMi7nP/jYaZ9hNw+GJARupcBfOnhfAtrlDYT5UCVb
bsyrwQd8rKIBoSmT0/pDfRZyzz8zPGWjwCy4qaXsm5SAgS5K8KdceQzyLZafmbRnsSTOzMnWJVDd
5LuZ9CzTJ2rUjXoK31DmzK4gAWR5gTDA6l1XmaqsgzaMl/wYV4el/q0GntnCFMl3nEMTSpgt1rPi
eyF/9g5KMcGe/vbXSbj0cpTdJ+eqM3kDwoVH9ydvuqZZGWyyFH/IZeJvB9se8ROExALMWknNrGv1
4qbeiEGKD66i34RFCQULTeTfphfZ+dlDHqq+xxBNVxoHNatWeYXH98Z7hMqC25i6Q9nbymc1jXje
oly/U5wBRezwBKXIH91CR3/PVFpzs1I2P7xmlndfk7Xc5ZiKhVLgxsflXjL1eCWMt7TGgRM1JIjb
5Px57ugDspXZn2NXll9aRFPVGYAFE0kcaAa6hBzAp1l0zeFUjqv1hjuM4/y5ixxR2MxuOtLD9Zxy
PVWqINv40ZL+qCpJD8LLJbSDhd+3JiKsNdQJnprafVTUvV/zBMoPuMlFJEWeQmxof1zOp+mYm8p6
Nr6gSmzUhHACB85XAkJL01CepklSqTx2UTjAhYcHow9gPZXpWUeJRRbNwyO5pyDI2qf57d36rCWi
7vrCes+kP2rxBQp2Ghpc3EyYAk+hUzPFoTgX65hAkAs2lwuuDJiKAeO5Ci67GEe+ShDGE/XbvC09
3zjSaMiUSCymHAShE6zyi/eMYCYuVRKQvAlLp49uNo96l3PoDC9JtGY8IP4CqUG+53EdKctf5jhT
2+UIqz4SFzsx+ISH9zCq1pzNMfKxj/UvVIa9hTtIcVoRg6gdd+J3tQir+yHLOpWtQPB5ebc4/mpQ
EAhcsExv3Ro/JNa66vZwOjIff5wf5R6KVS15qhnJ8JKJ3vG4HElWTDFv+Qx7uQ89+Goid3ULXljG
AWy/eB8JoRignIZysvnaFzc4fHR6quWNxES9v9yYkoMq/TwwNwVjrYHqL+Wp24omEl7/HX5hBu4R
rjIhpjlQxG4z8QFyg/QyyEhufDafSTlKGDrkwxBrHYeE3FKngKMUeXiZJNSaK23PxW9P0EwH4yIM
SyO5TidKxOReB7DWjZUosOXQPY1winq2ES6YAEp8JUlMMtlbDZqhUT4KM7zMbDm2K1QWR+qIbrfp
wcQlauT3lwmYugEnfPYrLJHYDjdBVdnuSHNoCV805njlMSqhi/DPGC32iO1gN1mmzmDV4gPeWzdM
NOJ9VZw7NPtcYKM4gvj3p7qxKm3Rscq6FCJpRTX/excnwfchdyIPgJ/j54z5UZOA4GZFUCW95nTB
cHnmcBBbAjs5U6C7lRnRYq3rz29PktgZfVOmG9neqVi/ajwYQnne1CiWSVR0wafZbJMyEsPU9Pe5
AXefksi6fE7WfpQG/w1KT/ooeVFE8W3gOaNV/Ip1VgOXjl27g+oDTSqNcS1QD49dsqLPOJaKQhcZ
7nuItgprfykiv2GX1SYb7XsYJbaNsyMLnTceOxe36i7ZbEFPZwb74eLHXSYpIQicLiUSRSY6JT76
akptZAwWZURYYKyG+YPufy5EGYCs5Jm7wGRTYRxz0EqJGNRIf2NQaKsLVsPqfdyWOIcc7N1qIE5S
4Y40Xv6g3EUw8A36VC3KWEGC/F+cFoHhj19pIiUH2oVJ73zkCwvm+12WdbbaNT+yGzqx7sf+oXIv
e/3+vscJ5K1y66MQn9vSDvgOfGOlECLIUu9cF9tZWRq3QWADCwNtz9EZD8WvWB+RHqJbtY0NQ1tJ
cl8JmsioPblwjGZWCZsppMEQbcY1ufSZ8dmWMfvA99yvU1/DC60oMRdCmrr3njeH0wMDCLn1Wp2r
VGPseK0pjZLncuskboSH4LbIweexhl8mLH0fGq5s/pu9a82tvknD2JvpEw5GdnW9Cslf1MWx5FLX
XsdUNFje9lLEQ714xTRHHtLuaXKBrf6V2PdpF2iw9NqH8CMzYSCNKuomJFA3uHBEN7ZVbnhxi/hj
Gc08bP+zuROjVqDnMGWuCfZut4BdueWguY1c8rjTRvt33r4+cBErR7tDTYeN0X2snVm/Jh/bwmy7
V1ze9jXlKmJDyex6owEvSNemoGo3LuD3BQIHlpd+wufYN/9sJlJfVadJZyx4rUVMR61BOTjSVwTh
WeJEFj/ixpiZ8lQrCBMykEN/gUypyqwY7npbElzuRCIz0iFBQTvJ8YGQoiMTYGDS5BBQQ2U3bxWp
ebQ07njw6jy9m0xuhHa6EwI5O169Xn2dql8RB0Y3JvZfWK4v/X9MxvZyQwf/CufLlzs8pVCVic+I
HsVaz24oWx4czqJGYHRmnNmKxJUYlstLVq50v3EZJGvndNOC37egOgHCi9bvniK39gG3Qyzjz/Dm
fC8vJj7ixFMW9vAhN49O+vSeysucqGMDKg7EotpvdQVGCkxng1Hb7TGHNr75aUdXIDKC0WOOueLM
FKiIrmA521AjpsR696WsCYa9Yvhhsg00iAHFc1R8Zpe3/92fJvzSVPItukxZzzhsvf0wlO+X/VHP
XU82yy9of3R4ffi2lQFFIIjwN6aOx8qvNCn09scuWdsgDhyrvA7GwPFqdGxjlB39aYO3G9P0MFyJ
40txmWn2DQxnjSkqRIg7bpSXihYFbvPCSzrFe45jkctfGtVgGYewx95FIBYii0rwAGsK3DzhuG8J
axvCKHigJm6zg2gQmRENI+8wcR26k+bRayU6fu6H9UvNK6qXS92F8rVxOfHUqghwIQQ48ehzliEY
UND3DeyUDP1rLu480+dJkqsE/V+tol4aB7ig4Hg6LjcZFOLxmi9ErMj3zxaluSFDMvwXD8+RR7tg
8+dQcBvvswGDdUPdUjR4ZjrAf7hiuEIiX7FraBTSR7pmE8eOS2Cu9zNKMQhNLkuuR1LgitvXaiv0
1W16j9OIMevffKH2CmD0hQEXvDsxTnGA/z1Ir9GcoHec5+D5yHXSosVNsuUc5dhwgBTXAlBwrZnh
crCwduQDSd7pQHezdzhMJ57s7STPl1bdb9sDUwDvqwtOnBrfLu2347GpdluIz6LXBaQzczaFS0FO
Z5Co0S8z5LngVsgHEivAYyDJKwFlpknAq9DdNFpXGuQgApnsMTSXQArQyKL226s1aBnFmP8668q5
54DfkCHfbS9FSSVPdOmoRvLHoT2RWJKP1qdR9uLo+KpuOKEvBo7NHVKjIw0WZHH7Y9fAKaUFjU/M
aXZORpStEbZBnflylmZt4/JEHk68Fu/X+bALhDGAozgVD7YaefOZjcIzN84mb7TAO1X+jETAYWs1
DAEke4wQGW/erC2cnOUeUC3/rb8tODoT+k4eFvkqWLDTM85rAwTnrWnXYsO7mi/WwAsfZNEJHAbn
7Wg36JC5AbEBQ+iaCoY6TBz9576mxQgWw6nTkTW86SIYZGbaInzAXZi80aO6kxo03mDGjWZTLsAC
K6bkfJR6vWhx38JtIkoNuEpMpCqHWNEVZMjFt7MyYt3uUyeIDUIzSKoFansdYqyc1yedpOMqnM7n
V5uYCBaWYjLP98M2f6xAEb1IOxJ5oMHZ4IZr4fbRa3BtruXxkxh+Sp1RontG1MBfJQ+QFyHpa574
hujyac2G4rpEPSrkqrh6fDxnO61rryWjvZRRks64Qn9jwOMdr0yIaX1OiuBL9I1i5EGQGOCFhmZr
ajSD9nRUnrv6c1bsCwjLD3tlsCQ43ryuIj5xUzIEtmpuKEkmDCJAfaDswCuG9U0O4dWq6hutrH53
m/I1ZtsJF0BCBZBLwbxSdQaF3t9EJ/lOhfUQmKEmn06HoCkPZx86URDFIRsoqzqmb+ktLXCoMlMX
BrqVuqG/HnznFcuE5XRljp0EU3H/zNDoDrfpg+WsZxspyqa3SewzqDzLBiJFYEoU6wQnrmcst5wQ
SnAlP1XDv5sXkDcH2VU9XBTKmVQQLoYoMUxGES0t+7I/l8JSFevfiChOlwAiG1TDsQNCk4fxmpbg
xITU1uSuDk5eRBvKYXXD2jpH0+0YnuNl5w8rSQwUgejC9iLlVaAy6R3rYCR+71luV2ABX3THoqZN
tv/elHlIpAR1i/RyKlSXKDIcXc14KslOTcJ5JLobpRtw+D00XO++yHbIEDQ7144QxKVqeyEO76Qr
9Nx/yyDpfx6dPt36AtVluT2sK2GGLi5D4JZnrrlSD93qwON4282XOegtvvq/6ktdqn3UBt1I7POD
dSB35zrW/gLQorZzO7BJpKeE7P2r3YTq9e7gl9aLNpAet1FwGguZfjzjIIsDebxPcbdMkaepzjMH
Yu0lA3xP6PWUPT109k2f4lzCA2CKQvs1CA+HPv1cQloTQF2pWuKbsiqF5DTbSsZRThtLwmGA/bhQ
FgZexGWY9TIh56nlHhmohqqHFiYHa+cjK5HnNMPR7pFhJGgPVN0Uagg7WsdfmjVnzQTRszqWaWyZ
f+LuEhJLsJpCgYeQPV19urBQ6hXv6Z9GPjfYxg/Zrl81WZrCql5Iimte2gswDAjPUyd1qqZPWCnl
eeybSBEVCaYiWu58n2LXNJxw2u2HyyK/vHHypHBJF8DLd08uy0N3vAUo8SDOJHdRiWQSuuEqQNg8
4/viFeb+1TY8n8pVnrWMHXmOa4incbGtXa+st9Oz61RbBl11mHN1BND5Rnd8UoXHQ80DOpYJPHPj
oL+zjVWDYdA5fsim6UfM7kCUpl8xAezMh5riiyF+Dag2NWhur9+xlX6pO1xV8VEd9vR39bJyJMex
9QVgOdZmdZtEa3X9ZI6Ad3LBHmtjBduYboOUct0JScMGIYuZlbOH5cYrmGiNt2atdBhBMDgjsedK
qkQe3Ijhj4mDyrCb+K/ve0fHwLj//DhPxG96GC6e89cy92WYvsJb3thJAxa2jSgDRmoAVoMz/OIY
e+NFVSghA4KCGzz9358rzFnvXGVDxLA0fFxp5bKLPfvTX6zw/gG+MNdXIN7TgmQP37Mv+pyKw6TW
3Bni/lYWWC2DP3BReYhLgm4SgCYFuUsBrWzp6LB/cuugYYqp5RTIGSl23eo4ck0Sy+vHKdJtCxI4
IW6HEI2cWA6w1hvpyRAl59iLSuF9ZFvKb8nMYqSUTrNjy8haHeKxthnh2uY9zqmz7neXZdp7eSHb
5sgvpfKpNLK8QWqLMDpbYxqgOIuH8eLY+r09cVKYk+ss0o5uo/tqdHO+3zc5bvRg+2ykdM0/agJl
SNIVcmWPhTzZKCNRdmdzHGu5zmhs2zITq4QE2SHggsvuHmcqDrLR25uQj4fJWl/m05p+NODLa/k7
S8EcKY5HFxBrHyalDH1zj2+YCi4zzMcDs/72lW0q62/YNcLTOT2n1+f1FS1R0B0k49WkMLI6bi6b
AS9dmSOmSz3WlxWwa+zIXKCQ8WDzK1rAaCgqx2MdaDjPIPMTQkfTWKeuOGIAiKRUnxzIrLIfq4nt
iv7i8dC9+930OAB2GU9efXIiqcSTBpiUL+4dwXOLqUKdCj0wVthnsSypgyKwWrire1QZcTSrJX2Y
a8Rmre8J43b56SXrap4fd6gyj8XhsZgNUkWm71duAOYHegZnoS5mKO+mZw6R89FuHhA3zpwm3TF9
8+gZwCnLFA5AjtHAGheTGOmpkJBtK+PRi1le9wqxAdcqlT+y3q0r3XqAfZ69KO8NBAh3kSHF/Gci
TO65yIy/N+F3DBOcwZDRQ6dAk8KoJG69OcuDbtNI7KGiMo5IBwkhmsv2sj7mbgTi9rqbjtVCMb2h
Bifmdmkz8PouuSyudMw6M6oxIg/yPthYT521nD1OfJ9tQrGj4vs/D8iZ3W2YW73Bc31RCVpgNt8h
EEIBrIx6Mn5XL18icSGhBoqTTmV8jqnWeyaWpwtlBW2BULxxK3MsWGA7wu2g9mfWYNeosrWK4AXH
or2gcMVcyzCNfIqYgZFSUHY093CAVo23JbhKBPNHR7pzQW9G2WRz0kBvACn7U0yOY+nC69YOZnlu
rUAmOlPy2Crrpuh3hkhrfWDWlkj878dwCt8IblucfcajpyFCFiU8x5iMBTrbi9EpBflweJsxYk3U
vsa+VDFqetRuKup+JbdHP5SBEa6q/5Es1xGB9/saUg0r8gnSZZ5+WLW7Ka+NstPYemxoCcrAJq/a
eT32x0qto4pDSmPv6DDQc2q1k1rfJvX/bXzz3scvROgJqpRr8nYSgadIDmmRu7R+zTgFFmzGazIu
/U/xgPyhT+6lErz+jg1Ca0hIvj1PoWWBRfvhNkxsoa8o+AjwjK7iLmVCoXNYF5RnTvYPxo0+D0WE
J1OalobHwwVegNGgCK9XqSm+Q74rJPlVNqIFiGW6QRXWwCnsnHyg6beYyWryJNagOzZuXWuJD9XD
8uwkJgy9fqZP4Pm+/xB7BHrgYV6ONOH61LNrnJfvkqR97+zOTvcEvOp5R0zEJcN1ywUwMmjzpCiF
7o6a7D4SCimiCeJdDlSUSIosiGRmtGIB5P70oD5bn2COu0gfF7oFtXCmeSMc198zPIEygulhI0rm
l1BeUwaZsBj/BE3oPHEEVfvDczonR7YGXq1H9Gfby5I0xM8JMfoQR+UzHuH3unQEhsuqD4CzFt3x
blluIaHSyxA63Yh85lK/PxcfCWG8wWZEa8FxBNL2PmQe2eTfP+x9vNnC0oFCXrw+qStwJiKq5Jqq
rUfXW7/nvj1at4/GdshDuzAkKKC0aSYqhKFttlQzFC7RelcHAq8JTq7SLDH+bVF0q2BOR/N5/NVP
7roXDWbcssYQsSSEbFlHT7bT12v/nF+qF46324P6aKIa1C34cxUe/65u9nk1CU8CVQ99tJaoOgzi
eWfOtbmwkKcPx3gskXKL4jeXumaCL9t3LrNppw0fhdoVZtOTbnOhoXwaORvaG6Yigut9FOiYNGix
FH91KJoSWXMQYbcQWjBFX4Wp20QX9yF2qLV66gYvm2u7bAQC0qq1qUQQLkuw4Xi9Kj1lFzrmw4Ho
vvhxAZcTXtj4gPd47Mh/O1TiQ+y6XYPcI8NZoAcrEtJCCzFrbFqsc/+GNxrw4JWOSkzNfycDtAFt
9YfTH9rpdPfLmyRN5Uf51uEwHiaHojyhtN7c0LocEB9CdWBFBer9RiV+SEOMTlMvMB3ilZ1ARktV
ijxjl72dGX1u14cStJMQ+m5x2C9mC1rLpROlbqOgmsCIw/W8R/UGH+91ndKe/gF+uNEO+K9bD5Jv
FcO5ZptOZEW5OT/3HYuFvyv261nNFwPwJ2iPz8OR/TytXDl0Dch0A2CC8njOr7P75ZDYaZcrx674
cr9VsBhsJ0XL5OkHcx5iNkaYA1QXm7/MPlr8JBArOE8h+Hy7R0jeXXxKKNtcv+lQFoJWWzGaTObf
bSA/5TX3T1VfMkO1Z6HFZ28/MSn0X1WcfkY1cafnBKXWIeseKoJSqx4cTsNnkf4LHMDy06t8jHUm
j2iWzWv34qjxxHZxy6pUUyE/DWzZYNNM8Cxjaj9Uaa5GaJqbsMZ7mV5ecVOPi7jSqRWp/kXstjIy
T5L41bcZb+17zp5rR0GXYAK7oQP0xRVOh5ISZYx5btz7lFj7WOoZ16pQSlcNJd77QGZXV6lIgsS2
13oe37hXk/oHgSx8fCpUIaA/j4vUMeL9EwPL3oQMSL40psIqfdfPFWORWk7oPuVMG+taiGbeycjT
87Uu5HVmuPgtK+jnxv75WOFHYpNCCobAAkrSCH9FzElFXu7np+SIKs3rms2jS08s+aDGyu6askUA
Xw/ZCAf+cpSSNAwKM38gBBiGs/tCXrmIuoDNKNGg0B5h/R1pGEUKwm51KsLPqZUunbGiO/SDo/ol
L/9ISurWJGP5BAjGUQ0OXuzfvknGqusq0LWANNietAiJiosFzg1J5WeyiBFSg1yfemRFOalhn8Qb
SXANOMhLxqWc9dwbZnyq9Us4/lVluWDtFpQB4MYOKNlJEIU/AEtRr3vE0YaEW7o3PS8zKIJxZJzI
F2ckziCXJI9S8Qh5Pt2DQwtJ6ILdrt3DWgVGb0qi2iYvgCUr8AMMy3q+JzvOKOdarUEDoLYm92M3
zFoJcoqeqywV9GDus/y2yGeT8IMTGOavibiSL6dkQCzTJosS6n1SUKhNTKkzNDUfHUi2pY9DXqqx
7U0Juh2pgdXgLaAOi5DjjZyYv3k0SCzzbGki1FQ//Gf1hctnztiHXkLhRx4g+s2LwtDrTSJYtrcT
mLEvQMUfafT9PN1v/wAy9rXRxoSuhq7+juR2RzyItQFaUxtvzcjjbuHy+iFs97Ezv0/AUzKr0KE1
IhC7OdnckqUkzsjSoxVBIE5RJAqQBPoH70O2mqzQYvDRmDUunSjEJFDM6NmasCek7MjtIeAW0QF1
v9mKXThs12YR0qwrVAAYr3TtIu/Uzkia+H2Nb/z5lb4VXDcvRg50KTYNt3XgJJ/czI55X5mnRvB9
/dAZ4LbkMAm64GCm2NWIK+wibYIQRaHZpNTFQDKjHe5MRW6I4CO68YyfaO7cXa1BhJNN1w3Exlhi
/IJuwkCGuQnxJ8LiQpLpjfifM1Ki3hdFCBbQiW7iFZcR1TyTfa2q5jURNmOPkSCK/B1eRZ2lIP9f
lph6/UYyRPTkoZyaxDgKqC2YZq0kIKZKNQvSSE8203zJnbkoaZPwAKT+Agddgr0ez0eD+aKnMfe2
UCp3VYen7dOL3MsURpPBWq2X4zDmQeMWqwcFv+Z3dFZh5tY01X8gO9/53vxfzIqCtuATKWv3NUnA
vKSxUOWSChp83SAcXZ5SiYn69+BjL8yGp9bPN5dHBr7KlmIqXJHcXtIJgroUwjHSr4zgO/cv6ONQ
AUscja9HnBYhnzxS5NqTThKSH2Qmjdzrq2jUVmc2W9JS86JEAqANCuZQzxxfsmlbC3tkB5dgbDXV
jQY+kHPeOGOIeS4Ui1tY/ab7RpPGZLjaB3CN4FQ5+/wE40X31gkxECMQq0SHVGwQJ3KggaEr5QfX
5/yxrs5xGb8rE2VTsF6FNuk2QujZesv1EtuPu5oCYiMxwbgP+7Vp3nv5ykLWc6oxoFnbTJiVdILJ
Xs/+eCGdES8bpi9XXMNS1bxbvtq0HevWjVbnW5OKCLejqSdgmSpP57SVmTdjnQ9OTCke4X01Fzdn
4cTTaIxEVmdgqGLNYR6tIlWoDaE67+cACgZql8shMG0XVp23XBGOwh5bh6RxE+9nbRHqmMBu/Qom
la93s/T6JFkixMcE5ADIfNu3e/QStGmFD7aYh+h5U+WRnzFHLdrBTaGoZCDk08Nwd7h0AyfP16UO
ExEQdmceAA1erJvvJzQ8IuyqtYf6b7UdI3xkGJxE3P9JyV7yNCQtoGThJvJgFhtIdIVK4Ptxp+dD
flrB5tmZsF1BeH/Ioo2Wxi1dpY5pHr6oLt05wyQG6BDynknDplOyP2JCTgRitywuNhpkbcOiaRp1
u81tjhvixmJcDE5FCVgKgRtbLhQcPGNrecWrfYAe3JwjQ9UxmeAcYuBx4b5OswiIl+g+8y7RkNKi
1I0gXavmADfkSUgIDT3FiHr+MTDt70Svcb8cTAuHqlblzQaZzz01yxY1ykKPVMWG2E/7npWKiLm0
o83jivfSZMj4FP2Be77oX6FZo/4un+IDZiWyoQwnMdp26Xt/kulAIuk+J6knHsAuGiZafoc1asLn
FZb/9rHikDIYs3+/tuPi25xGRyUf8zOdVW4C4fF+q1zW1lweUA5Q9tzVlcm/Xskf8fEcXfdXcGnd
HT5IxAXsBZGxiAGtBTdkfyTK7HZYEgGFotMYpPRrcEEfA5Rd4lECc60srql+ITlDIioQPqP0XD9X
PuSXhZ7ridN81GW48Hd3iP51e+z5SgS/g0aOq3UEl3f18XFb1k2D9mwCUreBPH/Iv8CH3/CqZ2m6
aJDRr29E1HSdJEM9OvsFKUkVXKqLEqAetSCTjew3rv3YPR2UnvaZdr+89Cq8HD4WNKwWuKcQNJoM
/WSoijhWP0sIIH2qtPOMjchX2UVM5N50SJbJ5/RGmkn5MWhH8vdXPMYlxY2Kn+ZeKVZNxrLhqsRZ
ybyPiA3aO0s8L1AhA+cPHfquAZNHmZSk9OX7y/nfS6XqSE8VQp7KXAJ1IzJY9jiognayM6tOLyT6
56XUdNPpUFkID5r9QQDCXXuKQbO6xP/7whHtCdFIfiJ2WFr3S2AdlLVPdDGbxzo+HrAEhTvWXg6W
hLBMB/43WB1w5nmAblGiVB/7hzb5XIe/06H2EFzzeVaVb3pTH2Nii+u7N5MzR/NEr/pblduB2A5L
I20dc5sW1x2j7humlFuTPdWIK84iecU+B7+UnhglWqBTzH67uy1zdALNlmYCXnBJENaW8pekX/3I
w2ZHjNj9ELCV7zLJlBN9IfFB8y2IUpXeY6zdCkswzxoS15rv2K5DhiXa7wsd5rZX7GzZ+43l6oT8
gIcv/4Dwsuhqdriz+kwofcFvXakLN+1Y5fjFZPwbZL5Lxjm2Ycj4aGk+iTU0ckHfWqSBm8Yz8vC0
YlPSvEfxaGh3npWiM1aYCGgiWuF/DDHFYRmoPjYVsnwdawfIKGUE2FKOdPn/JjJO4xxfTSsH/mmE
rOeVEaKenriBOAVD0xfl9FF8I8dvqYsiTdl+xmLTTtQ0EeDE3rDIHeh6FQvxuGZ7Xtyo/HoqTu1S
FISFubV5NZM6DH5eE6rUGXtSdU61yKJLkimziDCOswtGVrz83H0GMWgjtfzMoYSpr25F7HWrAXSn
0jM8KKTT3M1CnczR0P3/Hy09lX2qAnaB6HNSgMn+yxEbc2zvCagam6GsXgHAkb4O0csrNEzMz75q
fHeti3sDfE3CXKZ5VJVWGxqTavUUCMdaDrpDiHV/59mfseoI0ZF8F/ZIay9lsnUwGiLMKEe7pNHa
oT1KxJfQvI3A0Kt2BqSLqOMiPUdvZviZkqPJMS4pMQayMLqsWjOyIj6CgK52AcGK69bTF1DuAapN
o4jtmz5IgwP6VRsr91xWPcLDHwMv/Kj1iK31Z1ZrccxtD5/OK8XxBL252tHkSHMoR5dzTZWJ0e2E
/KHSW+852jwX9tcKfvRjH1MmclKtEC+yd2ljLvS9zpL88Gr7UNNGB9Y0vIqQm2r2w3StQNX9u+5P
SBcTd5nBNGKyOpY1smo8VhXER6GmdlnxTarL4Vbq0ucScOLFVtO0Teeun50j6qqZTAePB3KScufE
OpEHCAYBsVKYViKFszuddY14F3LRyk0ofFHic9tk5uKImZmOiUJrdUc9FpVaI9e5FuVlsOfJK8EX
wPbgehgwBEN7saeHg2TH38eu7aUzaxvnTlmawyzQLgwjhzCNbl5XiCCmGBEfJQROX14hqxuxREd9
0aS3p1WFcw/DlNHaeeXkmAjUox835XZHVEYBjjvr+wosFKmGpRS3DGtcd+/2gF5rZ9ObLBfaL8yf
iqq8gUvuIbIuOnPjdLQwgcYyom/+LgTdWEKmlHmSym9NhjN6O6jdlnbUIyerPFhzG673cit91ltt
GQZNNWpT6vV76nwR3QtT5KVuG6GeZqh98tKKJtvOIcLFpDKnZzpSLJQk3+zfEZ3RIMeCdgZio1st
DkKHshdt2DqDlrYWLloEtpfhfZUjFIr3VRkybeIgkdv3Ze+Odb1D9fm1QDIaYKaLK+N1saYdiXk6
Z7CKF87SldCWh2ITLXGVKLy6vLzR8jM3zRp/GpRe1V8tTCqqI0NJWuOz49FJiO/MLz1pZu9ASMU6
/ranjs8eu8Gg95ortNHLXyVgSdx7mGgSdJv+js27LWLUfg3uS4dH0cuMI4pf8UAEUiGc358GLOjR
qXEJYc86LYVeuniLgIN95KpGGAXGWgnefAIqZjTlqwh5n79wYG/HhW5L4q2wjRmHAXCYJGijgsoI
c+f61Na2mcu5/SWXlGT5jDBnryChzMk+vntMM7T7t4rR/Jun3X6Hkd2u7XjJWERJsgG3IQVEDnm5
6ye2fxpHZXMuiubNUrhFGVL1aGlbly4VhOwpbg+apoc8krFBCuqqLqtPQuUjlkmgnwV9HT4OGP3u
mk/K9+GMNcVozDI2BWqFuhuvT4v/i2x6J+KGNUHyg8Oae+lDyAMQ9tWKKarsy7W6M8NtisnVkLhD
4pHPb45v3DzWxhtu4rbtUAKjdodcvNixOGXFgtHLEtacnhJRME+Mt9HzP9fqPkBhxJpRyurjPp+e
3Lasxg4aAbFlsm+iUEZKkdSNA+XGDYcdFuqr56ofIG/MRZ5A+No50eqtny6HPS8zxcYQ0QjRH1/T
H0DT1i70eFc7STdQ2k5LdfDq6LpQI9zo4b0SvnQWBjMk1uO+gyskSP5NJbtfWA3nlt+PaA73G8cg
+sjQUwYjRwArWHfMkW4naNpGewMEkQ6wJNI7w02oFFxmXYSnDuChOQ9UsM59ZjL+bcvENuPZrdNM
4atQeUQmLwzn3BnYpw1fSYoaqhh23MMsk4beebwsIb7Ww10Dd8C9SPXyv7yjkUQxNAMptz/n/xOL
vdd5SxASI1W46F+cXidDkSy1ANDhqhmkU6jf6tL60E6qaLK25RtXmjQ6FHU6+DOJ3C1rDp8KTScM
sqwXu9crTl2pGsnIaRzboL4Utpg4DXDcXEXY5pOHLMgIDepI3leodGzk3bKDqudOEP9mH/1/31Yg
I6EujSZ/xSLEIiYuMIVIjUJmwiGnLw2467+88B2r9bPD0p2PwxX69Y/CksYHoy7ex1yeH3aHmsJH
eErrEjHqhsWmfyUNkCLpXRVQky19UN4x0jbNk0Ks/q3/nC7OQ/deZX+fOH57HaCac9TnPGz7IUz0
OsYmL6y8zpMqg948qn0DfTNevkc13rMx0p3xiyRj0TdexxhdOOCzhb0cznSj4NHVXRK+KJotD7mN
IBOKUWk0qEK/bRS+E9YG6+iIvRx3C6NGA8kwngcQ5D1H0iVrZ8v8iTcss3U/mJTQx7w0XhML5uN/
ZMT9xlFuoNnz2vM1u5u/PZ9oS+49KdE3naxyvjMqXkk6NRJxrcMixJ/y91cBHM9N9AoM6yH+I/Xs
O13gKAiw+WQHuUsd6hQUtk+UmJH7QlIhZ5pVpwBlwQVMkeSTO9Cbd0eutzp+/uyaVpTjXIUJJjOn
vOnahl1GXLbJnYwQbXM3j7aa00TJKe7L078pPVXJEqVGIbCTA0mjLABxnKPQqV9zdCjvW8LouuSw
8/ijbidaDwAZ6JeGJWLOMfgYH2xcG/f8KNR99aCPlTNxEoVxu3iA5ElXVkqamJ4glVHPy+Q5T/a/
FFF8fSCx2V9/RfMkvHPXAap3YXI27CqFOchtQuxLT0hoYUedj+SwTCFfkt/ERwgrr+mb7R408OIE
OgCMPcYneWAJFHcpwlQmul5G0Ekbtq2CXli9qgsV7+lDzlN2FNhIuHKi3mBpUw/jqrWgmexxDUYK
9H/8gbFEPpPZVKItRmqh9wuJ8WQ2qlkljP1wQWpYnqxZsLd+95icyegMA9823+0CUyM9HAP6fM6L
jigKy47DCdLPFB3YfSlsryStdOYpkiO0k1aPrlH98X1HgoLws+KPXVTaa6evepcUndvzH8n3ncHP
LeIQoGCoOmPDucPHjpMMzPqCtOB8xORRbyh8mMEnNxmqzV0wUH9Y1lRHxECKJvTBDUFKmhhdD/P/
pd37oTlPyeOl/KrirGkGS9JrAXgShJhYKKkUxP1Y3lzSfzOYp8o8c6B77BhoYJC3Z2aPfrwSVtPh
Uf/0g102HbXzOvM5yswDoKZqlnU7MnWM04hEdtr4AslXqinVHgfzrj3fZWMvADUZb2m7KU/TQrxi
XyUi0j5mL3b4saWMRFVggTdOV+1Uql0s9Cz06U4nUC09HhiSHJfi91GG5HvKldWZHnreW92tfCQ5
i+UMkHXQtSabldrVzKbY9s6jOjk4apwbPT38uNPWT8Bf2aw70gxYGNsc6H7gA7+sdUw02yMqH3I5
VbHTjj9SASHJ8yiUhYHLergrXML7e63ZHFcXH2jiybJcVA1Werx5bfLvsZYFEsPUIvun3HH3V1RT
QewqCNS2nCgi36QtXPNqjpdZk9/KewW9Y0uLxs0I0ZHscJsG5/RL3Mn8reqZraA4/Kh60fPYLF6F
UPxLv3ugLAQeCaXLgZAzLMSzeO+5dljneRE56o7o8Zi+Zbe9i2IqTT0dXAgbaFBSQjjtAy8GXmA2
jKH0QvsmODiTnhtO9mII2At/IajgdfBL35xtEl9DH0rA6Tfk5XAOv6idrO3GPYfL4os15KKDWryU
IUbv1eWUUJAOwZ7syxUpsFOm/KchAmy98DPe0OjZGX4PRrfiEwQaQhlEKaeBWDXw+Z6x8OAH8HGP
VSNY929f9/0/L14kp+/G5VABw8cLgi+O26zJev+zsVqN4kfEL5j6rb62oMLCRhsgEjlaMtdtxiE+
q/iieaCbCiEKGlM3GTRgCD26SKGP9ahgcUNW69wVmDFDKIGfASitHkiwZnAtR2CQAvTXK4qT1haS
giABWt1dkrFwb/TgAUP1xrXSGJyqiSWeFW09h9BWP8TzeecVNCUh1UqJsJTpHFZBM/u2/lsYohYN
E4MPZ5U/EmTPFYIK2+ReEhE0NqtRtoOizadzmMv0Muw/DdjMCvFNhYUi98WbSEh8uue5TpjpQMEk
hCmvjqajArYHAwPj1lblCggFzbPR7dXwd40K4VjxV3YDPvYrl3HRlDv4QygJRrMOIuGuJ88ZLJ9w
JPzShmFzGavkWgdYFPPJiOFB0FlNXmFbPfz7mwWJbPXD1di4PXeMqZwdSgaIcCyxTXaduKgT8SXV
DgFweZF33TiiPIEpGKWzPsOBfgsly8n2PYj8+ON0nMjhxJYYd16ihMFoZ164uCwhw3oiI3NecG8k
kj3fTsnT5rGOYZ2dfER9ouwL7eZ9M0fgqxGs7oOLwVPeeRZnOpdlWPiXgYi9aFox0J6TdJBkzEev
xdlPIcQD7KH2LZqeNLmhNMpFg4soxAzB32Xu60o0bKv1vv25MISzkSnagOSVTfr4NDYzbwJm33uJ
c7GIrc0pBH5MJr9jrEYejjOa3aUgDE7erH0wH7kYWqiAFjeYyNyH1py9fes74h1UoaZXLiRTZ/tb
gvxAhkP5IyNYxK4vwl7KDhAVPoA4AcpXsqE5HaJKd3U3pQItPWPjY+lJW/HU0TZ2g6vrOwjCVpFs
kV7remNpmlI9vS67wNyPonccHuhsRocd8gzrhIyCCLSDkY4Gts+U/nNM8a7eI4iDAUMHr0eCcEx4
iZTon7rmrp024iLtAvJzo5a4hH0ibWz+szMMrwhF5B+Kz0WW6auj9cVFmWKq2V9doFNnzqMAAdo6
AjElL83iUedsDqzTQIJAgWmIDpu4k3+istuoz0il1+5wnDdrQ2o8KP1x4ytPy1Ws38H6uebDHci3
fxcs21cfqiGpzMwo0HtrBEWnvP/PqOshWIUD+FyyK7Z/4REjBqkSqL/PJ6jO6SMXIq2jdOS5Prll
INpa20ZZYt5n8zR66BLH3nk6EWKRJ255AT9/ieL2vXaPxu+Ih39/xnaEcpjhWRXAU5VpIwdm3R+8
giWsn479oEUCe0sYSAeN8kgB4Q+kzGmILYhx8KeqFTFU+g6jN/pFm5mDzr5w+Lu560yF99xplvyZ
b3lXL7CZuTgvZ9DjD69bxeits75ax0ozhAyujU5IYw9SpSeyUPz8HPZFSzJbkaJ5+OtTyT8lFGKh
W2WVjHCTcvTaIeNqB1QITjHUo5TatDAa1PvvbGIDJBGZRp4Mj/YaegscQwLQpfXvkvVwsR7cVecu
TEY/xLpN7yLZY7VB2ZcK+MIgoPTBjK7CpBCz1S30tW6LDOVqBQbAJyBdTXGJtu5OPFiaS68g327l
z4BkNR84M+zUH3ZctZfJfEfaqm1IRDXHpqNpNEsw74BjsNMBt/DpsTA+lARhfFXIdRioU3UpwHOT
VtQelAmKDq+BqWTBE3/qX9RMRVfM1H/c63MqMFYRGpofLpujJ9flThYh6x1iTcCceF05c2mfyNW6
3V37EVUI4IeTKD1x8jwCK3w7wqS/Ss3CGx81TXK0jEDYQrEarXjb6ApIm76HWBqjA0PRTbDHe/kA
ZtSmdMmHXcI/YhXuP1Sr2Ggkf23lipmcsKryDwFRe16YKhsUZMwQwfdjq/i1aS56EU4XICs30KYi
MManUicX1sBfTYU3HmwAUWo53w+LNtO369SmqRht8SKgrJGx8eAAsLBytilEKhBBh7lZ9Mx28UZg
69HPrBd1rs8faD3iq+0JnW/d+sxyN3XPm3nSNCBGNRJGpV5WvpbS5Y0mEK83Pxt49c58W3xEkihP
HAkrVouaozZqw0MAl/oJGOrRxqU1M8D/50HfjU4ibKPbtMXnAA0m9CeDF960Qev1l6kiMVmIrLKg
KHbvGd+szopPJ2f82Tu87MOmEcarZFq8Rx9lL4XLgnuW0yaN6NFDvgrUulirT9/mudg5T7gswR9q
FPK70wa8tukF8sRNmDwAIg60i5Jz4HcjYd8X1D5wa2hqDCDlJhlQ7AtyhF5DrqxWUbNo07Pb+zgI
+y2PTK3Qr6jSUiOdQmL03BeJ3OAFXfROaDkTNBTXVEfqNVWOoriO2MxtuVtKja3Nh1JCpvDbJRNK
VeSeqR9Luq4kqSjEdHKl7bDbu0HEztwR5zhPmwtfz6gQU3c6N5WxMLJ1Sib3nH4x+fizKy0cf27t
8LfgRDTuYKD7iQ5On+9bwGPclhJfUGTlLHYci4KxHgmqkfZzQfAi0BgcUpX5EXwdNgpzoWMw/l8I
vZRDzD81ogpwZ4UWymT7XKZa2iRZfbXevp0Hk501O/deYArl1Epz7DR7Fpqe68ONV+Q/aOMquau2
hCjBu1lXHm+pJsia8lF/KZ6wtTBGchYfjmaI+W31BJauaC/Cz9nZi199LNk52ipL4rLL7+3vbY7D
Nn2pvWfOS9qoPy5knS4OVvNQsjAufp7h+8TrVAl9BjGzmc/wLNSTfTtkarQBJ3gmjr6lZNlE7i1H
kXordJcWNp/nwZ+L0sak9Xp0s6AdPud7He7k7VvRSn1G4qVAFlRZuTjSdaMcddoyPjf2d4pHDA/+
Gd5CBtlEeYXA8tHslL1c1AMSGf2yxbKSF1sdYWG1ONz9wGB+dwiK5wZB8yqaHrBeNl5d9eaSThax
q6IR3TUPok0TlL9218vWJ67wr1qD3BbtKfheWWS20piDShHLXhwENBnz/qetdqsWFwzZQLC3BQpC
14w6JYKDRiRmohkEt7TZTSjRFIjKRe41r+Efv80my0BOz9OyCkTkNif04W4K7P1tkSJivHAli+Vi
zYBIbvK0UbL1HO2nRnAej5MZllizPgwwrvuVcNcxZCa3uyh7BFO3KKDX2rBIwb8ttBZQZ99rWOxM
Hv10BVTi6tzmEnVEKbnmSQYW24t5OmE98SBVKuJhTZV1ZwfSmZP+O/WlbtkZauEbcF1BFNEviqiK
VRTbG5UynOrFogDs4MhUbLrjWo3afd37NmCnIWZ+OUZmm3W+VZrMOY6T1PRbXi0XGwft4PDp2G+F
VbEUIQVkUjMsZFb0Ibs7DT4NvY4H9tMMzkA//V7ryXv8ItdLRpaiOqpbKsxgvZUWQmKvjJspl9wx
7l7dcV7kX7parU4ib0MlbNWA86IPxdhpUAqOzolsrL5FHsSDj8wrfcwXktOvytWyPb8xyiJ4BO/I
IbhuVlfOdoUiyWLnn9pMT9AOMl8V6V5OiTyd+L0f1ai4XzZFO+4mhY5Woz61uLtyK4CYZoRGlnld
HFfjpYn/WmpU/BcqXZ6oEhGUzTVFlDFvp/QCrgsiNjQea3dYk7n0YK+yPHNwFWDwgY9CiN8a+C8m
3Iw1oN33cP3uBK0f/eR4eITdgMbD2rdDjCYSXpIl/LG/WV0TVHB7EV05/jbeB3IKvWKnuqKiYbHc
rU4CXiQc5ErR4+BOH2gqKjd1o9IVsHzIxxA6HoMZAMxYlNvhEgaAtKtHn1BlA7/F0mnZRH1Ex9Hq
AzBLt/A72pduJD8J5z1cJ9hoK2goIn/P81PT9gAKP1NY9WyXBEcTWgo40SPvDSQ1Yay9KmZQXOFQ
hzzPJ+9xsXYIFvhIDYtvy/9rNtvFg/dggVhpQn0utv2etJe2q06sbKon5Jx3kwDmjBlFBfgEqLiA
VUNqF2ifL7C1ZX6sxflVjVB7CO5TTBkzMuJyNXem0Hfm8neUN2lLuuNcdRFmwjcRz7q/NK3kdqsL
yqniKDWSsCapnhipm8DX7ERfIlJR/A1KMT58iXwgA7r30asIXEyVS+rX8UlQuwLjnRwE6P9kzxzP
Kwzoikmp9LPb8fWePcA40yUrt7LB86+4Pu+5EvWgXsCbBs3sGASkUSXstLoCwf5wJEtALxSkRU85
87/nASMLOP8ARt3vg2FE/kcOL3ZZdrV1KToiHHTaVbs1KUlXQAz9sNivM75OxHTfQci1HyotB3oA
WtqDyVtIvmpkswBg9KJ5rzDjEHWaftacJrvHGkoX30ZDnV9woT+YJI1Qc0TRK4uOG8TBhToLQ4Oa
U408Tq32dFUkn7B0S+xHzxbg1MH2RrpVqemweiodisO0qkRkWtEIzAXWxttKU6A19vkCv1aPj8Ff
5t80W02P7BvHbcgTYnVHQS5M63hIx6RDc41EgOkU20Sbl0DhjXZDnyV9FkjanVvmpdD11JLkY+61
Rat4n6eKSgrpDjX8iRI0bA3zgg/8ETz3qlFEL80wfnXd672A/miZRMNfxEClcuoh8d6xjjGgZwpU
wpcpTxL2nrIh8ciDhLppJErPNIKmcl0w2TTDFSkiGNLNbMZjL3IuuT3DANFqJK6ErTonDPWh3gQ5
iHpPdptNnpRiip9rD1MfsEDHUu1gvZ7U9C9rvfHbjtZN0JXjrg7ffaENWNI8NEnz+RGv4eOv3Rvf
IQdhQql1dV3OqpMn//K5sci58WcaoxJHzQUmDRdsLRUnYbtSGQw1xoViGKMLEhOkob4jB6YTit4D
7nQfpsc5KmlNYYI4cY+Q5Aodn3oHBXGNjIW7mQ08WGU3hZ2ziQZxrOfkcUcgMQ6ZByO5Q1ZsaM/d
WOV7JoOlcm0IUu7w4G9RiXJJ83rQKGDKhkMZW8Hsx0+zehD5sH7Nmg9oZMMTemP1mEz4bLlVu5fO
wZjUQs2EsNKWBSkRdaQA2V/haLoX74mpJ9YdT4aInrgDthQNzNhcM+1gjWtEQoW/nJ7YnwHmoo5f
0ZlhQZsH1Dvplf967Gl+efA2jWK/9yVbmVTnK3GdZ6gT84udn1quTOl6VujdF4YmQV+KuN6od3tM
Nan1DcHQqdq00J0u9QLbCA2bnBUzWbXRfbD0L+AVWQE6g5vpY2rkpNk9BuVdBUXHgmOOkFQjA+HJ
jVodnSRsgGDstR+bUiyU7PqAiLJUYqot/VKER/WV0i6bl34L8aczqkkt4SWsAmAukE2qw9/40EU3
qV6SvHBIHTKuYsgiKy44F1KdXeOyEEJnDmRb/QxOB7fM+4JNWfUkMmUcODT1FQe1p1osjU7HISWu
7t3TfMq2HNX2a/NL0JWwtmOHO0x0up8oVnmSfAQlJVbiZt2qLrCEJIypajzWinx8LAGCZEy11lPA
HiNma90GatRtGwAFJLdh9D2aM661QjWpz8d9DtoThC3J2RkXcpSEKTZmKALFPnDSl++ABoe8LcYO
9zJLoy1jdUh5spaPqQTAAnqSlwaTcpHNY7DaeonpnwDJWZWRDfIgdgsMriWQJaYweu6jw54/lV7N
lrMwsUlPC7uebN/sspI1UHBWSbN/HAq9C4FdiQrJcZRhxfpPEqlNucwL/QyHO0tPyu8Q5Ez19VUM
eNiqX7zbnuYdf2FfjWrsffEcbI3ERgDZndNj5Ya5beEIJ6T+7XQfkWJj+Ts8IGShhxoOTr63R6Rs
QfyRYFXJ7lgDzeG4//svkElZzm66tMxOqe2YQoJF/f5SLU942YYwjivjqDpd0MW5AKZWswrt9/9f
kh4lF1pAKJpY/xzJTE52uTNyvTLpZokMqOvtqJykQ/FpiK3NgyqUdCmqDmzKp3ABl1yKrgqUTL6j
yPzvfXXys7JwWv0uW/hs8/Yn/hv/ddUGc+ObqRH2w3iKTIfwZhww7sWfb7XM2Fy/1KW0qiufUUN4
DwRpfGiR3g1Q8n3gjj9cK2AZ8jwpElAhwe5OS+PkzPtSoxsAui8L5TgjuNhbyRP6sMJnTYPVBclb
KGS7Ko9hoKC8RS7sQVLIoMoOlh5sn81jBEkadVXnqnOhYH8vRw5xy2gDc9S5bdfXbJolMBOXa61m
Qi57eHat8xqR5JFEq5Gd/u+NBPwAM7OJr5T42RpexQbdTAx/afIbdmmwG1SqI/f8RXKNOB0CbCPF
CXe9dG+xFKHIglYW/gFoxa9tAwPZflFWzUGkkKIMb3icOk9L1LuyMN8TVVDOf4r9S3Jlgou/t+D4
X/R5Mf0Q2uN5x8EXIHsI/Z1PCuF1MZPY+YZWqHHIh1k+60gzsBlfR/P3W0yxXOvCF+BDsOAial6h
IS/NQ5SOrinQ1nAOEt8Qrz3mHFqxvDnfVDapWMx7YPbAlSHOZ+lnfKB6+jiJtySd8n/t4H3j4VCA
P+uIzqfhc+1+oCV68yu/NKA3H+z39XrQedBpfK/xGLnEyBq3a+2v+62wTKgc1lzd7B9L9ZZcxgjt
RXLiA9w20PKO13UXlstIL5wzOMbA0MRgfad3561Ie1YHnxtkwx260xXKl8aoxVGgVITNxckVUpOZ
7IrHx72z0XcxqyQtEy37bNZT9FgcIHAzvwuZKVua7k5vl5On4ShONRhMnM7rXgHAVsNdRQih+PpC
cUwHPLBoFlPXdJc9RcZbVY9RZfULhKD6gQ/ueM8A6HEu926uJVOB1vF0XeuJxuB5JuYt+kerFAg4
MRsxL16ft5rmOVRWdCUrTMcvt79abobfyWyv5c6A3KvcBk439u7WtSO/CA6kEoS9W7gxvTIgFppp
UGPEHH/yj0p5TSK1VaJRW8c2OoPe9iiKpsqClxv6P+wr9UlSt6L7O3dBw+lPzAR1Qv7PMTAEmpap
Dl0U4w/3viQDvt3fxPLJc3axgczJo83x/0CVR+UWUAXkgdkXfg1WJwDasfmO65E/3a1VgEnJzHaA
IFg1KXIad1Nx4bSWYCXP/7mk906pN0NRqY39uXez721C9fiTcjywfdausZ15V+1lLFbxdMzOylXr
SxpDbgE+l6i4/2XSMau07Yb36Kw7oC+ubwrLQqwTlYRb7v51b+182Y+14Pa467k7GG3ZvM0tIu+M
fGOejQTi0WKxwx0tMYQ6j4ROlKoCHQVFGH3NxDn1EoJ4N7TQHAW1VZgTIYn3jWEcerRoQfO0gnTZ
WCI4PfjpXxbfA05q/vOJhIH1+AWHWxqhnYQQ3or8bI5oZFB5ctuly2AoUFZ4vaqjAtBRy8Y+LLp9
Wk0hp+16OTd53qHHPQ7/I5lpoevKdqbsO6vjQ5QD8ouECHg80NUV6wFBhXfQT8r+UL4spkanneKV
zgQraSgvLICSMqlh4k3wRQE9xXuQRus6n744kZ3fC1DojE8hlEb5oLAzt7hJJZ8dBArRC/RGb20z
ncQJg4CiEgGmG6tDALqGasHKS8vWDrMgsg7S90zWNiw3WlR3s+keXBdyWlOoxoaL6tvsdesxDhIL
b4QRMCtO8AlbsUEjRKxK9+Kt57Scc3HK5XDDjZLUSeOmW31j2mK/hHOTzRJ4QvOVPh4JaNUCegPx
Cjb7+NnLfRU6F6eRlOuZUtRWVVGS2J2lIefyFjK6zlToIcXx1hDQhkj5whvHCPOo6woQBOOVvE0n
NS7mS1BIrTcVE378zaM09Fi07lj0dBI1sIbI3bNU6x4vir+6DZOeHrrKc26vkp0Dsgup/OhwtLKn
2TJKnWXWZAeeTowgfj58yUHQ4BNzg95oU1UvtOwuZF7OIloVHsVFX8Nr7RvWUxiKXvtK2py1aiWk
VU9IEqLkwTQ0Jy9XFIte2w22+4ef7NBW3By4Y6faCR1BRVJikYQj7weR/vP3synm+tfC/BnmRh2v
rIZnCGGBLydjXCviVa0Bko2qTDmzo3AKogzu0qALbkAwcjxGv8yYIneTKQ5f9dKFmOZaQG3vVKov
delye2IIAlUwAJ4fpMLaIq7/BOIBhDW5La5DLjcraqhemrqx0xZmgIiQso50Q0Q14adc9fFqeoG7
Q6fblQloKuwg11kN3IPIcQyW49HFMGBIR/bXm9HziSYGmkNFB5m70FpX0N8aLLeAxj2LqCdCLElm
rJ+LBuHcydBRw87BzlVtMwA+yXvWTKJK6Q7igmZD0iREG77xjOMxtfZeJD35Mx+quS8iHpOqqN/c
/dD9xAfdaFd6d7e9M4pKFOZv3QOszBpcj+JQ4IVRMWOgq1P2GNbXIgQF3lzvZ+wXmYpIOEMcBHU+
9DRh9LTxKfnGMlx7y+DZIcoE4MZqBhjWK1TsIM++CdFN1KBrEdvy2laG1pap7sdj+sGvohut/snZ
5IFEtW4/VlU0mFRAwrN/MFeuvEHsc1KxpZPXzeBFIwN27u/SE93IyOgpQtpUAV10ufCwPVGIdVYp
cC+HZw/XC8vi3wR3nGPmsg886byCpvx3e/Y1hz2lBwQV6LMjtVciURiViT+QS3PxfgihgLMnhkFD
4k8u6E0/b2s58XZchlsVC3/4R7AgHdeUAhVLqCCuLywY68dcWsTw88CQ8I17h1xFchJwW4wWoBzH
Dzti9DrWJL4uA4LE2xTXGwjP7m4b0tHommjSuvFrZU7mQgO8HTlvbZwhs1CedT9O+eac6GDawUsa
TLX47Mx6O3FcyEmnXRKkRV4I5MOsY7RleCk2T50QVYolOVX2YuQdQggPJOhjgDIZYMh9M0OxlmYF
yubECO+PlaWwo8m+u4qVrcnI7vrPme9BEYwxNh3PGcK6vZRleoQbGpv85tzwflBob1p/6r6pqMYO
VmSbj5hnp1k48iuV1eMjPWTeoa+U2vR7OSUhuOeK5AvHwydCojuGGg3dNwRztQUy/XNYOC/y/58f
m8IQcq1AU6I5wWbwYJALZIACJGhsVLgQYXfTPev457oUlFQccVc5N3wD0d3bsHhGW6S9VLJeBgl2
MMXbFYqvZ/c+zROlL09shaP9ir5OukZw37xrvV/1Rrm/5ZimzUmB5odtrm8mWxJKHeF13OhSmCvU
0eCwcIYDU/8H/yakoJIF3fnrUYRqeCJraI9dViKi7LoiYXHTnOP1C9WfNell9xYLwsvqmsPteGDG
yLPpRXYH0doMxbhD1Vi/aNl/9N9T2/yDvRD3LTUAgtil03Vg0V2BJ/r4vGZFPHWan1oZSnIf3/Lu
yy9MbMUn9lTdIzppnjXQaS98Mbtwyd0ieCYq7xK5hpBe7Pj9+/kL5ABAQ6fJdaFYUStkkaw+kHlU
NyZq/UgnP6PKReWfaOAbajlHFwgX69ahiXOtsqwPO0kvUqaA/qrQH2Qw31mSAR7p+4hRAFPx2XdQ
VBrmcTrX1W2fxfmMMoV1BrVBkXIuSE3ZjSVKQlnN2Gn68o6WB1ycINx4KI+2HSJd2iaE+LAbprjx
RGUbzmdZljZo0N/LRno7HAC0N3Ga61dFr8udN5W2QoOp/ZpNyQxwYFB9wxIkrJsDah5Nr5Gx7roV
NWn8uGwcN3z8DTTE2aOU+6eZzUxUn74s1ck5Jw0XoyXqq7IGWTccL2UiJ88oDXRp9ObuPYMR2obJ
CWG0KqxXFY7Hwt4Ofny1PGW1FC62diM8qgekNhg2Zjk8yvWderZ7a5HFvl5cfipLgMowcftK7GNW
KkTa26eQBDlp/ADiN5TyD0euq+LNM5fNyVCSN5Qjkdp4dHfmeAs3pWJmE6OOtdGvjqrTY/PcnIdY
/HoendwITB29wzvO5zF2WXix3hs8v3Lx8HTNPt3AfVdTj+MCgzbf1PCYuBvoddqaTCNyzkhBu5Xo
UA/tHHryiyT6xBZ0u1fCNMEztH9/xU2DpC5rDD4+sJIjUsykhtzVtCFxKn8Yc6PS+boZANvgp/E7
DbqEVcGZLXEWFlw6hTkY6dFvz0OmmMXhYx1kL1fwMzXaFINPhTJHx5MAOFmIAW15NSCD//PkSCeW
2lIQWnQ9MA6wIOiCcIa2Y8mmRDIzvWjeW0VsIK/AhyqlseCCnho8ru3x8sENvHlmLXjbbREuMpKt
y+V0BpAR4er1DX/uHbrsNO8BAmNq2fXP/5QDmebLcl+lsr7sRK0CLJRjerSjFUTZdWPTtb6SI2ZB
vz/E6xCsN0IvG93csbsgp7e07sfok2FiEbhqXToVvpd8WYrj2bX0JTQ4uWUn8mp0lte6rHWgKXXK
LvpzaJL7gEIhJU74B4+MrfK8Cznst70hwyqY9Bcb8abq96WDwKVVburFFhC1Zz8JDH03nbw7TMF1
KcC3i8oeoZj581S+O6UiJB8BX1kxuPmVm+QaKBb8iUum9AcH3WxxiZSGWH0vKpBXPv9evyeaabuG
A4eIZezWEBWIFN7rhr1lvwT8W/ePC9NrzEyuqx9RYTQ7KS1kjdJY5HtoY2NI5Il46+lt6AUK7frh
bZDGwqITM1oSFkvW8NbdkgMoNZGgiXq1kNIfXfAbBiJQoRDbN6NGu6OzMvBXRVW1JcKAZGlNQVsi
oU/WAQ4k9EYQs64FXqvEeY9T9cdWbIIXfwAPS/jzgKqqQtdP6AXFlO90aub7Y9v4/4ArXYhG3VpE
ZYiTiA2yd5iucbM/fzkD/7PVWNkFw3VIXsKP5unBalTzYef6IIvHAE6BDnJOgvOavdxtrVZ5XvmP
wauzuLn2vZqD5yZy3bxRBGUXtEFHJQoVHLCj3Ugo/ftFJ4KqQ9MSdF5Hetx6oMUVGeDJw6z4jtZH
wqOsNfLxKUhbI82oUVfJIz/b35unABf58LzpWkQYBNS+vmVly9XZzZwrUInILz1gVd/0kGsOwBu3
qA7+rLtRqKGAlhO5YV/7Week5ESWhoedG/pCGs4oRCXJuhAVXyf2QKDJW/Ss4OiWqSQbfW/7DH4P
zx7iK3eir5cswbj7qAiiAcelKStkNzqXEcembNdG/iUFRz2wBYxDfHJ/pCt57jk2cwtg0i0QHs0t
Fr/bzXqLHb5iCtDLudDqpi4tYYPDMeJjAf2MkYFQl+9AUOKiuogKC6c10swdlOq9TiVIo9ZbLhGl
oEE+qnQTlQOXLtRcN+8XGbNYNLYgCGratsoqXloEep56eLVbzYDD6BWHZbczdGCiewTToQmTAOBz
/jWTyYN7QkP7X+KBQtWWicPhXimeSgvRGGjtj/FFr/QgrDG3pdHDTHJxIMW4BmqKup6neWraq8/8
9gzgNPTKV3Q8fV83cSZKNPBEbNK4dasu7tCwzALII2PqUPoG82Dz4cDx6RExTvJ72BFfoTfNmp+k
T6e5DO6CUEpltlLMJwqWetA6TPRNdKKLLLa8Qgw+iGlacAB62Lbbers0AGkeZ6K4ZCtR0KfKTNg4
k5fqFgXotbQs1NX/3TeM75rxQIAIFT7wJROkN5pF59xvQHlJ/X5RrD+eXW0x6QIIsL84MXp2poxq
/BfV9uFuHLHtQP5QwR5Ku/Nxf35aA2ckDO40r00HSJZAiJdLE6mPQV0na7n1u7nBQoGVZa3NqQPZ
Yy0Itukn5tg9M5NOZ/3S2FrlnnHc4Ebmar5+2aiqSFlVIV5JjIrOKP15cCF/1Dkab2sfvhrYE+rJ
hi7q+FJ2yoCzVV0TbkrzYvOpWkie5Sbk2Vlaoh9c5kyTA8uIOAtmXkZfLDkbvMccsPONJh2wE3k5
1Ri73Lp9gqQgTWJL2SBzB1h+Mu+N0YXIX1dcDKyeumiBAHYJ3J0ENyk7LLHqd95NJILruYmTZzan
4OJniTKJsvqmPuEqK1VTDRebrl1a4GNJ2F55ZmSOgOuyfjuqyrkfyqwtm9YJYyVXzY2YdQ7xN7Lc
OpJQ8Ixg8Y0VL82RXvc9HPOips8Dia3kvs2xrg8W1WdZ0EBKIRTHag5KZ9yUlYJiEM9Dme34x46l
nNQll4lI2lZO64VP0pSnOliy+kUh1XkPwRrismVULOGQH8X6gzwmpmdi+AS257dK9dIiJ8SKCbS2
bCQodWkj4jnEh14vT3bOuhXIV/gGEV3Mq89/oXxbHV1pXtLqkMsDRDk+wpOcElq/rw4r5FkUHThl
CsAVNAWfX81KPcEqgW73LreGK10ReysBD6H29c31SXncRfwRhwm1+stGifs4NPMYGoJSG6msBTvk
T3YeBwpinHkaKiKeIxJOTT7UTXBDvZOMANXTW45s15fCOH8M6xTecGauwnlIMv+TxtgY4l2g0Qi7
26jPjDWsEgnGG0iNfpIv3jdQ6PoqMFHhfitNPJELQRWu/7SgDucWpqrVzwpLufbeA45xUNN3Mvpz
6g9k/ffaJxM3UUZ4+dQ9EL093xIax5CxKvSNhdaoij1fVHeUNuZYb7ljqEfaVerea/dJgp+HKyod
7/6VypmBHFOnCXFD6smFV07TARJvxh/xJpmd8ttEFJTcKA6eMmIwOkSGZxs0S1b+6yj0+0/0cf8b
prMFX2c13Y0E1RgjO5uIXKWtYcj88P38gSwVzOjdzZpwp5yl3DMa1HCAQiBpIQ+GsyEENY1DKOD4
4j3rCccPscZBoCwBPL2IujyfEG79A8vS+e73szNvj8c+RedFMGAsuiz/qrDeMr/FeNB3Bg8p9X1C
VswZCkv8cHfJxZ9JxsbvLMijMM6ioNbWAOFzvjVzuBkeLQSwpOi036VPO8mj1GmEfQ2JETzwArVL
sd1p+jrQIsIm7w/QWzcvglQ/3w3hSDJAXsxDlyI23rcxHY909jIzfEGe0rv3K05JbV8zNE8CTBxQ
+9z3twcBy/Z8sT2zAAGpChNtopIn5Ydh659K73/Yy5xQtGgqFNGSNtUrFQKQ0FBgK3GV+u4gP5u0
vbtRAgaEjRYV1rtszf/oiTLMpkbhQwXHlbuV19hzhHzYVf2R5Ff/POnQ5S+aMhOFbT222HieYMfn
tQm5YRiXn1Y5JnV5Pqy06S6bqq+orPK6uxAGjoRgYMdSIRyORkbR7O85GMXbttV9SaiX9UvyTTbP
uRuOMANDiJw/VzToMhu7Qby9eqJHtLxBQEAsR7u3UEtzUma0ydMnbDb4/rfT0TFUXWagcxTqzK54
oGb+VM34dV/PhxT20Dzk9aA2qrVMPoTAgeIKSbqIAjNG/lVJyFJyJA+8r+Wxvcv3ilcw+0UVhXEh
APMWuAeTNf+QX7VSfWEPfba+INPD3yiUbWat07MEMloDI7NuGsd0ePewz1TpKej6comUWTax0P/M
5+kOM680T/gO0dHdH0qxjja4L04VDqzHR3xiE+4FlBuudl2xcebE1aCebmbwYPpCJtgnqobUzvxU
Q+1wFGrj7ldhUnkhCqbMr2gV7Hqq14HJ4ihO5OjHqG/mDeeAj2ywKYdllVtQvj2r9Du+Yhar/021
ui1Akj/wx2IKU6dwTOgsZYnoV4tP8MjQ9GIVoyK3tVgfOEbifUy/9khdTOa7nJf8iWipwQg0ZlJ3
QM3iY+LJl8Q+Iaq+cJbICYU5F3msx/G2szvAOKtsMbgLoI168ee3ldvCeY+oBnxMIeOxzGpeymJA
PWjgaZkv6Itek1ui2J9v0S153W3A5WhfeHEMF2Q7H15ZQsoDFOgxb3ix950g2rsKvDwoP7tKZVzx
jusudywUDrPLmZoNXCiLzSfUlCPMt+Bm4aXHJJY505ncxBtMTmt1JTSWI15cox0VZyyc03IIv5D2
1K5v0/PjZ5z+PJa2Ydq9jIc4ytRXORSDCn6gkIDGRLbNrlHvLKjFYg5DmulC6TFr2UFIMkpGfE4b
zv48EYMLJwkTan1VQu8cFM5FMIfjCMwy7FGInYuEFsqB0h0DdN2JtBXTFKhB/DMKVbGyeRMmFjp1
qkX+F9S/PIoyMQwVO9poQOXdPWCzVzapvw5oeIT/O8rXXdjzMH5l62hzUU4lixh1ppjDiR/SYcmT
h56kh1c7Ct2p0vfTgyuzP1KbCKjjMxZ+KbXNqh8cdOWRKjQ6uexAklAk2v4hNGUe0sCCmsjXfeII
F/iKtkAHLNzNAi3Ihf2a3LBFi+mTqmGg2CbDh6RZRb/lL3duIwaYDmEtsPrZkHY4dkX9+cdjBDs6
lCcnhQBFh+Jks4dSykrHityu271JU7/XT9hh7hbJi3cJHwb7OXxJuq8If/qUy13/SwiTta6EUVeX
23fNAk+6E3UTC6jm+l4PZT70rGLtjEbJOzAQA2GPa8u9PRyJNSUV8ckabs2c4KML6SR7pYwOQfJi
2KSW/uT0TZXBsr4yxuQxNTmjvrPSZs2wyS72L7IPbfe2iyqzJW98zGTfNcWN6mdJnZdVnLtv4Ban
nuA1RK7gGlw4IBbcPqvfQT697vMKYN1dxn5gwK/rwcd2XX/R0WYznNDLmTEZr+CkxHNw1OQhLBl6
rOllZlFsgUGtyZ7J+GGO9ww5m8AQMym+BWO5yNITIW18ho8ayoNZclT6nw5cnOImajkHWTiYJeFV
o+grUcra4Itfek9I+g31Hn88djTNTRA9hp6WUgw5GvW2d17CGazi/8DTHgoksyuODXXDzTyCRNqp
0DidFyYa2uq8btWWx8tIa9AIk7kc9H9kSRG6VPg6PAr78XOu+uEmZ3CX64Vh7ksoeyyoe2wAxEY2
TeLZEeWUABPF4M/AizPR3vA+GVhuANT2tH77NbM4ZHA4uM1z0G+ZFSiCfbyFmeX9yprrPDBOYHrH
/NJV2TSCwXFBTfQJ4EhfHIKbbb1ZbWeMYeSOdUnu/1E7H8o/rMOchh6oVh4eDsGL+6ye/VkJ5/cr
C3Z2GJb2fiVn8cMGttgPtaAzy7b78xQRz+IZWig25Vo4vDdZpkaXDDZGmuM1Dns6cPEYyab38Nsk
hWAcmAxijECyujFJyvjQJ67QLiMTnaEypn5U4b2WKP7OjMi7fCBWRcasDm+0fUuewU/KawT6/5SF
3t/H4FqRIIw5njAF5mbKaEXz12BVMdjiB0s4tfEU4oL/D+8X4QUv76qVJwIsnUpidZOBEje8+bpH
m6+OstSu42WXoQ2jp5Ks0UpT6USqAADhaVkfNVBz3aMSb0Wfj2vAYvWHxpuBx/GTnT+/NfMCoS1M
MEwqk6tBluq7o8z1NCMyjfwtIToGoW8xhhjqwhrmSPAX/fuuEzxQHiRazmvr1Pcxze58EmjFLzRS
27yok2/zwOMKAR/AZpvjWTyPlEP8JvzzWM8DwynnL/Cx7MlFZtmAtrIaeuvb0kCm4rA0eblpRyuj
TMz9kCIuRZoGbJNhjo7Kyqp5bc32eiCKmeFhUcxaY8MDTYJAo5W3aPxOsUM8r8MW9uL3Ckk2KEkz
GW/+qyabPBhqrqBw6aMsAdSYV8XsO6lsHlrD7WztMBJWzcCJcCxgOumj/vNNbdTccfuRvlR4jkS7
TvYr9qhHYFLqDSlfarIgP4kwwuempRQnKyNqBfkYdO72UKXCN+4cFDs3UTDO6FJUVK4UwsehD4nB
mpbZQFrolHs78V1dtzMRVnfjMhL4O5olWOBH9J1QnOrXzW83BwHho2RkJLHksT9G8B0hQqmXpjH4
WtfSucfpDnGrYis6Sgjgvs0vfmu+fynvojHqZ7iwFD6bClfCnWuXDNLlt5At8wZS52ZUl4FvKQ9Y
ydRMnMauPMJFafoTWnVZRUdA13PUYjJis+9Wo/8ITtM8hSu/xpXXHb4jsfGXFhMzLh+KuB0LlUbN
lDQjbHu/b53pVH2HvcIAiMoskcUHLrQJCllSugm6QK4bUK463uU1IddL1T0eEe6mMsDWbLwc+qwL
sKzBd26nzqC2tSmmfHWn3zydX4X1rYX8U2bDLslJ09tVHQ0fZJONEpe7+hxpneSfA8iFxJXWN+sz
2Uih6tPLOwRPD1XoIDIS+Sj++2meq0bSK0xO7R1he3c/LrYcz8xYwWEoMKvB3ApB+rgGFEUq8GF3
KSXWS/itHo3sXkjSAnpmRa5fFXaF9Ax3GMBMagPXdMbNu1NrgNqXB0jq6tVcciycUbdxoCI88Kjq
xZT0dsj2qTX2j5HZkgTCE5UWl1OjSyg0iwGCRIQif5lh5T4eGaS8lw7pCOBm1Aix2Af5ytIYLr0U
Epmm1aGTJZHeaJpRZZcBWcKmOuDeHNTetVTqI+SKABGB9GNGmO3R77NCGu9MNlxA4qabvAnNhiZC
fK4lwRZXU3pQKan1U68MHAtNp0i/gdswZzpv40xLVqAagJeo3zqErCLX/p9mZxDMfWC8Y4zrstNT
07bBbQnGyGUkq8ffFvDI1NTzZMJQeJGqtOp5wAE2Yj0vtNedghmgV9lSIDzo9keAtbk3ceWnKxLk
vlSRdfoIAh0Fgkh8xvvjPeXD/JeRo275D5ASCAALwZslrHhyaKeWlfO6y7+XLffOyjQOrILIoAPH
4ilmsQqP60Jn86N78qp+O21BdjHrc8Ias22qbv08kCitnsEpiz0VeKQQu6t4iF6mucD8ztjMk8ip
qUAQ7KkPLwkOyuZHY/4QtxyMP1xiszoAHa98A2WgKmK+/KlwRSGaV2od3AAWaVBE/0JraMwR+bHh
3oP1Fd+SfY+qC9pbxlgyzzzdhABc7wRnfn78ZdISNwxZMc+Q52yDT4R01X5ZHhGcExXlEvsr8ihM
PzdyhUVjWjzvo8oIIfovXu7RFkzBJEggyRh6XvLRST5xpnJjrIKel2Cw8akARGJiqrYY3zruVB8M
8ICXgCh8eR0t4BvnVFj5TAluUNUr7KnmrUjCKZzqfToJkdiFNy29cWAYwWYohDgSE5PVnGJDm3F7
FmaDlvFTL6KC8sH2bV271wLMKIj99ThjJx8Sy5nRSUTSmcuSatJ1ayJURD5adOJVvVCC+mPuBMOJ
CqAOvfpzXb6Twbi9A90lcy/gJ0KsThSi1rVzblJKGy9vpbitWZOQrdorlPz9V0IYvliXsoJnVlVa
avg52MsqBAIlvidGA8SOnlxGiqbzCnpshkTKBI1T1Wr2vVad1xZwMY6jb79kp0Kt7QpFJ6ilUmIl
E8Fbvkfsdy+8JIov+C6dYv777yEfqZ7UapL5m0a+A4Ns0xfDNxMxgUcVRMYKMCaex+WKx1fG7Uf0
BG+CyDfAHRpjC3gQ+W4gRK63/WKHYqCNtBzmvU4gSH8uJI5nBZ1SSIZ/M2Tpx3Kk6W6oQbesyo2f
Zh6OWP1mgt6khDK3TIFjpBndZQKSnz2yExhh/phX7YQ1mv+TBXORyuHL/9FqO4UYXanEPScJr34W
2SYzf4gRZll71vAtHnS7u2iCb/+a7zfI6oBYPVysy+dRR8SjoB3LrIuycEHjkV54Jpnm/S8npE6W
kF+u80rGHR6Z1L8WyPWrBFUkA9naFnCJgjhv7HqN4h7zNiuHt6oi96DfddWBN0o0DwknvRXeoChg
m5phxkBNdLKGF+TkHw6ACfEHK6AATANIkypiHwrDRy9uPT6B2Yj/mxv4EHEqaiHQmJAmXhpNL5hl
B76qQu8q2c9uCrTzacaDyDG8Ib9KcegZkLNepgwpPJBGYiFKYflQPDgEC4G4dcFpsvT13sUCRnPq
pO3RjCrzs76bq1W4hl8Fxc7HsSP22k7pPBFSD66PMCvDzA5fOZHOns8U4HOJbOcahNCBT55hgiTM
9GNFLlrRTEFEsg/YJG0nnppq8VkzUHqaUrj4T5f6mFa1jqMdin9NO+XahGeOaspnulDBYjNBhexa
C6ZIIfYtYd2D1dluT4o87zCu+7YmX9A+7yZevPTPpDwbARrT0n8MRNto1en0BhsTSrPAtPjKNNY6
5CPRj2zmkOBgBHUx4WYzvjRFD/YeBB0JSYuPruZfVQP/KZdq1GFImpxmd8yM/99I2h/1gpQTZneV
3QuOJzafGVHld4ThZ8j2GP/lX+Z/gOO6muZ/d3D76fHbfOIjM1iLZUV4fnuQ4hStyCdqjxQ7sI0r
t7FsGdGifMZaoBSoThQ3dG48sJ6OCHS6Pd1jOoFyIsjKIhnEODBLxEE8ZyiL/fF50pQEzJGPJ9eo
Ly3Me9Xg6vKOxecu1ntoB10PU0txt5GEcEA39h+ZsMKunOT9eF2K97qDY/1px1+W1Phx9Jv3d783
giX0rM2g9CmxPffdbg3O+hG+gumzsHbL0jfCKavUsa7I7JC9WwzrTCLuUZ3CyB03M67FDovW3N1Y
n+p60KDEPt4gHrDAueXAtN4WBTNyBBn3bmu7/lOOavaNy0RoTsM7Nfup2QNo5Z3bQYDe7ZXvPelO
rUOoqcZwvbP/ItFo18U81zugjNmgdFQzZ7U60rz60dv7y5OZu3NeTKHBy2V2qdjVwkHcQNQ1MqXS
CiT572K+kiedPCpjM/0ksRkiYHE2AKaiDWudjsjRLU5x8IfKH9wU5UsqofaAvqXdjkm4dxg1yY2q
ncUMeYUOPXaZiYYuCLMNrCuPlep9Vn5vGCz3kdoAt/Bde9OSTS7ufSOVcGltTpHIDgZZQgcTDqlJ
ARuqRbJ6gAblOTXOj/xUUXhblADZvxjbPWoN29ghIL35DM22KrpWebQJc6GHPXE/Mb8vul47Kq54
4+BOegR7ZmwaoobUv/2BUsErl0VOuhKaK4EkW3JQi4XhHNO0N2Q7tjyCzR0tPrWXZ7MSgCLkS4QR
nTJBkZqVSiCnQww32nBSYwhALgfNzZ5/G/LEw+b1rSh0S/3y2jm4oskTSYN5g+sEa0Ez/3k1S6Rc
jBWZlQHVtfyP0naNLXB+t6ZlfeoPxBbWyDyMilKKrnXftYa8+9NXChISv6NkYVpxtSutEUzcReuv
FAUQ5aTBhf4vBIAE8tH+gxnINzy10hnsDoPvXHBHsfyFOSYj+zanvHTBm0OgRBlV95ZbjTGBfFSO
S8rTvOlKsyoM23qrlmG9THb4mH0eYDJSGbNQQb0AHpzcoZS3eLaR11RyvQ3fETxXGtRxIVyhRi1M
iQLLP7q7MyO3DldcT+t0l6sT5LQW1+zV9lNdMImgFAyD/er2yCngt12CN0WpNEV9pHKeUsGcs5oR
YJScXBzcm36duSSSH7InCpy6+fK7TaXufaaqJmKc96TfOKFUxuPp0Y2GPbfhG4K9qeywesnMYWy8
vhwo3PjJEQVXF7qlkda74l3WWAtVc+5oPH+ntTh80HzyLSP64yv2i9TYI2fe8yPMpkhzwZpkocPZ
8C3fqBeNLTgv+PJmegbQShbWsWCe5of2W/SCo1IGEOZ7AhHQjg/xjq+6QbRpEhAdPkOeb3Zs04t0
Hh3MW9Iiw9sLbLGVn4QXRZXyTU9X7R7uowyX9q9iMv/9YTY26FV0K9ll2zPN0GkcasBTI+1G4p+B
aVCZPABiJrRlFgioqwiWD72bYLP0LgRrAnkpyUCgWEaa6VhS5XjDpGUAOpzd7xATzM7fAcaH8zRA
2XKuF9S0SYAH8pL/yCpJj2qN2HenCIJd3gA5VWoT495zaqJfAj6mZWbd/gn+o4Ov6Y7VDCeGf11N
Q3pwkslxMKBiQ0x8QKxpLAmV49WZR7aD7ip+m8WyAHjGkcqJ/GtbbDPsuAAa5UelcMuxT2nnLsa9
4FuqPXzDjkjyg58/jIbrBYN7hc4rISi7NkDugSvXAYa7b3aSLfKdLh7UxpLZ9eccE/EJeK+g0KwH
Ji9mhVmdZn2d20VcsSwj26EeC6bssQ324+QqwRsF6rhEsSKxNHXzkXQGLWrTZbYrIVVICCdNUqcI
5v4OxK/57bwF1jl+ZREZKCx7tV5O/GLA01vm989VxRyZNUUOEmy2LeOLNGzppJB4ZfCQsKLt1Trq
hD4lKXNflIbKtkM2RqKdQOZXBfeLAxD40bv8PCypIfgbVCMcn8MG3Doct8Z6ncELwm9SyKNUAsmo
DCyZ0gP2AtZZnJ+U5DKd1y+nrcofIlJQQn2LbYBvnpnZA8VZguaPYXcUTjfA0zUuixbFZj5EdviY
00LKnSKjQYVy07HxmpLHUBn1lPGdV9xipJDMFa+fPheW9lavA1sWzVhfjQnVvFJQaTIvyYGtsCD3
ShsHL5aMxtbsEpUh+mBs0iXK5ZtFfqXgScSWOTZ07yi5+ie78ondP8Czj3AePmQnPFyZV5P7TEon
KgPqP7shuj64aQ6VRze4Lp0Z9azEhqAUq3z3DLiQLLAv+wgtVTHqEzMEk3Az1m9DagzlFtgLw47s
ofDPGk9MgG/G0rRSV0n+QXBp4yTkvpiseP3V1sJJ11rf4qg7t1PXJoLE67gGC+Fu9Ap0UhnHBzWZ
hHUtsN7KdIDZnNOOo97B6ZArsfxMGvbimCTBWSk2E+yooq1heUWMZD1NXeQKYoNKFYfP5z/F2WA/
tN51yaUHU1mg3CaxomHZMPAEDqC56LLIFQDP4fl5pZy4ZRQ8iQeSQEUY+NbYkuWU1zcDNonKZSYO
KJtMgIZOk9DW3iKXK5L65gBZNWqZlPc7F2ZoaV5aOzUt7r3hT7QJV5iC+cXLUZKs+zZ0yIMqT6pk
YAEwPfpN4XxVQLZQvXdmt018OaLBPcXYCym/1Vp44PszIm1CtMHuQ78QE31cc6lUW9pS6EDaPu4P
p3snjM/4pLfJ+2DYPlZmcNLevSjAUNwN+nt0H8Z8cOVZLVPQlzXrlxVPrUW+LDTAcX0wgza3/wrV
cYA+sxkVW3VlDHMZDQhsvuPH/XwZQ+HJUi7NFVZ5Es7Th2PbLlTHG7qr/MKgPexRyjWjqx6nTmMy
7zllSaSHZuVfPPxvMzAceX31g82nZlBPubyqm4XY7IrAv96Ym80ZrHbUKQFr8ctC6hNrR4kS9Vj/
EHSlvlZdOM+isyj7j+IOmRlKdKwB9NbocbvjfqSx3LQqkky51O+bWixZLUJenXfo9ytZXLDVcj7g
d7eYxkaF13NOBXVuk60zkMKSCcDAg1FBq7jyktvIPtyumdWpHQQ3pa7YlxaenW5NmsXjS9aPIhO7
QP3HCmkG71btMBefUsqlNwbl2T0IAFZiPXnbVgaJImUgWJ3hnV+n1yVTB+JRIOKli7ZHF9zu+xri
23jFuaZsyekvVRaS2vLBoXxCZiIC9259diKQk/gqOXkPmVHaO/k33pdRe1UT1TTZKWnGqD949Jcb
74ekuDxvqh1IZ4dThUIPFmAt6jkXbW/iJ2pr/YGiZ5ksCGOS4ERaGY7pzNje+thLq9Ppr3H4svK4
qfFpqzG0Ro4QmaIlJdWeudG1W8HH/QJMqVMrT8LZiGZPmRlyZqGo5/uWvo10gLKZf7gCXOTjZun7
d/RVN8wcKcVTuK2u/bPcIeUAgowhAVp7DWVV1g49z0KCZ/M1k1gks7qSEa0NJjytqKcAuRYoOfTU
kSuQldhxDZwPHiyx8orWgs1+M0+HUSKsg2MHOubWIKHM5wZDmTiFdkLfXS//9vOLnb2vcH/QsDNE
RYAkIq/dWEx0VLjcg51DvWC3DbZaqusrdEVvIm2ut0mHxdPNNOI8FtKRgn5TfW++q9fZuJpefylZ
kb8gw9wN57O/ECFY4pjvJiGx5XjC5C3g2pXpfjMEXpKwlKfHT0RPcFnuWoUAxL0Xbhvh5cUWluO5
Rap6O+CAQutJS7srNxo1DIicHCLFLI4xRi+qBIKn/ss5T2K0R46As/84INLzJGvW+OQMmpEjMBrA
/8z9vGo6uSsRREgGU6EcmsbLQZqA1yawQS+Efz6ss/Qm2vs6SWoCx/Fovx6tF1a3ik6VF0Bopg5O
RQF+SSRyXJ9S+//sE/t572wLICm/tVi4pnyj/MwOd35fzIQpY2PvnluKtricloFd3LD5pztGjyaM
suKBnaiyxol5Y7e4tg9yAKSRuXdUc+74B3Flk3wExkk5zezkp9TVBllktYST66cuTPa5I34bSX9l
HbKfk+5m7+S9TCeOJBNn9Tv7Id31289cJsVABpniCIz4jYneqRtC6nmTC02LMe9+B46+I6lw+3kY
mOzcC8xNmFxWqcNgaVKEFPCLVzvHgXsrL8HieuOUjek00e333qZR3MhKHv0LpAWIQ9XzvrQlesBl
ZKJh7tF4oyNnGDNivZvgSYXR7bHUDqvQzbniYz08zTUF4Bhy2b1GeW20P8GFSyVftGDL6SSgIqik
UVO32WAKFvAW6P9xTsotHSFQ+TSQjap6GyYFIrz+qcusXWS4o+FluigqWu1cjNoh+6rwh1lwz+Xu
jrULh60dSadwZ9sZpJ0BP0aFzpr43rqq8npyo8cO0wdbETKacT65Rz/Q82aroy5jDl+XRwJzar0w
wLgyqIZS/MMY33+366UbMT0W/79QGIwBbzjIqxLiTBirDYiglRkslSlRBfKpwl8QLK4EQgu7c2FV
Vv0+5/U+X8ItGXpMCR8EbzwNYh8E9VR+jZU560S5ndwce9h37owXlxLSO14V2dD+VwCUceSxB2u4
unrI7PXyTNHwOw7ARNM4bxKvaGM8UfP5lhqmQed85W6sSH/5g+XfddibFHSuwOzEicapJFS3XHz5
79JAhJ1KZM6SYAZq+zL771qi+GDHHAebwvfa7rez5J8ColWAbxSYQ9bJK9Y9LKYSODJVfjSe8X9D
+9MSVYGB0xIDkt0QuGbQx3mUNNqZyGupeWHf+5YeWu3OxkbZwnLiR047uK6SwiJbCvSSYkJCt3AI
+zkjJmBsMPiPm2zJVRfvQw9UpeaTWb3Bhz6Y3vG1GEjsME6fRpPS2OHSZW5hfvRG7J5AU4rc6VFA
wlf7coztojHq2ofcfc+SmWrRZwcxZ4dg+ODKLSTyrbCmKh6HfibhTIdJ2u4QQ7g7AYrgqB+PxOkF
57bFYfW24qvZs+jVjmND1qxlESq47Pyn2AmE/uGLvnDdn43G5+ZHe+WrQ+tRAKTWp3Vqa30djDSr
qPD3M9mMMkzi5hthVNnML5ZuKyL/WjHZHpfnNnHksmQbbYXSHeFMxAqcj8uesQ9xEdUTofLWDiIY
qJjbXDPrmD8m3FhaKGD1Zjw93ts7W86kxrdMNDCSsd0n8bNi5v4HViW3tWJTJAtHmn8sHPGLR05I
q4DKNEmngM2V8Y+BpHc4onzkupYTvTWncCJ9S18uIwcfjoNk7yWXk5x29BsNn0Dg4xWUVvUvlEUN
oJPstLmVsgUW7KzJdOP/XuCJziSd9n/AjpE96W48nCIqEL3t8W4axQhzXq5KpEdyP/y9aXnBV5CQ
GBGWGxbMFB5FEcMpoKhSWhFE3frSMhtscRbbVdO1bJ9kMKcerPhynm/nFY5b44WhHuJCH1MTBo37
nbN0/w2JpIrtNOf4Clf9ShWf7duXduW9NQv03wYS03py1gzsyeUegRcIl9HAJmcJCL9aT76/E1vc
dVPEUHJKDu0x7e++lzUaQXd6GsLe+H8aCs92i4z8tBdTgg8JDEC+gNY6rHNsLHHSviA5q4P9y7IK
oiMSuPoMGheCMv9h6wz8PQk01xwSzhD9sExbRcXGmt4MsYnmLEITj9e8i4tUI6dkglOIB9Cy056K
VB3tDCRG6GAPz8MTxSjT4o/+g3S40fAapwbLwheJa7M+pm2qFc+X+rGPE03Fba0wZWS4vgzQFwQk
YEQnNCFbdI0Bm4F4M9ADJMW5ncLoapg4toqMY3PDuui86eUtCN2glG1BsBISPV8a7DeGrSsZG/av
b1ZUoJIOplnyEku+OFM7DpnYUhrajn0xO4uTjsfQTlxMP0Xia8BO7wgSrO/SjRYiM/aQbOcpsuzd
ZZjGSRYSWkMkowOhizJ6FexJWroezqlPzaorNj/Wt59S92lBm/WIERTz0gJfpGzP/kTVYgnzbFuC
zA1pHHSC8tiSi+IWtgM7o/dsel2DKVDTHIppyCG4DcqoIVDDQYtKaeFHvz3qYm79efvUGAmIl8dU
MQjaI5GYhJHP0U5nZEQzNi1DkfsDofZ8fJXwiHmPax2aABJHHBpKW0syahqWHdTiUTVff4tBrrqL
LejPf8jIZ0NW+WjdzNpbphjjBNdhQpEMbuNShV2gijJPOZRswwpzgbsjU37XqwnVvnAzYfPZa2OO
dPSqAgSsVYh99Xclz4wbz/CgoFrjZ6tav3+/AimNbreY5p1F1v/suHVve/pwYasGpY7SqCpB2KgD
aoTmDcjMHCFsOFfZ3qrIkhdovJ5g2RGgWJAR8TZBFrQvYX/AH5r+j9NDlsk3JdefT4A7U2PxFzRc
/tTqJRc/PfdfdHjqo1bit+5SXH8n6e95kNij+8QzzVKtiq89HD0XTPPbUgJXrx/gI40Iqalx2hms
NkiFIR+Q2PIPg+77pBm0d5qx8/s8EhOYwR3PJpm4qC6k0AyOTzqjAC73Mxy9n4yYvDCf+O/9BmL5
K7dfWBGJ8nY6ed9F+6jARi5RKwTLIVhLjVratfSRHOKPxNAiS8qHAZp/kmdvEDMQgxRq0p/XX8iL
paeiWmU7/XlVitqY89wKmwx5ntfhjSES1niPXiwpEEiAkHTA8Oud/oC/LliWNdMk9wh8AHLEiX2L
teQsshnv8kkFAgd7gy7b4FbpjLc4lBWWHjWUC9T1XWr/rXLqpNVVd1AlcZmli/4grwTVjTb8+f+V
ag8EUsBz3XVTa9dp0uw5fqc5lmRAh/jsV2E/Ba7nOjhbvHVsCAkC7MdhFSFLymrf4E6Xf5U65DSo
vUcA6Hf2YX5+LYM3SCVkCDKtoMkfeoeDISSbzkVXlYLJu7hztVtW5UXjZxsmX5StcCp7Ea2gQoR4
pKE2axHoWb2L/n5dy+9BJf2pONQFd8TEfQS51eFPZOm6AOeYuZRTsGeIZmsoBBKMZh68cP9jzWnO
5hjrPCexJm5xj+CutCE5EDg04+MXb6fmo70X4/gpEpH4moI6Ne8qyv0B5c1wd2WcKyrCNspYtUw6
ncaPe4qVR+AgUzoQvoTjlPrFt/NcgkYZm0zDvSVL6dajEQKdqQ4X5oxLuelT0dmjvet3MVem8EBJ
TeJApSu+obVws7fGvcKoYDHBo/KnrMhz/Sg/5pcxYeVyuHbTldai1s4HtkybprJXDTXp+jB1w+a1
0NvS7Le0rmpFKwhI5fvct0gGbhSVhtFrgx5TB6FI5ErbiSLB8cg3iTJn89duW3/DfjCt/fh6H0yk
lSnyV5uBKsE47ADfqGk67EBFBut5uA/HfP/TVUjKNckMy0o2GKGB+Mye+c1uxkvClsmJiTdHbG9I
Rx7p1aYxW5RbfB6h9XTGSHvYu8JZFmAjh6qdR19TkmwAz1VoUjz608pIWRKuY/jdkXGD+/74KrJP
6Z+F0nNm27tzDjDwbIDYvZNhUl0zqhGuYqjyJ1R3SST4aSbCjJ+X31lBJ3dL5KjRMvW9xdPiyxhk
Wk0fhy6Q04JTa6Ab8xlgYdweU7pr5IwRRWnJjxv3xxq3pkPArXB/hdKt5H80Ajq3dwROAQH056Gr
hLkdmoai1TgHR+GcmVG2ArovABTxymUh6HolVQxT7A1NKS0XJ1Sz1CGf1C1JDKioXQxa2+VNQpbK
j32bN+HgK8nNNj8Xw/x6eMl+bCCyeDdrqpX0tUoH2SpDmjVMMYdRzHopPdqEtgnB9R45/uGzcrxV
XpD/b7DmZX1Yn+RfUt80NL7dzzGFDfL7mGAR0UBt2DGY03B+2YbfZF/+FN6FuzSvxPIr3UVGg231
qOh35HcVF+aLw4r4XRrFygIE+FRvF8kT2XSn3LUPY7zUIP/R+oBF0AAZLsOMq17XrZ82M6CZZ7Er
uI9PxqKD1KSvNdN83h+oB6y4rjX10aTIpFW5Ay6C+G4nxU/8IfEEIUua0kiwygKU4NaNgeDGwb/+
taaKaHXErlxoDXxahwIK8zR0qnRZGgyBRi02fef4AcIrZdfeeC2QB4qnXZmjFeipA1pZLYaJVtki
4FFTcpQPpmP9BvYxqCervWgWti2rcLKp+V2TjZgEg9xj954OOyIkExFKwiKsGdZFfue7EF8ltoSn
isaVDQ5w8sVCIKQbQNdw1aL+dJiXCL1QWsPDVaIfjbDnZvjlSpqC8e6BuINwMfbWY66s2B+EAjSM
4TLAqA6ibfp97LjX2Yo5RVG3yJgBz0iKh6lB8/ngcWvtwHL0n6CkCV931ER8A6uZOLToCf6lRsRT
vc4rIxQPg+TBxTjm5iSZe1/9dnUPZA6zxBnB88LCmI4j6iJi6J03T1d6Ug6qrUzSoXcMcwBmYtYh
7QoL1lLakZipUGAO0fyRgdIQ4p2ktURx11MgyKhQPlCn9SiWASwkiALLAy/U4omKMz/+Fq7ps98e
GxImjJuOQQ3NoKZy6796r7I0FtBqUB8KRT3KLl3KuiOX9HS9FHQZYvuGVPhm3bAEv+JDXSdWkuPf
RESnj//u/89/wu2cGlOkIUzArvziv/klQjh/CtfCbh2YNkvbsNlmZEuS99n2huyAvUkgPMs9cHez
d+28BP66a7tohcSOnJBzS+lIzGc0PAQtm16VNvqzIxxM3bas9ACs7mLawb6A9NgeFHvnaxiPZcmc
nGrGshuJRLAmBxdEuaDUljazEjdHblMf423QbexZwKCsQGKb/wl/wkwQf3pi+VPbr9u79Yl3Ur/P
disHUjD2MN4m4oHX5dOrQUFqPJc+XzJNWiwwIYR0izAZWRO4eD1+la7UMDv/XAolZrAUcGyZaOIE
wHX+THFfLglQfmVTuJMCCjQ9KFbpioxYg1DOCUaGl4NPKkDxzRctwyL97XGnlbE29gcaE94Fe2KH
E1kEOalSUHYAPG/9xbCrPmmBqPRbkAtP/EDuK2sKgECzpEAPNKAEbntjpdszQyqu/rofE0Ht2UF/
M1W5R718BBGMzp+17EcvXg9uYYFJKDIS/5Iml7byWFV4oYiph0DLi8/t0FQuy1gc1oKIN+svlMaH
kDFKkxoJnUM8wdxRMjG/48Ku+phc0MjYoxdd1Yvym5gz8ELEMEeKm5S+W5eE/GSgVK/rtdLFGVBR
Im4lXTilGzk9LzUeeC7zE+P2IR4NemcE4mkEWOWR2VGGdF0veYG81hI9I2nbc/UvtURJXZp7S5X0
hXis2lVyyzPvnArLv7cA8wQSx/foiwkcCl7+upqv9vXSxgW6SV4Mufbe+xsV/9oH8lyZH9CHkZDn
pYVIG3S4Mmg+oWBWfKi6II8Nwru6d10HdGGZ7VNWMLmZRN9FAz2KqRKKNkM2uLDhmsqRej0ROSRp
4Kcs0Ng3R8SHI96dKHFLTWua93JZl3vbPtYHkbr0h6JIF97zsmCPndf5oA0UWoGHWx40dauRb80q
R+ibPGWZs2GJDGnZYIOmLtyeQoVJ2/vpPyvYunGWEA10fAJ+/tf7UT8MgVqtbZiivXw8OhyD4NmG
M7GVnb5FSwdHsaN8Vx/oPKdtmxKHY2RUPNr9Qpg3AjZ+YkpjEsmDw//NUs0G2S+s9sfqMUPT49gn
sr4cPtXfnDhpoa9+eUqX45tyrlvqLI1YMeZNavE1r7LbQVEr6hrWOlgj7BibwOqZBD7Md7oJsVJA
MPQUSxshw8Vp7YCc3sodtghzv/ujVhuvCnFGslXa5UZpP+140+/AZzYXZeg0Gq31jyCONSc5L/WF
LgBZeM/xtUNse+S00Svebxc4AyZWRbZWG1UXGFKhEYUYcK8WjLpgEpkOXpb9eQeLkUtJ07WHh3kt
8OmbUAARSfmEzvCCQnsctdrO7AK4f6QJqgMuZmqeWul+ZVt3AeBbBEDU5/jm16t7sODS2x4PAB3f
vdU8nok+L6YfHeLGWzPBg8ZdB9d5omxzQFg2LE1gtrfQvFeK7eMYrysScI+u7jtapvQYs8O/W9Ru
HCddYLYq4icL6UkPL5/z0jFhSzMCEoV79ML0tz4eA3woO+Dpw6vbbYGzVtmynHVUG1cyi1emoCYK
0tlJ7QhPlilArGPu/K1Jzwsc7mQSpsLn0XotZ4O6E5GP4c+GZ+HHSvWHRjjj+Ovy0vn+diwVSju6
PtjqoHrFkIcV5JrwCCzG1/rv+6xRVD2ft9D90KqAjOhG8bg2UEmgUNdkKPIMJS7748DRlOOcC/OV
fKXPGsaNchvuh+ymghVjMrT9Zgjuj0qW4rl+DceVMdpZK7e3//djzdX3p7ZhoI2l7Oif2ab1mxjX
6BOaaG2T3/QoVM1o/om/wMpGx+wP11D76DCHHD4KXm3IovzVyfjijZLd2/1aolaJhLpTTlUHQVQZ
eunjupiKoKiZubEqF6wdLTQmGJwrBYOOS2V3bFrxERFBgYfi9rTQ795Wx3d96W89+ARkY1NW4L8R
jDqWYMoQuSIm0oGLracmVx7uF9psQ2KwssK/ekOMkaFmzdYzosyUESMbwTs2aUPbqORl49vFdd90
t2cFCK6mCn2YvIQAdlSTeS6iRq+foqs2vteyOhHPN2C1u8kO2Zn0jqc/M0XaRce+iIIISNSlXxxc
49858HJ1kKnNjbs3le63wyp6/QSFxZS+VL8lxpPAnI85+djKwGgyo1qIhix+xNPoDlqmIrOzvhYq
JxGDwBCH03k8xXJgsVORBeAzXP9phZ3tAv1ib0OkiZKB6akRW0hE48oJZkmLwQLCazI28QqYmBa3
29SW+TqSMcNchf8BKkZxAnjVjkIv49aordV2gEUgnLZ2pFatHr8TgWCDQTxpeoSyjMayJcQhTa+p
G6aJyZD2VyDSwuqnMc3qcBhYzHHNAaTwtkjQcKaIvrzH9Qy7VKGDVyWAK7dKgi1oNO6xkpRZjfbK
6npVfGJEXAoQhtF1J/CdYEI0aNo4Ie8gh9Jf84nUBasbbRld/2f6rJZ4hSx7eF6jTHWhQHD22OeE
R9g/p5kgqn9z3CoaRpFrmhN35KzbCMiGt9LduPobYNRcs/vr2PFUB2OrbiGq5YuQXkbhBqijOUdU
0PU/l77pqH4+Pu7i3skpW9D4pPPQ0NVfclbFHP/28PEkBMaWLEFVDLPukO9TjCNkXDD4bFt2LqAX
ZmdcIpof2zbmDYGY5AwT9gzed9DfZCA4luCZ3nyr4RJYfoHjP/H2BXL7U0srq4+OZw5iu7QDWz2V
KwoMvUbIS9LEn2l+AVjCygCwmdhxud+lQRLivX2kQ2gEJQyRs6Wt0kNLAfvFkeKgFRROPeNFCu/D
vsF2y6FTsbJHlYOZ0BTFFQcl561HSj5R4hHKLCIITpf1nuFT6bdpOk8XtHzDURnyQY04PR77cuBN
Wsi4WoQNDui0rEA0jpG1HY67ke/xUUeJ7HconBTpmd6+pgpkICpQ/FtOXbcFebxGZxoKnbKzKub3
XXSfnOiQ+Nr+WEIkv80iAZMqfqUU25kurJYHvSo+p5GGy+w2v4izDgCuloCGYXHTcFEpXCZKZYhJ
UsimcvkzZRv0Twu2K2cbjjDJRp2nrEDRhjHNqB/EhIBoZ9iLEJMDsT0t2QmWJGhRVfOjGo+Mzo7C
KzQamT7leLerOuk1nc/YO/3bChp00mv7eAf6K2sHd67Tw3SHpUic5/RYbiWC7XQvs7vRhix7WEgd
3xY4TPEcmMixoxpcAeauQvzxvgheki3PJwVcTAAEauT+MvHKGAuoeWX53z9Q96rHF/Plns6vZBHZ
npYoEfMIaX0IvKQaMcZxWi4+V7TdCx2KNa5MVqOPyIf1CSFGsrkIuulHhzVpRYH9VFeuMGHeO6Kt
v/3cu+lv5ZYkpguBmmtl+D6OADnpGYCclT54YrlK9eVUf/onFPDaEy0L35611KA0AukhOY+ra3US
Cr4NVFOxKO17yX4N8sYNXMkAn6FOSdUGYZsTN/ILB5Tjmwd3o+KDHVy8uxHxebKUJMac+8k16I9i
JFJco5UJM4LIxGK25kAcZW+HcbOKFeL85kOVdhV+VBNRBP5dUuv7VCDlozY58cboiMLWmB8xTYTU
B6e0akS+y2gAeYRsRfT9uKoYDqkSIZCF1Oo5b3nI13/6l1EGtpzplSa0YjhA8AMl+0Bv0pL0dlkt
TrprsLgAycEXwjg+ZiTCPgba7jw5MYCZZrJMpqZfdUhTiHM5cszwN8xzsco8wBBrknXioD2nmLeC
+JTMMyBLtaZ3rwz/f/ytZh8uB3PuiDGN4rOEUYr9ZwS8Fs4uqMZU8qnvw5n8XIFkID04dMkWGJIS
FwoikVU2qvUOXhMaYWrksYGQ3W8hIc1Mho2B8D8G/ugNv1pGDe5TryAyQs8v74OPFPl5TVQgXFOY
FA6YQA+Rc0u1YRNvUBMRAysVlJ/5GNvZOD+K4rkPizQTqPQgkjWNh6kxEV2iN9cO2I3myO2fFZyA
KFWqtq+ITiwFKfS4zMwj6ySwI/wfbowiR0PAIdJVmkojhX9mMtdEvMiH/DMveW2Ukd3rk2kWkz7+
mvsq5HHchnwhbkHcv9Paf7R9xILFXRAQ6EsEjIJ1Sc36BnZzX9vuD7fY1RVtnnZmvPlyv7cRrKNI
J+VXu5kcxKtfii5OTvThNGWGblj9pCDcdDB8TdS+oASpStYmvAQ1++UO3nghdqDJ6n+fTiqhOlgu
bkqC1u4PtkFS371I8QDnOvqI5NdICbH8m+TO22lOt+N3LMIcGhOQh9NCZBjwrJcPF53cI3/AoL/7
YfOig1F5r0QlD/KxiRTfq4a/5v5J6M0BVj83ajzLByDyStlzsfiUAM5pk1ISaduSIZZmfmkXlRSN
Qkfa6ETRX1hgEsdqmN14nP6eg6jcPlEG7VBNzchfFICJrec3aVvbjbI1i/RmXStbJdGYtnkgUnKI
VkudiBwrD/hLs6+mF19l3ePI3pCQJF7LqYwgwP3BZY5RPZHHLQ4GaUQtkEK0hc6cg5VHxPaqKL6R
fRSilZgUgYUC+JdCBN//bfnsBa6HUUJ6A/qmc7SmQNWH5KMdf+sI3jDNnYB1W+2kUp2VLQo5zYKW
9k5B39hsKIV8Zv/j5GjQjiRbGbK+EoatxGfBl5zP+6VIZyCITWp97zmyKh89JkQldKyAJEQTMSn+
NMuFEbzaiJKQVKHgaRpoYnyZkkh1pVTsKpNn4UEdIymC211SZoO529zGzSQ9+bSqVfLR2ckTBYak
WHiyuNSjsmVZ010PXppGHyHkaLmQkIxRAjVC06namcni4gN87mTW/GYtgbdc8m/Z1rrNbkmnC3X1
3sqQ2okP4eKxHixDXMCZkFzU0jrf/gYyVPU6/NIj9HqqK1pkCXuKIb7twCv7XFc9gmGN1pDN5uep
lPjNdezYCcprJz9QFWbd6Ptqe0hDJ0oyv9ffgr58VkHAW9Ca95ujDp9EjsSogMdi2fwZXg3crSHw
36VgnDTaOqb7Yj36DPV71NpQJgosKFGtIgLl65JvyCc8hbPlq5CqnYn2ezrpBWw2wES//zuCveIf
siMrW3LEZRNJTrexMB9NXk6EOWEdJb7AueREh0NSP5g2b7nB5T3kdn8jcnJbuBw5ZzlmbMtkqcsB
MlFqleVhwTrifKgFtRGmVdbW2Q7KPwrv5YTuRhTOJFFrot+ir9zJio6/grkqlWVW4sI0yUneRxUk
+7g9wWyfI8I+7MLvJ1OyzEDaijtyWqF0VweP3NSlY/tTvaEhEhdCz2gAMtfCY534N2GImz5wEZ/h
7+lYpVprM0ZcfN04RqrXnD/uxzR7Ei09wa7B5NbVx5b4ZC8b1ftO81j2tILLYnPfewnGK41XzJDI
hr3gjRVDC3z7dFEOyp9ICaXI+Og7BcjW2WvT2/LcoMVEouVBgkRvjLo1CQW7D/wulPJiY2WRu5Jx
Y4gbQu4VuTTc4L7ws7+hz8WMzd0T0Yvt0wPO3nQdeG5qve3r7Elb11iK4bari53DK9QzIz+Ngajr
Xf50MR/Vp5WsKVYD+txjkaexfTxnD5sWCMvYJTmabGyOQhyVhbRLYDPtl/Nb+sKaEElYs8wYZkzL
umimAHbTiLY1Y05UOaGLo3D/xKFSoaK77AE7WaNyyFYku1Sd42RQ0mfvxAzHNi8qCoktSP8ywMle
Hwpl17arNqRsdMzaOZxS2utzB36xsyr5Cu2+XRIAuQ5u71B+tpzhagJnG43NGl3/xizYZ18uvQTj
D2F4I04Gt8JYoXshwA7HGh1uol+RxgBcCE8ptAPvTHTB5j2Hnjp25EJhwmnwR473jXlIEDb7Owqr
rcBWEAwb4cKiosnbnuREhFKyhdw4pZ8Xutv6UGZy/FnooVupNOYi0Qw+xzGZqggjj5S7WG4TrL1K
ci1OuKaX7y0+V5Oqq1IAThJmlUmoatHJGdsc5mOxXmTxdYpkTIGM0oo31glso25PTI6YmFwf/H+n
/In7bz9o6llRBsZuuSCDJWFKap5JnK2KHjiARSqe+3XD//3OqIHz/IEFqOX/ymXvlJLY3XCSxqj9
6PFzsUQCnZpQDTpCDr5szdUrAUAbXuk7GVk1nox6NQfAHyXisnmZGNslqWGitVvDjPhRgwtAON7r
GrJdvM5FuUbPUAqspX8prnMfLJvKwIVfPu3BLK20XwmU3KWMq1Vs5GmmSCUECDYgGBG4wQDDf495
xE85pu30AyQIShH39sd1AWRLzDXgijBSm2h81EDCn43LTlzSsNylReHGpkcZLsuJcWZVWSnoHCs4
6xBZuqdEGLcQn5iQZHCIc+XJXMoPeEP1LDC5RWRFPer1kx6eMnaMpjRnymHzCrMuYdhJMIw56evH
Mc9WBGm11NmVhF3+A39MqnlQhII22YB6VKPGxTbyvX3WldcveznKRxc4H385Ozo3BZ34j5lHYjXH
4mwhCst4GgpAdxzNsrglG6XTp5uZCv6I7TSnOwIBA9pPQj2uSuJ3m/VumhwZrNv53qr1B6x/Ms/x
0seauJIkCO+3Q4QlzWJF31ctSFSW1TFTVqFdstuVbLgLcOcyE/D1KzKjh+obui9mbcNEjO/2lLHn
Eb3Ekw4b1QvOWKxqiM87vK6PCGdgtHTJ2NX0mNRwowtAlTly6Hc6D9yGJK1XL3JuItlpeqHFWKk7
q1Q3E2sXDaehqKpX0UQyf1HIb7oJM/qZRxSp8EyEDbvyF5I5fOZOfG8PaAMuc6i/whaDEXuVVK/7
fS6MC9HElhkLrR3J5KfvEaZDO4n2VccMaDObrKKX02VuTW5jSvlWwuudygsf4103aC/or/nVqvs6
x9neA7e2cV9TZadFTRHqPmGZ6XovBlo847ZOSiZ4GYa7HAXvMLC4T+BxDQYsieRMNr2n0zmRwcZP
to6xOoek8e+XbcTofrZpDYjVFopLNToskabP2I7NLzrhmubUJk69vZ201PetO5hhV1xN9kzYlQMR
LntEkFA/yX+v1CYXQHOBpiuh6d2/4SBs+fk2xF6NjsdgmmiLI4L+vY1oV8rdf3TYZ/wbuglgqAx+
dWdmbDqgzy4TD8VCDALYTVV0sFe71M6lEJMRUMw7HCvgbZSGICcUC5OzeV+uW0sxlV24q4PrOqKr
z2BFc2xDUoUudbCKBqcxGFOMLeEm5s4Od5NvJZgXAhGKSuZa/e2dRqSp348vCucBxKBDEp3sGEzW
y4XX1AFgmSi5Jp9gECAn0EUbBnwRiojJFlEzeBqcGfkuX5KXMsnRHk0KlXUnVJ10dwn3ei2b3yCF
YdL8XeMIb9GjCSdcj2x7qT5rrF348z2mtJDF4NtuB/dyZETLMK590wgh4OEmR2QlbFi8fQAanB9r
/X5BwgWXaxCI9KaLNQFz9BEjYzTVJKgUzHiOGGcWiqj0V5r7VBzUaJHtXNV80vH2vzVBuqeu4JEf
VskerEpDovUM7yDR96exf3L7/W+RSG9dcpg+Xz4kpicghAJql2c0kdVy6duvEClsATw6xbHYON9j
ZwmxvvztmXJZyFggPwnPbZDzd6V/0DMBYYbJ3CO264DUkjmfsMSvza7czBrBvx2UB29goObFzQqs
1tuRYX9ON57KyaM3OukcIiW3yy5qYi5WSC68o8b3A0EfcwN2UN8lHDC3lIHKyhk8a6nltSOB5d5G
w460a4Q0NjsdN2b3n4WacI/aK0yfQ/Dy/uvM1xMgcr6WVlnXQBQsyvdLs9Ee/Qdw39p0eEocXWU9
mdMFEMQMPJHb0r744kUplxdojjLEgtXl4CrHeiEziwkdLagLIoQSULMlczYftlh4vBD2jiQLfF2v
MC5Q3c+4/f7UiBhMgH6tpDCalb+KeZ3EVp1GfLZqii2TmacaM/IAvb9PCccizlD392h5eA9f2EEe
1KfNzx2EvKPtOggLKwMI2aviSwFxRjh5Eo2/lIEdBSux8j3p5YnW1M5c/1hmCOlrEJtZaT85ObF0
eMekR23xin5Y76a7GnrpELYdRfEs6gRP8O96BLjicLzI0rglf5NcVzGoSQ6npDX8tOv2X/W5zoai
xiJjhKGE+TyVRlC0xtuMErfnRm45iSh40r372o/4d7F+k37sTEiJhO7XtuOGNr5JaI19BLcqxJqm
X1T+zwGAlTZLZ39i8mxx9tFggBASxkGVblalML6JL5HKw0eVTJFrFHPQrnsLPONnTKa/WIzBTbc7
zSRsSOA2Lnp3y8b6y/jDUMqKct2ILZ+2kZJll22h8IZeGXUJao6Qs5FL9ekVmeLFDluJEAltHfZ7
Cu1gT0U+ZdyfOEof0IDqsH5HSxix6e8DUe1C51AgmWtNP98V4en8GkM+5e4URNLldHBiAKnAbfpQ
CIpqmWsJDtbcYMcCl9tLIggYR4Enbdg2ZsYHI9jwS5vhGOL2D/ivElIOvR2Lyv54kR5p/uqRPSlC
mFh79GxmW1SXlCxqcDe5/S9//o7WLbgMOMvhQ8z/rHnnPpBdepMXMsEhPwSpIEMXj9H+2/8ejHOb
FZn8EF82IdwrcgbUpPuVEWpP3YLOPTBHNsoNtcfHStyc4b+FXNSVxm6xn2ro4TVcEjXq7mzXKLTL
XgkC0Ph/jxJ2JWc+1k9PKiBVp73ECSBlLp4GGwrKjYuu8T09Iq5+UYUruf9+Ewj2ZigFeQIQ1hPS
12bWjD4RSaJzXOIQdI759Ct6gtY1sXPT6Gsez8LIArjQF+8Wb3hQhHvB92boFAdjJCiEo0j0WUoM
vkRbliRW65SrVfMSaw5/0rsfwDXIix2V58wxQTay05R9HfKezxd91uBeYGapQNHNnIcW0Jxa0YUy
bFYdp7XkoT3xMRNhl5Ix5tgdzb85tWMdf59hjT+7XDvfkWdt1ajXuAN4P/4ug4TWMKeLh6GkSwDA
6Np3YvY4Yi7yw9LVe+exAMxSaFRW0W033l+9RbQW6KSsbd+ndFIHXDOid1VTK7uM1I3czB0dcCOj
05bgfWDqp+lVhxTNwHZUnrbd19mDb2ypMtezBLWR2+FhUqZTGGxRyMd8QL8QeKtpLfCV+c9sLb3L
fxqGEeUXONgcQ8CRPeX0wwCJK3YBONUOfsL2fOMPUe6Qjy3va5tYjRHOcqJ8hF7PfkXobAuk2Q8S
84i61Qs72Uh0SwggK6atrwi3HcR9IKX8LdsXueVsoy6TZdBye2Yq0CTiF5sMy1cH/Wgd6Pd+j29D
sOrfLbQ8JtGdUOskcddcj0b1Puanp/Fndg4lJ+j8ne+No603JI9QAYlfO/5elP3/nd202i185xY4
qwRTpSVoe7nBu0VGoZHUSbxs/7Q3NivKqhrODvdu/jxO727nUQzIzNvwNQElidbdx0G/CatQqDqc
EivXqecNAGG7mpsN3OCWtpiIamrTkWlLaog/gaUhhrVf9B4iw9fjT77komhcBqz9qbZ79bQ6V9Qm
NjG+T+auBbBseTzqh2ViyxmHg0DtiBf29rB8fgLP0W/duiA+pbBXi+jSvs6aLli4+//UjtyEfqRA
CqCdkjSJkOUMy9zMamrD2GN1YrM9pc/3+p4s30/uS2AucZsDkPY16sdOBgRKv/FKbPPu/zUItd4j
2yoWjdAxbqHAQrugrGMSmJ+AGGLJ1FRZHEYmokuLYkgS3uGkKfOatiU1sK//GXbxAlBwkKhzn+NR
GdNb6o0Bze5l3J5B8SkhQmL8ZneuyjjT1V1lJbSxWDNYBfyyTF83jKh9kExxsNtEDAFDXCyJcGtm
koHPXNUQb+0jIdQ0Z4wXmxERq370Ot9Yxa0IQvMX1/5jalWsq17njOLfPptaUcvboo4ngGnhgw6B
tztI4kLIDW1ykDh3BMtdS19AQ2vhURjyRz2UpWStLhoFe9ZLW9mDLla6/DV5OiZo+r2ZuaJB9F0N
f0fY004piwHDQKlfkAsrhsx/NzPrN3jNF+YSc9wYNkTnwgld5Kd8/FfeWNQ6YM96A2KXCivkxCBH
6Q7jKU753OlRn0el+Vv1PCi84bK/1yu0Xmx9x7JXRMHzOu1mlvbWMHZ+JYEgKitF5Fn47v1Jy4da
y9QwnWJrhLGsF+fKoEvE8m620yfBt9jOmS6tMArNOckAp2uxikBF+3/NrP1PvwQQrSccABhFa2CS
xmDC4WxAGCBHoRTkPWuiTpTYQhdhXPJ+Y9Fvm2nvu3kd7HK/oNNZdlA5C6hz86phfg1LSuGYnHhY
qHZq08VMmamF2GKmDG3F1nBYqN/Oqj43qS54AmaRDs8vDQZYh8aSUaCDenQBEKybchivSNiktG8a
l5F26Kk6YIZ9gaY4sXFHremWkhW6XFQj/oHb4wf6MCdkIwUJiKq33imURRl/Ky9hheL7B3F0bz/Y
JuGfcCrsQ4xpv12DpZVzvkXvjU730qCxnJad/Oox1VGDRODuv+l0guVKe2YGzjltooe6rt2fcRxK
LC5xiFtTPPsZHMXXwlBXHFbV4d1WMPGox6nbnzYWYN0PrPsEtWCYMQCenLYw48Ck+Uns12I/YS6b
MUBPot1SpiaAdG/N/C8dSfGrg7JRA/zFAlu6PJ5YrH0QnVdYQVUrrgOMsUcjYnzyPn9gaz26c/ni
/BYWrAH9wMsFAr22pQWwq5YMpsGT9a24zd0vZPjWTjMReNzH0cnMteJ43mPD28YWrdYICOpN2I+t
aRlSLhz6Erw5Y8LJ+VrxOy5gYNKH8PBD3Pb6z57cheSMDa65wXBW6twk0PYvLmyuiBLi2CylLAMs
7k9BUDtBcx/Oa/taiVpa2G5iAuqmX7Htuq7dySxrZYOEOsFLnXCEG6kwG8Um9Lqm0uWx6HTICDRB
lLavXqUa+9BfCYvs10MTWmym2QwwvoyZQjXCAgJqySYNl32oQKtn/HbvawgB6hFPxrYFzBwpHGC/
G6fHvmoyZq6d1ANEHlxULyLi9DxbEQvuzv0/Ku/aSgLxVHOy/uCgBRmwn30okTKed27L6xcgBlAi
uV3eoD9H8/W3MVQHfTvIO8KM7tOCnwGNV4Ecmd1DEYS4epM3XVPWDqwFCAjHOkWbgyz3xraXn09A
98mbLb4km1yBmNMYQBz/kXRKzd1rfhiTotGJIsUrAeZF9Pk4c4+qPNzntgrm1kf5BxHnPhZ2fJap
DlsVmB3mKZuk8od2T01NGYjZZPU6yphNE3dce6cz1H5yaLYoOzQFpeYobpokdGp1PCURgqEcxFnl
JYiM1GWJjUm+2cu/JwbIE8dMINH5NKa3osxfQyuG1EMmjVLDMZbWdLRhXSgFB9WsRiKWckpb+WzB
HXLO2N9D62oDJNz8Cd3BxRXyZj0r5+XNk9PagdLBfBjM6sslbyh7uBIOi4Q27dzWyCXoM1GiTxYI
KFRvbgkRKqCzgcFdGvfI1FtkzPb9ydM23SCukgtzUGEkWwjvIaPmPx/pQr8YeL0KJcBqgG/oTyA2
nax+iPUicVSOerDv/mjm2KpCJ9/OeoFkLT7ipDGY8NAU56IlqMNprXw3xbi3TcZimWxRPfQBGBB9
f+kGH9YfNnS6oVbqGY+mdILHCXMSku7whGzXGYm/fLr4k3JNZGEmLyngIQeMd0l0LM//+6c3Px+B
UIvTXc5T4Qhpf9N/yqhq4fR9RgUqisnXnOyXQEaev62p7OIJy5B3GC6gQ71a2BqCGkD6LpaSQ8+w
heBm/9Nh27Ykk8r+zIXWJJ6qpN73GwcGSnwaOWOQ3jbO7+1+hkOE1LU0f1F7bltTVGteaUsBzPwE
M5rBmeU7Il8G46exoyMBx/wa2oRaRppYgY5b1hlRWPCZMBseAWMdVlCHBI1gnwUh4enuW0DLZBEl
M3BjHBjtQZzd4GxcWl7fiV9h7rYBsvziyKTbmEhz8WQ9nJDWzIViorHyWkH5PP5zDCiyMkTgVyca
Csg37Lx+R2jZACxM40QthccM0x0IgM/6GJPuNy0Mt35MfbQDAGg8++bk+nWtNyLZP3zr/e37JLbb
Alvkf/0FDIwNa/waRVKhTx5W2qM7f8vbKM53/5Ip21tx5sf41f8w7KzUk16a3wB/UVBJw7JJK9Rq
lz5bi9pWe3BYqUuw+7zfKYqCeA2/q/6yz3lm8W4sZNWh0V/nLi3N09njX4nAMlRdA1SHVcuarf02
cwLe2if9gavutN37XQPY92CO22hhvKdKgU8S1FjxecHpyCC+b83lzVDb/vF+BYKJUBSnixV30XOa
ZMgdlnkxA8qBm83b4X7KSs3jZR0dKeG4DDGeUyFZOJsFhjCcBWXzbsSrl8Fu8dLuSjgJvSwg9YO+
WftfsskyhqKdYwqgpeATP+QYqX/HxESULcwex0j7mGeg0QQqdPixLSKwHRwmX8b3AjzpiinRQSry
GKte/GwgXCReSB6Vn7k/5dLneygMQExiJfQgUge0HdMD7U1vMig1rNpMLrpBU5n6LVmF/N1Nadlc
1IkFGsjszW+G63PLbtqxFFfynsQJUSuNa+iZyYqxEmjHyFN51J+I/T0A5oTbsvsj9XEXwN+UBDov
oZvxQmOqg7xm6qgBDeg/h04ctcHViA7CkZG5AeAdJCe/b6/kBRGz23BZkg4qhwqIV31L3AMMPSlV
VBry6q2ApoHOLvxF87RJqnYsrG/co3lPKc6zqsrzKQvFkzugT26ZKSku38G0ta1xqCRcbPPshCju
XhTvAT0Zh92efmR/PXj1GzslgrMz9Tv/OwPnr3aMBuB9JdxlHBMuTJ8Kp+xnbJvCHHmvUUYRC9fT
mckxfWZ4jPd+VhBG0Uh/FndQ2rzELVrwIJU9SkGsD2h9HkxGOkgHcp4XuiT0oNItSt8XYOd9luO1
LES01/p645ckoa5Xc/Hu8cF00ub9lurISfJWXAONylF6JB34+791PwNMzNE1HjNQF2mdEsVB/IP6
aq3vtoTgHTCMWjmBrBUY5TvGBVzO/GBh1Hwv8+lldEUKT+jZPvyyVBivZ6vACQZ0F8H+4watO4M8
lBhsr+86Ns9tN01s3c0w+bLuBK5dfEv//PT1mXhdjQ/drlIJZGFDh94kqvbnhYH7QdjauOm/EocR
JYrTlb1lY345b0bdIpthmUWKBUh9UWCrxVzhh6V9QMd6Nu4GG+cPWXUbuhnZGES78bXg+2Wde9U9
IWRe7TYMba2tezVeUO4rjJ46aYfxv8CvI9I6vbfpf3n9aw92JNIPRPFM/N6zRk7+S6S0iPFX480G
4W1utoqhXjwA2sbn6lxM8BNk+QI+yPiP+i3PVKu1CG5HS6YHKh/uawpFvoa401BZqka3CjEzVoJN
/Bo+gOxqRcmhha7PSW4v3S2FxAnNRzdMxSMeKa9n1ckvBtO/fAdKB6IqlOgHMN4gsy7ytGEOwRjS
uwRRxwCAM4wz5MWxyrTRaFTeyy3TOZAIG12N/r2qtxdBBXwZzzL9a6wbKb/HlygcihErq23V15j8
69STYUfh5susCxwR9PBrsIqqG9o4duCY7wAYDqwtPB9/hW9+XBd2DYvyDbmfiIdGxwoAsAUq80Ic
hVQn9HJqkObUgeiDnjFtZqhC4Zx34FSjf/TLi9OYzn7Xi6qzVVcAB8BHNHJ7KMnB7OhdFanZNI3W
3PQgD3ehGrCXyOzU+2G0lbLuUXIEpHEsfGHY8fVmxPrOAIYXMqnK/jSwO+d/4Y72gSbGmdyMjj7B
okvpn+tMENgAa5BKolheYv4CtaKjygh/zFkOQK8j8v0mp/MsWRrDGcYWYOCLmuCCq/i1FJOrdDeq
5i6fogk1iMcgm+dR7yCdDBt0iHTIN2zfnJ0GwSy+z0EQEBxVkwrFkZYtTCbsLF+H58PP8BEYLWV0
P0yjVl0mQgUPFEwbZqwEx7dq8iAsj7RCSR4qOVdqpC2htdCe7OU5DXqEkjt7O5xsqNTLMNCaSf7u
yeIpOr377jtq63dyCp/37HGF8e7MW6/s00lbWsoVruchIcFSBBw9p4rXk7CbPI2i8OjXdQWdrpWq
zSZdEti0Vq53dxMO/IlrBi2iViIzir2xnvlYE+uU+T0H8JhNSWAYz9WO+W/Zgs4Ya1Qev22NpZJE
1Nu1a+a/Eyc+sse+5yJSa8ofJlqUH2ZLARRPhaNK7Wc1jj5JKvegiVX61Pvn4tml+XmTLEMR/amm
kC8/rk/ZCACTAw3h9VqNAvAhedWT+kkgstBce6Y3d0kuM0yFXPgV2nrAcnPgN0OVFk8NIWxaeJu/
rFSQZMERapc/4bJje/hU7YLtVNGpeYTHaoU+avIwq5WKj7HeBtIbUM+N6VKowJmMnz+REeR26VF5
P0w6WZK79R0oR0t6uNamaHLZLOIhZSbOn3uPfI0ujrbKLsoPK16ZBnv+n7F90TMW4S27ctdMtP2/
uzBX6OhlVeKSXnAOEd5LdmSnKbxaDef/2xk80aOjlUF569TA7xqgLhAc3N40UlVCsVSt5ZeR6GxV
cpsvM4+oQz01yGSmcE1BsHaA5134/w0/PHp/FuBhwmwIofmG74PoAG/HXEAXTiW08NUO87ixlb7b
/7/zdlSOjx2JRU8itlUecqJMMSr1yYQ/dFXP8xEHp+PoE36MuTKSyuURcZypnwKljF6iDgHPLNFn
I5BV8BhnZ7SncCn+e1F2PEkaA/fqgmiT+N6vQ4+22wXkN0UaiT91c1QoDPwye2pEjIvIcDHFQnm/
2K+N4pHe1Dxw7/y/f+hsrOJ2n0pdJpIiztLfLHL3XyBTi+5Su2wB0dxRXNznWQWrQjD//YrT9bih
HTXBN00CwF1dkPQFJXXFxJHRUmTYd2xsuSyIxnImKTDQkd26cfOsEib9ocyvwNPVN8qQQQ2pW0cr
MR3NCX/ltVt3DXtIKifPWu462znS5070ArkgVspWM+5w1SdZrkEkjogBNzycDYW+XySbw7AE4eLK
kQwNMVJg2JPse33MSWmoONyQkfjtXWztO4RF/sPHvJyQinsOg51K05CZ1Rf+yENsnoh8ec33wW8M
odT+pmFuDGWPLStLUu1rgbJs2n+lsfykyYzHwp2EIaO+EpTfcZ7XhooIeb5kx4ECSN6MCEBV7CRX
7uq7uDqNlv9QWDrqgO/tNUCz/N/JgJk+TzNdIWqbC2sz+GEr21Pc1jjL2zpH+GSA/o1maiw0Xk/f
gHNce5EMuNaGfQOoGHbuKpzRkkhsP4FQ0fqToczM5FWM5yW49bhaqfic1tH8TTrqAZoZEML1c/mT
VUh2IYuurdVxfoOt4Pt9cbViXZLlu+cXpnwVlpzVjkyUF7+FxQm7YKkU5qqj2m4NtzbXusl2hYlj
ArqXiAoZkt+Wa75/Fi7gidf+nX5xAryr26Qrgf8ow1l577GcAPJSv2NvDvQX1g3uHOM+mcF2EqCg
heVehSUj42vcFtAxa1ircHQnJS+E4YwpJ4pZP53016PnpLpsoKa7p5dLsuUq9rhCmx/PUGO79mxf
8qon66KyBC56xg3Gzl3RGRFj8gDakv0/YawfMa+cZAg09+1Ep0flaej+pgA5MgMv4+UwgBN+1Yw3
OTQhxE6UQyqKe35dY3ZxsSVIEH6qlmGtSt0z755oNyICOwlxi9LCTYV3BfYnSa3Yj4cBu8zeUCzk
HWJYN8mh9/0TlhRIVPBjirRWrQnOP6hZ6OYidT6yWjfdFqfQtuNXnwUtKof3ro8H3wr0r2Rm3zpk
dBQ1eVOO8LCDuDm7ghmQp3kx1KI8fTKCk62utjU/pw5ZkwyA9gShqNlREdDYGJXfn9xumqHGtC8d
H6k95ahrq4ph2ROyzHsPcL7U8UrtTWcTyrfokuTgWygf+lZ5b7ZSDDVGufUh2ZokqXMFEBtqihDN
QxsK+Di2siZDU+mr99SRBDl1gmrzUxhgRT1oNjYq/QzX+U0P7nuN3UCzkkkvkVcgAUFOlHraEJhv
YhO43y8/TMwS4d9gKxBptUxqyCFhaO4GvSdoPDWhWRUn5MX4oxtw/CEs0r8xejnfiiKTNoIXDWVt
bmuYUQAeKvIyA8D5/bL5BGwfd67dMUbqdD7/xcdPviLjqkygM8qfIdfOYXyzCuglncF3fHMN3LGi
IpgQuef5H8qYhHf+yZe2Mmp8xyqIGll+Dw2oB6nTS5TKk2F+zD/l34Qeac/HuvKW/Xlbx69HAKYn
Viru8LVMtLe//HXIJweBcq6gAzP/F3PE/TP/8Xaa9fNIczJcF4VptBEl98wGO8vIrsib59T8ACkQ
2H4HZs9bBORPHZPEfxm80HFw0K4cxepPhKQeaN7Q95wOdctg2YVsu2dTUKyhI4eVu9CDQhlX8k2s
bn2YUrbfAPfztSHP3+67MmCuKBHG/xrysFTtca9i1a4GhAvhLCEBD4yqkh575p5Uc8J7FgtXVoge
thXzwSaOv49MM2UXjB8IbI8gnXJYHT7hT4ZcIO7kumZLZQdz+wE4lPIm8BzjBKEA9k2z6US8tpav
UrLKigODTjdlYyZ15jlEFRe8a9OQiN8VS8lOgQzSWs6X5ufOS21tS4Srt7ncP3cZRV62xt2LA0bc
BpD6qHEHD8gyXdKh+H6iSbUTsuddboM8EZ13luJHXwIp+6P4d+jaoQqSK6UNHFKVO5v+BfKB3SGK
V+IYy6NlrkdT96RK3GbMJpjcNbSQSesvDh9u5vledYrW9CDUWIjrmtJc88NhoKOjLwgObw7Wy4fU
6OIAULgTDOHFCJBDlRcUHS1r7qhN+45iEG+ZLFNFiyWEotLrb78b9/Ah+wmmvnsGNBETHLbLFaAM
DfjRmY8Z4kQ+imlMH/Q8loihxPr3XStCX7+twdnGRf5g2qfd4lhZRxxV/JikmWK/dzG6zmc62eet
GzLwDBoaK4Izoe7/i8CyhGuDbJcIH1ZL5ZBWLU1PEi3d4LR91NCjfZDLr/KUaCXNgiQUrA7rfdYY
uZVEnIcNjKereGEoTcwfkgB+fqlMHuOsiaHwo2gF8D7LqtIqrdJO5BTafGcYQB+ktM7X7KtXU2ht
F7dchbaMZI6518XmuIi4vjk4EH9AlkkBfIlcF5DHNyDGL7hgZPmuncD4PgWirsVB6QxAuQDjTJLG
qfn+xsoye+laqKAuUyZJAoHbOEleV0dqMToGl8ZI9HH3gmhD1dtlNTnRhTnRjOHpp6IFSIwJchPP
j3gfFcLAwgmCN2HqS0w9D9Yu71sTvCI08qLQDjGlexukFiFZZ9oOvU1wAkXEowVGdcl+/k7a3vZA
O7cFnZOGQ1/K6wS+zxYM/v/4GhcAcWNPpmVwmzmth30W3PTIe4lqL525dLejXCzFomUEEWfDtrEE
4cXGENVENyvp4YGHqgOclJL8p5/GDAPVkuDuZJkHD/qTs3LNvY7qknQC44Gjte7yK0v5UQLg5wEg
YnAHfegTKH37ygSF2joWBOHh4/SE2Ge+Dr8aHDbgTYeZi0IFJY6eO1vFfHmn8amLdFuxki0tazNy
9K77/HoELoU5+4HfgjuKzE7CFnvL7WHzAcGvL6W2W7cPut78ouixJovBD7g3EXzdwC41Y+H0GSZS
8dwiElXkw01YLylF8noVqEgMF9wqDoaL34l4rwo2Afw2Jqeb+ZrvGOan2LZfeu1Bi9ZKyEVOdHdo
zXP/P/ekW6V9gU2hcU26DreJxTA3DMgiTcI/tCBDpFjN77+ZrdUjOMXLI8w2CG7B6tuWZxutMBOz
/H5utjcsSRiWNCn5cIfQ8V3z+5t+muX9xNVbhwfDb0jcOlzP8PBlMs+kMYoJaFef+1M84KTcJxvF
yL6Pru9l3cJkH5yK7MWZEO3aifaHJ3LTpYGObNPuEVPBl+Y3SVsae+isesWvr34zM4YC7aJ/y6MM
5dCB5XyLC2Hu4KNshbWP9K3Ux/Xs30U+y8zFTL3f57g+CMnLHVc9SIyQHs6zqzlt7ZAZCaWEW8el
gNgiKqmzTYrgVAoi/O6eOA+1KeIzEd8d0IIwBrd4ORAyHtKGTK4zXQE6+EnqYIA09v3q/48Z7mui
5+/x+MC+63fAdTVDw8RHMqGk2EG4bPzKNN6iys9Lak0wz0Y0hvnFod6ELJyHePvtWgkJ5u8aQzTF
rUr0A0mrO4mJJerw9aGY08gF87iZmbSeONVJ7FPWsvfGqaw2cUYCBtELs7EJRsu/t3MshfU1Tv70
SYQhQYAfZ0mjBvGarka46mWPGX4730nT1zU8lsS4hz7ZiKrban67ExxOTw6PI4zH/QOQP7ivHU1H
FK8SUSTj58laa4i/iyzAx6NPl6wRPRgtH8BKo3X0lR2R7BtQ9sll+2me3yp7znuXfjLDFhYGpD3z
OT3q0WP5mCQGrcAjgErdfT7K+JlnWCSG1D48DXYGVb+J/p1KULjpG1IZUzR/gpdyfMQZrDV4/uUf
QxJXYB9GwuA4iRIyxp217a43ktV0pef2vSys4HKiglXlkfiWpk96H9yfDxUAbvO6vYOU0B2DFYtz
ilAgsPaOhtR16GOKODd5zjRuIpU0rHuluPZKbvlV8KQ75PtgMCTNr/I+5WRTNd8ScGjvfqKKPwvi
p3+S84BXZllJPYWO8fTLJiqgGCYevZ34WvXBhdeCGrR4+g08M8uwkoD82rEfP1ZicSyL7sKF7Rfc
XFG1SkeKbY7tbvQqVt3QrgJzFfGbKg5yhOG83dGQ7kR/B+tkSqsbDoyXYCFRset2cUDjzxdSRILA
6Kbku4lGRdluPNgWm3OhDEeR9fCYYrZLgA3knlFPonP0ZEH76Tgo8BFdo7B5IxWtrFWQRrfoHLZu
+F4mt+7XzWrJuZ92+f9M7ArNwuFqDLX11FKnMICs+wkla8Jep1m8GpuniUwIVK5effkrCKEkW6gD
YgOyfQBNrMyDoAPjSTnQXmMbN7mSII/Aj4NImMS34wbAR+7x/O/1HNPb2GrwipSB8jJ8bdaSiCu9
9Bg6rMGFlvGYoK2w67AkYauQci6y0QmSFRPLa244xB037WGcWxLwhwaUaoYC8cFAajaLw/+TSOP6
yWp0pvIqdBjNEIG4w/cWRnQizG1dbbasZViTrIoIvTQyDbhHI6BDHWid2eqLh6dE77lRYgbBldR6
htRQ3qhjeTVVLiT0VjmD44PBz8RTKAn43ZWAL6ZOofwLmF1kInnBQsjCXNLoqw+mNOs0nyFOYUy4
r5oGJP2mtpATu9vSXSj+issUat2ljPBO/CHYhxM99klGYrr6E5zNmbBvtXCAmvs4Du8XcmMHdMak
b2Q8QeWWxH57moLo+pbcp19tbN8JKhm2vpdv1eajh55jLYeoHx6MbDunm6YmIEC1iPFTj+KxK6da
/XO/ERK7NU8ohbf32ciJzdak3UN+6LF2kIoz2QmvftMJ5iajsVAJne10350siEmt8IxBCV1ATnsp
mwzNEfJ9xupSA7tu9XhCm3dWApAhfEwkkYXcE/4R2Fyh52ZR7eZPl1ejwUd9oHLhS712jvjQQURm
nDxTzal5pKPoTl23sfMJ8zibnU5s0e8YXnjXSO3oSoCV32nl2UDf0kTkMyLlkfxgNAhnxOweoUdp
KWJPpRfv7FqctsVVjnjsKRWjAZjfBd6pyHQjqQG4qs4TQLqJbRMffeiO9rXxMXnrOrgTB2CPkSSy
CLSURoe7elq4iHkjqt+ibLj9XaI/Ae87Q1Pnerj5U8tIrdbmiyKXoBS8FwKAeEpyymND9TX9uIdL
tjANuZGNsR9XiZhXGtGqebBe8c66uSGMuuJzSmcPVJmBKeUOLZ4F4cUtK3wSOcBqeCpn/yolEr4V
ffU1SJc3AUxv5y10hL9HJ0j0sc3zdCj+m/52o/dTqRv0lxuC+TysVn55xjRt7s1792VCC1+LgkYL
XxhflDuSXSPGadE8JZOqJ1JlLf7DSNFoMrxOBJYo0Of9z6oEPmY8WzxpcavJv3xFVY+ch5q5Br3b
s6lG47qOIO3FECWnZcBCUeuTWP2M5ix1mKSFdKLHLF0b0IP1XGQR7kVfk77DxPVE2vuL5RE+3pH6
V4UjOpUOQQwNihUK9q7vyB7G6kvtww+1spvSkUOQwoyHkyUAZSnzJQ+vpK4EacVAeDPjdSH2nEbk
3tb632WEALn0T4NR3nGFx/u0skEweAdTFvg0OhCLwhBxE9pOyhYWWU1K2TOetMbz3rq/q+uyVL5k
RmduadcP40O4ZIUQF0K/I7t91GYJt3YtR9Vz+Bm+0JQMdZexqBnFcD9DQuANOFKqD9SxiQrMFvuV
Il32EsekBEXed4JhgzeB1itFRAn7o/TFiblWyysrPw5GbBG3WXoZCAWs9R644YiIimnbu2okjk6M
toSWfw9TcEhmGv64eyoGdKChENnj9163QD6ZVD9PYl0Fnb5vqKn+tofn4YScUYEmHTvxk78bj2ZY
e3HdabEL0S4DOy3Q89a2TyQP+wR2Bf6xHuo7+LxgUBLfbbBGBwT1j7uR9ZnCY9wqN/A7GoQxEqos
xaWJgG3QmOB1bRz3zK+WotEW0re7yFIvIKNjRuQ4503r2L9rVzYY0U8u09Pie0sabY00NHABxIXj
TDG4F8rjngynbpl+WbL0jEcS3LmNZaIg6wvQoh4Q5PUVHwYhZDtj1M+ZG0yd5iIqGALleddaDMjM
9YNWA4WvmyfakydEgQkDocaJYzSC6keTd2LUHZF1MDGpak7wrJuOJ6MsPew78VSC32ezQts1BCvL
wmA2JYskqpqMyoOHSYsNTikelNeI4/CTIixs50g44/Shdt+8+o14YLPxf0wc/LlIKx71aXTJSLzl
B0vZ7hyHZ+A8FMhLonaLPa9fW1EGsEHXQU7BPH6WZ9gs9yUTh9PKelEvL0gttL+ME/Y+dJKz69bn
77i6s5AMT2iqDExn+3Ml6tHMohrQBOAOE8TIAnBTQtnlIYnvqjRP3abN/Xib3Lzqt47ThlZ9tz5C
PcVOzwEHT0QzIWGaCYPqpsxO+STg0FTIfY8mwC+g9a9H/WmGU2+AQ4KyOjK5JKIL0TPb8DLqtkMs
/4l9nOnc82gKP5R+Bo2DPMzfrdVSSnQ2oOdhXNldK2vwlF3URsU12dCpzCdfYq/AyHmQngLQVpXK
LFritWaXvOAV7/+PiVnihLSwFHHFvnIsn6r6CKs03o1WDJPH/M8cz6Mv2oIwR4Ind3gDIzV5Sb4K
yLIay8H0phEj6laqpwvYLxFkOE9Ne9ttEUZYdLRXvY/Ri4+cBIIOLVyLjiX352Sl9u+PeK23ETKE
yj1D9gWnY4tKvt763pRKVtmKhPQ1JDHBMxLhgV4YvPJ63rpUe4NefRvuPPtJEApJEt/zZWrzGxQZ
KFJRYbdz049NTWthQconFkoASXtkiK6mO01ESVvJ7k11xWS2Y7S52f/y8ozyrpOwMnFa4dJmUJck
AQSfUBODRWKjvJrvHwT4Iv0kUhJwucJbqxk5G/W5vzFy5RsRxATOTJ9pOLIVMX6EeYxDYE/KwEM0
pjnLJuA58zfoiliQ1ruScRWgEwjjf17pw4i858mJuHLycWtYOnRvfW03oEYYWeEoMWhPsE4wVPVG
xxspDGFBsqKUk5P6M2t6bjyf7bu6RueSPO0sMp1loamyRSY8xGjOkNnVQ6hfbrIp9foDGhwSCXut
bOEx2HZzHe8v/Lu5HBshoHlm4byOJve8WTQkey3nR2ShfpBdYFzcXnqDK4qDX+yRsCOiwyc4VKPo
BWBo/ZYcb8qu/XITTudrlSk4MBmK+F6NPGqJ9zcXP/fqfxXAOXIHvui2TO8o5LJbg3CJRg2fXBed
3DzMOFCDkz05Ks7OjiAN7bwTT2FN3BWKjEL7WnqYMd3LpdwX+5k/1OBMO1yJQeJMO22M1pXunyxS
YByG/h5GdsFzYF6m9H9M0KWECmhSZ6wNSS9oVY+obhWPMX9s7sSW69ko0GhIPiVtarncemIH53Gx
jBLTXPhrxUNMLxIpCGEMiW62QgEA0G9n5WnhsUWum/CE6hxOa6xOdgnCY5fvb+ByjxX5BEx9rWhE
oGtLdJKYKuAXAJ2eEQx5sU1EB7xOw+57dL1a8dWCksXMQs+T0CXrSac3XAP+blcl+Kg03vJlTIoj
tvwUb2QP0GPX4lg0nx7YjZzxmYh4pe1P4zfUaU8Z42wscIRxN4l9l4LI/RCRqBXellMFp7kqe7Gy
1gJ+M9dYtWpwMFC/7MyPyohcUNb5t96F/8Eige7j6ZKBjBjsUx2HraaDBrN4ama0KuNIqRy03ina
i8kyO6NOGk9J/FmnCCCoxmKhYsSfdW5vmE8+6KeTDgEs0Ob2asJrFf0LQMPqKzK2WKI52Q577BYT
9nV8waUJt4kI7OOhwWHITWYz8dI3JYfnHHWcfZdKzfc1MzYcbMinwTz/qGdSxyinct1OhmbU9Lzh
/dGSEMPp3S9EDGBLMP04qd9Bth2apJqBh18J2t1YVeoXqDJtetHeYBy0+mmZa68Cx/8tZel7o7ti
qOyTwM7s9eeH+Ws6IdH6hBJOFCbiSobRlcAhF/k14uuOzI59YNOAYk/+JlZ8+kNFukjPB9hT2FpM
FlcvbB6WaeWQHXnBqa9oKeYZUQb+QYwxGiv1LACVuhxrMeOHFlcSDxaNOa2yqMR2dWpOxXIPnAu6
bxwEkumZQ4K6V7ABRQi9COw7+Gfz9dGYeawR5g0k77tzUwksrAXT7miN5W1jbtB6CllKo4uj+AsZ
KflvplrHRYHRfT4nX3T06OnngfRCKJN14jipjPzpM0S4HEIO3tcn8HsMenFBPkKWzJqTmI/K3Z3B
GnvDuVraOSQGrqIaVmk3+9QkOy3b741xygGLSSfX4NlMJxjwTo/y9gq1JNbRs4yG8oVrtvyjSWBC
Uc0humlAC6gM1qe02gTlc0PHqgSAVuYE2SV4PPrnncLpgsVcWY95Xr+BupSjalX8fBd5GErlqyOE
G7s9Z/XhxyW3QWi2mn0eyL724OALwMx/A2moOrrPFvNnaxb4FEuuT6M4fsKrd27kDia3vP39AzMn
uisez5ksUQqAfk964oIEAnQz+oMzd6hECVe7ajCJP2MGGim/VRaCHVy4aKHO7kHxszUWe53f7GiM
IiZrL+dumDul5pYon0KV18RI4lI4/mEMqooA1GWUW9rmro74dSXfk0KTCoAsrHjVM528wlqjHXsT
Nvg8Iebv9+iI5OZpIUT7fX6QJlspILTbUVqt1ZzGh9IG9Thrt53IPcPoDHac8ckDo2jNjKzU3nW9
YbbzWq0eXbTV/bcFiPuG+to5DfemTV+ysBG6PEpWxq79BU2H2RDUBHLzC/MedVF5ZAxXI7F7B7ks
kE11GUrszKzMBIPAssZestPWBvJ25eTNXI/AV4SmbzW/zcrQjy6ZF/I27g5o4SXfK65kmjT+BTU0
fg4m8qpBlegMNMsk3W6YbynJjCo+Cp4YA4n89sYoCaM+RNbVa9xvlw+78Gp5ZoebwDAAoEu/GpQe
Gzv3gfbJuZirKTm6QP8jETjPKx/8nHsUVfGpaVAOHMvrDOEmswKG5ZU1D3dyjTxKocM6BCnVuD+Y
gNwsSbvQ+B1y639kwv/N2tMdciXAsvbjutnpSukauyYfdUNFlVRUAYgrY2qPUltguO4d+pIpxLYJ
dgs9sbt5yz6ZoXvUoiwJG0EtV0AFjLexn0g3AL7VEPKEOmnClRmdCldICiMWcbz/nBo6zQI5HPRH
dEd4Zdo2lWpA0EDRFsRBhudnvKT+62utQ3rpBa73dt8fsc0Qn9/RDkGk0X/TR9kAlJyI8c1ZNuPO
So327VPknLxMt4X9a9HLKjILlm126gzajC+Q+sDKTubTgBzO2x8de5rRZjvY9lqvwXxUFbrhiWuI
cgKzTrOePHAGp8not+eNj+L+Gn7cQOV0BV4uZZt4VPNIKR8Sg7v1PHSF/Ibf+HkkAtkwRinxvebn
fOjCj0wdVvculw7Wy3fijKtG80kQ/Z6KIAaowX8lLQPMWVmYi4+ZVcBQLLfN/L/4xN2OMGC5jbp5
P4ptx1hT9X9qxI3XTBGRcZmpGC9XPZ+bxCFQiTyaxG7xb+jljNZQy+3XBDBn6m8Ea16mCK42GRJf
SbRWSYX/1hS7w5Jl5iN48OgnP1H9ZmdThPCgRCjUC/3RIMki60PIIPtgwL6vhYTUBcvG2BBMDZn8
To2Hy5KGEiofKkh/syGsXCbg6VCxo3/heMtVmZ1ZFzt09/lFL/9w1LO7B82aoQt6CQivwfSHeEWx
SoAGRgENJ9egxEHV0eOoSrGnGkoXWnFrk9mNuOKnoD9cDO82jURfeLpjHMFopUahYjW0AxTB3Mtv
WbL/WEFXYaH/LKeR81yB0Yu4kwZX5LZw4OLsXrHmyzV0k/CXrYX4H2+Li4h6FfaJXAHO1pr613fR
dA/aOTgOtpJRYWOlkDKkFk5bLTwTyP/lh8FXsXThbMh3VyTKv4hD2uYvF2Fe5AaezTUuNv/HsyJD
pV0flqNWyj/85+xZ9wkTHcP4OMoaffe24s9m1T6htQendDfOGMCUvHtUuXOQoYR6ZI4WiX6KPlEg
zP/GVFuIxVYlubfzhIVSuk5mC3HX5yce2Rx9jNDoqXzmNmUk25KFPg0LdQq8uF982YbbVN0NP8j8
m/aqFwiNxCpl63dyiCuUrXvT6AISffFmSB4Z86bPhTOaE6X60phL4pKn2s6YXvjBStwAKDma1cPX
xGvnJuCph6En3Bt5BYPuiUFf6Qk8PTyZYVatdQYK4fEh9ccCc7+YYeJuxQ1BVsJlNrLSqcPkuzxM
wwsTHtWrDowgxBVaNKqwoa+zZWpQA9p0ouWDpqIrPApgymjFAIg8SFgw+EQ+sFwk/de//B3A2aIe
2gYWcehpnyF3db9WlI9HMiiz0Fw/Xu4miOElGwnKGuQXK4v++wK7xrV21M4uACLnRoJqWZ4EzoSF
wLVM27OIDFFL0HEHWLY+y16jX9Fn6rK9ALYsHO6ThEv6mWLSTzPuPm9Wf4QdvRJaJ9vvfvcpUHrT
DpjUbzmwPBoVoXa5s7cf42bNuC8W4Ve8uMwHYCaeHUv8XA3qT49beyceKqTw2GqMqthaLx1aHE67
Vvu3kr5uu4Hlw5Lb1TyKXdW05yJ9rU23yAE8gzRJmDk6cu265Dn5JroTWV7UHmOPiV95dflAwXvl
kZBATPrE3whiTu39592K4WbueFq7cYY86Zwd9oG5628xySikwinNZVEeYSPQs7YseXkqL/qq2S+G
ojIN3vhlr8pf8/2nhdAtCvewCzZfHPk3lx5hFmbPtQgqTd0NbZUsAN1IrPXOBAHTQ59hR02NlHs0
m9QDVCA5EaB1gNg+yt4VGyJ6Klif6+DzhMGu3ZO8FJf3+6p+U7GUvLmZcNH63m0Trz2gPEHWhFB0
WU1xm72r87PnDFI1K+OGsj1QPzSQszVDKmNHaBUyTcO4Qsg+06CB3g8fL0sT9GyzqzT3Rw/ik/13
mZcSWradcYSECcCqSPEgiX/3WlD5tPxglyJ6hiUjVSvVEzW97MdFOw82D+HxjSkvKMSpkhC1a3VR
GTil/8aDouhRY8+WT1AkhGRwNR+FY1NKG+Oa5AIl3Ypk7KD+MkIjO9DXfMNG8E3JypdbYFdEIqYd
3r8xrM9/p/n0iSf8or4eHNzGrfrBepZrnQ7Z1vAopp9Vqg1ajAM8J4qSb+3l0xnqzsct4C91J1dc
ufqsg26dvDz4Jp+xqCNXNyeHUbdAX/Zmaorr1sJN0ptwLGYcqsUL3RgMpNxDruJsc0QGG2AL8ug6
HDDqdLD2G1oKK4OS20D+Uk0S2TS8kYzJgr6unEjllDQFa8TrMVpkTutywWBlog34Gv3J4ymQxBk9
2DqeKK0A2gA9huuG1u5Y+9zIT7LD0soLY61q1ugSdORRObbUmjhiIxV0ZTI1/o5sl1P42/Hadoq6
KJKIryHlOiUUMrl3wNTaumECWi9ca7diRe73eFr3/UWaUUcpe3HmTDvpIfJ0vi4KhMR4fAX/jUg/
3lUOGfzZ55esgEMwVLZjqs3B8mjtQs4BCDBJQbWqBV/eU2WEmsjSyVnVWnNsEr/HrprtH+aqZnf3
dx0DruNj1GTdJN01wiB7m1MINdKxnGimkbR6N75MnHwM/qRvMigVDww1aSwSRVIS+oYw2LEec0nA
vJ3jwtnKP8t68C3phfyaESfjj4xyBxkuf5q5Ipgj/fzmFca9iWza36ExdgDJiRtwqc6FJITJiY6i
x2a2vSiw/sfa4nVVz5DDYDWOAQXhB8I96qLdqX2ULeAuF6MNSrKytkpPnXSln/vq0BNu67QdKNon
N+nWWLjvlbioX2qhswcgP7JMPGieIIfe/6HEEkttJs8RNk8W1Uj1goIE0H1OfweObjDmE8Z9MVwC
4JQ1xBXxRdG+/y7fc8Rh9JksYKhfi7kOebCkBYbkG6/xh+gGOvKp30UxO7hCqtwAU0MKjkiieBjY
+xG3dKqvs4VmYsS/91rhWMMJ8OkTEFf639eOUgAH07H221jgfS3X0R32VgcsXcS227ITB5i9twxF
NHRtld5ctXjj5dPPpm64T1RcHIy5jfIg0YCMp0DR4ilD6Nfu7oWrcQ7vs1IoAM2VmM4EqTe631yf
lvgGyxdAA7Q+6VlrjdHf74i34ZTO1MiWShk2whdZslpS71KpDzqMsr+RlZ+eW7CAt9yRwo5QKvSs
t3dCEUZsELxdvq/9a/VrfSDR5gxzRlatxDGnwx/PZLisvSr8DSvDiW/lC15mxKRlFLSjQDMmdDh0
cze7Dba/zyx/cCsIUzY5JPGYXW6a9wOLLXo+Z2nWKxuiIXzPOSrV+4LO6pw/gVCk6VEwtWcoJcni
r+U1t3xGQTTOBkeumLj1MKqwC9fSURlapD9gO/NzY8sRdvRWPjklkopr4CRHRop/ku2RgZEFWrAG
JNzWsCbrWeFDcIOCa1s550ZR+5YmDcsv3JcbnHJrBFSnMGRTWYfNemYlQuo7Zrt6qw2d1O+dNR0S
HEkgGAWoOCq/NMC6EHSjV9VndAt6tuG7/wQjJELxZR4CfnSwFcVjWGr4J3q02WhrVco9I/7ICNXn
dYjVHMae4Q/RQdZKmE4X5yAQv2wwsOvrHIzcyvr5gNhn1PYRSMpr+0Zw2gWVK74dx/wA2kCTZrE/
zubdmQrHGIdv6jojod+wWREp3dQ4cmclVP2r0LGDJfyvC0hdj3+G0Y6FqhpXTd8GP576WFW2cRX1
GEKRAG5fWRXw9aYhF5uNdTZmvfYmAdNdPP7G2pee9QIiHH592g7EOA2a3ocWtlhMLMbDpj2sZaSg
2XusEXm9i0LudfIgb0Ow9EUeEf3G1dLLGY9KH05+kSOTc3IX7rdsX6LKKsgPBMkD6AUNJgK68Dhk
q959PTXhA+1injjA8lzC1VuhsUg+CHSn+2HhSO3RHDyofNt8COfU6RcOpNSSbRffTwcLavJO2b/e
ZEPQa9DsJq43BuyZTE1iZxp/W5ZRZJR6dAzvs4y2w1Pg/FwmIuNXsLZlTXKhaAQjD+7OYKfZKClf
5DAbyTXz+xdcnZ08noz4AsL2sUHZn6VWLS7S8nOTiGSUJGV0px2/6cD9zj7QhGQujmiueCab+ohM
QWoDoMbbl8pahrPENbSBblA1OUReEGPhxfouYDZ+xMQywcfQsshUcTi139dEsR9jetAEqs0sjRJ5
NvxerSlrTPlFEsxP3ElV3aqAAu7DRFIWuEpKgmRazfYMulJ/4vttV01fDLBMd10MX2we3yuvguSe
hBKSmgJNTMVpNuB0lAm/mmZoRIw7KZDRnivBK+qibDf78w+OWZiVNEt8zzOmDD2qJBscp/Y/cPcQ
RDwHt3L1wyxMUlRRmaSuEyJ+xwKUgoH/Rqz1fsijhkJQ6sBdUSmml2GTF3SkGPWV+SZAmHkB28KA
cZ5YaLEKMkEdxTAlzGiBUIlIoTvIX6y/9Tc6x/qY1DSX8DQ2yQy0QWC0l59LDM5XYJZMc9jGv+Ld
0Me8xQuf+WPFaHoaV0IBdwagKzmxHwBCxHgyXjQIz73vJe7NU4Oz+781mV7gUrR1dv5LOojKP3lQ
STerS2bSgRiS4yigLedUP6CxsazGaZprJLD3qX66klVZF9FZ/AwB1Y8nH/RJRcm0839o9bd3VbK4
Ti9Hda7JXhfMsOeD0otVevv+auEC6OJE0QB9PokQXyvdQAvkpVCgXQxJJ3mkIcCXnyTkoqM721o0
t/SjLwIsk+39orSspu8MylR2SO8IEqWu7xibPs0w879ko+nk+dU3Dzbw3bOHDbE9UV9FH21AMrlJ
Ri5QbArHpq4gMOQN5NZes8PWCIYajC1XMlhqwMCMO6j/mWgtwdNKYL0UrQLNbqvKqt1Vcpk3v8k1
gQoBYEPxlQhURURGUgOMZMEwQbn6kbAcn0O8IgamuQ69GQxflhHW6oiAYjMqAkS7y4az6YOjqLkJ
HHoletRUkvAYvNTJdwVNvGFeJhFhuwYGP+zo6rJONWf/TzBIk9l/9o8mOYfqu4+SdRcGpa0bVR0a
FKPj89OjxkZxMYI800nqRdKwqoXiPfI23eCKbRgVTxGG6fmqI8SaRTvfCGqMKS32y8RRfCgFsCDa
84eh++xcKhT8d6jjvq9Cd1NCD4rc6d+L5W4ibHd0DXk3XyDnr5d49cJUf/KehCIGuEAmIA4D+oT2
YPnQy5Z3oum3ng/ycXnICHvQefJetVERyii1vCe5UbMaAFTTcH1u04Ql81PA5C734PFgQVG9a2eN
t5DJx2Yziik/GNbpMTCeb0mxP+0gTvz9EdJ+yfdTbHK72Qp1PB+G4g/jZ6qkpeBVesGtv3KZSiEq
jfZGdkS/26H6mIaOX9VCUxQShPVKJNwhwpTzVJ9kDX2T6c4XTkKoGNJnRFduTACRNgfpaLNGV+pV
Y3BP+sXgFrUPWmnrtQLOnfELW0+1EBcFLwG0IuHdU8B7zn5qXzQc5DdxpyHws0ssj/HdbiApJyzW
MkeHBT2UBY56TGo4T4BLgabDkyEoNPzZs4Zj1GA5u1Jk0kYe2gDpo6T61giw37nB89ZMp7i6woaH
+L8QKOAvTjkqJGVxQLu+R2LpFTQQgFLpStlMwJx0w4RwvexQR1qc2v4jI5oxhuRGA1VUHTwWKo/c
JcEIuyi9OqnfS9NIdKFhIWaKzU/5K+f6PNUFqgxfkfBE4QaQnW+6vvubmKqJaAZsuploxmbO7bHx
Y6j+tVnD9W7BpBkWUMDTzCPED3h8kMk+f0NIaIQ/5OQZT2J+VaBYAPZfszVwxqAZM0wv0uj+4bV6
tlMGgEOxbK/xnOXOihdTQ/tz2+dmSmu0hFkaBnKh8SMJfbMRbm+yJTpyqcMaK1lJuD9kUgb2MvPK
+ScxlHANpH74PUjaIHiSWkZ1gl+0lRSzj8+Jw4fZ0py4LzLYeI3OF+W4d21+lM13l4yZePq56XTl
LOOCr5pc0z+BIIJOS6IRHGNywN8EJ7LbPY6dSUkr4sZ6RUK5H3RWxAhqjSpmejTmSr06nKCCr/mO
Pi92JSItTfhiVvD8pOeabrhLpokzkQupsQs+GoNZLK/rjbxpljNz4Th2h9kF1nQiBY17bdiMML5q
UnuimkB/f/qm/rc2vY/f7NrxF0VAoVv782hAkmpRI/eaaLd2Cn0Vwa27E5vGrLzRm//1v16TYWU4
gvlpGB0cWM5A7lFuxWQ9TUzymph853dmUEY3796xXTwE8xZmMOUhogfKIsEq85yZkO+S+mvM91K0
dEFV7MgmpynY3AzAGsUeYOXO0vjxseLwtGNVndq/zq/AWp6jnJxa8ESmYGAdU5n9fvtAlSwYg4Df
rzVhEulhNe2i2L1k0UND0kCPGRyv0NbXPi9WBpnS7+ljPL908AKIsQk3LaIklqXauOO+lWeZ0Trh
Ywc0K0NWHMtj8svngJeFB5mgAV9sU5lbXh/Wa0zjNQas+HFbdy2vBbBCsx+cQj9t/XQIFC6Djbmo
CcJTg3c4x5K8I6uqPEA40/B9JzQ3Pzil724sZ8frlOKCdqMsLs+FWFAiGFG+PQrOif0fWKOYMzlZ
E47pe9q+LnBbtRze2GOwmiJVGEkF+4xjk0kLpT3EIa+KcTWpGM/lsVLH1k146b7qRPEZnZ+5QZ8x
u6A71XyM1+zOsHl64ttBTmBsv5VAfnSQANG3L08XNXeV/kZ+8fPLwacnSpZ6dHzhlPKI895Ue3AX
eD32YuM9oJv1KB5caT1MglDMwQlHATl1p7+p2UcTVbjyWj0KYPC6f1aictz4NViHQk4fWe3BsOK8
YSbOr2QMK6S8zzCJAyJx2udhbeKFwVwvqHA7mplqmoBQbZsrypSUucCco+tIu7fk3/zVNq6ZKKBz
14QxP5KmOX8BXVuco3Fcdt54QkcySCD/G/HGOqUmSRobfQdnnFOdXX2FceiRlkewoH8stha8056Y
JUrbAEqfzut69EB1NBRZ4EMNX0g2ZSijadFqm6HXrEfd/ihv66dwNpBQ8/EHW9MrWQRFKvwdmhl9
MRTFiaVxFKLMRRdCZTJBEY6eoP+HNKLwHyotJzmGPXHrYo7uW+htbjL/fbmixGhesYIWHYb9jn36
qLLV+rqWuHXyLq1nFKK7E8A1zmNDI6CnoNm3IXnU9IoRVcx1JS+mu/a87cO1ifgWHl6y9mOpeZjs
S0rKr6UO27gfFAGQ84yIVuPeO3spKZnQoPDWyfhFIGETmtAe4d3BI6z7k7QsPoJpZ/5ZeAY+olOB
gFf/9ZMXnXQSXpgVULQqkr1ek4GXyFi/fhBa9OVyaAtBwXZMfBMaaklEdu86IZ3aTSLB0W8s2hxM
796UDXN8O+FBjkx7+zFsuFoYB2G6s553daS9QeJ/eGj1xfi6vA80lIIhMrjv6rqwGJp2U950Ut8S
BW/cdUc67BLaFxRI5C4RNPPuoMGs1AuWSd2IsEXYDu1Q0b5IYL8I9aHRLxpxYN6w/q0Kd8pAj2fS
PZnui6puVjF4jhfA79oy+ejPguOYQzN1BqkpQhlXU5E5BIQWBX4Ayw7/UPMteg5uTWO7Q3WbTlX1
7+PCcfz4cKnFc1oVM1rKRPOcihNFdBwaGUzxJBSrSL6HOepbrDXMugC2LJsBelqXSMX0D1Mxp/fK
NvFTuk/EnKeoZVlLU9BdFnUSIWlzdYSgFncse5H57jyjCXtFcOSgVfI6YRtGfbfPOdvTERWmcRIo
OA3oFnryf1J4v957a2IUfY+rItcEbmV08qypybnRQ5Uvc5YTXxm8pLjYTfFq5Jayulja1q4Kl3U5
UkRpinyocR0JRtuHO+yMTXFFn1jAZL+r7q52CWbtYP6DLI7aPr30YvZUpxaALNbu0IFyFiQ0zdHx
YnEU8IDbxXi1IK7/Z2+YQDtBKVyxBgC/hCg+NJyPgkqIa4S8Co7/qee0uYqTmS5HMMLfjw+o0Z3Q
dfBx0juJmAlpMLkF7W7rb5gBEmg0lii5fSkk7feZXPgSbOWdm0kz0l7vIjUsHRpkmhNK3Oft/r7n
TrOnhlZJqzlI1PI1q8EtPATPSFQ+0gF1y7iJ7nPvL6C/SxxC1fFfP4YZ2CEjJ00k6UT554J24LQD
WCIIeqBhxC0A/4jgeVg2SKeuPvLcdS7/SbMQdchlNWsE1d0nzXfFw+fM/C/k2Ew780dutyuiunRD
1i6gdXN8CWOumYeu5RXGbG1I54fdTm/xExWGS6knt7zjZaz0HnSrgy/8noMj1cqdclukERufRG0m
EGqVcdJUY+dVgQQ+foPSDGusnY7E02/vyc2EVc+eGL5H4BKDvUB4WthjHb4SR/B+cCYzEofIvUsj
ia2EBT6EhTvzDm5grBXom+7EiBJmtImXUmftc2lehH1GpKX21B6s+FN/QsBO86lplAeWeGE3lvkF
+g2yh2mAO2+56o7C+lUNktQ7/hohAy7OYAUtXgZCuOKpuIKzookC16Uc9dt61Aik4Po4iuXuLM4Y
RVYHhabK8bs8ZBbYJLoYoLgleMzs+U+v/xrARH2i/pfJGTgl4Dg0HDugdx1P47m44me5J3IbAVc5
Wx2H7h+CSis9LObJFBN3qM2sWRPDACaSILjnkJYzN6d7zn6C1NA8wA6psFqy0K/1uw/JuH25xWW2
ay4zZOlWDU/m7e4GSILXEPY6TY8ItdUm1lvPz39sGxYdM7RPu9peyZCOIPBI6vbDJk67DDNEVn/r
fkf66eigSRtTnwAK6/KPcwOUG140SyR4H/sxEZA9KIpXaqwc6nulY7vhHCAgz5ujngdXz+vuOJdG
tsnuoYJmi9Q92BY8ZQhw2xnTCSCs1XCwNp4hSQXfBs8y6T/tKePPn71pSTOa4XeifaiLt76wIljW
k83X9l75iZPRLz37rfXpW6V0p2XBfRq3C6AvdjnNUwDffXrc8NKodhtu9sFFB+YUX75lTrgVt5og
Hc4ElIrvGlUVo8QIHAm2TFSFr81sJhtXMyaty6SOzaFpOaOURbOuqqoegk2GromZr56W+Rda7ZQ9
O+1skVoysTI2uGEz8MBPW7JHwTPN8sdPuDkZ8YC7HOo9t8KGyV1lJhrx5xh/EGC0bUrNKHfGZ3X+
g4PtQbRAJ2l6uqNMBIqUk+ITmosj7gchU1ChhU032mGzIVP3Tto7s4LEQdqL/18BTqsfTvVMtiuw
bwmD8arrdK1mQtzXZmkOkb9k5NufiX+ATdI5PgFJtuFzR1l5VzFh84gkBm2EsPkftuNuWWZ8E21U
HTQnK0ZYiNxOCVPj740HNGT8WeHThhVbHsDew7k3raLoREWkcqrRc73WNFsqvvu5j3P+afyNl2M1
81NHwtdvRHIeX0qbPcX2sSwuI1BAJ/f+fLSQS8Lhy6L6OpSsqck2Qm7BCCGdSnCJUbp/vxgzEOg9
OoVLnFPjP7h8dbY5XlBXUJ1EMBh1+pZsbqrv94t6c3/vnGDtktWkb+IAOoobMIYOm2AvqHUFjbD/
OrEIMZVtWzs7tr5FQH3ygdvEGk5Uspkdzd9DuG7rW1p6ZbM4Vk9+GwdEZv94ojbQTR6Rs1/ylte8
rCTgTfMNje40ddur1QPVQftuz5XBtOy9OtDaQKDa1ZvMOn47fLQ2xprYfRibrPteyVpyDTzK/KjA
FfkooR/qIggG9/2/ULpBu76d6xjTYPXMGVB7oOrQpgPlTQ8OvUYBZBROFMdxc0v+IAF7+JnLrZN1
rtQXp1neSyHheADm2a/9Wj9vZQ/ENXYqy4zJEfurYyPJMtWTy1QOOnMom7tlyynR7UGJPArr55To
64TzueGFlOQZj0uJTYDO2Olmhrb9R+ZpeLV7av49BRg6FplogiEBOoSFwtAIxWjN5XQ8HBtzY/qA
tm1+AH7yHpF2efyp2jGxTHJ0Qz0/uyb767Yzm2H35NHN7tu8327C/mzKkoabD5/8PbGPAHAigpBM
gcbu9yQaG1eughSySCjL92yDwZuVYocYtcS/02GeZGM8IT9KYKrS33pb2iMciKP9XBb8hCS/genO
gVCUKTFMdKg4QL5MB5bdzMVc//8AgJQ0elznNepbvbwYg5qxK07X34pnVPgZY6kfng2mTKXIdBbf
cSomIySacdJjJAnsDRnKbu9QN8F4DaB6QumjCRu8qoK4If3VR8+rmhR+feX+Om0GC7UuxJbrAx5P
JnQkxahtBUXHYyUrdOg41N9kQnMpYsv5CJk1fW+LHCJBCRpbxb5OuMYwrmFBXumg+0/CXurZPRPv
Xg5Jc76mg4scM3omcQ/mq4WW7EGbbBXwOkgap67qkr9ntrVdoQJkb7nC3ueaLiC/2jA2xrCAL2Sh
f7KuS/PuZf8EiwUXHezB2LhyDeJ1NYGjGhE5Puu0gcQ0tdObVCjCdY6lnlMI3Ck0ZygrqOn9MuLD
vQpFS96PynpjgbTLKU7ntHZw8vQNFZGLnSpheGJCI7duvhDlD7QJGkmd0NWDuz77Lzcltv41IEMF
ua0nd8vOhiERJXKdAHl2b/mD1356KuofHDvISq8SzjbksEAdjIpRCVcJLbQsRqcpbrwaONbqiyHD
/OKrB/hqzs75eyUno9XXvdFtboSvYdnnwS2t4t+8113ot/qX/GgfRW6TK8+tRAn5ETMZDeMHnDEy
tVxTd2ipiGpwYFb8IviJp0qQIBGhTie8kMY2VjWkETYqJe5B9u5OnsCiOjT+JQK0cm8Nez2xzxJ3
iygeJq/oHOYrjxJLTixB8eD+Yr/gQey6TbVj7oqghK7jU9u+CKEFaWmK7Z1FWq4JapjcgdBBrvW3
xRgqVdRbECCBiO7yF6CcbF9qtSmz1w2jrcEw/SgWArXtDnfJ2eMcB7K97OtsjiHZYTdTMAD8tC33
W4nLHzk/bzWiawfDZw/AbkBLav+KdJ+l9NPDhRHGrqF5vvC+iopGdfSaeF8gOIQgOqpcd8E3kUWq
1mFT2e9G2TihOVUg1OmjS44tXkFkGinu84kivquI6A4N3j4xi5YZxkkx3Dhan+rEod3Sgke5xGDu
CMAUk9oHppLUY7v/ryFbhEX4QUeiewPMYwby15kWyP7VnYOqDBOJNaO2V744dQxCWTmAaboMMzBS
uu54WgTuBQicbfj2WgviHvk6309/cqcDP1Jedyxl0IxPMu56yOP8ZheasEABNnQ5VxQpRBbz23ai
mctS1aJhjC8ji6tihzTlxoNSLmtEBumnSrX54esplw4CQUYWY8yhqoOrbYnnRjbgGGKHcFidLITn
oOspQfQ1OiWK07zGUSnWJc5mYjFLEB4X1EPH/cnAiDC7nzniCuf+AQ1M34FSQA6iSwDqjKLvrU/N
nmVuAOpMPrNbNggxZDJ35M+ojN8GfowzbJ1d9sMyCGUk9Pgp+DqmKMEvR4gaOAoyGdBbBja0VB6K
2kPse3vZ4KVMEG6m324c99a6RZXtZWIMsVkl8J0Ec5aTwfenwdCK/4iCYdb0PS1f1xZBjdrllOtK
/HklJUhKBd+Wj/p8bHBY9S9oQgI1OJ2zEamwvjBgAL9vdUytPpcq1HAsBG9ulRD4lQnXNcq1tswN
OvAkz5FqxDGzlmmP+KRU4E4RMnpGM0VTmspVDfLUQCcTWnZlJ8NbP4Fnk+0fVbagAEt9olwFVzqV
saoufhucp5rSmCdv8isszNZy05TfbF3/PO3e3mqLYtD2BxuJgoiuSaaXh2dIh+7+7x1iN5Li+HPQ
EAW5UT/HqWe+IgT0PZLKEU6xlOpbDLWB3vEFijMvw8YPMZyX84hXX0daMioHbEhBLGTRvXHsGpgY
DiErwB482Z7IsyAdTwDDO8lYIxUDHAl8ZtVokZHv3sjkVHcl9Q6lxIvbvIiyVnv5DS21rScMn2e3
TR9HxW4t88lOaaBcU6X0fWHRnmrAkxQJm0UECADbPyyTxAVcIl7lNGG/LF7mTKKSzQQQBY210yOa
meb12Tr+LP9lYpEKI9GBTWaB40TEGqhNuaCkSt6ceAjO5J6yBlL5+cFQuqgqthpoNlE1I62JMw5y
LjkUWTJHxae57rpYFA9pK8z8rOR2Tu8qSJw7Uha+dlz7UX9oODYejqDikqKu3yvVwV93kLHnO2vZ
UqUTcOczQ4gIXBX/bippmV/8w9WKCSt1SY94HIsZvs4q5xLCWEVwsn7asRDT1FNlHa46RAJSTFEU
nyMwh2hxXehGvFO1BH7yKW6sRDJQc/mkKbHasVMOxfYTinMNiWa2SEDT01HFV7k2I1S5pF35ZhsZ
5WUyvPZvsMAi0XlrTX0M1YA/AnxNSzcKQxaf7MMWmFR2QZ/YoJiL6YeuOvGkP1+LEXQp0uvmDwzS
bWwoHnBp11mkWhc1kWzZf3FpyUHn6SR0dTtOA2HuPDqWuAzRYwL8Islb6nuTzr07JaMJ5IwfvHEv
ZkJaIMDu/sBYr4LZxcHoSQbhrqxUi/TUX6aA3uppMTiyUE1y7LtNjFhBxTEBD8ZtPozdRW1J1hVh
gEUCb/aiwFz8bUtxYypnslJmDYR4ERsVjUUoUA+74KmDIB65n8+YFzeNVb1oVZtrWnP7oZJcRTY1
I863NV0qEVfOdtln3r++wuaNEepePW3NbPD6IuxiPjztIlwAwW5XelQpZUP6+4p0LBxBzzj2PSsI
AH6guIjeLsvh9z4YwIOX5vRjircdFh+/TGMdW3afKlPN7b9wCXirnkrMFopdY7veTWMn61q+Lbb8
pU0OYorYc1YtsfUgf/iqOecYaSCJ9MMl7v4ItsLFVCTpib+xlUFVJ1WJ8JEcLRofQk44D4XUcvmW
63IIwFhmpHQL4yJdZgiuO3EgtAD0AiNTnkNomMbrmxcHOBFWIyaTn2t9izq/xdxqldJmRgyETC8b
OC79xjj6+qouCLWJD49LSSFYkBNLT7SXFPLTbmB/kq5EqquvfLnp9MalKDX8u4gsf0woleMqnxr0
80rApyk9SnEcc0kKEheAR9uZgAmq5yeK/ou1tmkPcHBAmMRPBWd7dJGt1lR1JsxQwv8ed5BQu9Zn
WpVPFhvAI3g4sy3L1LrVML2uYJ3IuqX6S9SkZGi5BPaqA2NPuPelf0H5JXqkjNR2n0yvYiXmbKh1
lrlfJIuiJ+A6SkVulhWl7Lsy0vLUBoxocQZTFkkKKHJFtE92K2Y0IpbCsmcioIj3FBVdDoGNWEhQ
F+wlyZ/8HeyprpS9krcZr2ESvjLg6nBWfPqYP9UvcObLNzL908JYBZG9kfL3Y5LKrUF/AhE0Ora4
ql+56v/Q3nQlysDxMo+CGGXdQuS1TsBIZkAw2LwRVM7WUCuF7LTPWixjPSC/oM+3l1r8NQU1zuc5
nQDEKHQix1PmZxXaHwlY1NRYiSHtni6LdHBXF0J5wK3KUb26n2vf55mQBAdeQVh5yrusImo5U/Nb
rZhKm6zmx/boVLbkSyevek6hBJJxjXdmh9vpr858WZjiCEQB3opAVgjobd5uHnbRE11w4OJrzcrs
MmRp3Hh7jnXpAdTarrfj5O4nCDAD/3A9zWTtSeXPbSZHYxet8XYzik1qlgH3/M6zkXjkSvffOEzE
jPdGXpaiGFce9vaRU8HGTWGyqHASRgueL6M+VIrw9WVKeDz2BfQzF4ilmt7myoxkRmh21Yz0BZ/8
uC7SwXtXG1WvHML9fhYjuApY9a2SIESHLZ2Laq2qvlbA7rhvTpNtCyHCVZ1No/P7tbxIS1G5XOqN
Bd/PlS3CNEjc/A94OG1dHAMcHTjCgLVx3WMJ3gBnwprt3bnpkvOppDcdoP44o8KrxCu3iDppJszj
jTJ2bklKzs+Cr/iQkUKIME/RLetNDvVRVLaVAT28a2ckaa802RzS8INl9ZnXaoWFtZRCS5qAkv0p
qVQYWrZycb8Befi8keMl2oKVRWI/t8Vo4ozdYoiGKYN00i3jOgZU3gN9xdvW62VFMGmgv4+3J4Ou
Ln5fNkfGLbyCEtk/isC3eVTwonoJvaGtfei20dVCgjYA0REEvvaCeMTgwKyb3ObOMHgW9Lvxm4SO
66+Jx4Tk+qREDzD0iJDmFnJksaHBv+6m70J6Hv83IUcStRhnJrC6vUMmoSCgMFyGqKvjokwuJdLd
xtZtIdsgNhTKQb6bVwDVkQsW/b7jWn5D+xKdipPrj332cXymNsMDYYsuJK9v5guQBfQ+I1Alk3wd
zdoLFJjxxQcCzjDu6bfMseV9giZL5LD2TwifuQ4UQWLijT2qiVPEl/2kNRtnR2Yn0+XGNnddYIS0
fE8MTCAh9eDAm6qqYMk8l5Uv1YzMVTzKh6QaxOqywf+TyszikE4ec1t5gYBYeSJDyHFOOlEiWH1N
nHu9Z8e9cAsk4mOSF4/XL04fyWs4ScdStzPD80m9Jk9YeFyq3JVxNo1HUxf84VGWvX9dHLJonFPN
7JxpFxDkjqrwbiA5tDpPM1+LTdDyg0m6JqE+6gp88wcXZvi8Gnq4D7/jKl3mXJVQn2Szw9iSKcp5
boZQibGiO/knr2rEW/m6/GEyOsdBvhMlgFetlbSDpeQ52pcHWbR3qlXcDe7ih5o6v9onxrIFQglU
9AyDXaCeCJ1ooi9ODhAuXnNFtvRynPs3vRK9sC1px8gBMef71A5REETRfcPMdrq+BZNQzDNZS4xl
BqsDE61v5DQOV026hwCbfOASRADuuEeki66sVMy5HXEWC0lmcqcxgikzZXlYFsSwthD8NMtdv9a7
jM86NNYv+5eGxruqncrOm/p6iINAAoKHojbWnk9IUlKMVMRepsIfXKr4R30z9TXcx0Oa00A/dKRX
m3v80YaZGPaf8DGnhPQaDB2ZBiheRwg/fRhoshFCFtTjoFGed2167HIiIQHzCz8Iqux0OJsdiuqt
EV6rq1SbAoqa7o9FZ4SGx4nYxtMaV8ERGhD3wV2039jPrhrpK9ayfY9AU040OJ/YSu3xCGhNTxw8
Aoh8p0vFNehXcMMjW77klC+Ey0P3Hl9o/XISuFqleFNkWSefCZutLsLGirZWJkEkUlryRlzVC8FV
G2+lhCAV2t3eRAEsAyPIy8UEL22B42Zz9pUkJB+tyWznZQrBtKUdaitQP4GVn1taKPc6H2i4BGrd
ZDI+fi49N8joGsNrGC3qaLml3XBxIF4Z9c/YTJxlbaAVffC0cTzUZORgYYkblJp4SUlGtQvY0Mfl
4so9JiuzluZfXK4KhOr/3cKnUq44UhIlfUFFrppNLTOiaKdiJqQCkKJAiAKlwMhN0z2NLc1fUcVd
4gLfttfSq6qgPY+zme+d3jDGnKWdr9qT1H6hr3ww8P5shvuSHzweCmk3Rgb/UuN9QyUbClOjHbAe
sIuMgDZw70bAUfzCPsT56f6o1u7RJ70BCH79nzrHsIZwANhy/d4lK/amUi7a7ihz6JUN/6bC/qCm
cCGZEISxwggnwJ7SigCMAc3hGMMFWBSakyS5QbCW3D0CNSOlO+RWcrAwdzF9IkIhrDUTuHqpjfv/
lu/XV+kN01WmmpJclYnpZBWX7BzS/LcO9E4N6lSNmF61cZ7g9sr/6T3mYE9kow4wUy0aeiokLJxW
lJv7hR49+xbJiKNkZfHG7GTIN8cV4zrLeeMjn/Uk3KTIj2kih1clENghKcp/xsPvnNYwfLbbF65y
ZJJELSVIiuMpPR+aNYp06A1slAm3s/NWkgTYnJCOlqJg/KjIU/5VhbZtSrxa1wS6sM1fVMBLV0tZ
ikfYbUpKqN5LEJCX2/ndHBaXC8TPqhGq1fK/SJw3qSysQq4LHQ2gI7jjp6Wuj+9US4H6M9ICicqw
ReP57yKHP3n3LNuBlo1CFVCRWVHFRtN1Auki7ckajVYd9EuK+lrZf7mqkhoKxhnJExtg4To6h5HC
6mxAU+DRVCi9Ux79a2cglwBwLDZJJ+Df1Zw1GNF7CGXlFEc28tucnwXVrsiy8BZe1hhy56/JYzg4
ZtRKo4URNxqaoxJX40KU56lEYyy0aAnVsV27yfKBOYMzxkwdxHGMSSruKg0ZOu1ONdG5Ax274lIX
vdbUsNrgZi4Cxji289u9Cpc0onfEL0ryhfgn7auHKovWM0GaF2zJB8fiuqdJL/MmyRUsTduVsICu
wfS7YqurByeNm2Tpk3/kd/71qhKjFl8/UjmAdIauHwFufveRG7gmFUUuOrsyWMze6KM/AKak6H+P
TNqEXeeSHMyvP+Q6PUoo6rzMk86V0OwDTpyf41RDurff8FvIQydMg6XYJnHV9C3hKVOn5FUq9f4y
J49Q0ibZ9Dr5Dj4Y9hV8QAKfYciy6c85xgrAA+Xs0KgAWY5N3zJlUQAWX0yOfsv065BQzCNqb5MF
DRwyG/UfDc2mvNGkshg4RRXTu+8SpI8VQveHRFPJNCmrDCm7qgTveddM6TsZ6C554aFFy0ZyalBS
y5qOnykANenESzAWdGYet1Tpx/wOBMfo8sUx6XFCtvUTCp4zhac0MCcQz0fxQtTh5AeIR7THYGQF
UrVSDP3XpgnKcRunEaxI+G6MYTYN0wLxho+OpXgQvN9y17k/oiRU4wL2nZJS1XkiM1uzxcb2Sz/Z
SMInQYA61S7AxMkenwz3XJ4FnM2F9Cr4KctNS39TDT2Q6Kwwx/JgMX+rAa14Jk/ap1CHp20ofhHx
6xbaydUsJsL0qYzekpM+ksg2n5oa1xs3fWTngczMPla0F8l20FohGTr+A4+WAmw8ZIU0V4AnjGjI
7b16kSVezqVsX6tOvo7ujhLFTkHckhfidNjHjKSo67L9TOMwwhCJSiA3TY1CK+R9eiN9gDyZ/gs8
2LtLaB2Ggi2qYZ/h2Z+2pbxD8U116fKlSkxXtfcCis/WbfpbU46JHXQYfJWnO6CWhg72O9TVSDUR
4Iq3NEp6ujDbvq6gdW1Kgo655MKiF+DlZIfkG9a/ZneU4E+EVZcP7QheGk4OGPrfT7OAIscZplHc
NQSJQQsGESfbigx1h9Xf8uhJn3stX+WT/keiQKrlNm2Hl7iCNTTkbL6ZAC7q5aNsXLtJ4O7YkUnM
0MoNMJbICCzJa4Nsjk/KqSkjU/8Ns5/WI4IGfvJbFeXka+US1nOjka42QolZIyKFsdI/GHuU79v6
AjQNGr9Gw3rsCeLepFvNUgLmn2y165fnQLwBIeE4JktUnBxsOOuAkRX8HRoEW4ANAy1kB5amz/m1
Kr8FewWxI6xwglBu+3XKNMe2yAu3bDHSsdLt2uSC5fdNGT04OB/c4oZRM2AEu7ls3LZV0fi3FzOK
Rz3dQHOLqE5fIlcq5TmU09pd/uQdJl7QtpiehOnxbB5n/7/baeZu8QUgQd/kjuTxZND0H79OMuTm
Df1/hf6DVbG3ZaOpisokjbzeXSWcYOuhf9zLqr81DJMoZSBt7T9wpb0oPdQ/ctI4jTB4S2BqlFGy
lbV6eySzSod3+NiNphOyTfzNpV0cVHT104gpCmqjNX+iKbfnjWb+zhvHQdkLbgjhG368hLBGo42F
p/pjvPvPDCCcF9tg60243Uu//UgVvmkfBIiyXGkeghNZ45HYhlUx2VnOLlb1rXZxqOGr+ea78ISP
rd0P2wfJs+82SJkudDK5doQ2PONoz25F7eHZK0bBQsLe7khY7l0SbxDRxpPvsXbZ2yUr/ZeHT7zr
qesFa3b4QEobYVv0/sBx+70qQwPcSai3Ewz7HicrFaIjLaWKIlfP9TTsAEE7E4lEXGTp5h3ZeAHl
7jErIM0h74n+tHVdhckX1i99doX7OEwhl2buqPJsaGbGAJUdJ3ifg8N1u1Z+u0KrmSjhmDsdYmtB
4j8l7GiaZH2aeDIQB2rCChBLbD13Tj3XUvuD9TAB1nm89sbVeq8X6JsG3carkaYAMCN+qrbP+BmW
wVEEvavD4rYTmQTd4goQLnKgdZHZpINSBnUmRopU6E6BY2/+7A+itHHwfRVjGX4R2Gw+pOR5YYLT
0OgsK3g7g7fkInZjE3LY1wWzF90GFiD+t2KXqJw5VPtNn93sh86+nEKDtVvJRn9bpiFt3y4ER8p+
iZaY57gE/BjLley3RzVHCpCRgCgcCm9GDItq7UzkK3zeqzr0e96IXiQZaqsDrC2QgKNvgds+K0sQ
a5jCU6vpF3OssWoiyhXWLVO01CgtRXyvQqOwceW6NpPXIAb6B/nkTfq/eZIrRny+amvC8jfcx0zy
hkUacGN7OTUKXBS7SODHA4me5UFhmNti09nlkDUfnAymB7DausmircWzxA9dcQoXyGmPX6iDWAiN
zCCBr2WULvZObbFXZnUg2R1wnOibrf6DbyEORyHgw5ChHKeyo4N5DT6qwyoeDa/WBm6SIyjnyDkD
+bDEZXmvOCVRpb3QRHIYQ57iLuZy8fXk1bf58H33K57MgFSbqtVE8xFNZuKDMEckWpzExkHwacV0
DDiwKMw+rSdwpgtDkydwtEF5kCTmU9HeLyE4Nn6twgesekZuk9TsBCINMhq1OV/vi5a4tdRNA/wl
2l42oPBKt/P80Tv1A7F6nDM2zxelYD4f+3N+qm9uKfS9d5oCIraTbwjBA8r3ypD0f8XBb9MxonMF
8pYtsebUwqpLqtAoxDT+XqGHvklHQVH7LQ5DAQrB+QcsrUsN8YFTs5TGe210Y0RqOU07gYgP3Lyl
tNeEyg8CvmLqUnRdSNRVzGVVxc4LURh+V1CROYPDhWPsd0m2CWmxF8JAsw0b0LFlRezsYFVdwUHA
5hwQvm6TB0gm/WkNRK5Or893GwBGL6BSjc3WHdAJlUJAvCEIV3PqGnIqnv+C5fC2DdS36X5UpZvX
MNQIxkST9W/NE1En/sLb1Z1aUDN79TXvmoBDENmbo8vUspsZJxDttsRwZtisB6ETveMv9gDCwLJc
WkShczoJWnODqA87hPAjpsmYj8Dp0LUd7svUV2nBuC/YmsL/qY1LNpDnJrfWLsPjHva6vMdldOoy
J332JeRb0TMy6sUa88fCZiJaz0KehoH+WK63BivwhXUFgodl7A6k08vDC4fLeYGMYmngXyVbYaYH
e1jesKdwZ/gFFn+93gfzcuvze6Zo0hh3+tzhxYigeoAzS/CU8XBfAkyygqAQzrx9MkXbP8xHQKtm
7jiS+JLpHA2+fawO8ebzvPUKGGvIEIC9UNTD3yuACNsICjVc+pzUUsOgEUKyQ7a+S/41N8LnOrsE
anDn8kVCGdKdi5YFdbef0gogLQs59c0LR8tWITFlKAbZG3/Dl1FVf6pO7IseLUkMcRjQh2TUCAUI
BCRpbTM1tmajUUVdwLHN+dZxmpbK0+sanlfaup5PjVxQD9lVouKnWxN9gw7WlPzg9GJaLU+l++TH
sYCV9Iw928Ardn1pSJtZQqTjGeCeku8GgcL2OpZLhu4PKKFQO7Rp7+ev9cteXBBjMNM0esBXFlps
99T2H81/sZ11mKfqJV5qMfqPXxNVoZgMUc5pX2v0DsOlOjNQdtNRHwOArz5Hg5TWc0oZDof8wpnZ
QCCOF7elELuuSl9wd4HKrIlWcGowWtgEQNx7EzQtQdhG7yp8jppzlGc32W9KMupSGgXkou+bf9RX
CVYtL8Yg+NrSCbwymz6S2Q/vB0u2uJVgoPlU21GzcKw05SZidyl3WAKPk99bceucdw+jyAjHwqKT
/t4sE0T6NW6QfSmKCxkja6nIlgztzisYZx58ZVFPjTCsOtQ7dZRk2pdSFQXOTSGakezF0gZl4pac
66iHz/JLdWcfCP70hQCIoAbiZGkLZFzB/l9g5lEK5DjJXikkn1JD1BgAa3ZKomN1RQl/q4ON5MpM
cKEj2uSxyr4SOvDOeG6806we39bMV6ziUSVgA3RkZnie4G26/lk7q/NErRfjYTe5QuCZ9XJlX7px
45D4iuaelQEc/J3RusfTemertMSmb0pcMZTcAqOglPnS7dnc4f+IO69ssOSKBPn6hOzFkM122FeZ
xcJDUB3TxR8JB+dz2JD6ymWNnt7ttvjfS/ixtxFE6jwTRqFqlVt9v0NTPKTspiQShO+iXS4FXW6i
a87jo8UzQ/u37XJ1QJDUktKm0rbqgBoXOM58J/QTKbylmcJR5JhUlRt0rXApj2H8Y0MFV4NzsKeF
PuwxCF5QlKDarSpGhtUugF84/K+jzZJs2KwBkyTSb6d1TgqkJZwPkXf+6cIZ7K9VlCIcSgCONCgP
yFMUN6Xsvj78dzuQmglYeccnge6Xo+bz/vGxHPp2DHkyxW0Zpx69g9dLnvLAN5XfhlQEZ4B486YZ
fc0+Kb8eMIs04cklbphpxUWFUpR9eB2E0cH+NAZURmpub417qNWI5/tROiNuiyK3njSGEafgtJ1/
xemg+Kc+Ps49Y+/Bn3dKcRcRwFBsaH0A7dN5FWrXtFrnylNY1Uxq3D2yrmRjGz5qZMTgRI010RRt
NiRAgqn1nUMpGM2YMzayWQCsimIcB+v3lqytvhgArPyv0udAH85aAxQWK5OlxefgtO8ipmE1n7nd
gail/yMb9cAF41bYaeP2l1HPQiY14IUKbBO27G6Zn4v0MYmkK9TiUgAU5B0xy2EvKMWD1kEKrWHB
5UHesH9TbE1LVLgYaYkDlnqQwX+yUmMRunMtg2+2zdq/MGwSFp9HK/2h3AaoN4DJuXif1jWlJJ7x
XqbC44GaLChtI+pqKwQazfNcre33CIuSbvONwTA7InyWbviLkn9xCOpTkm/SQ8xC3UqAZkVjQdA7
hSPikWvHNtzZEe5Za40HJAJdy++/csLT9YM4Xg8YfCboEN/I9rRCTVYSHofqLUPs9lV3gV6Y6GlX
Kz4M6mIA5vrElBVY0ZzqsRK9PEqMpHIC+kyCVgGIplclQJ18/nOk06iezBC1OiiS/tOZhUHEWqoN
WsRhoz12VPTT9vE3WDyj0Qy+vKQxXPhtJZGoazm53m5Go+QV1Gf8jlPgwhh3ZZCj8tfvTKwkt5s5
+MtnpSy0Cglt7roOuRxMJ2kA340IOeEr5nquAvPO1QOBDimB5n1iT2NZSVKY9/xwcnpV3Lky+RZm
Ejya4FnEJwY45YLNLZzQ9CJHw0tF/CDF3DpVq01sLvD44WNfuhpRov6wqqf/GwRy8dBanHKTw/Z0
xL8EcgrSPnRCZz5B4YoA9SG94UvA+AnE2uBNACPtNayVck/CdcR+wHrPI6KA7xtefILzdiJ7HW+z
QrZWlq+zMrP3hYHQvPYBD3eva0QZJm6fYb+GLym0AYWUDF1zP188pX2RhxxwT7V9idd1GtVvu0pP
zhhE9fisn/jeyCu10rbV08tmOZCSTbOnF0iuyzB+NwSRt0utrp0BsiNFVfodAcs2TqhbuRBuroy1
HPLFORRJGSmR2yXLg6Yge800GWDgggM7DXsNsiGqR0TxMzrjLD/EIlKmC4CGBlLHxneqc+Hh1sYl
5NxVb6K4mqYuGOslGUCI1eUp3Eo/xvW1C6LU3fGDK6hLH+1dI5qWuIaPIjr0XqLQ8BTuFfRzYdHj
U68NixZiYkB3DmzJ50mLs2bBCMH42TfAZ15GBJGW3IoNUeM2TVN9mYKOSqta5Xt5q/BdU5oVYb5+
RO7L2vP7Y07W7SCqbh0qDMzIYJdvjGv5ixVP9UMUKEKxjl4ohZmffp96yEAprGE+vRGi1IIm7gtm
ga85Pf00o2OJt8W3Utsbyw86j3lP41/sgAOyK3ClRSdbpaEhtBn7TnZDVbk6WRjJE6mE85R/hKk7
03hHirmN+gTttr0WdWEEW3tKRAZoBzN1t1ARRvd5Im1Ta/GDe3YMCXa12TiTqnsn8r//0HhxsZft
kU4GbwdsUIw8/Xmwwt1lt5fLnRVAzWeQAnrYa76bTxQ6/8FyN221sYJqzTdzzDwFEfaKTkDABrGl
GJ3ZJZVuVtK1sQFpZEyEvPDBD79QFD0ZcDSWd6JSn1yTMgYUtpIcTrjEoXWzvYRgsbc1xho8/aI4
0VQqSdP/ufyXgBrE3O0kH55WgKDVv3+ipg9flND5Kh827O3KYk9nrtHG/f3poNvCjKq8ahRqWSRJ
r/p+uSxj/HBVUIF5f2DQB9o6j1esDuIILMrAfH/VzJUYfRXd+qSrDnLi7wWR2WEHZFnUWt65mAw8
/YIV7ZUA4xn9rVMd0KI6q2MqpkEZhHIDW9P/hykE38G1lreiM+SWdPDf+LMxUVJBK2o1UEgW050/
8pTC4R5GcyKx0TILjJQUyEJZJQ6Wt9P5qO9sA5zbadO771mLkECFebai/EgM0LIH8UuYcVdeK68z
Hi/Gq2+9dDMUC9NUJ2WAXnKzJ7WQK6J42uYWSgbReeEH0eHvqDC6sOKSalgHCNzG3qwXPo8cnrKy
yw0qcFMzYJ489g4KTJdSAfDOJGu1bPdb6wwLEJ45Q5gN7GJK1aEjCAlZi1je4m/D1ttzahlSQWPI
JCvgfQjSDNQZa5KPc9lwLtUEq2IkZS6lsb6E7XNYRbiEJaXE2GfRuopQ8QMbc9DHn4yvOFu6RfLD
A8j7GICaBekEsFH2qUapSzFmDjtP4WC7/HacPuCq4h5s0cUMBQlUDQnrCQ0bSUzAIgY+4m76+Iuv
lqSuLksXVCgnzaKUDEjyXh0QKwHg8w37Jw1BznCX738qrFCQP5T1ZlRMUusSXhcdJD3877F8fNtU
9mijBYiNqyUfLF+b99NXFuTtejjB1yyD0Yok0qNcfhzb5wYcTEHfWzRoEjsdgcw8cto9uNr4FkWc
+rcAl+vZ3pxDXH95JjzZ9ezfTgM6NVLphrH3Ah+ZJ/PGLZZt+9oMMl9NssMvlueeDtKFpDt27YVM
JTKWXJQzZbMLzZtv486X06xAnmm2nDKV3aONzZs0ewz8n0TEQcsKkqm37Z00ABywFNuVblVj1rIh
kxOMtAObDg3JqV46/69szBR/Cp/8Cst/Lx/kwfbhdquqMO6QfxkcEFONDOMSpReSSzp8GK9FZ4F7
1ms77uaDWbFze3djFZEAmTfP0tzQ1I7Y+Y5zw52qWSRwNfYXUtVSoaaouGG5tFXHn/yQapjQGmLU
WfZON42oxlPMoytc+gdVmIZsYEqhx4v4lyx4iVOx/OPzkGPzu9O+xgqdLhUdOEDmRigRsU0jhh/b
zoXsxc6PFmGGi5f6Kaef8C9+A7vlq5e9326NJIlVTTArsu7Jfh8/ObnZk6KzloJi9FlP9bh7WOf6
WVsjDSECQwDA+ZlHKhLZw/YxxI3LsuQVbO6WHY9/yqATt9aQymIfGBwMU7enUMrb4L72zkZiK6IO
N3MFOuxcHWwayc4eK4VJjAf2WDXDIaEre74e5zXQF2C3UWvIIP+BbXlib6qNC+YK5867SgW379/B
dAKwC7K/vo5CZEzonE2797cujHMIqo79FDvxEwvPNYEatRx6nH+k8+hWSxvzAkVwew1q9hs2cCQ5
oLratN48vk1kqGfmtFep5os5muZ3tMbyKZFQO47NwmPoCFbN1ZZI9mnLcwnl0C8U6kopeevVWgqc
S0L2mOnqjAoPl3Puwg2iAW7IOIO713+Z1nnuqtysfQQLru9rw95K34xlqCZW1ZkWUX6w0/YmK8ZP
GF0CYPvNUdw2iWdcb9jeWEwQktp8Swxed0/L5yfBbrb6FLt7gOpo75JeZc7tCAKDFfzhdNv6T/7H
KvxYfKzOWpeJ2XaAfy+J05+GlpBDUoJ1VFL5Mz/K9D+2QQfOSoKVfiTbqO0eU2lqLrs4YHZ6dID4
EMD7piKMYT3m67KkNGUbAmRyHexj4bHfiJ1ZVLo72ELXnJNOd3HnYN5J9fPWZtRvyOPO0xXcp2l7
YBHDOzuCmpbY3fi8mgxsXGTZRXHY4nv84/R39Y4C40si205D5SJ2EadNTtXSk2DRWKli+RhanwRn
3oBPW/0Hee5Nli6NniQ4linXmk2fkXl+BDsSkA9lczoxQxBsQgE52jD/o6OiQ9K6PZL54c0h/5xX
HWP9QInrZCjii3/j75Ssh6Uj42kMnCJ3zAQFu/U6zJ5kEtnu0zwCX9aoW4Fk/oim8SgcJoqiGuGG
+CAlgA7EhM1jxaG+TGMHZIBN3SJjbsMtVdiHQfEy/Ggc9K+5nBGdLSVaiSyeMg71r9x3I8xxcWu5
EwD6unjp/wV80MMCeK9xM/Bzm+4XUbyk/X68kbABvepRv+T2QwkxNZirx5cuuRuLB8678+jGGEzy
rAAwwqO2gCKDXENGJtbT83/FonLahp4OGytpotpy5YKAfacUZ2KJ2DXd4iDqFYHMOs3Mrr0xcvBI
1w7UbMJsk3BMnPTZv+UOlYVrqSaJEiL9G7v6NMfutaT/1piup8YB8IE326LW3XYWOt85IEVrX7BC
+BAXEXU8VrqXluLo+f/kKwmertvrr0P3E7fpvf/4PyBeLmtAUs/8a1Jys1GN5KNNfQe9u8zMCPBy
UczsUGim5cqjoFVz1VhNQUld5/oDIBGbxuSXnD7dlL/2JkNpDIqhh5wKw+/ZrHcO4BYPoXX2tvAP
YjP/HnOZL+6TUxu9eTtpRYRCS/v4OkBFXohaJt7cncMMC0cZEWQL+qXIGPqCYwZU2DX5k8Vdhrvs
44sg+v1QHuw7HCqcPbB0R9fyh7FaOujp4Spzwfg52P80Ff9svh7HtpJBVFvKo1nzyf5b3YgnV0J6
d7N/NmtWthSO6HgvHWd6fC0MGhnhhoVwuYUltWw4ijK5E4C44oYN1LHkd4PBiBhV18fm3pExB9Y9
ayOnXRweSYQuv2D61zjnndJFOLJxSFBMzs09XBEOuDtVggN9J878+1VPvjYMxwb+0QGlRyTuCLIW
tqc0EkwupjCIGaEM5wZKHFt8KRgi1gdlpIRQ2gH9Aual3jVPXE3AVeHsxLX9HYOO7U02QXzGtaqR
Pxh5ykt1yJMVY6hA8oDxMholaSFu/4RBaoroWpsIOscaKs0MYhLyEQUoEEZhIv2NraMrWDmuX8uI
7c5gUfkzhMmfaJL/jFYUY8MMCclmqlGqxtCGhKQpJnTiptNkns2aYFNQFSWQpmHIi61TpuQnrQOe
Tyq2U3zMrMs9qSlmj/ySZzr11w7Reo+YtvZk3T3bjvmR+sAOlB7WpP3JB6PaZHITaMieRqLfjS9T
KFuJgIu4wzseGXvfVxU//5kt++kW4bQrVwIOsCRdMg8HLVz2p1Oixj/VairsceUyD7tl35nB1yo9
pr6NzstfoOHudkx2qZ/ACedjx3jSwn8lFSSu7lS80UMY3T/P3qquOCAWtOBBYDs5IyTMyqNYJi6n
OZbehw7JbIc+YoSlQxZ/PuTZhrJ9L1pPfaDZ/gOf3R4bjNeUz8UDijWKM2iJ1ob13Zaf5I4vmusZ
zT0YSIp6Dt8EDcZL2oxA/rSH3aesPu7cZEMFVDhiISARxJBJc0OTlvuzLvIDqnEaCualI9HqC+K4
u2+YKmKN8sAkRxOZqXdyF9IQQUZs5e9q+JbokWfApEC7tZfsQiqD5Astg95DzzRHUyCwku7iuzlW
avFgt8ud098AoWLh9vN7Tcoq0sqc4Kk9JP4tGO/9JYH8WxDhN7YJ+CWZBf1hbAdAJnrETozs+cCn
CvXoFH6qhunTJt3DK6qivx46jf5nt4ikasSyQnzclgcadfcctz28krm/yC/YxyMpnCT/KCZaridB
ACy5KURrQBDsudXLi0hNMlHEi6sSqn1K7hn4S79WdBfJioLZS1+CI/2TjpON1JWYg9652CGop0mF
qZBWzhs+rdvwW1mmopEt7nbsBfLsDPII/zMSKa3vjzs9YyMfTjB1wFEg+F0VcvZbTj8WSsH+Dmws
kyDB41hvq+chQQmpBNFfOQgt7C5+woNLb3TWbKR2v9Gq4F3wVtbY19Ph19tkA873yHYIXpCzuFZ0
ipge7Akg5weVQt9I8vO5ShGyXNQKFGzM50VTMOuGK2VDDa8s6cvD1zw6dVMRcoEimcUCR0XUH7C8
71fikKQso66LSCWH48CaautXndYrnOBc9FMlvceLVaQfLsBel6lcmBLkNp7k8hmaBnyo12UhS+pC
thlhhkljM1OEtuzML7eF8d3XwwIG2CQMeyoEM0+UosquZVwB/0wNm8/rtV6tRxrCswUxO1tpJwiV
T6gV0Ti0KbiczJ0WfLuG70C4CRixUUGCeG7jr/f+yhMEN+ud6L4ywFFLMDusZq9S2b3kbhaczGUc
X/LiDZxXBN7is6+op2LDQceiZf4qDE6nLWfkml9xS6NXZ7WqLa7aknx/sWI24HTFzmiyETFdjqb7
cq/OqHJmo+Cumf9HFN4RhzwjyTZf4/3g/+lr3v6Prm8AemxUC1DiIq9FyV+JB/YTVa24n2pWz/U8
bhSg+tj8lIklRAyg+56lG5sezc0ml2pttUIIsvdtElSyTgNGiAU3pEyT/hGE+yDaWNXBQ9JoWWjI
LEPbW9xL896dM888/nUKPnL/erSPkdfGyC/0Kwmkc90AbndB2RF4himknYChBZvifuXfREWvSa1a
pQD1wiiKqmZGbFhyr/d1fd0n2EUV2LSv1TFmP6JzV+RdIa2WvDdWO+11qZd7suJGFNDWVAv8alKQ
btIemiXg9k69p2bnMMYeqY50CVDJ/2UR0y5ZRmMMXA3OozgvvQaqHPXY6COSjgHFGD76OkjCDEmR
Cd588/WruzLYqCAmDiL1K9bIuxHzQb+JORUFMOFE9FfMJLcz/AnoYDzisivIvfDJhU9RBtdywhuP
0pmDlUYEVL7Za8/57QWCYI6A9znH4z0IwkpgxjU0pCbkr3rDK4axvb1DBlZkTsgVlNAd+Zaal2Ng
B439nHwDo7PGdkQWXjX9J7O2Xqbe2kQh0J9MvhToKd4ImsZyaD/YtYn4+8WxbG7hxHxnZP1+HPUv
kdsrJlW6xMymV1qfevhrEiSfR5E3NOLIqbuIYaxlLB2ZtyWi6FJMn0zkGyMK59Zj/yjbzTJvZ4yu
2oO0DSAGqWzz2wc52Hq7p/mEQwgMbNUagLQly9PF7u5CiAhYkKyfY68tO0JyCpnDg935EJetPcrR
tHklNBx4ASKYp7eLFZP7UWQ/tdTKYGVCMLWiOs3gD1CzFqKMm/5Jrz9CtQjuufZt+l4IyO1XON49
gxsF5Nq4N2Ez6vv0I+vdd89u5sGXR9IIlrBZHBMem7sbCq7NjLLD4arnoPR0dN8TaGLkcV8OiU12
iIgOxrrogCKNOyOdhYvQbGWxJjYcjSnbQMDvdr9mCQMrI6+hFb5T38bcVRD7P3csP0sLf3alApBT
Aghhj9sqBvDYx2ISr9dy8uNfFIAvrR9CfcZbBZrZXGeq9Wl7o00r47UpnvtfqDYqeJu9hAddLvRS
Q61HQrcFOa/ZrwkAXyUa6qgCqgx2v2lqjMbZWIr+1+5HcJSO5JMKH9+YGBIjrY6jTs0PtbMFfeOB
T8nw4q4jqsGZsSFc3SqTfTAQCQIOj7a613ArtPxjlw4eO6XhNLgGURmwBpf5U8vCHR8L5+hW0GPF
Off/2mvFbV6EhU+l2FSRbvwdguiXcDAVWomBJL0L4p+3ynUKmoqYRFP0XI9DI8jCDR/6sYVKpfB+
tRE4hcx1jmqu1S7Fm53AO3bcC7VN8ujMzUqy+rN/dRAq55AXDUSbYSttN+2D+eyelLOpSRW4T9PY
avW7kPbv4OVIvjPPvlpjLHIT0ugugdp0lw4snPU31G2/3Ns3jobH0mb+DXSaArVFnVJvLFve+sr1
RcHF4iKPaPJMOIz/8d4OrqK6HrEV87dSl/BBk7kBidrxCCVZSKOLQe4U1xakvzzUU03ijxqyqCGu
xQTNKvYPVqcOLdYfx/S6W2fvDAlANC9+eNIolFo+RwPdUxdFuNrnfQwTpKdnD4DVTlY5XTUAcma4
bndYH682i2xUHAzdbK2TJTZUAz0MTToWfxoL799kFf8/lbIJBngum/PbjhP+U+1KT+3E1pZwLT2w
wwi6KQ5kdNAKYZOkSdD4tuASu5WBOhG0taUsa96vTMsLhnV/nUVvq4OIjNbA946u93w9gmVR0kvf
6/IIPkx+LenA9uumujPIyrtd0IarVbzVHYerD8W0INtSREzVUAjLxMBHuUwfDkFIj00PB9qwhR8Q
O+GgGTMaEXgIR+mhnmKsokycGIVf9PRiQ84sHghYdTWtkPwo0f8brbrv83wHCuN1QHKreacZwnC5
Gt9ue2M00yE2KBXBthQC3pIGxSPzS73zK6XMoJqN6vkFp5yEdRVO7gmHrK5gsSYKmT+BCR/uvLGu
qEks+Crd7AMXJPj9qA0QzFBkOpYHd/WoyVbY7lo3pdVjIrp6TCVo6M1klBwhjpR8yTIINlgAnThM
Z6leRR4dhxQvH9sm5KBqiel2U0fJtGYkkvEyn468bHJvFq1ppKcr4q79gTbft/pv4kYbQCqNTzFn
Gil64WaLKTLQiTMNpxVHcCEfpW0mN6Xd3mV8BCuf2cyzfLIj+iKnulY/pxKv0WXWizy681Kha0RD
kboHO9V7RHFCT8/Gqk6Ww5TpAkcutXNHcGqPsexqA8AKZyRE2JQADJeX8yXVibxX01dT4jPCyc1Q
//12N0772nwYLzAfrnAEkgQbFZ8q/ZTjbppjlu+nHWciYJWk2atHgB1aAfHEk6yfC+LTYaiLVSFK
ZVAaDIEO6Z17Dp33FB5vCsLzS88cVLcHQyFuvmGkk11REfz8/9NxuJGgaePsCeAoJTUpkADVWa6D
O6+gmVe9IBLmvUTE9nNuZU0az1ZjUFSTjsi4UIg+tmgdYwpzVVjgfj0XICTPAAqG+cDkllb/FO/T
0Ku0Vzlusex+p059vQ66MDe9AvOyPbXBnQf8tPeSHO3UCsCv30T4TOV2Kr7zG04JwLoILCKrArRS
zImNy8nF4DD1pCd7MU+SIewWXLLiMrslRtuVFKygeQXZa5zG6wAHLligYGWW25FbKHTJUg/0Vgdi
qVAB74MF/nWjyxdWVqIDJTM5KlHN+XTGRex/I4hw0tU91p8yIUJhiWKCDwl+Wq8fez080UcaYURP
SMlPNoeT7CIF+3Ye2PCx9nGhDgT5yATvo8hBHMNTYrjpFnIrNL++DTT0i9EGgva7EludXy4gsHHL
/sozU9HfGQoMm9TcWM2vikwaWXxFZyjlgP7nRKgKGzJyy3stW7QhQ8sFAH0lvzO3LpdzqyH9CqJO
LN5pTTegETSxMyov+RD9qDhRUwRuus+WhH0Stp0hh6wuEAOC3jMxP5qTBb/1wKxWo0nTlyatttvR
vnyyEQ7GPSiVfFf2tPPJ9aQKsOfgpY9Z6JbyqvcZmiM4MfPqBqbW4Iln+kDpjKVsSWtmhdd6S4N8
wm+w8H5rI5HjgM6Obgb+wpYmmprKoy6aDqQM74zhryZdC6+BTH5F8KWjSUC+BE8cpkO/NW86J0OM
d+RmScUkGnXL+b2CoCURRO6zQxnSmsxdhjtMdP+aP8iQ20VwwZ7PL8Q9+dYhv/GcZjnLqEXpRjdG
2+O4LURbwDWr2oKfjPYJjkRM3+wFEkqTb3uSz4tjmNeDeUiAGh2kSPCgdhWxJqu7MtLHigXvwED7
hn3BV1yCcjM/LPr8WeH6ODHMydASdgPm3bJv6DySskZXzT0bNI7YF9U0huXSXq1CVLvlyG2eSu9U
eQ1fbhvB3qAvOyD6NJOOsZiT3sceLiGzXhn1g6IbXykGEyu4foYku1Tzk1Zm/q/fg2KgDau8OJWv
/8iYWmIqk5okJkREve9PmHc/fqsUAMeeC1ZoYD+8Trgp3OXmTwB/FBZ3nBKpx1pmiYOazYGT7hds
SsqzMmRCbFN6/kLaL/XYQKDVvpUXrz4lkiRxTCvmkkhoEmhIuVH8jF8tLsCGVJoTFqKBfiXLIWsg
Rmw+3ky66VVLb1o91ve6h+HomLKPkfsRghIyqXxKruTPMeX9x1XNxfizm6ccB52V2VWuc9J6gVzr
hJaLe4QKjsOe+49C1ZmxSSC2h3tLamctcmSUjKRGarPGtGtcw3BmsL1vmuHOA5eVquS0GhoJWgaa
/HuuXqqypJi7FFc5SiMhSdBPjRQQhYRxasgDmZRylvk8uPPZ+M4UszAuksj28YuA5bCNloY9VbJl
Ughl4zf1fR+wjR7sSoAaGcaSzoOETpT55iaiYuTC4gWdr+1IpuaSd4zeZWdBpVuPoZwmwHCX5N6a
IMiN0CgoXhnHdsPSvVW70xyPjZbZkDucksKgN27Pfxjsa2SaK4DpZToPFGs97Iodqmn0LZHp0Ktb
eQ8Zo3pPJpzUxZPlbPyC/Eqddlo9GuF9PdfbqUxTbpyNUqaVhJ6qFQkIyo8Gj8C4t9egjBGutu8C
D/YE8ud7sDxyyj+jlunuXbEzHEVjp6nWzeB0xswjh0r2YXnwqjlP4GAeevxcXmoRJ8qje8gwZ2Rg
KPBea72uslv7JAnE5tsxa1Dio3lWqW3K5gQjNUbUIaP/7RxHB+GHgBsNBCY1LxO+xPbHxVirB3iV
GivgivgHFnP0RA0R0jCO2osUY714HhbcC2/xdmLBsP6tAzJPITcqqBmvC9tdahBuZfmSP94AG5CK
6KluTttP+ZdohMb4tKvbdQk3+RqjdBGr/cM2C04hwwd1Jekh14fHd1xs7J0/qHUSjAkQexHaSCLT
povua7yU683yX2Jw044Dgb1F5BqUc8Ley8cXZPTw4DUBustpaAyrbpIZfeB8OgSr7yipXSX4DqGk
fRpF+mhLvu68IiTWNqCzumU9nykbHG4fAI+iCPUwRUf0ZWtOPBggKPxyqx6p/2aPgnVj2GJebvab
UNqnjmV8O0Wjj5mUXqcQ2bpPcMyHwkr9j1ENeRzEbsyK4slEMXmUv6EhtFDr9/nFBTg7vzH8iTBK
t+l+UqdeN6Opyb5YcuXiVRCQ8aZIUb1M4CmZ4NRV8qmAkZarcZW0zjGaTgTI8et2d5Fb6zRWYSmx
9Rv0rmwqxepuD/CBO9rroh0D94O5uO4WDmIfyDepn/+QP3AC13+X/ZYLYA2iVSjaGACyoTiO59ZG
kAqEgcSQPYsa7g3uLkKbg2GQQOfL3Fc1r5ROS9wnUKH0Ws14B0z6mzlDbOSIrbflJIKApJ/Z/xB0
SPD6+LUePzy3YPtoB0ApPDecFbdCbsFuG2aD1mJ4Y0MOKVCMI99UXLscZMDmfuGL5jhMIRpF+rXw
zJyrxsFQBrdBLmHMVayp3nzg7l6fYa9LBCjdbY/U+S0GxA5/ncsClGs2Mv7F2TvQoQ2ssje6K6HO
Ohxbmbp8OpXmGOOshAzTgLQz37jpIyFac0T+JJcHdH9I3scvLrpeCbpW0BE6vAidKN9FR39bXuQS
h03UZt70qQpffUgVSya+L1VfbGp2+f+u3mTtt2e7S5a2fFu6Vv4uBbiwQwWrfqjhpCN/dEE96cCF
PKSvywJOI2JbhBwni+UfZ3LDlEs78zrtOx8pNU/zBd7CHhEHgm1lCw+tWe+ll7nXwXHgiU98NRuM
OD8KvYS8uv+LWJN2b28/Ri13fDXHUB3+FV2Mdf/mVoazwf70UAK2gr0K1zP7whCttkcMaB5vQlrO
qoqTtprkD8gCBiu+8fSaags29ADfWwV0YrIiZ+wphaJ3p/Uo2R9FBn6S3EeZD1mkf51xogSkHJVn
Vg+5jmRvbfScWEadEfi3+iRrz0oaAl7vIM6BbZ5luzjxXtvXzj30m5BttwxUigtvzV699X0wfvE7
h+sRSvgM1sFx8AXpoQHQ1AN0XaB5137s9T44SDx637fjHwi/GrZDRVzIYKJ9lTisR467oyd4y5QW
7aItZqcafsNgeAr4Kqu1dYZGRm6GMsUa1hdAN+62E7d36sBj4MI3eomW6BXpIP1SxxzGk+qPbKyW
oZaonJN2r++ER5M8BuxldshqK3VSZZ5GhcvWJRtVtI/0N/PRurImzcc3bbBsQoa/71N8L6oumrZo
XR3T/BV+wXfXrViQHLDxnc3oE03FDGAeGioxqaG7rc/t00+aMfSDmPhk6jwcVcnC0EYe9m6/W/1k
h60zmBYAoxfBU43B1zIjjmaz5LlNgQxJTpJzJ+quIoM/dsPRKQd9HwmYxClme+OjDRp74TM5d7rO
9nEyS2vNfWYMq6hs6g8DdrwYdOok6xIqCDKcSfg1FFWbzKqGr16n8dmXg/tSr1MjP1yfTm2xDpyf
+OHZx+baiI4Sw7UG5MZPuQd2NHZhRXl10anCAgCQBDtUGmJruWS6IdcO8jjW1DQj3txRRA4ahRQW
t1lfkUl7YqWj5z8+F99GP1kEWHkTRKB0Lw5sjrKDpYNlkgqCSttBO9HKPcQxaDQKDFoMNuRE5yD2
6pe2uNz3rg2Ai7+mVFwfDVXHb/Q/wbGhfkO+k1KrWg/A3l8yYca9dpz23d0vcCcK0SQpyFHEkSTf
0B8zti/dIHjO8on0pB/u0SVzWGcqMsPlrPQ3UHKy9gxUEoUWMhUle7heTuxQz4v/epOfG3HvFFp0
plFFQ5UazrtG7fjK7f6I9w3z1aV/F0k1mUX1OSSAXkDhrI1eB3TIdkCmoPGiOWdaH0VN65qyWZNX
MUI9qkaSsPaqih3f0TL+jAugOFyDJF+heCFGmiY80sdG5WdTq+0ZJlexyNYlCWsg8XxHjnI0ZGxL
h1RZTOFO2yEe0h1LT1P44coLyrOCU8a/NM5dGmHOd7sOwrT9dCKokP1TJ3Q7cYn0ZkruUyxQ9jNq
oAeISyV5+2O16nLYGJFtphnmg8lxra44stds4l4HD1qDVZTooWn7V+8BIjeOFc6luHh3+h0SzGZz
HBfnpUkIFNtCCvNA5Bzy7S7nussnbLvD4vLBFkLnthprIDJt7ES6l+cjWM1KA9Ex1d7BzvuhCtQx
VAg/Lcb3O0+5S84wMwekShTUILbJ8MykNgfiH9QFVRf3MoXLufqpN6AcnSI7xx6O/DeAWblU3rUO
JVgizVHjq4/MN+XyFH4NNXTybyDQfk3ihV6p/YZU6MvAn4Ow5lZI1YUJ5/MDgCa7x9dPHy8i+MJ6
zUSOSjGw2t+/ERxHT7H1Mkan563XXHz8Uy6wKvnQySj+YWqaEqiRW2G/G2H1yDOmLOiO4MLPdkA3
3XZ4Rm2G5tn7CMq/4a92bNRzhObPJKwsDnLp8taX3YOt1ij87WdfEoj5ujoDbTFQmDbRkGbKIxjT
fiVwbEyuzjfIt8As1pCypS7cklPP3l1lQ0ZLNCljGuSTj5UUobgeUlBJOtRjKEw8yIf3gOHvEq2O
mReJq21BsXnNrXUITqRGMqfLUydcV7wh7LvYHHqvDQaweOhIWVT5sJgMHCZX/cTPGShOv7koN1bx
PJbCEtngWCQ1YiixJ2ukwVkVRmNUOPVOzoWB8Ck1ZYQUT28oVaDIdt7wbBTmAGp56YDhVjW4dL9F
NmKf0tVbj6iI/bX1B78apnrisihCut6Id7rO2v5k4RGckZ8ISTrgM1hgHxYXLFiihvjJq7bHi00U
uKTHQkix93H9R1qSUgRtN9kC4Neb1liZpYGbTwicl2kd12cJnypuMDrAxzWeCD9LORqJgdpC4FNs
Polsl7d9wMaMy/tZKGo10pyqKa+aouB35X+/0lVrmrFtfe5HefEeX/4x9gmQ/zspg3lCLh7h3MPw
OLrSf2ysgMQpDLupWMjptUx8jzakXQ555qPsy3fOJQMqRpN5QlV59lCg48QvBPXmz9B2BcjoeTjT
12Io6H3LL/k/YDJrWKgm39YnctUcTCzaXHV5pnIxTWq6Dc+gf7cTXlpFU12aqFn8hGDj5G18xlkP
vGYgaXJyvLxu0prkuJCeR1wpD0CG/4ZWFu1UGW0/8OywXqGcRwQXQPH2NRNJKCpHzUQ+PnVintTC
rQKkbI9no2CERk2uiB8/O0t4J40bkhy8SrxWa4vKe2qQXRNLkGOrMjf53+AL7mbpfwf3IIFG5H8f
mTgYBnGBVR8f76F4cBm9Tul1//gm2ftdjAtdJZPyOZuyA/K8AfALiB7eB1gTlxgdyskKfYuEPR5z
tcemgs47exA/bIFeer4Kz65aAL35XdarUbRE26rQlS0cEreQtdrpEkJPG5DTJ5lqbOGw1a+VU7q9
1DMj4m/EJBg22O0ZTdv4OOXQdO/jmnmT7VkSQJA2w32hSwkjRWGSs5q1WSU8fF8mAmPDdDsdPy9V
wkmEOaAADZ2Twq5yaFXdANgTeHxxc4oa3AhDASESpX2LeohVbORtKyUfjIOADjep6dta5pyyyvb/
ihih4OkYlrM1olnpO0JzcP3BC78Y+259NaAzUFDAxkL8pzPSTsnajZqDgAcQLv+5LETMwq5T843Q
qgdbpBx+A+blhPJg6wN8CU5c5uBfR5DdW8tgAIkQb3FFaisb3ncYpokdxz0T3X0YFMK+/aydVCjS
sW57Gzg79YRN7whrAIFXYEUUOaj++Vanf+Y4F6H6n57dLKyTqmDcvdcY6NWn3iVmVi3KlujqPS2L
zcv1ZKhyQo3Fuarm90TtzyVr9MMS/z8ZackxQgVjA9F8f6FeN56FOUTEGsFC8i3L64vHiCj/0dfE
djrFc7LZ0Ip/BXbea/jZ+2CrGfyUGaDJWR4dcTTT3WUYVciwrplOINYuo5hIEXsygC/rYM0xBJFa
IM/bRuv/PiWyzjaZ7g+DJN0X4wCOh9Q+qEtGwR5IekzMpG0cW6RczsxKdslgYkQ2sCeT4mzkLc3/
0VHfUbA89F5b3xKF1iLJJoqZ8xgyeQlIsIK4jmJNjFNIuwyaZf04v3Wm6h5YEjxRGjskOLvepZ42
lZGhxl1FSMtnGCLwrGa/3vYB1yElFIWy2Ofzuc6MdjzBbB8uxiH/G2NANl+z3paEgUlHCICN+nml
1quBAjNVHc2g8m9aw962LD0B+f/At66+C4hYZifqTsNwRF/p6UBwZ6yNmQO16R9Tnlr9M/LqsPlN
RoVYt/h5Gz6LMnwAppeadtnlbl+li7nDnzmUSiA6Q844h2n/ROl492dQ8Z8Zfi5jItnHkXGgTi2Z
JOapdra7tgZTslnPGbsCXhNnER0sF6bLon/1WCKAwBXyL0Tpu2eFlGI6ok9Pt+7bqFufh6wSLxey
6VxAZkV7HHC+AhzcLScFonT5yqmHmxNIprorkDNeCpIjXeAT4tPXmXNQdMuql3LdTCaoAjVhNqGO
dehmNC2thwPDF60+8qel2KRKtWPlQJOAOSX0oHO23xtogbvtYYPPrYdmMYCvPunGZaAD7AFU9bAd
TZTYfOeiKpGJbIhfdSvKN7h3VshR0qX9r3DMxwX3Jj+FGf89hNCMKZLZjcYmPvADRPWDd74Wf+Qm
TxqrkAulnRyQ/1Jkm+6eiAAX5uegfbcni8YqHaV+R/qjAyHn/TT8ExC/uY1/n7EvjYblcDeDrjqL
5+dWZivGIzAJBRnd1/U8l2kjMhkQNSPXXQRBFSqUPphVFzUIWuzegyW+U9bjCUn3lo8zE9C8i1LD
zhL8nZXLrZd9prdG8t7RwpIsu9O320xOvkg3aXj/iS7HdF0OZ8ujxh+W8BzNu7xsHXBJaThwORhb
jHG4zGzTiSZvFnrynyIx6Kv31QXHrCo4inLGlBDcE6EplzjS+iE5B4XR+FEGprr0nOXkeJG8MYop
Ky7NiM2cq/MYSo4l3Ko4tK88VQkM6myNTrPkEAOGptYMxlHz9ceKLhQLAwv6Fpq4goaFFNlYbhwa
zl2Dbm+HoyaBi9BKx6/nnL+OKLUiIOLnWerp2NHhFxbJo3GAijHkNdfgJCu6Kv6eY9cYobe1VOPY
MeNHwb0WOwgvPk6jq2MpulTUIB2VTu4SG9BTiz6bkFKksndV8NDfLBc/7Kchq9kKAZWX/A2HVK3p
vGZuDX0RpLki/vBoNZUmN1ehmDU6yHi/LF23f6n8VuaGp8pVHCWgil/+q/+1FnI5b5HwSFqRDbKD
uilB/B069AWrhgAcYiraDN85UQ5zSaRIGP25KSO5thu2z/onFIqjCUmXRpBZNO5xNvyr7uoUjk1+
BdKDy2w5Qwnm/Gdf/mjMBPDFspdnRojtwVGJtgdCvW7UKaH9uA6NlOdfkRjTXplY0mwUBMBIcdPU
l0F6F153bnTmulFgBPCj+NSZPjcpjXr/LaDzeXNA+auuJ55XeeMmtYI2KMKOz4mx9hakpZAEyQ37
gCSoiVL8bdB0ULpG7qXW5OFBTP08L/hNofnJSGLSoCnG/TpTqqjp75p6tOvjD6lHnkiKtuNRQpTS
5/iu9Lydija0yP8YoRJJa/CsCwdgTCxg6CI0ykyngHIcpYGg6INOjuMsVEjq0x7Wrw9OobZLqdvF
RoG61CTq7JiJYh+KwvkPrF6k01ZPsV6FEgGWRXMdXKwpml8UC80CcUmfGQAefKhNXXNAJ9kmRVIp
d5AiEJ7GasifKhys32XzXpWG9M/JM9dTvjEPMzF0hEXyD0RRyKlmPd1bmAKkdVtzecA4/qca4W40
sA8AXAEbMCZqcfApsRDcaUUb69avDluTBYrF7zyZSx9mIedmJnfOIeDRZttxq1YptWT1RW/aPsyJ
jdBJCXwXtj7aMkqEX/yMw4lnGH94XD2wgZVjZlUepfOo3cqfXbuy80p3Gb3XpPbGvGXTn86V4gDL
5yZaunCoNidXx8gQC9TkX+fTMGHFeTWCc3bTmho/5R//Gb4ggFOCLSSIFpTRcPJ+Gzp2AYMm9tCY
b5SiF9UQ80IQvoXztcgV+S4nkFs7Nd9pr/ST+SzeVzBCckR4fB0OnAfd0Gch3tq9uHT8OXybmo1I
Ob/TmXyVsnBskh5IoXNj+rDBLoXFnk2qwm4rNzWxEjKV7rCKGRNiorJDvPpKp2P6xlRH27oJwOPX
kCWZVf5SeGIYSDdI/gqJlpKVu9oHAHY13XhDQHG384qyZXXRJLFMG+DojxPu4DQskGqMDjZ0pJM0
jQW30gCGg0+kTPYWOuEM+HRpApwioXP0kFmyIktCx7nf1Jq/ZCWXj2YcZ+OjOMdI/wXp7XvVa3Ph
B1SJb+5do6OWkn0WurOvBjylCxeXMQFgPmpOyXvP/enS9WB/FrwOT1NQMCDMaHB7d/XlDZJob8EP
fTW4mqrKzvvyYTSnHFhJXUqVoXC1rh8A94Nwf2jHlMC/bETwwHYcpHcp2wLGxzxOU/fr68JBw+/8
i1RSBtG2cx6sap/2J0MeC3jQ+u/cVWReMhtrI/5PzVN/JkpRtZeuLYhvv5NrvTi5tg8KjUkd8Hya
uY6LH5Voj3/ighG/EeoSLiI1Ow2+1K05p1kF/e9N8Dk3ygXXUzCIMOWkpIznnzzPSZODWbOVZNF/
P9ZXjfI+8mYnRfs31ns39iVCtzx/Ws0uZ7+LYoFnORXt873E48hOUiA56NDMOSmGvw12hOiQCfIw
4Oi4qigo0LAc2vSG2g3yDMr4DTURYIOZ6XPbC9GUKoDps+WYhczvwSohhwTgbkT3TE3V/r5I2CIM
aQw2xfXMEqZW0zJ5dttiCSdy3k+R/2c1W88cbHBrNpJg4QGiz2utZcb8jgKZdL1BnracE5NfsECP
oqaW8eO6/Gz0rgEpoJBA/YGH/Vu3CWiv71CZ1XR70nUjWoEUEyYeOMeojoubofgexSFfIXeNL1ZV
M9ZIOzxWU9KnkFg4BFYXKrDX/56tjSAKRQfEtdWa9pzsLH3TVycmNWIyqXFHOTqEDZHW8mMUgj/P
mRZh1OndwbtaTHpm0IAU7cWznLJULpcYFx1Mgd/GmtGWaZlxRiWErf+jwzcY3dpfEvDJvXBn6rfh
SzopjXt9BIWOFVjjBetXHJpdRY3l0Wad8MMYA3iUqzPTK3rP0LjrIbF/5HEouPxxBvRSIRhpkT/v
dI6v4t0TjoWuuY9zqBhkY8U2obgNVMFqTgCUjuqF2ldfja7poETdRvhcHz6iMnkq5Bv2DKVpgM1j
QnKGw4U5ZOVK7MEbxH5lQM7Cuudls/JId3QS+X6aZbSa/M0g/rWU3DjmKw3ryC1houv6z+I5bJC3
2jdScQIefUSCf/aM+OYbcKQfZn+A0cEieQdwOkxiHYj0Rz2Rckr38DU8bKvkSbBfo6tqTiLyFD9V
bc78WmqiyiKTcQFqyow/1WiDR+jWmOSIfQDs8wl/gCIAXCvNJlWtLf6FBa7oMh1tl9yS/pIFkFXA
rYXrxG6L/Af6sVnhY7ASmHsoKzLl4secFd8AchMUpIe4Y06g3fgNMH+NYzjVt265UYduiDqq9XWX
6U0hDXICyIHsamR9rRQcqcxQCzTDT1UWiHt7SVSU4DAAVVy6mZBN4DzgJggE+tx11Cjwdz3yexFh
io8I1QsxuOAxYVqMLSe9nuGYEkCjrz+nbDk8c+w4OAmpxfdI2mhSP0w8GzyLTo8FCARMRdsTvdcg
zj0fkXthmD3K7QdFGgBNa1JWyHsr+RW4eTHC31H5loEi7BuzUSEmqSQHKk5uxRZP7kK6lR0EE8P9
XoQQhLAw2Vupi95ORl4FeYM+hmJUu0iACXITmqgVl8WKa0Qe+AtEM61VeTRS0lPZXO4QHeNQlwZe
vBVGVMXGgBIcu55E/i9vKFY+/LQIXSnf8qk/mY0wdYQgayH+8deC0e4bYGRjrKABExcBNacEr20E
L+ak5v58+5Mds3lYJbQhliYZ9JdXNTvO7r9w2vrGjbL1nTZA7VzPVWS/I16VvN8gLlu9qiGmIQYV
nVsWLNv0H3NZR4vjQx9YfY/UhCz3INMCHk+NJdNrqnFeQR6Lt/YqYowjJ9sORH0d8rP/fcXzWk4P
6wciSa+ZCuf7T2M7oKrz1HMoSjpk2VVc3P5FmPSdNGlx4AFO3bi4GwKLHzH3rDxFGuaWToiUOoCU
mkGFhe9PL32M03iDlZsBspZHlbtN8PGdkNr0HCKQvXMnMEsakvVYmN+sEfrDh+EDUgKa8KKwUQlV
SmARigSGXKEr3dxb6SM4lyhWsTDzajWVuYOaiDnE6OQDBSRVqVlF59SeaZeEpp/erZFHGUWSItjD
K1EnLEa1MkQJCg654n5Q0quIreF+eBpRYebNaCcD4AxFLBEu2vbGByrvlizD/wcPYFK7ARB0vjzA
TfuNN533DhbBmSvEuZtLedvcYd6Ls+LwhoCKxk54fXq4b1bPwvujUNjCmUbq6nj/af61W+NzpQz5
NLVOIhM1joRy4UKqTAA6SQnwUM/bhszz8W+YKe+TFNnBhKYZBOIgzivo5ZiA0+mqWK+4IDoEH/7s
az1RrsBqFFkN59nxmFAWLc8ptFxFrHSuFAIf+fr2H4LRQXvsYxutP2zvsx2S8uAwERLCrf3s9ws2
fMIORZNYZa9Wrl0brypRhpnuvlnvluGaLCCYpn5ta8dAFKQX4pE5R6yZyOErWyk2w1fItwgvtvbx
fUSwknrjifSkQUMGAOO/qhkBOhbkyvmAAtWUghshBd9kEYQWlpOmL4BykaPskgQRuUgOZtnhbWSS
J6wz/W77IfVjX+cgsmw2utgC8pnmS3SlFtzXEPdkbt5Bn7HB441BOg6k/8LBwtHFVCorbZv9bFCp
mfSOyUCZQ0GKfeSaYV5p5CjAhCrZD0Gze57zTc9yBycSjJcRzHYfPV8oueOJ7i0bjF/p7uUViKHP
/bp8Ke0BZDTgkgCt+pZeAFLOKXUIPj7UHX1h8QErsJwlkwTq7K87r7QgQGsJRhrIC9byPSGwEHUP
HnqM2BejzX2UzDMM6MmwBBXgf+o+DvUfhidZMBp/75E34GtjEhQW31G0YXm0HKKg/OwH6Yslg1Fd
dHl3oTVnmkjWXG5+745MurjE04uJ+lcZ2RROhdraJSo4wvq2bfIUleopThDcIFbLvsshLIMxMsh1
peTKgH1QTDClU9nXr65UvrFbbo25/K5G8u8plE3gFneP7xzYSu35aDbU4KknKBqtJMnN0h0TzHTr
mLnznX/EXUOHeeBxTydUtZcEWdXLm6PFfGW3pnOIUE844ZTSAFXzb3qfB7MixHbdpwckY/vuf0Jn
NPBcimW4R12H30EuEIc38Njs03U+XuyBu+1LtqW5T69seg9yWK4viNnA/IDD9q2yaiOhS0OO/50O
wfyYzDHqXzn4vZAU1egIXe8hoaP1hAmi+5urfvAT3L4QsXvYyLF/4cmEgxJ8atQtQJf1KJlXXyMs
VlPwLOodLSDBYY4FN2yaP3UVinfChf+5a/D73P2J9J8xNZpkEK6B6vR/zp/LGa6YHEWyjvB+I/z8
MeKVIIS+3HbeHAukU90RDFNd7EZBIrkkmjo8j+5dy/luQYa3bOtxzbdMinokb84+3x5bGYvDCiAP
shiqyR7AEORhqXlHuntzUiWdNlfEBcKT9xGJ6tXASffGSPGwXae3loccQQlOz3l6CUj9SzqzHXJ0
sjuhCyBJW0ckfVAw1SFPo9CqDxLFk6Te5Hmi/TFtaqRjEF9s5WK1TzkKi5sLqSE9pOO6GuO2zGVf
1vyCJk8utjzKK06jbVfhN23eUlp8duegso7FLdk5DI4fvl4q6wRncK4vWmNyv8XA71bHVbwOv+Zu
E7cc3ZjavO4LmHVqUfu6RI6O8lCQgZL46F1n5QR6uJ989chfkJBxwbhq05PuzFgF7NSebYKgKvD3
ZKHY2onCP1CM5YgQ6BvzUAYagBY+LuVWX1svuY4w6ZRdsVjDcDxk/n3sQttLvaRSgrknFB7vDUaM
8/RScmIEoYJf8KeFc5dFROsQ1Ed3GAbSyqVCHT0MIw9iGp5OAkrj9Q/ZkDPZkdvvo7FaFJzt1oVc
jQRHvG4PxdxX2/k8r5ekCUqPet5Y+hGo/hyOwqXw7wynSx32snZPHyasWzAk4XqCcS40iaYopUym
58F1P4ZttTxMu7nKHr5UgNh5HWTYAb/RYECFLqBoCxGYkOaXQfdcQ4IheEypR70o9oghGw3onXTE
RkLCkuSCw3gyLQbcMCNiWi2R2p78A/sztukkdHyqF++4Rl3pFIXc05nBGpRdkFDgwUSDXfWkkQME
yBYFpjhkEPszNS3eDKoPU2+yl8DZBVKSecHcI7aeqvJGbrq4jl/xmHZDiDDM0gjXs+VE//uDFZ6x
bDdLV/bz7ks3CN1fJdbt56OqdGUMaqA0hjobCJ6WU0Yd+YZ2djgRVHqr55GvMPwPmWQ79Oxyex+2
e4F7Xf6sUNnytYK6QEHB/Lx/mivTKaxebXQxyKh2gPumzOWQmU1HOGDPv3/R/MKHFP1hiiuSYYGu
pBUg+DPsXzAxIH+tpD4+ketk8my5bJZ2BKFCzj+UH65tPxPyrpj3KbmzpilSYtob3wYJ4awE637U
14q15jFqbqgiYfp2sZx61CiiGi8UYkuH43HkroDmOtpsopKtIF3jlCfdf7GQEeQeWH/PaEJaCA+h
mKZaFDViIQsbgccKmPu622nRBimzwF1orNwOONvr+vZ7rMhb3zhDx1O13hU/a/y4mCTEJiLvnAbm
R0PGp22Tcfv4MyMknvn3kxFPHPOChaGa3expBLj8eI7MRYZuxNK1nWNlUr+/QBplofAXxUmqe/jQ
Qp56lRpa4CWfoozkl31XPnFTWhYAtWM84V0if9OanabmacGdmQEKRang9PJGubyPlB8lgjjiGPvj
B+ENLVBq2wxhaPq4F0jsYObGCwYeerYFsiL+MeMkOicCVGwNC4YqX/lqVusY0RaQXtwHoMgD5bj5
YVc4mL7NkdXaMADXhuuvgF8HtM+eqic/yg670/Hfzxmh4Ck4kQunvO9PilPpf+GJtfCc5FBDaFxR
xhbrPGgxt+NnaoOzDWrplvgo0Fliz7ip9OT8nVwkX503MNzxgmWvNuGhYT5Sqn8Ih2uYKcOioH7t
OALsHVoDTe8GAmKdG/9IlZZVRPc+J7S7i/dqN7TvJ2DLf/q8538i+K/Y3jz4HAACWCE6hy/0uHi5
3b/xvog+fTAOkleRdkQYgT/Xzj+7pI+roWrG2923xbNyCpu8Fq28In/TYWvbjvgQZwQnygYQqILN
ybaUG4Z5CiVly2Pi8SS1tAuMfIBrxrBApTtg0bNBRZs/BzBSO0jaAIJyy4o2sYkiBYGwb3WZUZjg
38UcAHecNUBpLQ87Uz9NDQWKnnNnaQP/NhUQh2SoXIISpO1A8WetBaSzVXYCA4tc1FA3XB38kqnE
i+is8EBv9WDMkH0H6B0sMcn6bXRHRbcXyDSpc6WMFTpuQE3CHvh5u2uyeILJCEchaqnIvKVtDmNT
n9N4KUOsPO18iczIs654QOx/zylLth8ulBfdiJJRBKRpUyeD3O3clA733yF5eQJijKTv/FwWgBvS
QTC69vYohcp1+SIcvtXip7HUNMs+WsEYRVaQiwGTt1MkgH31JO2F47MtpiNzs6n639Ez/MIyDKvE
EhpawyzDB1R/qwNGVvHVu4g062fhHgeBp3nrhPirQuUI54swaT4GXn3rGRpiJQH1fdbqhu8wRwAu
DHxrr7haeZ/xYGKsF9VY0gqc1xRFuZ6JlG1DWt30sQ7pPNAZYhmqsWvXPNc3RquZaJcqxsqkAHAb
OmRcEzSUNmmbq5kKu98jDghkc5blWB+iPgd9oqQl43FMA4RdpSmGgOmM9yIs5BRCaIlS1sh4N+q0
6dNZEWkySSCrhWpGZxC0zH45641D6ZdC8Lcd0l7UNLVuNL9i1oj8zE3u3sc9/VqorxWa5oyThEzp
r1WkD1gl8q08ZrEf4w6baE6rXj7f/HK2SrU2DiYlOg23n0MdFFXgoCYUE4qPUv87y+BG6UEyu6LY
4kYhLgcUrbsxWNXJmMvsNhdwed7FM6/PdiOHmIDlTt0+ow5jbQelY33puf4BBVPlWcqVLa5bxpky
or15Qp3Z4NjMK6P07hEReRAJoMKLlZD1I8ag1sqnK5kmw+0DQuV81GdTCrMfSrRlTfHWUkinx6E4
u8zZ15g9KJvKrwjA1q+H2rpbCRonD4J0iijyzlHq/L+LzCjyxtnBEhNjC/nsUSJK9dJcJlEalNlt
8KjRP7463DY3vRJsjdeGG9VE0ngNyunxcfPnD5mxRD9Wy9q2NAPP3DB3ypxGev9t75mKRxZjGYvp
NOJafEgDIA0NP/YPCoii5EhH40a/BDvWz2IkSAKxKF96SgFqsFIUJDuXEkWAyYNwCdKiSJk4sD0o
IzO9To5FJMdFc5aDmz+C+oQPIV/qd1RuVLOy3jz6rNOk1YbFyy/aZ4XCGJV4qjw3586RZZ/nxuuq
p2WLYCK/Ms7Rnrwl+TfT3wBBonGqTsfvNcuoJ7n8g+NSx2Bj2PBd+QFSa54HuuZavhj+rhvWSDNC
/0Yi5X45PnNOjlL/wdKPNbuJChViqqu5RTWaAmGkY+DrtgZDNEor2BW3uF6rgrYKhpe/NAPLQvHp
rfdpT5qlADlGvO2dgzWl9nok6OAytndkU7A2iasQ3vQSAa0nUtuRePSgH1OiRyqElb+eChJn9tGJ
2yUTpLzZ/MZLyPF7Sqze9cW3ow51bFO/pmOiDmjkeLM8e1AJ+MGQBZE2CM7yTIxo3caxC/VyPau2
V9NOr2xVFOFP7kJyYgxpFJlAe8/t2fR7QP4SFTsxdU4NsduANQc8usIN2Bipfb4X9jSF35O4oOWb
ViGiKLxDIKQjkVgrdj8zGg4xFdpIj3cS40dDQFqpEcdKaVbZ3zodbvK0w1SoLoO/iVNUdAlN/jOe
wLFHqpMAd2tjfMGHIrqWa/Iu38saUABovDrljDe//AtdeVZQZgrowxxEhBQkVtk/A7rnQl3SFUWY
/zGUQqlrQezUZsbKqgdEjwDqYJu9DRn13iiSycSu8giwF2zoB1va1PkQs1f84I1bkXlhFZI/6V3F
piasP6vKnfUNzH0SqfA9Y4SzS21pGk3+LkSfoPMw1xFwkG+aq34HG/jjGAy/HY12VX+icwEzbqsH
r4hoK0owCeA6CMcVJi1yBk74GSB/JFqXlvcSzeE2BYV3CcrN3v0WfmeKBAzxrrOX8BmggPIy+V3e
0gHxkZJCljfNiDHNRExpAy7av+qwl7KnRXVlKJl2L8tXGCWuUt8W3i4Wtz9zUHeEZ7K/lfwTkOT0
fP1j2i4rLeELy6pNZSvW+M+nQ3RGQibMJL8kLyGhIu0XaYiBDtEAZ9Nh+Iw5s2/Nvwfw9GDa7At8
axZog5nPy1yv0Aow1GqxQJ9ZVofYNeMnaHQcE5kgrCOCDlA0qfBy4AY48hcSaXu4szk7ehvGmucw
Thq1uLyKY+oTzAhYrtpLwr6sicQvQy5yto/aXbdlOtyi/FcSJLo5hyXdRQh8T1AnxxKyG02pfMu6
KdT0Ku+U18psY0aDCljVYtFZIZqb/vpP8G5GwCiuYtl3iMnHrHKNMkuXH1vPh5le7JYdREOUIJDa
m4jD5k52U8JtDrlxsuJyDF3zCuwORG+WNQcUNjk4XGEsb4kLVX63ny6XkHIpbis/cKVdEmQb1jjg
9RuRwESlvzIw3hD7wAmCnjXvtDQrN86iF1CjcZDwbO96odD65iOyQcfzx9GTJEdm/zrB5rak/IL6
fjSpwW+VRnzPOI35hA6pVppiMakyQeqxmjNcPpUbKQou4tdZLktGakeCYnvfnHQNSAj942Weok6I
u85XBfPd3Z3Wh+CAcB6Dwovy6oel4cu2dZbxV0oPBMIV4phcn1EqV8RkdKmHTN75xx6633wNFIDq
wY9wKI5BSiLZQxzTn+x9kTr38PICmpEnFExldVhQCYBYJKXu9sPpjAIb+HZy/B3ENyVh3+KI3iSM
MHnSfejOXGJAPezg5Jw2k7e9861YMrUb9b7WgaxNEfvZCccrbzBG7VVhr5+eP5NIIKMWm6wbluEW
JtP2umkq0F6GZ8Ny7WHR914WHqkNyPnMOPo7okdnlLZfiFoKaYsfuGiu8BrVNKYOTEyxGPWUxjw3
TiafNCtgrj5NJ6+HgL9W9k0aoBjzYHOUcfojKpadoNvb7deSfvBHgiXmM7IUX/0uZzlivv/IP9mS
cNS19nFlP6TOPc1ecMCtAfXxSghyB/MkyfRi3TniPZU44PN5sjMkex//3QUVqblNR8R4R3H2kbbX
z+w8mjQq/QAgVscyPDFoUVtzGsQWF5R1S10d6GHirkXPf13M4UM8hW+tQW7Qso429RVpnRlFCmfp
Ooa1Bsns4KTz0q30z42HuKdUV9h1SPRaQMFirQjQd/e/h3E3qZzGmNMVQHYyuSE3CJWGPXXgykmu
rndCnfovP4gA8UMUp+b/azmoX+fzk3bVIGaTt4Q7l5M60pO1PxCrCarN6uitrYxG5Y23xIpyp4Uv
fGx8OqsJAsuE/LGT8tuwf46FgIbnR4/t7jribXBk5RivLMrwQOuoEe6B1zP0S1NNCfR1o1/NtO3I
nzvKibWzBMRK1eV/m22JdnjdGIiufxF+Go9RlZAEBO9YzzRM5S648PrKxU7HFP8eGz5XrcIquhHC
1+nJ46jyg0sI2kO8XZmCcd8bqPdQdOip5dMOPOhFw/tmdUEiq5WAn5tyze+fssRwJqZk9j2iGavd
8iiK9I1MDmz9+e/0qTX4mE/vUmvdA7EgLzr5shN40BPTSJP3p8E5AwS+LYF4ssQvZtRaOM7NbPjm
DefIYj1gJCfioatLg4EVwgvW6xjpFVvA9CjgSAgk5Bi9b93/6r9nCUH1TVssIw8aszpCcfKNvXkB
GWnJ1cOaLIPxtpWRywSfYtp9C4L50mufUkq25Mp0sXdlXIbkohqSz6l5SheXcZrkpMVXP5rLLxmG
wKzNeLcLK+YbzoQGevXwneAg30CwvNaH/Z+UbY0NNLv6hcOcVxU8WvYffhs9OKcMR3rvG3jJujw+
ivkqPDmrqOp2EESoBp4HL+IWJH19SebjGyz4QggQP58rcFoM5ZF2O2sl41rKCRsfS6c5l3AUQea8
4Srjl0kdPkydsKV8/ixo8w1W+jVpchGO6GJv/YzX0aSU+gvJdUykOJT8TpH2kTT+0pokGmfejzel
UCKS2iBFwFmq8Fa19K3CUgJ5XuZNIXYtvVL1Bw9vhqufKV1DOrNTl6GUCKCjm3X2PM+sgRnhUZmx
p6qNBlIVXIUXEHLSWX4vrDbPPFtQGUtMpyh83oQ7KSTPsL79jEuWkEUTM4PCsqhwljB25txRxsqu
k481XN7v4i1YzgndpUII1UnTkSpTUsQzOJooQmMgmXpCyw7FGEP7duhfTPa3HvE0nbbVMYgo6Fe9
BSlgvKH7XPpBZIILFWyhlxkJtFudIl6c2xpgnr3OSIv0KevE76Kfl2u/1SA3RuofKxABT6x8CHiD
lXoDtTR16KDtlvbk30R5Hfs1cM39mTHBpE69aqGWxgalxystXAW05ZuugbGzFONBIe79BU8txfwH
LhPM4I6DNW1vOAfSbtUlyOCCbRRuawQ43M/eYeWAZcgb3jlw7kKbfV2LCxpSt8aHXvDusTNTIutv
QM5QmJJPj4DsZZYIdZ/AF2uYtHmP0pUOuPFX6lQwK1mzGdhUb5Cnuw2bturkSXl8js/QwsWa+5LF
nlC95Ll9CgpLtdaNacQTUGMiX8kMLUvjtaSaHPZ69r6A8RE50qQPKxcban/hzpfAfWFRO4yNobYL
lINDcj9GJzuPMb/9r3ed17ixQw1K4AkmREbuyfkvrfYJHIjZK3EEUaOMERsV4n5xEMG+Om3o8/1G
/wLiHrYMWhiQzmFD38F8NZUg+2gtTYJY7HYML+TTszhE0Q6bwFCS/mxsiWX+lk+UYwHd85cJNQTb
i0tVC8ki+14lTE+Q5FzBsPsvBL2OX6FxCFjhGqAbBJwZLK84r6JlgtF/LsSf5N+TyE33XJ8BSJzm
WmZ3RNkh8DipT/4i/+tMu6kA2986XKb+mJqs5TDroCDOfnbf+JH4s4Qh77mleO9eChdRMj0UjqFY
RFKus5N4gwfM28xF+HF9SFbpVE2zKjgSePVS9ngMBkEc4B66zn/Vzgo8gcBrENOE5OE6jcqMmtqM
l3wPMkmp8W+FTta27n5Mht9ok4hsA7paZxCFSpdSMlrCSqG4ZfSjUxNYFHtC6ouBY9vXgOc4paZV
Pmp6/PbIURu8EU4mzJ9X3aUH9LofrfUhlVUiXhNQs+BpM+IdU5Zn+QFgs2mAu8NbcISXPyCgiKnr
9VsOE6UkaJprjd+97OoW4bLtcpolASdn2dFeqoCU+gwjzk88a8m9WhhTH1BeoDElXz1J0m5oju1o
wbpQWOokbfy83N/zaNsHODsVF6zQFBG0/pbpSODcsDIgf0D9jm/PbKCH7+kiRUUnff4Qi3Janw/C
YRS8kZA8g93D/5bjPCyJE1NJuYpN37VkRWZGsw1/rUA0XqUaeh5FcwRNPf+pKpMvchhV7hHG3gx4
aLhBaqfxOJfPoqxp533KVIO+Wr0rCTfUmmlTd9SnXZSEtl4beOMdxG67wnyi8yY9zC1UhDJwvP7y
jmQICyJkhyWULkZPawJ9uIxo8Jw4kEXPgStWqq6G1Lpaug6ZbLtoxRMTC0djDzMg7T9gw59VFrKb
us1f+ZyPhXC8mMVGA4IdQNL+/G6XvdixpGA8X5CuJAA6QyRQkXL9pjiNZDjWY7w6rOyBn9IjXShW
tS10FrTIr3Hgrd+9Y0nnDyHuvIcWZ7Apq12F4qDP/q8gIWOMcDY7eYobB+dY5tlL2GUCYisZ3c8a
U2Fz/wl64bWup0MbxbseqZK9CoOCnknnUAmr9mWPkyP9qKX/IsI+lVzmpQVd4qc4zPm2yxOEnce1
BnJvna5aBRGeZgi/Mq7aPoWvmwxvDp+g+p7MeUTl6LwIWirliFYYuFjttmFj9csEKFznukzEW9ea
qsb3x3+2w6D1+HhCY6TtyN/pF8eTISo1YPt7pWKsFdpq2fiYVMkx7w8TNt86r/FZeIwEBMLJC9yb
ZtH862aQyi6ldAQnuvrM1/WXlwoLasFCfTkxNEAXH0ACEJay7w1KZw8+8Qq7S+vWO5/og4N1XaUy
/poRjwfPY9a/am+RsYmFfmmHXaG3v+qDvTe9KeRBIuNq8X4HBu6y7SGE9UuD+xVKr9rM4fcatcOv
Ifaazy1Z+xXQl6gL/eRBy+3XqIpaQOwwdVEh1T1x+Uc6jAbguJZh+OyZN5nhgERhLmGq9XO68JeX
xczrSt/RDqduNFc6fcG1BJQr2aom52WzNolQ0YC8TS+SXyLEHrVLd42psIJQzoYele40IddLC85w
Zx+oK0rY/g5C2YekAenaKKy21PZu1SErp5CPLkIozLJM6jRAPsCNV9vobD6tUWELd9edxub+OoSk
fVtSzqrOtMaCjwAFqEovfqvEyGHf36J7CbHKLGwzYHOs54FfeTviosaOadf1LalN1HgRZJhHCZKC
1EPYbvwxJ8kOh4FnPgxS9sN2ms58FwmaFqL9v4R+uqabvC4dMDtyZg/1YFU1U47jVrc8k0oABqU9
vbFIfBLTU/4AT+ikTtzN98SypeyB7sV2Xl0Bkok5fTzL7K8uJNxghKixNPupThQvjhGixXxxwZLS
45M32vQ2Cx+t+Ev5YQTePrk0NFWgyFrYXjAt3QksyyuaC1guBrgpUKQLRC1jgnXAko0I8no0E0ok
lKQ3svnpB22WZzZ2yCqzK0ddmlwgB/uEqzVUFfUeeop967W23D1wNwOtO470sM6KYztTJ9PAKCfc
qTOss/aUOzYPzKeKgxTRPlT91q0+pHoMZvMIJIVszE2zDOuGr/QTXvxBlezY9gaCq3RrhsKsd/Ht
aoJyX7ISzDCb/x1lcSwKFdnU6Pj60Zu4VY+8eCZN//zuFtYo98hdwBNqbTjX9D3ugnLi0Zp62qa6
02CutTc19Dhf6COoENWqSFQQcJU+dJkkeU3GbQH6qT93j/0b9YOlfU4hjU/433UAFlFfYvmRfq8j
E9+eEgjUe8W06AkcvWhXzIwbkKOSKhMV4FihMCiSYk6Nq+zPBeip/MSuCDSQsCwGyUhxR6rerziR
0Nn2l3dIjC7iYSatT2zSlCq8IOm52xkPOXZnln+dLM5JAmIMgVJy4Gs1PYtxvhVvVNHI8A3VUHW0
AnJYTVH2UhEMZgrmfPEQkfo//9Ms9b1N08KARyGQfz6j5Zt4Uov5EoN5jaseUlt8N0BmTToKI1x3
/ZuGQSVGkzf5+1XakbdanlGTFmCye9Fv0hXDnJ0W15s2bGir6GF2VsO2QIJHj5LnBCBwoHKmAfV8
bhFEKOfaWUKB0YNPcKO0oNR1pbNP9PC+2G0ku6O6pjtn7ZKAnt24ZlskRzOdfRceJuD9x9Qh7Wzq
qYFz9K56Zv/w608MRLuOy0HJW+4nFzQjWBJQiF/42O0zI6TIM5ikmMwOt/yd0lehkAA5zgUx8fmv
+LuQgfL0GqXkvm0WaHh/udyOhD+m2Lg7GO9LHUgMmhpDXxb/vhPx2Gz7/DFUicQKkhRlmznE6BGe
kFhuxlCpbG0RvkMfjdtJ+7joUDB65stM1dfY7XannJsLdJNAUUWXnksgFljyA1GoWBvmCw5iFx/M
/eUJSi7ogu9oghQ+5Y+5CrMVRI/WF/OEqlK3mWfbwoNEzUiFQxm5IJymssX/AlBIt7a7G7oxwkVb
Y0UC1I0CnA+6oQQ/sHjbodfIFROBd6LROMmu7B43ElOzoquLogHAtAl+exq5vDI8vPqIdLV9PqKy
9gUE8JM4UEbnSGO61HY0CX/DDlfve20YT072BYWTMChOwgLdJX2GvMvBv3PaQAPLv8ZK9QsuPwCk
2b0H4gytXxhDqFTaEqu7O17abg4Leg2kGKWCCWmNWn174Ge6SuckQgVRWXncyRNE+/Ve6afwEJqp
vM4o+pLLecmprKV6iaCw4KQKnc14+wLOe0AFhLuSeY4O0madLTIZXk1FHA5p8UUPDjTj0sPzdcWD
1X6/OHAtZ2/AAGaOb36Xvt8MNZxrfM0MgVwjmUXdBL10k3HP1vHo+SMdwjCbDt+nE/MP0Vgj9eqr
UigZzOnLfA67G22v5aonM4y6LERrEqSBEwivZNM53YjavgVcsSgtXErcTMhli/gPhLWIvc06Ay17
XmN/P/NJIQf60z50gtJJzCK2ift96rrvy9IfKYmH+I6PGnRXoHLccHYi5cT8RFxzT5IXg/oAo0Sv
PQl+oD5R7oMryGT7soIhpRUKagPqcizxPGYxQ5XnCdRYr0G6LT6hfbX3re8iVeIo0h7n5TE5hAUv
CEWg+0uWis0dpa4ThPvoFYAqxENxJ8QMr1TgQQpCKCUsd2O75LyOQM7fBi5oKyoYBtrX1tIrmJ8m
hTnX7A5TgOjhibGxmwxBXEAbku8FfQzag2/GMYAfy4cTDiDxs2aMg15sMPFMJuknSJ8R+C+qVOBl
QM7DrM9Yt+dVyHmNoFAlt92WjdE1ROM2M4vAMy0njNzIoiGgZfjy1YdrYcYGG4pXS8+j6QDZMnnL
LYq0knGpxCwb1U0vNkakO+zNFBH60lEBNWzKEisBpfnLu8L4PYP/MvOP1wsFIPwZWz1XBCqUfyny
A8uG4ON3eiAC9aVpWpb9na9S+TJz4hVJ8UlBgOvCyXpqO2Rn7jtlucrA+BvWgOCRCHn6ksWUV+1O
2AMD/NCPY0V8+X3HVPZbs+i5Tl2dVbaO2yvQl0k4Ropd7k4olWmB85DsvSE7QEeAnbQOX7f45DoM
oYY5WorjQgWCekVmtEY8cLdb4+y6lbsAKn4wzk5tQcttRVYvdHESpxqeCqlLI0FL0S7IKmnM0L4c
kxXvZkptlFuOoDP56zHfbuQ5eGcbEAVCjwUOUWp2/XJlBZulbyHqn2zfuvSSZJy5yI+Qp2LubAKQ
Mff2vSLSKp3pH3yVG8J8CW0fP7lTwgBuV6ux6rYYX9kKfle5Vic6aLhcDoLNVDJHsse1FVtm6cdv
c+JLzLseV8iVmXPwZIFMQinXJskBIAuxo0Sk2BIPk6fG+0mL2AN2onD/VDPQVFe5wjvp7oGjiD3O
gmJPkJm4x1KwC38sRcUTlWj5nVWV20yNRFrDWScfj4IOF+OWVryXUzQzlnQ0D6as3bZsbC4dIm/w
sQ1EUGAfWHYqdeg3rXQAhav2cfKhxEu2l47bsMfcYOF5+8rGaRejtEYBSu/worlfR9tV9G0W8+9E
nNSJmjf6+b3zUwb7j89p1xAexfBHkes7mKQOGKOvv1l3+l7gss4I3SvyWwmQDV+3FN9a3nNVi5J3
ITynUf80LtdmxuxGFMW7jlX74etMQw3368mkXJbb+WKgda6OlsiAgiF2i0vlFXTr3a/vCX7ZiLta
oTbPECeU1+p9ctDNbw2WTViA9i6KSD1RheM/tQf4BW0kd0V3HoHMG3P8xwvBsdhnGmMZqQuavhx1
a1WLeKXR1mPH6Apu1s4zy62oWvOC5Njn3veRXyb6L+KHA1vYj0pR6CNlEsCwgB22Itr+1EZbyslK
9Uw7n70OLRA3yDUtf3qELHGnansOglgNoAXU0CAdOZ+w8QZOAKnV1wasJIF2E0zzCGAheth5gD1t
bDJD9BRREZdXcENcF6khOLYeASEQMKUBb/k6PfsscyXDsAOa6BFQnqqvC1Zxhpf295i8xUqp8AcN
tRm+rhDAoevYP9Sx1O0tJmvzcDs9wXXRD5NxZimq4zJUAioryP1VVeys1IaGS0qAnGo+uMwGojJA
0Hclkb3YTSaG4SF5478hVroqH/+6DUKCukw3NYyMRjepQnPUWJuZFifEDHK8RtEY7eQ6bF1WHKUm
8vfcpfFLdjJAms+jOyo2VkRz4T2kwnKhxsf8wRVmN2e8UdARI17KzjkOe583ud7ZacqNDq6RHYrM
RZmjGNdoBJfv8ZnJ6UAjg0dpH0Kt1wC65MGNIy9FCaxkf6rnBlm7pWcagYsN4kiEm6tQiQ2FbzQ6
DFbxiUtJSflh+Rqo/NSk6b09o8pQ08s19F7/HkNN8e+0TUzrzIx96aYXJsH2KSZjGWH+7PJOaawt
VoNCE93dNQGGBDCR7BT++R/aB1WNsNAH0uv+a7oiatEDttSHGHzfUvdhkza+DABnEP15VEIpWYUr
ziIfKqctAI3E1zUujxP4A9B4h5N4PxX1a7PyrojbAk8x3ab6WPZs1TepupQSZdKVnV3hO5pcysU/
d0tyLPYWExlzEi7GWXCuBb7iqv/TOKpFN3PVV2XnTHQU5a0/4wBDiR4m4g82pyl8RHurYKq8Pwfl
vUq26z+a+fcPecP1mnwYOEbeaqAKCTsYHVgqQfNRhrdbpTm/5yHTqK8Y87vf0qjo83rOXAnHW2ut
OmS1NIWRj80b3DvIOjYLTsP3ZUPcx7aPlbXaZkl+rNq5nyNcFt4elGE6EBkqB0eLs9+F8uzWvupN
Ch113B8bENyR4fGOLFUx3BDC3qY++NCbjqpOuxXDGSqPlyFXKiF4eeepRd6kpFYIau5cJSNTvX+m
wGSt/QF7gwrD+lE6L/+6KtVsfqlvgryBdzZs02gUJv+UUp1Ip7e6i7CDOstxbqs8Q1CGO6Ea4sUh
OrZ0XXhiUXZz4XWYbywlP99mS7YfVrZZNbab+vbsdhgxnFy3ByB70fPStdv5Mst8WCGQ3drQfqZS
AxTWhgV3Ki3BNcirYegRiYqHSsjo3Ipz6nlFCCvWD95bks+0T4fy9fdpIDGgIwKRAQTnLSiI7yC4
6mbhXMe/T169RLLyVMlGURgTWGpxtAIE24fKIgk79ASTggltodRyG7PXoTLmICi67J7DNSTmGytO
dB+lFwW9DZKNT0jnFntvpObeMusnoFOB43yzK72ATZ+VWSpxsyV2vR6nmdCKpDg8FRP3MEt4J2PJ
IatCLQDGofJVJlrbqTPWoO9Ul18dfeOc3eU3XQEAk4+XreG1HblXBWToBApLrMzAjcAsE1M7orq7
CNR8tmxoENeYP8d6/Qhsg8YyA66IWUNl7BceDsB7Qr7Z9tceZp0JSzh+zow8FvE/eySKogLg+7ul
JQB0M/q2xrl8NEBr4jJQnEw2iecEWm+VixJba8aFZ7CMjArGyWEyU2F8ykQIZzlA7gsnUx1cw3Rp
YyAJi0G5tCODis9CSZDsLIehZXr2t5g2HzSeTNgyEWB8HRg9+1naQYXDTVzZD+Sd0p5dOdiI4rFM
S5+sfDMr5pgUtf0K6X2PCRCm2l984LhL6Kw8D9oOq5P7ZIP2/WShCZze2KrsnibJv12aalU18svo
R3bo1f+qWSacpcDOjK+8LnMY4mrh12bb1rP9Dh/6Ahvujwy0yOVOF9Ogszw6UTEV0zp3c5YVFOVz
JL95DyIMOqwF7jPYe5hrqd/xfoLSaBvkbkTilW13GqTouv2bYsz6hNezm/xw6H9BQONUzqWsiFKG
pwxBC/ji6k3zF97sF9enzffSgQg29rAvSh/zEP/4D72dWwyDznz/eU49ZYqZdzt4FqGTFoLdMYV7
zmdyP4l1abjdS0Lu//e3+uHLIRklmtukUYToIkVhlRsUn6yZD6oCVWvnG8FF4C8991qDh9Usa1iP
TPmuJ9qTh7BLUNm3+ffg1BTGwrvTF5H+ATMMS9kr8Xp6hPG+4iACYddkgLEUFMMCz5TOIWQJR5Ak
eBZJUdNFvqHlOKPEiwm1JM8SmADDbSE1VAn55ev0IDjhcciTAxOEZAQYJD7lFlf8IZFXYjyuH9Pj
/9FPerzcOSkfq/mUCs2P8YtIJkbKQROVoW8FDxa57+hNX/loqTlkMso74xX1Njb8tBcOyXLoJAJN
Zg6LL6xwF4gfwflhACtfSwkpX9MOPNeD/IaPlghV6I7Cdyt7XwIRdKKekv9NTroX+cdYWNBJ4FJI
9soDvYjFi+MuFfFQEofvRwV2hNYex5Y/a4J8Z0g72h8QV01k9TKeFApfzzoQQ026drUljl5YCIiy
HepL8JzwwvWc6aIiP5nBWvj1qMx7DOqGSpA0NaRNhUo1XQsAF69bIJvJnDJ0n+2vpIPQDenNu3hg
ycLW2VlStruO6oHaFyQGlUrsk1tt9d6DC00zwrXGd6+iH3+2QiMQcMw1f9jUQwEN8ps85HE3XNKs
d1k7q/k7rEy1AQf9C2amC+2ZWn/ZH0HP376rB1PjlYTfj3ADKW1ml4Qpb8x49fkqm1fv/hagZ1gQ
4zCDwXKibs8XJXA6gqsTUMSVOcvGgCddpI6qBpuX8UIRodEMnf7chvIfQBhlU+m8+XMmDjlne/oR
levpHor0XMR3ZLWsSCCxoDPftG+3vS4R0bh0CDRDfc37gQfqFq4u9qKdNGDCjUaMYbWYIVB7VATn
hvgOnxlBg1xSvMTMsTt2skW3XZaOccyt5R/ReAnLEYpSjikbaIA7Y4pZWvlLM4r7Ktn7W8/rZGpj
XViHJj5+t+YgJEFBKlMEX2CcYtfgtAglJDoEC4AuInQ28mIBDNYmn7rxj179T8A9EKrbm05pMhbp
UbQFHdg/E/xHI+LFLkhlyeaqUreL94lkt47KbaD/0GC01zzpeGVNqzXA34qVO8F51OXuWPv3uFcV
YUldKzAZbQX+zjh6GwJPVjXcLOxkuh3+9Aa41VbmS/WI9r0JjcCh7bM7xjhGA3UVU/KV+7zhfaEt
aFOad5aY0zpgMoDqnwwvJkdyZT3IX5TYbEvVZ1sUXDjf56cbnQiYgVJw66oi8woz/Cqn71NAC4WU
Dq4mXZWgxksXBz8u9XOlgiDTkNElzT43kbfbOAXDnewWsWuA0jMby8TMW5BGt/b3wAcefs91ECYy
sZ7nrRlV8GqIvhavhv0o2ByCvf/BD7uOBuu+xrhYNMZQDNbqLS3Ff/FHl9BLvs20j0UP+CD83Oxs
fd4GsGiWoqCQODafTW6KpxHOpcK2VjXOlTWjhDUm7rbYBlCfd3SP6oiUhF8W9htd2x0EIi1BBJCv
UGyYGQ6StRPKgdT4WXTxZJhurgrSh92OAVXkxzmREV0yLQ9KPxKhm8aMpDfMMcIuuY/puMkbBb6z
wME0zQp/aBtFSKc35/+psETyi0ygFIkhA9vFCkS9Lq05SokyPGmfZpkZwyzMSK/RNRol61KBuHJi
vIZx/x6pcl0cJTGXWoytVWv9/mqR1CeCBfT0UkeaoXMuAu9nlEFeHEWvrBzxy8cfFyPWNLrjICna
3ruhUu7Fyuh2pPgRcDP4b8Fq1gv0hfv6hdy3onkj70GCGNfL+PkttvJ30ezWcJD1zAKWktR/8GSV
Kq+DL3bjgTOJuU1H8Kf1HUYwrUJpQznUEW+DhwNArv+KLX7YA0JbU5N+GnoVy8zMn628bfYhWfEm
sEJ/U61pKl4jny3Eii/4RZ2tXyjGLYCx6zkERQu7XlqRcw9q1y+uTHhmYJwGBvP14Va5Ruam0jPc
RkKxkir3tY6j5NWzZuI1aN+dWtF7rlFDYHWWwdiV7ynUO0JR3aFCamf93Gx+3p1y6+6GupvMOhxv
kvNAvRXHKntufTwY6rU3ftyB4E/yYQPMFl14RuCJ1w6L3EwcYSSg/zPQzP/fXasR0Ixzzgd2boqO
9rD9hMslQWTqe4E2Sxc293ry3tt70LlZyGlvTWJwGL3qmVOPJlXqAoDgn3z+nRnLTStdCSuBrJG0
LMghXFhDr9AC1flCAhs4AFGO64p2j1ca3t4lyz8Av36dODRykxjTQButt1jTq5N/sAlMa/GJasxR
i6Jhc19sDwIKKzJZ0LrZlHab+0W0ceuq6HqFs4t4r9m6VTfSh1OYsY1HnkRqr/HsfphH8hlwVWmL
WvDdqI3FCe+gfxpCpQ250F1OiVYPxRU9/6AXi4sGuBNsjNSaFmhTqOTB3DMlXvf/gAUDxAWEtwCa
Oe8tMGdrFqDzbevT0wUt9u1bQRUx9rk3k8pugzvbV/TJ0TQOepb2BAmOvhPVBtXPatHras2g3rrY
k2PvGFSHXiBKYGWbioR0WnVQgqs+bhv88QVah0fS54oiG84o3OGvKjs/22KiKhj0rxL5PVbG0NJt
ya5UGVyOHyZ5AE4KZdKvpHcxcTSzNA09sR08fori7Ba/bIF+gu9emTA4ZyKgDeRKIGDWNaafdf2T
5DjPtXGAb1OeGsEbDIVbDLkwFsSID62ArCgmW5Y101lcd489TGizZb35hI3LcGMFXrKFU7/1NrwJ
VWApsaFyx/t/gBRFGhhelPanKbSG/V6s0f96nCG4wRNuGPS74KBu+9HaDM4eRTs1bhRpkyt1dFmN
meH810ZWHn5xw4usVJChNCgUe2NODyaZ0SZcIMwVTO9xRtYrm4CNmTO2hHbwXYCefgyySruC+1jm
hlGD8u0pbNKLsZ8oiQ/dtFoyLbF/9NdQMppyWWu47H3rOD5P4dctXlLeok6ZcvSWnsekG6Se29xE
i/nfMqA8vnXHfzqtx6YFX1D2H/AKeYCqaGMUMuPAcPKqCgNww9/Urw9sYwgyuLL4tBix8FOwr7UW
lZRVEds2vdlJ0zz15HFv+3t9sPV7leAfh5S86EhmdQqs4WwHN0PmBkhI3tHcNCugXAElB9AZ2RlH
7K785r1j384qD3a9sePPc7pZdugh1HMa5+ps5lICNzTP5266gbaSp8p9ihfgk8Lk4wyHFRTCbUfO
wz/cWCtA8K7/8Y0pFDOatdJdIO1wmSawx7lEi++cInBYujPcfNkO3VOBaN+72lwTcrnWzbIgEkEd
4cs1OqI9P7xrFo4mqaeVqOk47cSgSnpRAImDQIC1pWSy6qCibBLRCTAQjyvWljTg32U8SzcXFfBs
rM5wZ4yqAZ5wbyCVXV/0zM4Lt4V122DxjL9NSNXNVU2U2CQtg5epm3LqDGeJYXvgP6yaSseavaeL
Kjm+8jIYiRNB3MVHY4gPEaHVfFXIo5iFzqUSBVt2EQOiopPdtN9pN+9qZzQ55hWpKum73UhvFTCU
48jWOVjw4DQHLWYc5mQ6xZkb0YUl5en4sRVnocAfpnbXKseDWhJUCZGdd60FPCVvXOuUWd8vyMJ4
2+zmfrRCL6ntFF5HfdrPudcyiDnkbqg0aD4VEfh0InzFZU3T35dsQUa/u90UY2fpjatV5eBvBew8
57h9YR7lkalzrT4ryRij8zpsIa/KktOwKWW8/hY5JPecKsuUhTerSvCFeNo+iSvlehuKpFdHyPAj
tkzDzS4PXuv+FCsmAnRyMKUOVpaeEI9CwtZCzapd2pz3vDx3lSiPsEiAo8Jwpouc+v8fTe96PVPP
i1uPmGEPOWNy79iyHXy8akFihetow16VbJWJDWl53sDI7KZ90nZjDRc2YYmj+Bq1TXhB6O70XY/P
i0rHIZMQrxUAgwAUu9CKte9G0h4QLwKPZFm7BNYZKJDde+IhbWN3mX2FRw87X7ocXxd5bhBKRWuO
GR46RFldDCyZgCeuqVAui4nMiL/PhUOzO3G3JfUSSaSZyvSOxm4GGxAJm1QP9ThTArgbwSTamCuz
3InnTU472f421TuY7L/N8/JpfqhQDSWcdJDpa6DKnq15DkWi4PU/3b3qdME2x0IVobupJH6njzp2
ZeAAckp4DCFwFWX553S/Up3Fai5qdbkaIc4gQKmyPJU+Z8s/koR3LpLvTUPItoY4+bTyr1LfRLZ1
5eZtpCl8lZI6vlNuxAJTjZn/I13zJNzWbABj5ogMqpyFuntfJh9VSR1fcNPuuCiKLfPaJQFsKBts
/2Qzkdf2aAhjvkd8nS9Ft2t9bvoWXHFqUNELG8etQ9JzAzzXAx307FP8n9c52RyAiHlDiQ3x16PW
rH0Ti+dONOYhn2X73V5K/6abHF3hQXlvz+4TaalfNm/HAKtLj9zqHlTDbxz2jo9sbJ2gA2Fje7ld
O1GR8TRs1P7V0JmTgXahYz5FzQYNosvHwGQU+2C5ekVGgNq0N/ZHAzH5tts9HiddDvBx0eP/78PA
QyBJt4o84KfOh7fo+rpuFc20kshi0rdluqXV1yKLMBBDbWQDMqx8tE/W9m0+Ww3M1r4QUCsHG1e6
SfOsZOfJFHBSYTmnmUfoX/TZHXQMqYhK+iv1w1yjWhdfl6XOknRl3n3SeDtVFC2XP/SRQsYStUL1
kwWoSnmwCuv7DxGUmOJWyr5v51RTUm89+07i+bTBgpY+2kDvuARe03WIXvCA2sN7UfVS7GbZNHO0
u/qAt0rrxnOLpBIMimeqPyLbZpobqzD7NLbrWwZdvjEOMDguPBWaPaUUI/xwjP6u4zGdqpFo7mas
HQhiIFnx/oaZ4Nn9MTxlswJxmvy9qnF/5sYeMWXg8nkAK2icwKdS6tYziTiTkTtKJF1urvdWEruf
8xqn4Q66zZQ0qesA3614luVmhxGytYmsKYt0wGBlaNui+KQZR9aZ+AWUZ2baz8fTRtWXo/KXD2U3
ZV7WhaxztnO6bwDL1niABwl7h0YOdEvgPl7heTrh8idKe82VqcsxDH7+Dvi/cU7VyFliCBKW8acO
UwoVZLMm7mSxpW3hVdWrrZp9+E3LEIVj7X8W1sazKbgWIR4LxyPGdwdxzLq7BTHCmtNX769B3QJL
+DkXkMF4UBk+pHxZJitvIlQ9Bw6wFs1gJ/zq59PcDERCOcxhDHUsbzgGInHSE37WgyuEGYCyGAQ5
Hh6N9PR1N3yqOso4JlaciIvc6ZRt05fdPxwOS5BVvrYSVTf7puBpDEPQsPkSRxAWehJtN6GbCciv
XTnTHdpTOPXzgrdgQkX0g0c4mLNGX4f7pNfx8Bc6dTJROruKLO7Hk9F4bVDJ/AmIdXe8VLUyiaG2
ZrjEZyeFKcMNiFByIbbg3QAso5wk8uEkS8PROclzB+dzTFktPyN9hVbZ6ZpBkcyICElzq1U88Igv
yXmqJPeSubW37yDidRoOk1Cn76u6f4QtPsUY+EEswBPBYqExQ8DJ7DQKEhzGPqodjjAYP9PsViAc
4ELN2ijQhpzKX78J71I/Vr4MiPrX3U5yOyyaydiBy8WxmLkgIsWUnAf3lp7KaU9LHXUWWmGHdgFr
zoKPFUJNfl36STZRxp/MJEM+MI/jN6DL1DKfpqq3Y9mpxxbSZBwjWtyi4oJBDN61EjRDXTgBiYt3
Wf08j+S9mKMkQv9Q7RR+vrDK8v3bSx+/2hiuhfQ3e/P+J/y4SlsEWN8JqZ6iWj0Yg/Kj8Te8DkVq
KYuQ7hfAxR6tmhFiKCqjeF7Mf4+cv0baX2q67gStgDH1GBwTrWhPYxxLA8ibM3B8CwcpknEJ5MWb
yUaZ2D21E8jzQC7YgAfciK2I35y9cMGlaDEODAOnTbMUnVoPast8DHBFM0/0wk3KqF+1TIfuqfYr
i7ezhOiJ5PT6TL6QF0zdeyYcCs4NlvE6KtYsHt5/+n7/l7OjdN21tDnw0dqg4nUUkO9dWj0QI6Hs
H8ePMyYCu9Bn+ahM4ySuibNHxUB5Fv39qx+pLk/+k4IWXCtBfRlM7wvdEcZ7v8RHVRXPus5lBdga
KAVXZz5WFIydrmAf7OUUCzG6EBoMvPskprG0El0LrJivP8zN37O3Lu1X7xdue11EibD8qWh5Fs/w
mm8O82vHBNFFlc7N9BW9k15btW2kqB63T3q/ToFAVvujKQYlWzXW+OUvOweQyZiAIR3aT/0KD5ZB
uEdFDrDtFREgYHEKm3XuPk7NfKpsyE5oV6Y4WzKSAlbftdbXv2HQcoxD5dHBmojR9wIuHv3jFdE3
rUj0+G9d8sTkHAamheNL/pDZBDfk6qI7bqMouVyBJabAPhoqLIK+Irza9z4QLABrtUeAATYQFupg
jBSfuDYSjp1VEYGnnDpYtCJCIt2XDVEWjI55CuaxwJRKKMWOQGmccPwKA3zkkMeoUzqcFWD+gnby
ySQulV85bok5MCv/EVhks9Nj5TO2OkxW2PqULoW6hS9ZmeQd8cHq5+NAxYA1qf/etH42cVQnnZdi
Y0A0o1+rMptTu3WGPHacmKOgWCBWOFHSE+V+IKm6GfgOysj8ey/NAWNpcmgyIt+6D2VTOxyuLsr3
HNRvJC3pBIGK+K09Ac2A/RRDYmJei3utFzgsKSO+w9tkws16zAFqaDwXQiYTDlqbk+if5vu02Q5q
hD2Kp2+griR55skTS8ZXdnxlXXqRaoIrxCfdff9iDGNDRrgPJzs8IZJaitlL2ex3GK/JA4Ld9NzM
Jx+OUsdW+HQkVadTNTcPJ6OKgxvcWK9pojLE8yNGMTxTlL2JOYgnMVz2ekb2gVq8aNipQd/WvLEX
SocRcO94V+gzSKMS6tYLVkiLBTzVS9SVagYMvI8tCnyfo5FWYE5MvoUi9am0QkjVuqY9ILWxgT8X
wNBZLCGJVufJJrhNhoYuFCXO2i5oM09UpEUqtvlfugDdQuwYHGJGnezakfyb3KHIal4QErDxypUY
oxbYHAY/8ac7IMFHoQZ+5+uToxkZsvF7FAuqWAVSbxqIthHyT9z7A1Ci0AQsQ05v022XMthAIK0u
SZQfYcpp83gWL7eJmB3SfIdU4ulhMqLM2+IAvwv6EvP1SnWjY0/tTGJ1fvnWDyQDyiSlIP2Aped0
Ukzz7SrdOXmKkE0MJNZ0d2HlXV1y1c/p6xPVqWvHr3u2eHI97kxwmQhAgNauAGqFJJbtZ8odTxOJ
2kT0z+1MkOn4B8Gld91R2Bcf+TkMKo1dz4N5oMi103xFOwxUsKlBB25jqTw9JxRIh4BzTPXT0SA4
xBSpqq4eRFRD/F+nupVWoy7eao1rryE3131YpF/d9oVAdAIZET3bEGggSZjDJq9Hodee2lXg/Jsx
77OrhmlMaaADHz99tbniE+G0vZyutRxnrLwXCUjHNncqGOz5nilxal/R4+T6hbvotPcG77/o/+8P
JjXPwrxmBMlh2QcBI4Tt/lcytHDoZYPDXsZuwhJLD9J+4vWfGiaTdoyd8GQqSkpSs8ity2j8OJ1V
SBVz9KdaYDnp7fwbhAUoSEgl7Z/WBfQDuwSSOwvdAE4M/z3b/V/ESF5hAekjqTz8gwNftNVhmc4T
wsXi/6TQz1acy2ZFS0kb/QwxtN6PlrkR65/3O7whg+FXb9Arir7VJsSAM8WpJNPS9ncy3Z9XrWtb
5cwmj4RTAbno/7NdboT0LrzoQBhPN+O3i5SLg4rT8HHGVzbM8tY4Q+P5DnAfxbR06BjauXyaF+7X
wd8yGsjrsvMFUoJ5eC2PmSSVF/sw97G7R88D8m9EtqRiYly53sN1lrTViVpTSfDtksymq8u57LGk
whVFeWDPwgQ554vzhu2TyQlWmbqzcNT1O+ps8AEvH9IvlFP9BKzZstV6cZdjxldG25FqBoj7WXL7
diyMNTxcarRJyIFY9EZrTtlVIc9SBIZjbuKYkQPZPChPIgrH9jNmqCkRpCnj8PSWShDeJtmyw7d/
rTIwSDwpqaTbr1mhJqnAxw/AYSrrToxEwpk8iFxbOPRU4l2L2Q647MEgxikHy2RykHUPuo8gkWC9
R1OxEQhiO9S8KnJNMdwkKQnSe5nxSV9cnsEzryeOSv9qrvSyhyN2dSlKAfJnSuGU6h6s8LUPstZ5
+5qaqBh/AC9ASOJIY47MUL1ChXiE5CeKyzLc48XeTA3SQD0dfJfJRYn4LLKMXYWd94liNhjD9EEo
mNvnTTGOJy0Zhs390fNYqt+bUf8+tq6ii4Fw4BpjMxiY6Bdk4K+c5Wnj/FnL5AyQi8lpbNJCsxRS
81HAinQrGjSicFy+Ga6BycLMhai99+qPt+94kaWCdts9Jh8QGNl/9DshqJy1swoXtJGe8tIRA2xa
kUT+xnZ+2nqqKgAuXtsIHQyjnqNcU6ezJ3NJuUnYMn7i+TZ6E9XKOhfVaxdA9xTBNWrQr8c/nQ7Z
IBixiUQqN+F5emVUhr8PLmeVqpaOG1GJ6yzmPTbnHU0y5yu0daGXC6XRTg40t2JLQvRKWuLT+YQE
oCqEig9dZgAkpzeTC1hiCIypepjZmPN5WWHdQcx3j8Auz4LLE4EyrPTRIHFi/K+Vs4L9phXaKBP1
uKH/PkFRCrankLY8bFIP09dW1uBus+ApOf5332oIsiShmVUeEmm9OoVv/M/17poueB0+Wr41uZWy
yhQONFQDd8/QeSkJ9y7xmnK/0SmQcvIXAEheOuoOefo3RpjzqAPVGz3p31TfhGDsOYlGeIbMNZ6n
SAQfLmayUsy9qu9GkClSvP96ZbyZwrEenwTHrdr2qtixPQSg7Oksnt5kS+cFBV9S3QLOUSKrSLLn
5xomAyDnsDtroNxxvm5ubzrGqIVCn1CquyaENTOrPHmiO1C8oGIwNoQLjkzrQ1TdCfN9JUFrJXeP
aPlTJLF+S4RLclOJoe1fBuF5XfKUsExrnkZfpXBkYqmfKcf3PZSBPPB9vQGUfBjU71UjYC2ZH3Oc
4ZoyTwD6GzPp9Tg8/Mhp8zZFkDN+adPuNhxUx460Bji2IVJ/KiB6IgApVQt52WvpMBxS4k2Ki0B2
Ter89G/7c4+bqiDckv6nnSe4MKUZAv+8Rn0D5yX3ixvBGuoNwYow+99LcVk4X8jBfEuTAVywXavl
PfXrVPNFSKk2YPsdVDHoM5Kk4UMZjkALVzkUTBqbwKO65AYQugnwSGX1388Z32ZCyTTCSqK1WV/b
hjNoOGL+v0aCJyoCb8YfqmtC6ch5HVAhPQKarWIgHTYhAxHT/VnQDFwtQuacVyZLo0jFOcd6L5Pb
oF0aTa7uFec8S9YlppWkU/jMJoWXkAL3qySxC6NekuAuIAT/83MRrSK1MAhFPj0lxGkCq6rs1DVP
0RVeu7na8vbjNv1QYl4uRJnEFh6BlnCSxQVIKQYZTcnn7F1gCnxWgW7KHCC9VCWhAlxyfy3Q3ZUV
hqkPjT02iyana+ReIWeWat5NKsD8VOIAcVrz1/MNQbIby5MsnsZsHloa3PnD6CQ0+uAddK7b9Qkl
VbWi0OgJOJZ/JOSRVFh8it7gPmUbgwwDelb3YDlZAdsbL9wf2UuL6TD8+x3rItRXXW7n36PhiCEj
S9WEq4PBTUT1wu7w0U4cQGibTsX16OFvO9bCFTseFMprFqKMPe0/BbdeU2rNPplnkvIam3j+sLqY
C0cFp2UvR8o8pikR7NdT+yMOND2Uo3G6IvqyLIBYuGt5aLrwN71uJEXoVtp95KUyYN3k4Gxsxay9
T1bA7fHMURZVFV33nghRjCzLtM4PlXeFz5NxD0Zpn8PD4tUgcMpj1ZyPoTdXttFYXqBbIXG+dDC2
U87eyjMY70wrScNR9DuJQStGgO4HHWcVEMMnQqFfuIm/mU0LQCyg4ChiaE4YdWqb2tsgXENEa1Uq
S80PS5+rj+ySVhOrA3ErqfLho/yJcsiFZFRNSn9tOa6smL5jYX80SZr8r1Bhb4Bn31rZMSHToJDY
bZgKmmkDlTQLTf8xJMB4w7wlxF9Zsr9/hSi59rLFZUndmpmMzFGVLhtjeCrSDL7mWp05cQcLRFRJ
75Sms15JSDXslfc9EmumzJ3euL4XPdkvkQcWS+scOzPe+i+WFEwvGY5w8jpjLLnL+7C8uxJ+RHfC
B0ufbvRTsCGhwFzesrzmGfXx/g2s8Rtp6d4dg6NSXuODozzj4kb70s1dc9krdAsTZhIJCenYYWgB
YJLOiV/PZB7QnyRo1uPCJtr0njfhUPlz8425rBwJZGkt8pQdQh9owrnclxObDkHIjTo8DC/aAeOy
fLZlKbXbATBFENM/zYk7sTqRTMfa0hWiG4KY1H9LeVLH+3YpGdjNVLgrlSTiq9UhMfN6L+JrZCN0
bluJtzpUlfaEkbhYNMJAHqKnARO8kSWUsocVaWhoNFN9VC8PAmXQdBg93r9kO6FNhhT/OZzFrLUb
eD0Hg6ErxII6jB5dvI5r13cCJC1l58Ax/OaiguwtE9adxuOaNMN+KghlHOdkLeDka9M0lN3A2XLB
7tARR0C8WdTtTf8Je8HRvdikyBn7J7gVAHtRV4GrGhvtDCTBL17UuffcvLoj4RF4nQtVmPfKp/b8
oVh+w+UaO8V921pLKK8yD6P3M8bfxb06EKa29s1GgjnbsBAcmMRGVZ9+1BtxuO69NaNsYA/rf4D7
iQW7ohS4UQkImG1YIeCS9evBM7RGuxENzv5qXS82i0XmYjgiFD8JV31A2hczam7hlOUZVzWs2ur1
Td1XAxBT3QLToq3Qp5FvIrB9dXipSBe2nI/B6GF6OJ0bCL/Bqsgmo+1Atvq3XoR70vIV/qJQlz3M
3JWUX0aj0yz4caW8YQdh7+MJQqbe24tyK/yfhE7cEzvtCEzEPQouEiiW4rsQU+fgqMbYJn+EIjtF
RuAVWsMm2sqvJ8PrbMrdrBB8V3qgn6IKFiBYxm+Eqw9s67CjE9OAZf7IFZr/LGERgRFFxwzWPnXw
+y01WFTDOeDSac+3OdW+nIC2sFVWmEHQE1f30I44PRYZbZI3QpKJq1GCPq1ylEKGuQwnA0DY7vJy
jb9iQVVmfxqg0JEjGVw6J7H/WRtKI5KINnX3BawtJY8VWYqvsaOV3rlhSknzlG3XKM19bgL1PmDx
QPBVuf9F06x108EJ/KIjGRaLb/69U8lNI8VwaU8C5EHsiOPepZP2fD7J0MwlTnytSxQz3vrdKDnS
B0EWwkI8+f0GTUxoVfY2Fxykz42vBRi6x9qg90nZNmGIXgWURxsHrAyjsj3NCw6DliPDF8+a9C8S
9HPpdWnEw/Ht2wVhgZ5u2M10iCU2xA80dpSrrxvlkEbq9BEIRGcMf415Z+bUOgd0SqNioMeT0wcP
LOJaVdapMz8hM9eidbHCq0BYDeSS/I1PzxglxO0lrDWiaE013RsbqH/AXARzwVClrPY3csnt+1VW
dTmC/E8cC+yTgKlIi5FXQhHwN8uqAhRHhMxFdvkjk0glh9ZCJsUse758EBLdzLOovHOIVgiu7qLK
C2aq9i3Vx93v+clPVP/ZOKpvZ0C6qcln9RyxIW5uKM4O8aNHhwkfryYQQS4ALkC+AMofPO1R8yVK
lXnQuhITpL6VQfNE/IvYWGNHk/ArXBszHiRibqxiEaorgjjdN11RjXKNnWl5XPl0hVMmu3sZol/p
A66N4StvX3zia68WwG8Hjsv4qcOmRLJ+3iyGrTuLEJ8SbkYmqMRwb8a5JCt+kcQY1X5t6CZyzvqo
rMXjbyezYVoI3nHkSmEwSgz3lpJulX+BMF5ECUlmECz6M/GGcm56fcBsUFIR5b7STNX0QCNnzgmb
THnY8UPA5EXnKFb/XV1UCd5Ax9VEYJrZJobR6CmuL0FFANYSh1qjD0a71lTPjMeWD27yLEr4jAbr
xH/JvOKx0kfZLzayfXqEYvbM5kW4AH1E4BXZOvrX79jrBLB+9vzEpWWDLA9Iz4zRHnEzZJzHgqys
DRcbx4bpNq//GZYCtqKWKNGXsAAcl1FcN7BFDQRNQWt32thCna1p61GXgmkOzczLbLHC2WEoTMi7
T2KPeEIOp6Snoir4faWa0QVByzhKQa5iJuwqYSxIqEq/oyf5uL2qu6I+GMGYe9qdO12II8a1RJpS
G1g7LpYE2fixI6ZxaloYziKIp8UvA/9Zknw0ei5T+aVZBybiyRuUieLf+EFvnB1eDdSMySoTbcMH
LehTMAErbZTXHYyGrqxru0Y+iaEOg7ccyE/TVBlIWFrjuKfEMO5/0w+omug2PHCxf09As11Sy4fJ
41x6zPCnGeErkEUuWHd+1sqweMsRzXAUqHzMYNMsuHxBqAnQk6Kt7p1a+aDK3rpp7Uv9viiQI+x+
QO6CQ3+fTOSCof5Aijy9RxYXNuUZrATxgYrMCW2Mk+aL0RYEJUXWJ5uEDMSyU5RPAGgJ2hcxTreq
XSzGZYeRYsoeHiDLG5gNy0ThRXUGD1S5v7DOyo9qHs0Y9ZlvUHGkswBYPYXSLI40MPFGKN30ASNM
+VnGIZy63nfG+bAgx1wHzzdOk+HB8iB38EbBprXVrMtNpGQU98Qh2mahyb+SJED44/Min0HZfIbU
Q3Uu0wrhYpoVveCYq6BqhrFnRB1I+GkxnzP+Lre+nxbLSapMUN18hKoHWIJWBnaFTB7OJ9TlPJ4J
POQyjPrm3h/BVEzZ9BJgFk5ZZo4jDcGUxIGLoTnYHAbCJPECvBDZzpVBFlW982Og0xYG2/CtS066
hbwK2eVMwpnjjZla/6ewR8mn/MFCn+ba+lebPIDkSbGkeJSLi2i8wex9PZfYREx7K5fc0bPslEWU
T3+Izxv6Bxx2N+NvBhceSUMgouIlyWI253CaB//7QHZLehFfVjug4xGDg/ISm/BanuWuSQucEWoU
7ri+Gk6RhbyC5nhxtT90xiRFyEmqb279Fu+KLs+f+mVzBAZ4laytrKc/oXB7qGAZw+Lr8hrsXSRA
4BB11vOfo+xUR4wUP3oSrtH3SZvoQIjquKk86R2SkIYpNdHnlwuS+tsqBNTEB8dsl0//GYjISQCg
gihb+K/yyQknTxoNSxEsPx89/8lEBzpCRJhy8l4BnD6SRL1Tgiic3iT0BX1CVzEbXWQYff+WzaE9
vj6bi6YkO0aOlx358XRgWoz/t5D4+DsR8hUJSoICooUDnts3jlXb3umyNFJJeEvFm9jfonmbM9Wg
MprOoc4y62ys6jbOE261FeQdaHgWSFddDH88tyCDtjVYGeS+gUnHyf2U+2+fygk6M5rz7sSuegl4
dl5Pxt+QftkgVwDGVXr0R8EPnJkNzCPkG26SjNO5qZHaX7njxOw/z8L1KYjZQzwiF4PZKydg/Cf6
kyKj3602pIk+TS7pXlFU1n27/Ha/PyX238ZIhnyR3GSpqkD0b4vDG8PLxMlwwqjP0eiPCeFaYp7f
MimHNd6GHerI3pd+YD2pzBMPArldSrg64HJk++0UF9dlI9Puvr7aiLgp0AspLKG31BXI2V+N7++h
12Wvi+R2c4BnzlnpE8Y3PgYwBdixH6SQ8CWYOt9CLgcWOGGtkXFuz1Tz/4umWPHKsu3PpxTCmqD9
qyQnWJDadpnZZm7TZGcVB2aHO21scmKYuyrUw4ggGBhxpWTo6TPBCaw518jhUmvUfGPNAuGlxHaP
lvWBd7HtOTLLBtsOsSwUJnYT641fSqrrYVj/gkS1aLIm9R7BIDkxuEEDqKMrZ/1fATfeGoxbbKAf
kxs+hRGP/jfwFK9cggUWgx3aBQU7YdwCeqlBRyf9DVw1W9AVI/muJCGLM9rQt3rKTwkhFuKwqVs9
pXw4jkVq35rlXUHZKBcKSyZpmR1pQlHBPuSPGvDaME6Wzoz6PPmOxhFH2qu/XLoU54MIhp6metUF
6Z/vJUUdsAJ5JLvSBCm4JgW5Q+EGazEn7p2Y03P+/ylmcIzuiNbrqJospo31K1oGxrg3oRSfZkm9
dd1rQ7cxgemqmYmOteDPCizrE3DIfqTHV+XoRkSTMc9bRkruQrWrAtOhVzQuIMh3EBkDwF7Xv/6y
Z9f69PdxKTJnVlxZVHe57DvlTHQHPGRHdDHTa+GGPgtWUVG/8X1cZXken2SlNg2noVreA9QAxPmm
7fOJdsHEDZvnRSLGr9EvzM+gXmYqZ8y1+ut7DeOnL3l9znVl4a33YHGTDKyJE4IpjYBLN2oPBfg0
s61f2rjtZx+xO1xFldg86r2tngobirGnqr3gOM24fOX7oX69TNSe0bO0Rhygv/lpkRM3JUy7F5Ap
Cc8Jb1nFGg8wWD9NrGljcpvdT7r9IaKlyGAqvx6+jmRvA3ZYTPr6CPclwv99bkZ3CwbdMtMNegVp
xLlakSCgRmu2j7kmFR7vsNNtI0PV54IboTAPMwML8jf7yVgY0qtIF7VxMJwJ414g143e0EIG//kB
L8LIOWd96SsTWGEjc4P1KwtSdpBwxfYcRXDyGSQckv+xY1rTP6ydwMmselw4z/64Yz1JLJbcGpKh
axgsz/uneDyBAb7IFD0zuqdorZxBwQT74rGKsGUl+5gjjMxA6cgzGXfS7+B2JBBdLxx/VoD0n1z1
FsXbjPUe9LP/rfHqcet4oPzjxvMhiOI31MMVq6GfJHBeJ7a9Tm1/fnkjN2Y0O/iZwSRObK2FlNxi
dr/jDPBgzOPxwtdeaWP+9QBXVkGNaib5P1rQbuXnVVFM6WGWQupmfxgHYHRbZaeC+AT/SdPdnh7B
pQ++XVaUu+0Gsuz/RXzw9kSabWWIVNqeBsZORM8H3IdDHQPl2AqFtHdMaIp//RG4HFW8AK6iD+5S
1w5RqMa3T+l1nL8QpxHRUpE30ngX8c+8ba7atEmOjUfXhcbYGlYnTpkjrUrS2VUVzSFrwmweQIeB
s7VsbWIoMLAO+rAx/fwmFVnH6MOjPLAqDtLTkN+ppgAmlCqRcG6Hz2Jrh83HbeNZsFGEb15p4Cqu
r3NB7mUwedJKBTjTa9yLfFsbewLyn9ErW/hm/234ec7GalXTQQfINjohfNIU+315SRffJtkjVKll
5hgBKjzjMLLqXYTggB3Q9kmtM1YuxkfVZFl8P7qOkGy1Bm3TOVlkxGWv8JO6TmZCVJNY49EkCT4o
66EjX41cHs/AJ5Nvdfs79pobHqelIvgKlKZ8YP+irhKDyfpBQJ/ZSpRUScWw2vweRCSjKdTNHkSk
/m7wxBqUoVkmuhVCApWRlp4QHm7ktknjyu5Olh5GHuf9tMVtG9EmgXoHmgmOrQXMXofVCx1HextY
pFxH8buuuXP5kXgFJOngqzTVKUQWiAs2VXzy0ljFpO1vra4xrNRSdxNLciKLOeSGXXlikab7IeIV
jTx6G5NZ3RMf7U418B3TLkcftPWJDH8N14ECfmlY/oWHhbF88lDqi3aDMA03PjGhSzUOG61BrrTk
H5oEeCFqtrZxF9/gyr0Z5fqt8fgTcfmlSHqGX9mDaQphvyZV6ERf5ulgc4SB251t7Vq2bMPGs4ZI
rrnppTTVo7VZ67FyFHdinAhgrO/16DB6cHRBD6cnp6eSM0U02ZVUvluMFp0kCWiHFjkEecgbMop5
Zjser4KPajhOgcL0ksD29MQm1AUDcZS8KafWUDSZw5pPXThubUvQxNZskLpd/FSmhSzjGNJ88vxV
qvkxZgVYJ34y4PKtzyn+GBrn4y+mo86bPzPEQr6ldn1Y/N46FEPMileL9hlvdUDEJ0P+dzk2Od4C
GGg/IIMCQx7Gqy0DWVn7axhojFcEYvWGGE95vKF4AYHDS9U5vt6ksV2FgHdRjf9CJKxB2mxfyN7d
/qe2yWivsP7imBa2zi16C9GKxrzD+QEFzKkL52Wto0H67q8HE8DlBTJABPX+7Yi9OZFx8Bg/93kY
ZWv0HumLn33xbPNy6arUARR1/TE5PjPfzH+WYjWbt5g8/h15XbGclT0NuLjuVCz5BO7+YJh/KbhI
y2bIH3RV9zKAKgmqxEK+F5tKv4+bBKtPuoZ85PuqnC+swLUfn44HpeJPo31OxtOIQ6T658zKfUhR
3NQnunq2BqH3RORTrzASH5VRDiMHkZcl0vNdhZGwtOSK5hCbeJQE/0YNfi1NO06X8msZUJLuF5+g
4y67tFEXIjDovGCPBbC0bp2ihxW2Ml5JpPXbtoEu10OM1dIJKT5Fl4DnQTtZ0AqtgnhiNzxs5ER/
J9W6hfqkjllM09EylAT6jg7Vj8s5CkF55RVWa70pjXUINIumP1HFoq2RBu9yAu8s3wRPAU6fRTCm
lh7iVNqBRPm5kY/HVs9oddgeUctzzKqNHSaPIL72lo+rg/uDMTvo/HyNwGWQ5hYZTyZKUiNLvBYc
0pczWLgpCDbnMAQakqLAIYtFI2gDwZo907u/UShmCSdAobPt8V0xPZ7AySvEBIdey879MBl3bs/a
PiM6N+5+s25JmFzIClQ7qrJe45ku/BYTs+FC2yeTbXWZAT6mLuAinb0lS+F2oX9AlZ5LyM/BwZJp
j1ihvClADcjsR0Mk3U6ynXYaCEeWNa/VxK/lxTdhfwIfyzcjoDkoHC9zt4+m9PABjAigV4DasROj
r2MoOduGgyaTUS/rijQYzwuQuLxnF0UmcF8CVpqY07cmKvE29NURsTdHjLjrOD1H8/vCwdzpLtHj
I3AxxR7Qt73z6eXiUM/4ydg+vHArYYW+tckAD0WYOjhyWcSk/fLc752fn6F9fZ0BjuTgIzj4omSu
evrYOVHmJWuEuzEWuQQLakbSaFHqKQgV8cILfAoUYC9tdH2LuzaCK8pWiMfz+EWHYvp+X+DZJgKS
H8WFMyzXNBcIS09FbMTDKBZ5p/4mrmbk+obErs4Td2ljRUAnZ3S+v1spIsKGXJ8PQUZxQWKUrgxW
QuuVdhF7A15HdGNyUJm2k6+xsnYEaLt8IfL/xRhP9uiLMfLSft4uKbhr12GJWFkXL/VWAL7w6Kio
2KRnzODo+OAGt/fZddgmO2I/TRyHuywrdkdQTzM4Xhi9KyKLJK4805KB1oBUUisoe9vhcZXxBXkO
jn5pduqSqH3EhVKX+2NsgvtkIAx53QJNFMGCPKz1Y/wNfl3wBAQtNrfr2uFvs+mJ9WzUkQMEpa9v
/lKMjvCq21S9ukNYhvdh89Xq7tre05z+qquQ3E8fGAKNbN5yi+ZKg4xaJSeYT1WzcZrXp5PmKD5f
YWLrTJZwVm6z/oQZkKUjZkb01ZIYyU3vzX454wtr2LlX3TKkRVcYmyxyVIOunJCZp6N4B1OlW2BK
IF74c6Krz8LjxUtGzGFUIMZ/eLxC1r0RRFHXnlKUeySIBCXCmy+aQREkRR54l9A0n3aGZtyVtSIn
jN+tarRNhHFo7aJTQOjbDuogc8Yvd96y5ATs7PGVuXfirS9Sc/INX5Vm/WgPuDjZU+ea6/2AsmCj
LwF5SFvjG34XDXeouD8ZK5t27pD45qjTE3mNn7A9WFkLnc7P1h05BM3CkbP8Tp4pXNSCQkwFFQmk
Tcv+5gkuiUO4yAU14UidU7805vppLfLyq4+dh8/vDiBkPx3L8Sr80zLmiV7Hnp4yYZ9ArrIlWGr6
n5oz3FmPWVc06dHZmIPdmA1/8vrghX+5iIPTDXijDKuSXkAIB5EfNI9wS5S5ZMKqKApZ81zuwfSp
5NgXr/Ff/UEFg2oKQQJR+zZx19vStZTG6d9GJOzSg+5F/Su3yxDdrslxEGFk1ryYBxfO0ymBQlsD
czci9n6MAeZah3iHc5s6Igs4y37mWSmrc8LhpryI29z1NA2L4Ch14BZ4h1rks3FRfWDEIq7IIZW6
0zjqh9yAAc3qDKFUrW51iVrhm8GM6OqNpc9rBxXvqythpXzLftYSJBOxE546/peoyLvx4DO5nleA
I3iV4Id98uIEt4p/QU26D8a8n63DuxAPgIxhZ4xSyaH0yjqiilWQrHq4NfKSdR2IX5BzbKTk4AcY
ghuZlXxmVlRzxuq+VLOA+31GCBkJ+383XqjAa+6mwdMdPxAQb3QfZ/ywoclSKS3BnYQMB44lG1Q2
4J1TB0owWfV+ABKWVNHiZDKfD2BBJlTjaBClhU8X8Eb5VtkuXnyU9IVkkhHHyu20kHbj/XmSm1rv
9wK5hDWkbXNYqdVBxLaW9YI9unj3Ik9Auv1aOOUOoUM/mB+JsIvXfwwToERPOHVp+SbSBylt9tLX
3If+aZCa+ID8NR/mMaI6MDxargjYZgP6HHQ8vHOZ6sZOXjk12BD18k7ENUpEPc8vCIHXnGOZv6Mo
OkVasl/ig+KuKuePk6dzKYpFl8gz1W2mBlJjyElTEpc6evlMwY40jaBoZYK83m7wcDBP8MdxTnXg
uUM7Cgc4KTafUdzGlF0NngMSC7SE6S6ng9G0KU58OA6YiU9MpJiyipcxR/NVVo64fNmSIlN6USFv
Z/MhSw7+9w7s79MD7wqOsvnffwvZCOtHfO1pAFR+XZVfnTPN1BLNerS2d6KD/K7Z+yd77Dtgos+Y
qjJGVMfmMFCNuTp0rbpVUR9QUwVj6pOLcYtDYbSV4DnNuWiaAfZ49vJ0Z1hztYO1F+f3GZct+0sQ
kVKDGYy2dGnzB4a1gp7MkaU74EpXBzumlM8faD34zx9NyBu3uGu1klpA0UieCqSDScmlfHJLRv4Z
hDdGD4a3OCRNlVHKCfvhjGE7AOFmLXmWqaeE2tA/y6nGBa9IYXsgom4b8chzfwosZlGDVrtk5OfE
Dt7qG0+lWVMjbDVYu8quGWBoboLmQrzN/ZvFxUp5kcehCIeULGBs+uPgGQH5gNdjL2abkqCiyaON
M0UmKo/YqpjZiziOhGC85XdaN0Vrcb+sWfN0oMTCXYXtAmfmDR0u4Vr70OL3W+TK+nBOnlVjFJOv
HtDr/OZIlPtQtVx3cezPiHhvnoG3cBc+KvBKcfVZJ8rCwOD4jIFvsYSKbSoLodfRMijNQjeKZ8hp
0FOw8gl7fQN9eEwOdY3j6vuWRQSSoXeuNXgTiW2j0ZVf1NJWd/JJnbc2AjDadzGDnpNoZY7H6+nb
HjcZ82MDWTKqI/omGsk+/UlwHGqQxFL0E1eaD9V3DURRX5Otq2bQqCCZ9Y7Y0mP89lkl5rxflXv8
K3ZjQJYZSKgQsKt7wUuz3N04dhIbQPka3I+QQOYuY/HbmcGyZxstiEnf7Og096OWxXpSC013sx4N
IdbNje44vG+KOHsBceu2MeVNOxNDQRwsG0+Kt7c1vR3e8hNJaDe2y0zdeMzzTUt5gVpoRSXlaPFa
gHwEQ7yOwcuZu8d+HT5M6P+JgEDCk3ENk9+nktN5zox23OPia84abi9UrJ9nByiMKqC5YOFexO7L
3Zs8q5HtZkZUhRL3WafDpQEzXSx+YS9bqL60ie8xy81W0RszyKRT6ipm2zFbZuh+pBaiuTgJDqSJ
l6vWuciSXsLy9uIjzYI77g5G0sBuvkg9veItZdasOou1Cm8k9vHsN/kKn/S79Ifs3DwQk4GyWsoZ
n/jFGwCrd2+TqwgrCdbePC5lTI/VYkiag/SNN+kKjlgaxdm2k235o0YGraPG46oNLeLnDNdj/1DG
URWrrmBoq4TSjTLteC4UNolSBYmMhIY41M3/nWXc8haV5rz86Pzhsh/HI2tDSRmEDJ4ZwdUjjnBt
Gv3uhb1ixVXOXHivu9Lkpdvh9U8Umw5qgSVc9B7roMF2oJDYU974kTWvB0/sPNvjUG+SolcCRtAz
v3hAbuEXipWSO8kHOlEB7Ax0ZgCl++juYRCg/UiWhAXsT0p3YR7eLDdGdqUeBLlTPr0ar7N/S2j0
5A7TeKTzmZefZ4FoiOnGAEIL0fyk9TU/qLG6GxXLJ1mL6D+h5tHcJ0Pj+r3LXY+PKAHmE7gWFymQ
Fi+eIDm/8trh9ZKX6twEM0codHwnzUYxEsyZiX0HySyhkAn9eG2Fg9AmzeZGMN5Cek96I4J1/YQX
qhZID6j69k2AeJRBfsMY4xaOpk1STfmkmAr1pM6ue+PKn2ykySYcS+Mace9SIdo7s5tizYakkxf2
UH1+avKe6hqHxkDd5Kg04hBitYouXviyKMzOKrvncmJFZ0bw24bewWIFL18nzypZUtES3t5hlq1G
AU4CzTtXwAfvh+M/86qnbINWD9visnKm8gJni8Poj6OcKuQrM6ClO6hbKKPVkHu+lSuHNW+dqvzz
kttLalJt1y23YrPMHARtejI/ZPd5tJhpsQQqIZnJVp402SkOqLl9TwFpg6cI2MLRBwUxvJ0feumZ
mRmGLH8W612JulAPYrhBxLDdrnRpcXNzAe9+1XY3jZCZTs4nfIFH/b5BmiKq2BPxfHOLM+NgHEMm
7sB3yp8x3sOKqsE777T2SuQaBqm0v2mcM6+j2OQm84/cyfxDBT8Xf6/HYa7NyZ+pcGUjXfMjOK7y
Pr7LQzAi1hzSh1O8hn8uHmLKogroZIJioiUOiW6VPVUHm3IXEKgiNWM5u+hYlq7O3ukW8Fy498mX
aFE0C8aDp2WOPyBYiEBaI/xwaQ5/G9oy7h+tf2Cm0n3vW4IWG0vVbMlYszpkYd2geObojYhM8Hrc
3cdJbHfek3mJKc1x7spT2tcc/j27ga/LDwgl/js0AovS7U5tMPESAiLko3EZXNZ0KU6eBYcmHmbs
cBcmSQMRcQFzP/1aUV0YLbw8UzF0wLhhQnwE9qEq2qdWu+IzbDmv4u0um/tPYFRI6VhvTbEf1hUJ
+wHF7UoC0LE9bq8bYjGNBBLzuOZlhLWPhe93/WRrN07yznbc9pWWXqk+8Gc12nxLdGEpQaEyO+PS
dhibxr4K5fyInskLBqnUcRcpYGVuTUfrChWx5YBBJxe5tEgJMCgoJfttGTwVlbrY88l0+8MTJB19
OwDHh6eKtu9ApEou1QN9saMUOtXlvjLihkm7R/mqBWZmUSpIYHU0LdZxbUxC8KqEtE6o2ryRrJED
F/DniB/F699PKJ0dKfakSIxaLIQEPMaNSoJjO2h7B5IcSpSw3lrC+icGI7x0YW4lhoTBZck3TfzJ
1+4IB70jT1S05IUWh1mvbA57ZgndWFsaI5EQiOe0KpMLaAlWNVFFxa3NvyhxnOoL8ycE8j3DE/Iw
AKoTLtmtQ34xCATKJw1zz49aY2ifMptPyN+D1ch8STAnunQ1a76BqQIQeYDtRIElYeLJNtrRNVDI
fls4xx9p6tuk+cxf5BM8cjkFeiz3geERzfx0NXy6lpk4hORkK4Y/ui89mWUGs0IBdHRjWL8ebooN
L5okzWWMG94QinKwzxItZdPoT3V2c7uqWpIBbapLk0LwWYL4PpUjXiSmxtt6670dsdpaOL5AHy6G
9egS1nqizYXfRjefelm+AxBpKK/sU4e7PbVl2IQ3/fUaoJxZhUNYekxOoAnJUvQduegCXyBYsmdk
Bzy/9YzKo8NM+vqUq+8/dM3jRl70UJn4LEzKJy8eU/jo04QbRDqF32VJ0+WNqAcrSsRO/pXtdkMw
52bww04ryZUgxAYLGklX6ZEvZuNFOsrf7S2QI3+BvU+3vRVlWkvkB0tP0le0QDfCh7fciSuoHrIU
dqDUU/RYVWLIKcC9hGLyaBkUBV93p/9oKBQEWsQaad32ExCVY8S0UgLEh4/4zAAJ9IJnJY/PeOJZ
bB3kxcMqSfOcUm5vNSrTU3pfUUfhuCxmIzUHJeb2cpgw7yDi7huhUl8rtaLtGiahpqS6ukmyqe71
3Zu6CR9r8vSZIJNUWMTiV6XZrANDS9mUNbcY2lYYJsEcu+u2k+R+xzBAmIZGRZPzdC0XW7bNiQXN
yHyO5zZClnB3p1zRNFY70ZkV6DM+eRre68vZcglmxtoUM2weuiQQNXFdC0uaYBHaMyc4a+DRV/G5
MhhILsu9HUEP5P0ilBNXSzth/K3j6OtEiq0OKDN2W/gRqY1OyndXH5w/+ebYjyeMtXOc1h9A7HL7
bs859JEKiiKWydiqeQo6tir0AQlvxGoyOvHhSTYXe9ia7Lu9dSj2CoQrG3QsXBOGPXZqKimtL3Le
+xYFevOYmMdsGo3rziF0JOcjioG3j0A59/oEcIKjsbpTUG2692NWNrM7JCxF8eIbaVe8TleD6KXA
FKoVOD/0iDGT/MBwOrWqkixhfFPBbyDqAOj7hwvHhDT6nUDL4SRnenp6cb56a3KVW4+jkhsRnNCo
durCrmID6pVTj8FUaDkqnrJYWAI0ocgQ+bFTC5ctHyON3KWsgCT1FOC6IeD9TfbmWJAquT2RrD44
KOTgrBsb11fRkjevCSLYZSzYN1qTP3ek+6rfxoEyedYrfYu+1xGFqp4NWSs8J0sKS8gTqHv60TPk
nuzikQm+NYZBYykbwuFqSefLZWH/LLDhOL8E5iiDyUDCyAY2rK3/7lNCPfWmhBXH2DEc8o0ei23v
zdLhZhYfX7pZW5t+LdAVSqxlbChRwoKZqT1ltEZmHEFCI4g4Ndw1plmeo20GX83F3+vOCmldrNRo
HIMPff/+yvOwuTcVfDpQh8pqqXUB0dyNoSMuKGxIcsqJaQ9mqMrYjzXc96O2+tUd0J8kEDjZ7bUs
GX0rb9aRfD9UVJ6VFsf/ff2Kyzz5SgD6mQV4xRDOpvqONG+nCSnQuoowMGRdkDFOGvsv3emI1F1k
OIadGL4CfRXYPq6369nxDGqpLZqaVz1sWcw9AHTCD7NqYg+O5f8OJW5aeNPsUj5FNmmOczv3QFZ0
hXRbL6iMAvurymteBf6C/MisEbQEi2GjzNV95H9tboNhEpIuKR46bdd/NrvH8DBzpIIKkqe8PQm6
LckK//biT1deF4a9Cx3A/Is8Im3HIW4zH9kDbAWWPRkhW4Ndy1ZDv/8Eosky6wD8Su7BR52aQnEY
t8r/fPUKl+GJ1fybNUvmzAEKgDEO8PiXaI5CcUqthGzqyoMifwBCRL6/GiPE6XXn5LhZzWzWUsh+
qDQSf1PfH9Abjh1KbtCKaaJefxujx5993CpAavXpkaCuJU2SMly5SKWCiqEPIGsfdVb5axG27w4L
AeEB6Sg6NFFv/W2u+Miqtp5GqNKkbL5ajSUu2MKEGazAHoFpOKdKRrtKPFIQXw1HOQcq4iFfJO7l
2xqHCwtugZpCyT9ntTNqPCtpmGMsBxi0NHiBidk3HaCzL9dVgrd0/Ck2s+QKRuZomOON9N3eLVGt
OtHVC947DjTGkd0KOAZy7E3b11dsImkXDj1TGZXHmQUJHyNsg3L+yuhb08VOTfngjunPMNdmf/QY
LFiBkzgHybKsLLPnoFr5d4/mamqVMuUr6Vs1M8XKXu0LOv9cPawyceU4qR2jezJ/PC1wF2ZlP0Ac
GtCytdDIL2AQ71/ON1FIJDrRqnVd72bNqcqf/LwMkOycvFwweYTalzTO7Nf6trndLOVl5GoxDOE5
PNooCGVSD0qP5Alo9Ru7HWso3B52tcBbhIrxMAkKdKVyUgCPvx7LX5Vhf4/UbRCu/OOWhtTuw9+x
l/8u/BfC9G7tvj5EOKZjh2xr6/sqJ89ul6NjK3hPH5ppv7kqofQjLR18Sw8rfHprPHjuNnmvg5NL
HYvqBe4vf/e39ZErf7P+rdflSwgrGucrK8NN6fa3MWH4/9BNXudQErznmhqvpUod2ZIhlpABREAh
vdpBrddWQj2WneFSA/0yUSPdZ+qUGOP+s4Jqy7xR+uC1r/PaltMjH5qmnjr95dkaDhlFUDcZxX3b
dbGtjc72QWPx2pBGM8zFjs0UJJueBw2hp1B6b5tWxS7okFH4RvkkbRutXzyuCD7g5M2B7z5lKKz3
wQn08QlliP/vW0UW9/39j9mk7tQSF38sO1++C8bOgeKTDbrfD12fv9PUQg73/o0jKCz/YjD56l/g
Eu9kADAiFsUz2JawwcHW3kxCk684e5/1C3/SvjiseTzXGFVl2g4mKfIXTAzxHgVaFTYBNoxmt7Ja
pvLABNkR6O9XE2OqjpeFQ/WbqhbpbrYtDuTqvdE8S0d4RJBCUo3/5o4zAfXddrKOy55VrSpMtH9l
sv5/VAa6edXytxi1QIi/6jJ3dXjXgz+q8JSJCzwJQ6uCFKbNOI4pfbRKY0mH1WtEy5nEho+Dhrp4
O+583ExWtIPKUjSUY+bFbvreHpKH1sQfrtrCxyoHOlNaWWjmoVMfjTsdAg0zY//kmJoO4ZzAGQIQ
TUFBYC3//IJYOHUvfn6/+zeA+KXnfQmfkcfM7bK18OVjnTxlRQbgpwRErf3YyImAcigjwrN2Pf5b
a8glIw3sqmI3NvW/a4RZLXSxks9z78IxWg3E8xkKtpRhtdH/+VuC6zP5akMzFDgEiDz2GRnvgga3
/MUTnUrG2WLRsolryxbpnQpVThxANGsz0ZbwXCqS0kqHXNnYsYR1ghef9vR2HTzYQmo8JZDnEK4O
2voKFUpmb359ZNLZluXaTKlvWJAMW93jenOixs0JIiZDMX0kvXk9W+BVOpLO9V6VEj6uJm4DTl18
24f1XpV9/ZfcB+3BDvjMFPh6ushCEkGbLJVm+15ju1mcvvivZVY3hFPqrUJ2cYgXGbWyhg/7mIiJ
RsCCtBYYMvhFIUkMJH2btpiLx1IWMp3Nun46PiuLzMcCiX7wEz85mB8UejvAsJxwHYEjZaYpaIM2
gKO3PlbmB0oEA7fd3kdDJfUcu7QRX7e25MajLYoyMXoC+PYpwC9hOAfPSsydPlXN7NqlGoL9/ykz
Fba0AsAf3fLi5ylCwL7yM48uJVQUK0W5vOR51pqk1+v54rnFcgSTrUJQpM7DePnt2nHSRXEYr5hO
CimJD/iXldfFXtUyFw4MVrmgOw7AxiMUX5Wx5nC4b+gQGdCjIXLDVFgJWxDRf3zc7sDo9b1SvFsA
M92EpB2MAVZXbNranihi+W77urq0qcCZjFZdgnlwrUopslRZJ1nuvI6GR6cAXwGOKK96PwkRq8tG
IE6W5UG/zBO7K2W1xA77mPT1BFjDUG36aqDpVyZbBAJGKJ6uOqinOR0WSVV6BgGnVNauwzyPBTYF
2Jg06gxCQHPLjGcGPpgJ2ejFJf47pLsax3335aUvPZZiyfiJTsP0KvT3ocCgB3Jn07CqJO611Sbw
XmbJhZiJ+NivkXeKV9gkg3x05fwlaYDW0S1hodjVF9BmpEzQgKy2U4M2KvEZN4zihfo1pbTCyZUI
asjdTLIMHjgbTzzLRIHtjm1TZzVyweJbs/E4UzKjh+tz4MDXlp4I/EbPKEwKlQLUf86MccotGLL0
ELlbXtk+UT10ssxV0dCQKej3iN8RbwvJA6VRiWI4l8GZ9LT7/Wcm0IRk6J/ifcaMO9Is65vHRqE5
xZ0Y4Vd91rHaJJNttS8bUQEULac+g0ZjH4LUYXEONCr3xSQ3GkkEl6HoVG49RyVslMcJjNYcboVe
Iy6qu1BtbcvdwyAj61Z8rf/bz+hNo2p8+iarGmffZwOL/iSL0uo5T6FaeBaMtkyxIpmOxAUkNyis
gjiLKzl/DoMeTmi4AIBbb2TdYeEIDXZSj+fhdoF8aqSWuR7gla0VNcFpMeUr7cxIQnndZqm37bCw
g8j/2uaKK6fDpnwOonXSbFMR6aabQNiMn8BDrYtsWwRHf4x0X+9pPpe1Uul59GQSMO+lX3NPShDE
EoNJao2Z86E6EcvUAcu+/fBNJnqAkK7RisVqNpPQ/oBzd7rANALSmj6moGPVy9GRdzxba/j9zEBW
7rJsTTXwLP4lCCgBR9MPHVIHBYOgMUl4Ivgb4LWepqQON0yxk9MQGyB+jAf+Ayf6206keN8DZyzD
BWmGCoWkFHfsoCU2POnKOXqGPGfC2sWJAuMmsMW3GabI1ATYfMlXAPkykMulKP2fInGlMEGvla4u
EI+IpQjt3X9g1xrVBgo9vG/KepzI66ieQR2UcKxUtWqTOfPfvf9qesWXKqm2dHkCcH9kIr/HYbRk
mIzs7icXHl7AgEC2/nl64f7UewERu3L9yi9icI9d29y2wHxJuiZ/sfmdv1quXaU5+dsSUryRkxVr
ri9pZznyg3mD3ySjtJBiXORvHkphsHLdNfQqykTOFsODBuU/SKP76M54cMmnvizZ+WuD6bNpPPOx
5vwSsrwNMTS9xRvlp/8VUWvi4P6kzU59a1NgY2s9qpnS9J18HZg0hOfDCKgkNjAys3ktR9M342Zb
a4XCz9d1WUG0EhogGRruw09EDVLmZ/yKS5FxLAS2Od/kItfwdxj1siDxFKSSTRD9QScOh2KleC0y
kTo1LckYZTyVFLa36kjRGQ5dmwckgpwmTPNpn02kXnOpapTFM/9BIK6aZ7tkuUuUQQAIJchbP2Mw
Bw75p/r6+RKFMwr3b1fJYjv6ZTRrsbwvwLxZ8cc8KNe/6O+9YDktOOl38TLSLGzHJNASIEv5UPLw
CIRL9W7k6ZcSruAcyG0nFSFUD6Kwvk4SBo0670k7XP+deEHfJCDE/Jr8U92HQyF4H1ourB7aWrSY
3B5utIClPhkolQzgIZtoIhyIXY8lfzmuEqx+mE5m7T/okmanOFIwYgB3EEwqxGLdpcaWsEuTNOl0
8m04G6CaDMhQCpRlG9d7d2+5YoHVsQ7kneiVBVl1ITKBL6fmmFuG4zMDZYATdp9WF1HBbRD5QFCq
CgofBQ5YNrVMC90Vj9LCJQLa+SNOciFY7jbMHbgtIlPilZEb54R7nBeAg9gkBmylrcZM0fD9WLCm
Eoy0QhJdhxs8r/q5J1ZgSu48SkLtb892uHjVLnMgYJkNimEVDwaa5zOvwEmExPF/QKG4+Yokjfk5
BiQeDwNtuSLZRszVB8RiyzuV449rGZR1FGgNXpNerLiRUMnuz/kBqSnamLtkQb0OafK8meBAYXJP
cE0+p7rs5rrhPtvRXkj6ZrItQdxtPt7ZJUO95csXYl5/W3V4tmimlvBFEpmT4NN8Lvca2NLW8Y+n
BIH1Jy6hwFZHT3WaegP1fh/uIubCIa9Me36UClOLJp0EtjvOvCUBJHgyoyWqfPROEXXI/97nqPQF
fjo+HtECE5wPpQn+EQNajHI3URK5gcSBD26+mP6y8Zsh3CY/4UkribmlUzxjnpuOKulnQwdAFZZT
FhomP6UlpbCsystEVg+++wpRMiKOsYKawoxY6EQu/wKb9wyk1BHiCHw9P92IQPl3dao1UpR2rEtz
0WyLymSFOcczC8KHEcslDz3uAU0gZvX56+9SvdPlpdcAjLVRbqz1EX7zylBbenefq+fVqa964kfe
c0a/iL6o372h5SKkbp2KISpwykcKoeYhqcnWHl8qMM1BOG6G6/X7vPahUcVqb+2iyP86iirGdm+t
ZtXtWJLLpUnK2WxIa31tlTLn3zT0raQ9X/shkFzIE9kaB447dH9KqkSPsbTTdvgf+RNK/wZA6fY1
LNRMAx6P+6yiiVthPEtaXKcdRSV926SO0+umT5tTVRLIty67csfDPlA5rYKHWIPFPpVw1mQKIY0M
AXXW1WucgZg7FDKz3zR2LhRiLsvNh/j2OuzC/2ENAk2XeUlYeOPmIBXPN598yz/gAU9bllnUgWtF
dZeAKZ/EJFk/2jkJ8owYhLSEz8LbIl6+nz7IDshV8n+DnLEQECwBYuvKr3+hRnc0+f+GaD0FJmWM
ihAFhOzpE6djjXln8BH5pBfzgJ1DG0FcJWOdxYjD71JxBsjojqcvQVeHc2VYVXKm0pxElMWYr0PR
kQQpkUMa9j7WlXCX4iulVG9KtMtqeqdva4mmwowKStz55yWE/cc4JEBCL7prgiWSYn9IOJZ+lO6S
31g9ZoQpCYml3GLbEpnp6bKjvQp+Lt61DVJ++RXM+Iebm68nLTSAj0sKc7TNPpoJBshtchLBU/Ed
0wpukrRBpoRDJ1J+Va+3XCxNLS+7ff2uoyYTVhFHS37O48v8BbTfSSZVLSUOa4HsOHTq9zPFESmc
gNuhCCORbIouFktYtX8nF7G+PkDXt8Yn3fylp0BekUbjhVXXQYkdLE60xya5mLx3AgNL3AHvKbxW
oSe/hB3hDuSf0Uv8fv5ahcw3I8W86Uh8IYTYgD2t+YY9rx7eM2JPxUWgxyLohowfR0PaugLRsABo
kknttRWXvbbIzIpz2shYFkBJQ17ATiGzKrX25WyB/KsOVprEmCdQWUc/Nl7YnAiu4j378g2p2VOp
mJN6scyKGdQe7cKSqnjnapkW9EOVPiRWafH73W47KDyQzO7Ev4gWayTxxZLW8eYoN7hYdG57B7iu
IIzAyIC6+qomhkyZ9RNlpQM6EOdfueRxEs8ytvJrifFVQOlKSI9h4xM1qMNY0tOCNuNr4dVIKQVb
SEG9uct4pwm643M5cnrF6jnFFKI0Brt/Jbkrp6S3uz5alU3QFdCEQK1Yf0/evCoC4iyhHMzdKLRi
N8HGuLUMsvGyjw0JKB9rWU6dhbk8ZtfcWY+WDtKChXDIp4C5cUgF4ovaB8zfNxJPKuTPs4aqosAD
iTM8RUYJS9rqkpWZpSyq+3JNtQ3NMftCMWPE2K3ZzNdzhDPLW7t2bvstY7J6AxJftMEggY8/hYQf
LODCmtlRs7TpcNW/71Urs7Sqawbt07i6HhlCxzFeCBrxP337trvK/oHmPUrPW5Z4Sj4AM39KJ5eu
4cxJ5FcYHhixmGu/5PCeryOuSpCKzClf6WB8i0pvtslAhyzakr5XQUufAC6nk7CY2rSs7PetapNH
i0/QZO8Z+heN4YA75fRmlfbWeFJGk3HomItRcpXdmW8PqTtgse5tc2yd81GeW1xfrkxOqnqC/SxK
VM1+oeGLKWTYKTqJS8GEiM3J0JumCsNGHQYZISQLEuXJVnUaVYnekAzOw0vwyPQAAm7Yy7H+Orsb
pp/Cab97OG7Inc75BzeK9UjEUuvz+owUQgvE8Vr0aWvFUoquMxhmtFnC7UKNxO7agRxG9ifBp7QJ
Rjgh3CezeLMCxhtixFh/ZJ2me6LfzAA1+6kmZuexcf5oLKBdbRy+uKnmV47nRxUoU6AMPYi1hHRL
6RUWVH9FVUdlM65Ah/vaE6kqTkt6ik25rW3CVcMY51u7qmgR600gykGLnYH6g4aa+RxBqlswVewz
Z1cAgdJ5EYQXjq9G9aQDSX9EB65P5q4jTj1Y1J5EfSJWtJ4M79fo3yZAGOFe/vMJwyfx78dETJkM
BxGNaxJeldrY7AcE6TEMAtqYKa0ccpJ46GGGjNhqF7NaEgxGNL/S883FDVVJFO5YYQ8TcOPO7h1o
SlV45NO/znra0XaN1OvE/+vgmkXAx0up0p/jkUxL4Pa24pCkiI2iHvLLLvu6ukw1h8XAnZTCD07R
aqn0WUmU05H/gfBfVkvQSh8vNvhc2nkFzjgMl1ph8ObLEdeOyG96+ZiB+okuX5k6BZC0EYpYIO4J
GjzP6G8fEKca97UfF+SrZOAJRumbzLSSfApx4llJhGfPeqZ8leRnAYULNwJJx37CeFt2brEhXqt6
odt3/VGKd2QJgYbVaHaqMT2n9d1u9IkUZjGLUA7nlaxB62+W/YYAmJ7F352dRe2L7KrBayqIrps1
HErybT1QyQY52JCHKnpr4u8xBfEmdMoHjsHwaYmanFgnskIYgC5NVgxmXGzfHkIxUnBCF3zKdgkt
pIQc4UyJd5tK1X0XBzqcc9zNWWL1bvncA3uZoOR1HLRa2apFob8KqufzWZZvoULoXdIiGI0KkdzL
B/6EVbVL2J83pu5OqrujGGfq+V/Qw/rn/SSuk+0KQtIdHWfY/ShAnGn1PGnk10yMyZ6CgRC4IsMD
5dgljT6+/dl1zqPVaeqVpCIdOudut6ZCkbHx1wSGal5t7P2Ee9rc9R1sNt2ypL/+/0Ho94ctV15X
HgnozjFPdcU0msdgjaTOtzOFPLPKudso/K06m0niZrTK56bRmPxXLJlmj/pwNmJdkR5fJSD6pFfE
soqXCTXuGRVxuYlGzyC+A3tKZOZUT3/httca2pd4Sp4wdAwGES0XY1DDxBUL727jBFot5j8zZ9XF
w6GDHiFhQ9JBelmdcNMU8hBcPROLZfgoxi2zh90wGsYJjGw1tcUS8W7s91B4CMN+Hmsg6Pe5mlSi
4nuzbeiUs+7JlQMKJ4kjcX07UnrcNmkPI46DJdyCG6+CtI/mUpL8wAPkg3KWxftLq3crJXZ6Cqud
gPmQIF55zTyzaqnLsWoxy4Dflgxf0c/I1w6Sd0Y3/58qMB6H3O7E+j01cCjhDi4PMoKIsA0706y1
8b8olqTeQ81jO3iZznV5nTPzbiKt5LwdJ8PO7ZB1DyqoVqLP+v2aZHKe7m4816NmXTzycl+JsQio
vqDpsgZSvW97264VHdjUSIi5EzNJQvWvXusNJemfnFXX6jnP/KwU9HRbIw5d+2WFcJBUtsL1M1ro
la77G4JkaEty1CJAsJowDctCPnjceH/SIwdFDBBlcMhqZ8LFMzNOYW0eU4O9Ee5bLEShzIt4MTCA
2RwuRbWUORpE729/CGd+84cakY4coLrDxKKzgm5qXmbTwQ/qqhQTq1UMMNpxd8NEyBwksvGHGgIT
ztSXJCjZSHG9XPeMvdvA4r3+tWwa7klVY8E5SHNzccgWdYMGmOAZQ0mWAnFoca2qhXBESchNWRmC
2cZ8DPEhRSsSDFwnO/O0C5O6ccIg9yd7wQ9lJZKfZHR7eU74kdFlfKhLY6jqz0L/cHW7eh7/ebEe
IVNnH0ATJCUJUVqZJjBlev6X2g/MuQl/uk8ZezyVEI28g8ZGgHo25Xa/zh3A6vzaR/KEHbXLRmQq
Q6zxrORdvbf0AuEiqXHBCIGgxQT0x/yDNJs8IiHw/ZJUwiZG8MVXBIOif9EeOahZdD4TRGNNs/c1
xK+PLDakq3kFSru1SR90WQ4Hjm/MBc63YwE7Nst0CQytXRRKqaYpJkoMTlJO0CH+rYfw1esSndcp
tNULquM4j03H21sgQgf6PNUj1/eM3EQiFIcM5rAPefuUeMp8z1EUU++sZwI6gI+wCJwvwW73fcXH
eHp5ehkZ3dqKoAepOGRwkHdSPBT7FMAHejahvj/kVg9szJ1I3IGkKEFDqUR6bL8a+63IYuCsxe+9
GF1XIR67+fLZrFRdqe3md0cIP9WjZLTHMrD52/luWBu1H27wnikqwytVfv3HgFZn3zB7wfFaJhMA
zvshPyZVPbkdkHqT8R5JOiAbv2i+SCZOBJZ8QdwQAkUaF/JKcGUVhNs/AQd7yEIGJnRyAixcLPAV
De25NxUpAFKtTRqhAUOOb6upWoVTFywuXEupMLEVgAa16TIq/AzOaWAo3Djy+LfG36hj4tg1gTKl
pujQodpE5u1878j57daPLAGwN7eh1yKCkrqxVYDUj6SQK8Ugv+TjrYE9OhSoWs1J5D0lSVEwV6df
sajVT/0goSU1ydInH+vX4fZ5nrXa32Jc0C1KthEWttAy6KRNkhJjfyNoV+8AZHOyyD8fthGwJJiv
hnsMdBoyyUNmlPhg6ZpfvUtHLF9g+6qG+TUgfKiSJdpoue7C2KU03DayDX2DOH1Rr4OQwVy00qCH
NvmRRXo/+xdImpaW5i9Bdc9QBoSb9ppKomDHtcpo0+rs2hsVSEPYrMb+4+z7YwZCnoA5NtQC2dCv
q3QXsFyhkO73wag09OfhoiuI2VXO5n2L/MEBcfGmKX+0mFfwNUv18pCYqshiEPhYJCdkVCR0dZyY
70/x+4kFYafoo37Np7YClt6WNRMBtpD6eROiCtlqMnCWCDeU388YlO3Wez2L0L84FMh7EduKRWDw
d5vT4HLA31RULF3A9C/kwR1AQcWMH4CDXohNu8I+MCVEM4JcsJNW2H8tL4capg9tJTn6ZsX1qjxQ
3RKZ8twJB1pSbZ1ZEOG4vmr+o6bCG7KSBUHcAZkfsJ1p+eILVdO2KwHHK8EMgMFwY7GR8s1zVcF5
nXlkVa9VKFmm7wmspiKyZSRE7iaFB+AIvVhhcDPq3cey380qUAd6DISDFelIZBJV9aeY+cv7x8nb
xJ9whlFdJ5r8usznVU+fWi+rHocScGPHEHOWcGKjOF86ty2o6FeF7NmSQMoBOIrSHRx7FaNLNu9o
NA9ZPkkJ6RUlR0dTRB5SEIBznyRuBisyr8DCT7vRusqFP3pjdT6DqZjoxCZrWJ4rx9OznXZenIZ3
5OJjk0dAD6Hotyx831DrEjnJHA4N8y0oMliwE7TrfuajwxLG3u7D/z9oszb06E8w9A43uVbtDK99
FI2DqI8HXBcvHQzo6sfvaxeqhaIYJ6SgDe39FDh/I42KNAfUmfZSGd8oqVFPP//dOyp1qVxL0lvf
+aOZfNZNdbi2slv7aKhlpr2EzlPf4icruT4AqXL+cKnmCIKLY3hcsqXrp3s0nwsCU7Q3a5BBGe5j
CwKY9jE9fpJszvv7VV2f82epysanmA7f/iAPkKSPd/K5F64sQhxXoKocBbAA+Rhx0/xAydIhW0uy
8019Vy2jEPPcNYUY9skt7jK1MtWB9AcEaRBvWLRB0OvOdaZp7mBY+lhwJf/M32pKLlE2KsaSLBlH
7S3ca+owlgnEtLLGelTGxCzpbgMtZvV9yLbxZGHurreEtu72RLVzMtytzgnFib1eJw/s/umHtzz0
rEMmUa1MY8zADXmTIMj9TTYqUDbdcLg/QRHWaz8ry7Gm4vfMJPvo+flJ/rLcREAcFYBbkWj9nGr2
a7teU9Vxh/CK/4LLOQ8X27w2qT+91zDhyzcxJZk/eLuZZaoKpuSDgQR284DV4wAXN0LKZIzCwLcm
rnLEV9e3Egpyp3u4nxCnC8miUaAligtfYJzdoB3GrM+76BsWfI45/NBfhlY0oyxVL7Nfy51GVyvn
uyX/gLr7gFObTJKD0fo11rx2c3Bri/aG5Pi4jS9HTI8FWSewkdSPvVtP46n+sYXMo3kJ4/Tk30YB
pNX7bb5cFQjSToYYSlMxrU02sl8Ck9XAUiAOJ7HxyuC8k7yBURcYuVH0BoPoFbL6324mlzT2vS71
049xVJWXZM/Oi9hmi+6NZFHgMQFcJ8XRMAchj95hYNg6M9/QfvirqvnPpF2+ynE37wYHfwjcWXlR
2aMKh133PIofx5JtJoIzkFfTXMpzI3Jfal98KQEZh7k3FumvKHnYLpezSI51xTigPVWlAPu0fjcJ
BAQ5ziHLc4gwBppzOkoIR+MLORVDErvjOPTL53l6noQlLhJBqoHwz00MlLsQF6Tc/5YK9+OK25TF
u7oeUCw2AuiE0DgrC9h1KczlCrwXvDyblThvo6wwv9hMQrGJSJ8z0xQYHFuPQkDWt5r/OQsxiUk1
UggsSzX7l8QSPkJMYo3+6+Up9lV7FW4vF28ZwzgP2htIJymzjPxaATsJddoc4lsCaxghMZCrsEig
nSXDMj0ky7d39L0JxdjKeC6n1ecZ9TyGaJ07p8isGg01PEi8+jrVUSND7p9sxo9VbG+MW68gdjnh
wwQUcyxsaI/PQMu4L19LckFYgHQD0juT5dgwXvMR2aZ9Q8E7POrrCIodYlf1LdPtIbI7VURLoXwZ
e/xUTwWaiCx5OmuDyzIyeNPaT+eGzETmj9fMmqfpR/PqXo21/eq96GDQf5uh+Kh//1hkdv7lpCzb
AVWAA/VPHc9RWd+jR3d+H0iEZQ6T3dN+x0a+fnDdRly9YQzKeMnGqsTd1JTMXYBO2orEg4n+cFNy
rLPcNP8v46vk3lkeR9kTTjl0Q4kEvbbcCPeGU+SBbvsT2PJ8lNSUWOBPbMyr5iMq4eilx5HA7uQ7
23k9t/qj1SjcXCCd6E92wGWgUeNXwr4ScTvZDoSLDpaLGp/WsGDTM52sJ/+fpzcdffOKhfZB3xc8
6u7UkOwEVgLwKEMy8zhrYAj/JIaeyM+HaL9mxaewez71BfYnYfpCLor0KquM0jpskBdTiGXKNRgU
83eXHo22ZjbPXqS9HlNLNxvSOK8RvAQKOXbMY+Iisnu9lJA4Bn6/vZUbdNRWAZOjv8zy9jCBcLmE
m9RJCgPppJOD5GnOlJHpa8muFAUQER0I7JTdGKiE6nzZtCqsMRlaB1AHh1kTfNEr+6G5db1OoYsw
8XP4uSYJtX3vnrtrHynUF4AHDbkk9cmAuuse4DmbG81vGmXzFcYLcV5GAYCvvEC1dAzqntrBcjWW
qzSAkV0QXbtcDlgphqU831+oL+GrclOj7BCtmA/v+QCNQWt85m9JwKzNqZkxIe8GElV0Nb3yGIAZ
r5+B45pI2pudPHtWGtPn4fzw8oc6OH9UwotMHcdl/T2P0yTBl9DYFCkTKjJH5U4wMUNQ2zuLLTKN
hskr4fp87f+iaTOBOABppH/PFETXs7hL4REDSiy8M/zwavGQmgjZPY7GjFyUq5IzZ1NjEohiDd0a
YvupB5gnOJi2yLIqHOvSIthfz2A1kGraw/gbZH3ZC7sy11j5h0p7GjGvkgXEYD9IvnFzAYi++rTA
CGwylrhdllVVV/p2/pxY3wkHneCxyWx87Yw23jB0xqJ66IULkuHdC7kZgs3zuO441A+PtY/pCejq
DymoMWjy4L2RBehwPEk7GY7s4oJvDCYxqVMoWXKQOhUOq+gFZGsHEp/XpOydasOKT5uKC24z/LAM
fo25Fgo+nFQ5pz/NiIcAqpHNQZWgHgnMem19+x7X8LdUB6w0cyBVifgvUkzcuBRV8laKXuMQOYtm
1uEJRTusQwANJYR5iUFVP4/TzfhEkjw1OxAdii+TuFLYnUuHUWqGn+vEv6MOoglZpngbHnyYTuZR
Tgk5C4YnNe2AJBmRn+tuJJSnO88X2EKT05lzhKDNCyjGxLuf+2s6bd4WGa8J0m2pMJojkjgTYIs2
iA1fzM4GURLAWNUl71skQO3eX96gadyLlfhoY0eNXLJCeNiZqY4otb+Ht98S5+JojYCgCPV6F7Qx
b4sSODUiMdD8OML0QFUI+DGNqUPpgI7lRqObrlNUAiEzlCRsQ0Q2XAkPed0n5UHcywehgXrI5QBL
2KsdbgFXbRcd4il9rzNJikDCPqBnzyUsi2lU2m7BtsB4zzSkY938uK8Q0F8QPfob+OukZTLPvMzA
GXPi+ZSpXcsiYm1uJuIeTpPvCmKqdtLfcc6MQ1wc3f19iAYiJdvsGm43JIyq6wZEhi/vA+/JhT1M
M/cs4fwu3KM5s0mtgZ+zQjTHm8q0I8VwP5wtYfPWe0ESYUZSbMZK3kDuVDqh5XMQJq1uK1paP+Ye
ABIIlzrgmGl/FQNbRpp3e1wJDGD9pxnQLCsymPnEabXF5s13zUspk2q/1wNCKOlO+5Ovi3HeRUSa
15UNeW4p1gcn8cYG8K/wf+E9VgVpC44On3V0ux3SrtiSU1frAuV/Zb99Jb7FsY2cAEbTKnp5QUN2
Jl6v4tqvs9PjnIU+kQ/Cio16BdnZqwUzpx4knw3GiRIf9e/4PB5w5K2uK0m1C6AVShlViw2epwoB
KuT+qUhjsMhsqgUrn5LhspEBgKYnET9uF607eUG6USeHy55OVz+IroEJcJgcyCUc/EDsLzgBcZ3p
XIZws+jfFcxzCpURKv8/GyeEk7rLjcYddPHy+QauntlAm417G49sV2s0tSdkXkrIpUtgmJdjMTng
O6XrLuXSdesZ/qmHrIwDtHCWP9ELABSZvSh+Me4OYpQBucUBLhxB6FAO8ZYGu50hwXIubyttsoDf
yHAEuHpQnRi9a+vxzebcFvav2MkrfmtGBGUR1U/grwrd2UBnivHoa/EsdNsbDGcctESl7TcKzrAr
loNGR59mz8IggiCYRD04JD8QdSQKrWt1KGFRsxrNnEVfw1TDWlgtYuyjwQUvsKqzWn717XkR99C4
EKtGD2U7D8HD9t06RfeOvMU0q47DM2QPk5FICaralYMVGFIzmC3ZvC8eTNap/XeoyyAUM/+WH/7/
DdhGkHExgniGfiKZyp5WaAcC89zksQwFOU5v4ImHOR+DvrtHsD/ZgaHb2BZlBeqFgNhHJRjk0NTR
nmxMgnaIRqHgglOZUBLk2k4mjQQF03cl53w+cN9vVQPsUd7LTSn/ZaF34pz3uF5imK/b1FbJEM65
cYiDBmbJ8z12NErSvFNJ3I8kFbx6w1bo6eG4GbfkhaE4GLYt2wdk1VVRXKmD97KAWuF/tcUMS1Po
GuIIyoiZ2Ca/X0yPj1+U9acR/SGGbquTtmq9+RwjEpTuv/FuOPopC+eCJabCSwq3z2W1DLrcN0rJ
2ms8WvAmaloZgDx4mPdfeeNSepMFs3kPDfy3V+3NnGF5ri7Q4nj1HLlekjeUxD27hpJpvL2t4AhN
VmRhMC9FSeCTmwMLpyWdBh9cuF7HytU4j0sXn70lSfr6JX3OC6RR4DD0Uz068DxzU/rZLzCS8zFu
b7ZSfwEkIHcwDdRt5vFZkFDCTxHIFJQlBzsEBVcZ2keSpn7c/YY6keW9h15op53i83sDqhvl665w
TPgMJLeF527lYJc9hRnS6B7Wp9u+NZ8eXUeTzmc/Z8+Ewk8+bEHC5dSQoOVRIt6YhtpJzpyuNCIk
X3nZWhALtDkWNDjQKviSVGJItRDKDGUP7X6NVWQLbcxWlNPHmIM0L5c/YCkM5UH5B48xvyJOuM9z
I8bdYGWFr9W6C6z7HkemEGKV/eqc03qLHp1KpT7LP51mF48/1XPtA3baHa1q2sXqSRcG+z8Rcdce
1+9MrF2KbeDlKsxWgklILYluvl2HAPXuHfxnsBJDBjoaDXbtF66IVgVUjmmm+ZKrK3OC0J64ZWCo
sA7JlsGXwPowDsLXt+zFH40j6IAC4WYVqmxwP1n7cMkIAGCDqnarJ8bZe8Ilo6Hgv/jAsSkQOqZH
o0wtfz0qa9QqxQBs2OtmVBj9sbXBRmZoYlTde+B9xftnyScLWQ+VDKwjMq4HY8eachiURvYl99lT
sY2QmhLFkXOTiyeq/N/NwRtbpGhKh0idunBF3CjGPKpCPyHsYAO6lSh6G5bPDMgq7DuLYflS0q+L
iKuwNX7t6XymwJvAOZDaxcDy1V/RgUZCXo0aeBpP7DG5k0XD/eKLVs/YVLr9briIWR0iJC5i6kqe
9C4a7ALB91BtRfy+p/ZkWb074RQfUe/Pk7lshV5rAzTlwajMHSJ8o5+F5IxsdICZ8cHGbqlZNtOB
oKpHKHxBjOCR2ZZspWwphMB7iks8p4SKrgTuKwqnz9v/WQDf7s50D34Ty2dQgTFwl6ArUQ3IiRAd
iIjlqwCCEzP70myjR5T+JdVhI4Y7deKhenwxEfDk9ifoknK8+armCAGiPqJayvCaJmMGZsqV8bYz
2kYn+F699B/QwQOrlXhV2e3wClceOiKl7lKt9DfpMgUxec7pfc9r6s7s2HmFdKDSTe9WeeNHEdjk
u+2Fz0k3KrqmYrB2wcY2DiDlMe4WusT2p1Sgeb920bFAHlEYFGXD2IDZgMyKrOubUh0U2nmEMFlq
a6BV66xjx/dCeW8oajWCqB/h1uTCuGnx7NF+rqCR9SJJmbUxCypnQCx9AM5Gnl7LLQzJjU0NaXSm
l8H0R/roG5lS8PJN6UPwadbzv8+VSTbUmQIu42yQTmBEC/NOQxGqNouj9OC76/jvaEs39IeegXko
IOrdLfuI7Oi9HGTynpOiMy3fO/LIQNQWpphzbvCFqf3h5befvIHMuRJVVWvW1DxikikT9LaMVG4G
gSowqPoNclVcOFGD5GGFyBiSG8gS7tzg7dAnCulExURwzLACV+umu4ARURrtcW65vN7u9hG8G3EY
Zps85M8bLiZYcEox19G9uH9P6kvMYH0Sng2rZSHW6M231pDGZts8Uoe91ryzBjjO8IiEn3T4Mr1O
enJc3mAcWG++JhrzhIq4qeMHNH0SDh2tn9kVSwLAU1tGKUK7CP2kvHxKdtWJppAlCK39QHEAky6b
3vywuQ+2ifzA5zRcd0szS2eu3pAy0LFXyRozGjRQjy1cXoPuNbfMr8GBuGRH0bUp9C1Bem9T8RE3
EZVE+3QbsIBXCcxNeBd7Dt3QdCk2XlrMzKlIBSVmZfkZzZEJbcrmidbp6RNQoc++KOjQ4bR5hCLH
JEBqTFFzxLtwTiPqNs4snkhgKI2AsvF0HrwPXJbp84JOg9Qh3ZXE7XlgXdGVCs2SjP8dBWnp2oD2
eXwakop7KHlbkv8vnNYPgjmq1pja77WYtzLeowhc2unZ90wawWCjfHFIHmGWz6MxX0NtSqh/Kqd6
bB1AoDGm4nQWe7ndkdaq8VscfYZgyXbrs8BQSAGsNRMxgybkhrjyYXb00So6mC4MAh9jubpDWvG6
0pZ2SRJ3TvwLGn0JXrhY9FZ9mlp+3cLRBJYkvlpvEtym3pqLIXp7P2pv5iI3VqgQ0qPj2Jegr4up
aXkcIM6UaOt5F0meOAfCTg2gvBHU1MbhXiTPzNxq9TSYY+Fao1pYqeSyaV2IygLEp7LBLK1hOt/A
qwoyMuF+QkyaHVp8JGgOA4b0/SfNWOZ0j9yi/HWM0RxO+xiDEj8IW4+v3J8lAQkwQlB28Z/ux75n
3x6w/Gmg0OibwhxiQ0OMYfihwu86PTmsoiAHfLyrr+oBWlcSgWwzQL+5gEWjy7sRnEV/5lI2NfLC
rCcFHo3e8WZg5UvRo6OPDBxncdhGI3bt8lewhNQtIovrhsqsse3ScKIjNj3rTqJfjm03SN15S1W6
v0bpMCNlBIRu8fEWbK0yhF6qzZTFclUCrLor5EB6vNwX8Pu2TLjEoxtd96EjVkT/gS97tEnuZOrQ
v5GLUhFclWIoPUpI30ocwfkNx9DSoihTRat+FFtymrxBYCnlxsuiqaY81rjPDvnnfXNg0ygWHJO8
VGVtNkP+GCqjDx0f5INtouyjHmcdB0EJ8mGRerDj7kcsgnrNBVQRRIh69et5x3mE3IJMJ5EZaaOJ
HWS1MhKJaQdECP2qiTVuYStghzwc+iz0zEVjwQUml1X06hFCdaNHOOgSzXtjXFKadw1iCCUixtB9
+PeGQoB1Fhsnk2mIhSYYxTyQDPomvD73o0XJISToV1L1B1l3HKIgLDmK9er3r8op5a2/09pxXD6y
PZjshuUiAStEatKmRC6BbPYDvpyNQYoF3PeY+eZq4WqfkTrPX0INmyIYOo+4ZuziFXN2zX43ahph
ZT1rqbQROiejcLJhNDuE/loYKOCrZ5HGKVoHF7wiN0Bmge0xmQXGs+aljLkmpf0hmvsL9OT9maLX
bqKyfOcs8BY0lub3CfEfCDQ7Ny5S8xi9QF7tIre3xAj/uJor9pkBRDNkgK+uLbzuvKoYLx/xCU2d
14i2xKrBOomfjOarUndFrZSwLR0NyaNsJxcsKpjDPRVnd0wUjCSgdfatw+6+VRx+nEpTCcyxHQ1j
lKql66to1eQjXNDn3izRTge7ehZwYymEWypqSBsO5+oJdoyZDl9MN0roMDy8iM2K4GgdYzbqQf7J
KvTkb6FHLk51qHHJcL+8OQTg9GffqYP3EMrxT5UKzgo26/J6URX24q9qeTB15B069PF41POU0240
ucgN2YhA5IKdxpFmNnV8Hgrq3J/RpFCfE6VumraE6FIW6METGBBKioUPgSvXEzWG7XFHSGW0Izcq
3KXSgASE6ZHpfqA4Zq33dj8cX7U4Xp6ZLN3aGyI8aRfGvy0kLeLpzXLwY5iyTsYAkFXUgYKc5x7J
m8+Rcw3VYLxHaUA3BfQp8ZF0EnAXQ+Ocirkac1PAZ8JmgpgLOhh5eKwLlch0h/lgJpNImooZRAZX
XkaXqKHWiG5kIknlc1l9bqN/ESY8vh6cNnUrb4SLrS40wbhcJJTVcqyCVfMkPlwh0nB1KnnL386r
op+fM1aumaOMhkvqsFogagSFOOAYDENiAxX1BHalJ5FI+MXZXBD3pUNph1WV1kBcNCH77++AV1mv
WJoVQOFLzZ0ps/7WOfBF/AAM2z63ExNL6/tw08FTrqV05t2QxDJ6JIKtHn3Ll0UpKrERh1/vPwyY
JkZV+EZPTZCAZrQii6ZLMtqaNysdzpIw+sAQTanimblu9YwoB9/GXcn1xJKyCv9dIchPxTfn32CU
0cFmDBskztwpvBsihs1khZrE6RL9TBNEvyo/xOtMs5V/MokSgL5K7ZRA9c6XGYzj/nWux8mUN1v+
4yeaIBF+ySPMtQuk/Y3dYbBDVBQAn5IYjTjRtlk3bqH7DiHtnw0Zl32BBjBvK3rgNx01c+8MRdA6
hnVJM1SKhSkX+HBe7fsUD/t7dR8kpObTMYIEDHCpbXhfTVEAZPRLu72IwjZon5evaqQk6Bwtq050
j1tlw8pQ8i6W6gfRPbWEyP1zmrBWPpLthRa4qnXO3Eka8Sd34EkBuWJR1uSJ1C/Fwwerj15oaEoz
58Kovlh+MqywdKnzlDnRMQqdPphw0oZqSrFtM7dboDHyTsymOXAGcvEQOL6YIKyyQHHLMfJO5C19
C3FFhI/NUnJi8ZOdHVhmiLTRK2zSHVq8vRM/ApbBzKqkjw+UEzgXC0sOiyi2fPvWMeh7rwcRzs90
5H4kXFJM+EmYjfp1mA9DhTF9iu+MJFncLzhYtt9RnjyabfbLCJZIqmJGa/hWvMTqU3U39OhY1UN+
TsvwQep/3KHMCNsixGr/kb4C7OTRiNzNSp8J20OuMh8mTaYRdOCcUNO6c3hqBT5qTlS6KUgi83eu
5U7aDz5GiZVwFK5mSFVRNK2DkRstxABv8F4oWRNldq9T0unJ8aWFM5JioWM8qxTd4hL0MIhfUbxn
kux/Txjd+CGv1JZcjwtWiqnHa7XIfAIzQMEWGabj3cQ6E3EXh5jUtYanPtxe+sAdTpd2+hiscqZV
njqK2S2gpPEzYxinA8QZMJcRC5tnwUbNSJYzzORBWXoAj336HIeofgqjdSq6EF7HmxPyaUF5V7tj
7uogLlJ5jUIRbOa4X1wshjsFXPBJN7NMs8+ZBTPy/L/T5CDQZgbY+wsW3hUKVi94Y2jsAobrwJaS
v5cts0DjxGJxkJROz1qE28gL4OJN+sZvvHYifXBlCrBrOt9aScXETVmCr8aBuUowTuDzbfdky86K
uKz33ZDWLMYq/rxfEyWXwgmhRU7egFXAe1BAfOZFiXTI/0yU2vvtZ4C52yJnxnR2KoM9qc1/6s9k
dAGB9ir5Sok+JK8vFJkJlg3kf4HUJGGEH1gY8RMtTMlqK5tqCEaevmQC5Q76qJM0vRO2Ez6zYqBI
jOFClw2tqTouz5r/pHwyo1bsIHXexmN0/CiwF0XcK156jtfh5TUeneO7m8Y2YIfP7xvTO/QPGNpf
g8Fs2tGlLIdwVflk8laoLP2ftai3FcKhjMs4zCptURgJ4cKhltBjRgKHmrms6AmIfwEcZiyCxYLh
IZR6Kmucqbh42yIxObMCtpTlfA+VMiyY42pjcMSuBpBe3L772Ol10UW4P4NxyJSvpVLltvo4wPwN
r5fcswn6aGh10QoIixZWMA5/2kv54f10uvzCdtBXUcdEgYJRz+CRWj6ce4QgUhZlzZtGCaptTUaD
6AMEpYgoQzIPneE1zbvnGXfPNxcjP6p8LBG1tqvN5rxS1dRz3nYg2ozErtXwByXfwc3aTxc3EKN3
7yw8HeFG1YfM1igvwphn9J8n2vqEYutVOO6FObUZJ5gAH+AKLUN1v9QA78v1CYhX+JMQVVI+PTrQ
3fOpHvnSAoIHKeYFnglrYt+XSyXzcOtMVDU7Md0+C7gsCQoN1XEAcDxvxG3DSLRm5rBYkE7Ec0s7
8q+ENx8531AFyzlKa1cx8zFCyJMRvSkYlkjOSPdlncBhsBi5bPY4ezZgn0osPybp4mV+OEWhXZLJ
TCCO161B1JkPx0sjJckFMRR2dpqMM/bRY8sNVZg7GIGRea4DaBYvJwstR2kO+taTqw/qRPFwJzWN
uEPaUZ3rAt6OF3kHTpEaS9QAF5ilN468onR5BG5tKBGVTrY1iFWt55Jtj/SOJm2JriUfkTGZM8uH
sPHJpsHI04lwHkZQsZmnIzydRPM8m2Qk6FjFqRC7ajNK3+Mu0mN+1C6PIzvwPARPHH8vANFbgYK8
es1Z8w5WyC1fxKTmlfOT2Eo6VKB6qH/dT6ytKXH0wBE3E+LI6qRbj3SA6gYQQ6SzNUBnxb3rivzs
8GOgeL0JgHqCLe4q7wtP0FBtPr07uzaAqQ370Bo2saZfsFgJB1LsBPt1bvEd2tmWSoNvBwpR5Hv2
AuNJlYxXmnLHPVr+qSg4ayOWqdbuFy93zyrKK1XHchTn5oS8VAN3Em37zI14kE36bCX+ERjLmmcb
d7W9hHgFHEh4FbZ9TyqDEytCxHVvQj/HtALVCcTQ+z95BgmoB18NFazmIthJasaG4bWcMqqkBfNZ
SA06qz0mBQy0fuukZYkh2ZfOusk9khZG9d8Om8IT5uEb3UXdpG8NBY/aT22qFzJFpOxklHqmtYdT
kQvTyaxG6pMDKcx3b4Y77VhZgXdyKNYeLfQuUo/G5GydTdOZu2KJGeFm7waULQXhTNkHMDt+vp2v
Ovv1tQY2ccZD3k7/LY+HYUX6kEe/QNzdjtwsfLC4FzW8dny8yMJn1A3E4xJi5N9EMhdZmG/aMRV7
Vt8NII6gPoPd9uebaJKgLASm3K+2q4INoRrEHiwgZP5U77pXxVLwI+PyMFI6YUoaJqF36JLVtNm9
lKbfF8VSiFiwwy5BPS/x8yxgFlFxAWN1PypYM6x7IXwt4e2/s4q+iVhbsMZl1afgNgbe8KUC9Ce3
e+rpeiyBpQd7QEoPbn+ZBGsDNeCcytNAGd5Z7XdPPxwpncvuLGBaqPTeFgk3atoQ9mDDY8BH7c8u
d6DrKT/WTxlTYfY+LSXrB3VJaHFn38kAg8KT4iUG7d13IOmZdYRnvNusJVVasbj5DUEZiFWYiw+i
ob9s6PlIGS1FGSpXDbyMW02W+7ek9YfB/kpvle9VOGvy/nov1rUrxzm0XgTjJaqv+6tbnuO7NQuD
SqlLwu0W7hlTIrI96eP+c78j/DAt35cuVJe2CYDbvL4fgSIdgWT2ljX6Pch0A96gaYYUqITwt4Qj
04AxfwTXZgN1I8/CQtCP26HJ4beiB/rQU+DaAPl9v77xgCgSudGzndoLCsHbfh3N2drbuZOQ7vZH
Gz4Qi4IFVw1ixS/BpZqI5jip09a+yftdLwuyROHMiW3IHHBUuh3e9hz5O03MtoLFx1NXB4rncv4k
PT5S7Jt2J87OMigrNahiV46SsJja/8yiTnsZdIPsggaRPe2+zxXdFNl9vsoXPWKEk9rqDlt41gPF
j926ljdg5kc+HxQBTJn5ICGKQIMtdrxcK9FglFMt/FifdvjLrnWcZznGJiEXOSIYUjDuepSIT9qO
UbTRwmU/qktwWmEyLLHwSERzL6YCbXQMCfhWsVsuOPAJlOr6VrsJ0Q7FR5hakMK/BSwaEPb029r4
AsWfGmJioaDxIx7hlWVMCxG/AMihKmd+eSDA9uBkyKG5kFfozW/qtHt3Nzt6I5ygHw2Wl6R/UfIj
NGkw+5KFtSJ8EwAgTVrwt8RE5Or9uhS7qxH+JiCYfB19dFh0XYf4RbJjn4DyZ/EFloZP02rijMk+
7Bpn++M93DF4O0MnDNJbRNOI/p2sbgNQ+ijiX4s2DDzXWwfK3XY9uzbev7oiVUMzET7/BZlI/DDG
NG+/WRszWOjPINfnAcgC3Hq53KaOD4sY5j3Z67ipAcGrny3t7vdM1KjtmOE+ABW6hKzALPmlSPAd
g877drKSA5HTp95/XTUyQl23rxItrwjg/ZwJZvBt0RWi8ByAoQwPMIodnzEhF09oIs7fbqUFbJeN
tSHIdY8EA1FZku+7URaRgt+ROdzlAjbVweMagCdAkrtT8fV/hr4MF2igcQmx9Qab1hFg102OYaI0
xsYKZGp14x7PIwYZq/0MmgkKBItgxItEI3wzupOWHe4KViaHCbw6wuuDeb7o7sBFgsFFRp/5/KcR
DDtFz0ON0ckWqR39b64jUN5Q/ZYpZmRyatanXogOnlDLDR2yKNm/p7E4f5Vhu9KlsJjwi/DMdMi3
qb9GRMZ4X5rtWQ56f6Fv3dvGi8gFZ4VPsTt7sFGawrNT09OR08Uhwns7GIbNquOdtP7wI4+xw+78
9RivSTTG4hRnb6B1boeKfk4UPamc50G0t/meCsnhgNevXH1HX0ANKdPF4i7Gcnt6XECirQwlvj+b
ECTn8NiNip2qHi254YC945JpwCrs5o7A0ukEZDjV/KQSnKsqhqXwA/bKGF3SI/YMtkPz58a51QoE
9zsmxPHwh0l5RFqw+/0GF2VxMyECnxdQ79xcQoLSDgEsTD72Uj3y4VxmIzXn43YBnj4PfHBsHmCN
JTGl596CfsDq16B4/WzzBYTrFPp03fu0NGzk5tXjVTmB4rPgf/Of0om5cDMbSDPC/8P/pZjTd7vs
K2x8zdRx7+2DvZgrJ0MVaxbrGI2ZYcBW9Q9Yp6Zhh0/rrZGyAEiUaFqGZ7zKZUou6ssO25Q6UcOr
wjbhn4TD8L1NBzleGagN3k4/L9LEGyBPgSpvNTmJJ5p2dr9teASCjWCaFSyHTlXReIK4J1SrDET5
kYy6XMrFwecn4e6Kpm6kWnzmM8vo/AQ5bSgbQjvMEnlVpUzDYYH0eJOU1rtPWlO+43a8NA0Ym/Sy
+3YLxYuSIHjuY4JhcHgA9SvXtR9mhrR6ppN5Cvxa29bzlNBRKyjVuZH06EIvFbcfWP86d2hDZUoB
ux+KlICJc7Yrg4TMmJBBsU8NTaRFLaJ5xuxJylsEtDJvTNFCszIVbjnOIl3jiu0qzqlynF6hZbtV
teV7CR7lM4KIO7eBaXpjPd8G+4wQcwhMc14H8v7L57qdP9MDwt0dHex+J+hvDGN2lzcjfKiQ6b+S
aULAigKCFrmmH2YBUvwE5FvLyv2G5YjG2s6ld3XRboSOXBzyYrAo5vOiwspU1zDT4QfeJH5FuXf6
PQE1+un9p0VCIKxEYqWoG0n87+W7U0r++Tn7tRq+a+5Fx6HpsLNQAL4ydR6q2BbiDLEEmQhTXj0P
WGExZPogLTTNvJ75Uf5iMiKIMwtDj4PPny7da7oHMeMmj45oQXw1YYym8a7rBdi42fr5lhd1X7DX
sXEiACv8lov/QlFfM6ipeC/HKieRJf8OFejf0VbobJHISBEjy8PV+bHfNkK0A15gRYXxF/qCvvFH
SzMc+K/tUBdDPMnY27OAVGE2lIrz2ZzEooDC5m28kpkSn3at+/z9NsFHbmemwrNQFFldsEEsz4Zt
CBLQuwkbKBOtulT8O0g3SQpmVhKgDUsEZq1HA90nux0nrayh4q4dTcaOBux8WMvAu3EDfEn+pW+1
zVsTiXX9Le0zUg0OSyXcM2Esv6nhemGMd4ESV58poZzARe6B8xPSla8CXDLViJp75mBCh8YZAzIJ
AxdEJ8sWL0hN2xS0vB7qAej2UEshNdnxPuYBO+jHSeETJ3Ec9BZpoSWLgl0C8O+2uEHfX2Niubmu
NcR5ufy21cqGAiXCFj5xAgZldRprYu6/cAnYcVB/Nb2RaS4pAGb3pXc61sJu1ISfAQIWZrYmx7w+
8fL9WZ7Nh+LpWe91JcVDa2VG/mvdKsYoV0bydebRxM5T0qVi+7kV8vL5U2kKRlViOnVuBZBsBpOk
sLYw57GnckCZ/lf6nuoUgZV+UnU33ycX+6tZPNN0x9e+7VD2IE8qTSJE36GxopBrngoFcmbU2nQc
SZ6Y6DO1DvA9fursdFATsKE/H46RRUPfvnJcuqoJR+f3geEOkW1SM5yNXa3qLiLeDWciiFsIhJXB
nh8vFQt/l3zwUQJS+XZm618wv1DMkleOI1Lr2UuHEKd2lw1C2g+6hv0E8r3sYq5G76ctoAIcNLZF
bFGBnkyW3IM6D5W0hgvJBvXcBtuYC9qmJbQT23S2+9sq756nAFppOjSmNQxI5N1tMTDM/XXI1xMN
bfUaHggdJNU91XW2uaaH1n6vpMlCT8qPufwuHiiTgYfTDwSkO1iyhMAza9HIrTEh7/nBypuDXGKn
3lUsx4pNNxc1gqj8MRm/H7V71Ro6Eg6BkmPJchGGHPwETVzR4xGNjwkY3cHmluOLlc2XvgwFe+hs
yqmKusN/fef+XgGYVImarDd+A5eRCA+t9IXoHZaaQPjVvGGvCtdilAGI0K6Tdo3F8PvK/n/NhHqQ
1aR7vWkPO8gjE5hR5DHPmyStL7+C7sqIcTL4AxwbUXuR3cpzVDLkWxrogrzEL1sxY20mfE7PozDZ
2/aPsIlv12tG79tTfSEmeVtxPJgqzmmIDzFHegVJxnZ9zI8hYtby6x5z5sf/cqKvTLFoGOQtkGyC
9CY27NVjIe/DiAZW2pa0kDEcwSwl3Wyjs5LMGef6lAn/zSILC8q/WSCFxjCB1C6KyisRwvzE2cMH
ELacJrLvGAzXOxEKaHZaRlAQIWNtfauGsqalXUs8AqU4CA2uoMHO1fsJNnAdDJE9DOPy3XvPUjx2
5is8GqdQe41bW/OO2rrWiy19iTCi8rIDGf54zJo3bnwRp42b9Jwhf6iDkpOkz9xXRfJLS/j7Thkz
2qYNFEZkox6iFLBHrQFTb7ArqFY9aURToJM3EeHrNdF/IxUjkXYF9Rwl02u4KxuEIsU/A0s9ab3U
ZEyhztZUylGw2AocJcu+h7kyO51DbSFdAitRZnY/nrtX0+ibHQb7kVqxw+jLC73ez3hj4WuVevyk
XojA7DhssNU7Y+dXbASoBD00VTQVJldIkHxrY/UjoqR/6S3XYy2MlaC7SGZmOHpZlCFaZU6R0nxu
XUz/GUiU901s3BEHW/yTNwQN18Az8mA9JCu/w0Xj9KQtzwNB/G39HqnP70k+O+iLOH8QiJKP2EIW
ye0v80cMCKLiS02kdCi/8+PC1Lxp2e4K60fd2ofs5wrgeAFOivZLs0JR8BEiddbrjEMrXa2V06LW
0ETcNtZrPYJfXaArndEYuA+qq4w83hyWVNYr7ff/BuAL3Gh+MOcnepqhvDr6H9xZrJr+k1UK/C2k
KEaH01pPezLBxHbuCHW1xOids+XO8/6Gt68XV4d0don/5RSxtXg/l5NchWvO7mlYAbWtBLWquR49
N6tbZzBYby0o4L3eoXezxRpqu7h2FvDaEG6XuDzGnyTIlQRqCtft0PZgiErP+uAG8CnqQtKOC9/c
E6rGO0UBWsrq2XYoCeH7G9mqqnKxL5x06A5emb4GBrPIN/mS7pbeiVeUWtW0kD5zi0e+TPVm68dY
BSJxHCRZG5O4izzmzdIujaAuuYOyuRR7bmUndqNt1osZhPhRg11XFQ6LVXj3o/PHdApnFunoHNHq
0iuZVUfQuGuSsa4pBpUUzcwceW5eVZI3H4s/lnFmH1lMv8V34u8vO+5Y2U6nte4guxyKhWYC4d7I
idnlUIq/fgfAGbpq1V8hfK6t+71dYbwcpiLas2HHmmHCPkOnkSPofvE3t9a8EwB2rfOq3a83+Wsm
uMIHWBgXUADQe7DDJjqYzvakwZqRmskuLmrOAUCg8N5Dh2DOiXf5RAvQZNLgUsYM52/6Eqt0xbhS
gzKUXiGugKjBm8tWDgos7GlCUlK1qPqLmCrZnSQQHywK49K9QvymKNIXL0CV+/RK77DGiraIn6oT
oK/+kreIhsE7CPy9SJVlTy2yQNuqeRYecOErYA3xOeFuKUC3LDy2xQ3+8rBJrkCSzx8ghqU4BGh0
0iBlTe88xHbUglO8pzi9QktJqgA5M4lI0RFn+6Vb/4ycfbi7wkg8NxDCQ2jDuqLSmlocC4LpxBKh
JqlSSk4oDsknHIn8LqAejyBs8uGoBEvwT+CUBmqwXqLRvkNNv6cQvwh++KJa7hxWT5VSlmjAHZR7
12aIWIN4SeRwJD1dX/k3DIsjV1lBO1GTFgONFwb1693fZKbvKf8/1H1Atqk7hSMM5A9rzO2Nnv3N
1F2cUV6XFfrQgR6S9oL8IGD5wD7SiQaARmzTDF0iJscdZHx8rXKViblcUYEr5Sx7CZLMcPzxYAvj
0Xn/+GeV4eetps92qPraRGMAt9SU0+0WpoQjdn//8DOYXQvZIfBylbCGUhVwGo7BdEXlap/ObWw+
yd7RggRPm0fKDCl2oqTryhXkg3aeOSQ1t9XY1iaauO1GodYhB333lEiMBnlttDYd0C2A2OnI6/7E
LaQAXSgIjekpjEsj255LWs+uEoWFOLyTxUDX+IcsQOLkR23GmFDAtCDSy7+mGi2siEC8VEYPdEi7
mUbINr2xxyHXMQvkSvhkGsQaCoWhq8lt/yvD9QOEihGJAgKNS1AiTZp+XiiyutgSGe6atde0KTFT
l0Fjw4tGaV1rYmwoqTJ83xtbeBHuIwwtgdN4eQGBhGGRBsXTB8cjXnvkmY/lW1hHByuzTNX0rXOO
mSDDbuWbBj7K5mxLtK8Sem+QP52L8VD/tEdGkmvYYCRotKl24qxPoU+AAOj+rnlKw7qf18QCmV1F
GDxOYlzt3ExWgijscjh6xIWqOtxUYcQRH9J+MIvW6RqW4w4Oe0vogjGwpQmTArNOU9n25Y1Blg8f
8cyaGmOivnJR0Ohi9bNCUAclhY7PuHwgnPHqCLQofCPKvo5USGFVy8EdIlZIGotjtpxlnCNnxAQS
48EeUnrxWUrwIGCeHcjZtSKjdUyPE+tRaFCtGmXUSeiB5Zc7sTWoKfpAud01F0oAJKWdx+fOIQcX
UaHr5Z+0ry3ygTwx4zMpv5e+K8+Gqcd+gDJkv40HuaUvm/wGxej6HCamyHEYZlXaWJVLwYeEIb/9
GTH7ENoa0SQQfCCrMJtHT+Kter7hDP1I2CwJYTUl9hhZcBXN91csXPoiqrcGu8wPKsdXXViEuhXF
FHydFtRBIa6tkizsR0Clrajq0LMTxjWNEOFu4nbg4Hw6l9MysNa2SV93cDnWMOErv53eGZ6jk0Vj
ZepGfm8aSk6As28C9Kcsnn+GgZPjwwflBjFPe8RQ911EH5koyfSl6/dv1z97NgHn6zJYZQUnk+JI
M6BimQ9hCRRl6aTBuXILX1DKicfkOJ1TjBU8gQuVBI7qf3J9XGQubUhAzneC45BBxXjadQPwS0DL
lH786ZXEyGh8oU//5oJnfBb+r9+S7fOqBGDyz3ux5sLqgae0JiKX9txA7WPhnyEMDmYQ4Y0oSEag
PoXCce5Gp8lwcMNdTKSYcNADlWhSMTzjmC7K6DVARBCcC8gDfTxiPx1J5uTNypUvKkt5sLi8dFhU
1qPQUyu+nDAEnzpLR5vdt0jPWqsksfHjYVrsCAwPq1uEjgvMOQv0p3W1wSFvXU4mn5FUtmUc7CS3
hwMDAZ0E9XrQurjRhKC6bAU4SG/didXb22iibJbOjPeKwbXmwU4dnAc56sccGdy3sChf4bedRrVs
UkV4fL00sKtezYirWWondDCm5O4ysJ0lHGQ6xS9fMdxpRZ2WtCVWMuT8G8DYZfHI3eyJxq/cEbdR
XYdxrkqZQylh8sH2fE3AIYC56a5S0wA6xThpd0csSES6XWp/lEFadI8WZGA/dXYd3ZvI28RztFUB
1QI6zBvGoxV+mT+O/eh1pvVANpliq2mnf75Ko7nVm/TDontkJctpxZY6ozLhaRsdUlihJlTBRNGN
6lvteQlPMiilxxu9EvnzJKNdyD803AqhlryVg/xTl46LAAfXnr87U05iTpyDlEa9mskdKYnceTiE
DdUKlkY+KfEW3lFrc+38vKX7XOa3uM1b7VaVgKiyHM/ENtP5dC/jyyE2/XmJ7VKqeKbwF4PQqPdP
nS9gHIkcsHE5p0IbnhBaqxgHhAjNvBzeOVJvnauBZ4VRSTPCpf/PYY5hYJDTjlNA9VoZHn8/NAXg
UUFR/+s6cYYtzlEV1JxNXDcF66z+4is9/NUSbhnghT18rXIfGhDvuCyaF/RCg7bCbZ0qy9gEGAgi
3iuN/wEY317sqEOzFc+05lBbqISqw5GLEtRe3Jyo7MZnxA3/QTahEA57iDnInckdPbG6TAk7CCMJ
6FtU7mc8vyDHQ4yS0D3RrKrx6o63apAArrA1fI1rK0xeO5tDPj/A5vmfECgEctyW3G7OHrMJ1Trb
y8JPpDR92VEUMygGJzgEyap/FOhoenz1qOV0nnAuEm/gryFRMytuz6o5mg5IzkdFd5wz7epyMqI6
MWo7XRx0okksLY6oBBbDPqAaQvP5if2MsYPWDPYYSHNzD2uRP7XAxuIomUPfbIERFEkqj1cncc69
jcGWQMEqyI+Gw74BgwNODXiFuCu3wpScJFmOM57fVhr+0XAKzVHPf2ebKv+PjkW1O6jqEbGl/dmo
yYb/Kw4XOBB2yJa1Yh2p31sp3IRo/Sugjwaxlyh/CpDJRNYhgAQOBGJ/AWPsIHA1TR0e5l7Ilxh9
f/4uPo4vebSQ+jjnAFy8PU31U3KOiItg5lwDhMAK+5QEPJJTdpGuDlJHqfIKc/orqNs+m6jHusCM
xhFsMMRm0CL6/z5mlDC8l/T1QF1aTk2v6p8ocCWWhX26ir1xO5i4Ym5UN5A3FhaqOcWNf6DlOIwx
vtwsq97X+3hhEqTYi2O2o4jLYv56o31YNGyPp8MReAQTfW8FpLCWn3dqt8HbprxqFbMmo6zL51lp
h4A7QS0xNbWfIJgSykUdXQdoZTGzONRfvBUNxK24ZGVH0lsYOYvKOFLLvDOfXXjYtAnMFV7QAjBs
2+HDDWh8KqMrwcUCFkC378pDgoISlyjBpTVuSl3jQSJmcbofIGYzq5Cnh/gmydXOz2pmH1Q3A1KT
joJuRx2TIrY3AwCIJrEgEOCuYCR4O5uLf2yVzP/wqgtUhD8hDFEoG6hNAtVntZrEZ7j5cw6SDoF7
Bf+QkthC2IlqtNwab/nVhRombxaSkQchuz9rvAxfTRl90hYf0GVgR/efqLgiK0OV7mk2broHOn7C
2fqz2W3zPoEnf7u9EPVUcLuVDwDXQ2QTukJWpAHlqslzqoE8OTp3HAHWjAXW5WAwrhEAZEegjyKY
dii3cEsPlW0WIDvWsWELfL6jpQJts6RDHVfCb7YtuhBNor1/bsg8D5EQNaElm/Ug0HqcpErvHC2Q
biksub0IXkG9mp41YAwQEkyuW1T6vakOOwe4qJPum/DvoNs1Mr5OYE+Txa6zgxSq2xLJOzUAqYok
X9chPUmx66oCsVYS7iJ3dqlw2XLxhyCFCZHnlkEuon8OJfGtJHI7p0788x0eRMdSU3loGp4AQBRF
Vx90RP/CNDLoqK5XzomwDDSaN4JXc5HqdF0al5SF2L1Fab+83rtdK64HmRk7LHfq0YlcZfGah7hJ
hdjpJnhXNIhZbv4+UHZDrc0sanxsi9RvTK9556qw5/AdrWi4sfDumgTzM/Iw+WOfP86pQ6Jpv3Qn
qG2E+wMIrjjOOQlGHoPGQV9grRn5u8YcJp3CoBOvwaX7y0xNztpdmaf5XGtMhkLgiGeO7oWFsFUI
93SyRfGebLIMI8gyywfePAaq/niVoZeEzgPf9dpPnhS1xrEMKCm/GOTlF5J568umL3zgVIYWbp5o
fRFnalyyKivv9CWHRwupPAI1ooCHTTC8K3Rwyv8sBZlWHu3c32utZ8EVi6Dib3APXEtSq4NAXPhf
mvulIK2AogGFH4XCONqy1x/QBBvCsvGjKVtTyjAoUrTtwtZeAB8p7hIE3TJVnPaAkwcqcZH6/3QM
LljPLUalpzrYvkYIgY+z8ila/ai+yxM80zhVDS3v/8wUqNlHqTD3BOEVpLddItTb/vC9gyRIZvHG
nep1vYGlUwUlPlHRn9rv6C9Gxm+dCGXsP1kkBwQLOF7MQeh5tgxaArOtTqIr2/VnXN/mAcCmUJb6
0Jo+pgtZlS4fAfVD07oVISOLLIFUrPvNcC13KCfGUdQhDHKE2uPM+H3mzGYZLA1tED6TZVfCMp3+
KK9HJ7uGm3iL7xz8U4/tPPNvYUSg2eT1v4geF93rhyLqSNZw6+GikVOBTHFBcNDUrn1g5NPMwl0b
oWVT8lyf7ai/cfU94ibr5QD6rbBMn20BJHVY0/xmhMxMGVcWA/LlpSxdba7sbpBNFR0ptNcNuQkt
yu9OkGnxF+AF/i0ntdy6wmzsvs/sK4BXc/APPjSCAhmScI2/ywybDgdFFRscgJFfVa2WjwwoO2yz
sL/oIQc4MEfMUyyRIR6tcgTneeJ1wbDmcpqfXHAVV+FfR4TxLgLMDt9xHKhR3H83g25voo4uS4yp
vULTNHXZ9nVJArd5UZ+TKI4sSIAFxWqoaVJ75UHqs1Rx0udICiIZtifh+ZX2Fqt4VLxPSQWdv3pQ
UW0ndil2xrEaoO5uClKrJ7H0jEcXZK7UgBk52QZpFg/EN3ZRsC98xcJAs0CBKAA4RWBSkSvXQ16a
Q86fEz4EScFP3NCUqvwkIZpaiYgpUOOZ2Tr9u+43b1BXXjHFP9RUNR2cuGF6TdaILtBts2SZo4LX
K2fBxfJs3pmT3qNEw+RFoBoYqWyNdCdeTNj7elhwEdCQh1bHQhJSCShCPcXzWpO5JJ/BrUlHFnyZ
QgcIKxrSWFN4hEFsAn6L3DxhphWuTrmto58L1LlBPcx5n8uAR/5seUzbJTXuyFmeLNuMS3Egono+
VNdxqReaSsXe2ZTTz0EmC5fRbUMXCCiY2JrSi4uy9ZblZwUvWE779HZ1NfJtjFgc76uwwbsP2TzE
Jvx47CuXl6gznqeo+1Lmjp+yu4y5eREHAjVmOguxeUiY7Oyan67bpUY5U9/rPq44JNcKa8jfVuZu
mbhjuIyBePhtwmRRE8FD2uYcashuy+hix2SMWGI/1v53R7omqWvDwGxqC4Txg74h65it/HVktOY7
Bxnt7BmIvmu7vIhdXrJplgDNB4LNNQwM8X+5Kl0aicsK3rT1LLpsMVt1wYK3tMR2bsVGZhP3CRO7
3STgXrLZtJtFMXfBHglsDkZmFix6X5nhRG1PZPpQ0DKDenK5gaOE2So60TrHI2jwJf+L3KSdgmoD
ZD+ktqAMsl33vXKcc7M/X8wnli3OLrJ1HBmaWPAh1pW+Zf5YuaQlvYtXgK6g3ZYSwDhyx7e6+nF/
tw2vftT8+S7q6gUX6X22qt/UVIyGH/p7vowTGsgoVc5NO1wtUeFe2nLBlTULST2xxSKNHqxirHUa
ePIuP2afIgSY1mjL0H39TcK63nCjPKvVDaDZdnr8NlmTkqiDc+1UEjh0Ba1Ou/Nnv1PXYca6H4RI
+taCiegnw7J27ioDZdPKJz3IRN8YGL1u6dYwU6TsDXvo6tRNYBgi0X7o0r7W5M5brCd7a4CxOA4b
ooYn/za7zZIWO5yb4iIst1NPlQHn5tPqZSEsOV925ZmzY9gWdmqxXGV+FhoT1BDvOXSfV7LMr6Wa
A/bGSorpdC8DaTp9X2/iAJCJwSmRyrovVRsRMVTdEW8zBziPIoXIIip9B36hcQHHZfmqWMMsYWet
nZX3AO6FkijKXcarl0AcK3FzmcaUzOJWlOnTRfN9EqESziVX1W/yhJ3Od/56KSs5c8FsmvPLpY8q
+A0qTjl9zMjn7mJh/OPoSmrOWYSiaw1caG/mgDqVgrFGbn4kLOblNZaEzDvv9I/Rgu/JnyrRP3OC
se9yjm2cN18piarNTrRgQnA0W03zyetDthfOX4yxwifWE3fdGyOf5+vFboEjppS9RItqK4lPSChJ
77LqME+P6vmUeHHN9essREFR1e72Ie1nyRoFvEXOmSzmf+phE2QFu4wqdT7HSinckBljww/JJgwU
JSPjNy96jxyCaOOSCdwKB+MEAq38JngY22rDO0S0TpthLIyZHN1OvUNjVQf7iiWvLUhVyA0lbhKK
C3uUyzWBdNLcmqxh3NSEdWtCZTxHPC5uaauDAuquBo4XgYUWVpHszJaxdN/rWJaCQfoMtYz5h3VJ
GY82LJoKY0uwQn3FTlwVnx2uTE3Vmm2eU/LCFoBSPr8L8KDaCwapKGd6+Uqmlgn0tCZMlU4pwQYq
0K295mnAr9O0EVA4TvSMT/QOZtVWQ57mrIy4F0lcph/ubr1Gs+nMOKUOQGj/wwf9nBDVnzO3HzdW
9CgZ3w8X1pF4iLszH0EJUcjL+w7V59A8S1b5S6kpmdy5gE+8QLaaYElFMiDSGeiWXqhSN7NpYp+I
dIsveQxoMUYfEP7HUxzx1c98YnaGY38PMbeglRNOPDzpbR8CK/V65RtfJdgELK5JeWH4sVHqhSeS
Ano/rHE4WtwjkP+bMRs5P4VyAJBqBenV+8lGF3kAGBiKbqe5LsHKP/5ZuIC1CrOW8msH7cMj0ehv
3IHH2fY8c/N42K8enZw8sByKwKnaSugrcuEYhLiMJOr++o0rbwK05GOyyvIojPucnlM/mMbV2TXK
dfnJs+sjUCFmtB8kIN2Ga4XPn5A8g5+MC+DOMTCzTNwpWkVE5nwBx2iuGRVkyFG4LF5eGlKyFe7n
/pGFTmoYSQUB7opxhqutuPvB8G11U5Dvkr2if01Z9JZNzlNBXA08Is5EaFTvhLA2f0MyjurteBlT
xERs4JGxd09q+hC004Am1Rk5cAPatxex3ORfrIGbfdio58O98LOtdFpKSBX0v4V4C/uDIUAnZKXT
7RmUgCMmDR/biWVLeT5zJBEQXmwG4kYA1SqZoC0c7gslvvvVVK1wEMeW/1dQhoY2T2zBrj233aG1
E3tHknIco9gLeChicdQ4BXA/zMARHO6S9aF1wjCX2YwRZaJn1cwsV5fQ94EMVcgDBa/667Jc5EAo
6tIIG52EINvRpGlOu/seekP5cGc7AlwsUrOSMFk0bWZN1rY1xuR6TPcgIlScu84ziDFJGzNfrs/t
j88MfF9qPIkRq3iW4qyoNq1XIHFYo6EyoEipzVld4hcjTKqkqWYp0A7HEA1jHMS0jZ6y7SnvGPFU
u7t3R+ffSsJih6JR5Cltt7QtiyqFNKksdDOuad9AiAEHXAOOFl7DmKoLsA6q/f5JOB8Cn0p8agcR
2EM9OA0SNXD3DsXg9p3HEXzn0rW2Tv0dJAq85STMifSjA1/OLPZXgib/uLOtC67BIjvl2zadPHxw
QdKNX6sB2LV6I/AJjI0mq6D/gWAus2bhXUJt2mu5DR5syNEIPoB9KSTv/1WacFjXD15nPIKvGdT4
KOxe8zN7liCOMPTvL/Z8B9RZJmQlsqTHNI1kZZe3zK1KHOUFaf6832NsxR26TgUCu5+a/DgmOA+m
SSjHCzTdONSPYpm6m1BzA4NjOr18W3cftKvKl7hm/soCZW7BmzH+NbwjXlDs5IVAVqo3MWCeOpIQ
DREsNdZoLrpDcjH8DO4sBlrKcAcfMKDsaciwBCT+ktdC6K19NHQgblNqCH1YjjDPMLwcAqBGsf1D
UeXx5+8OOExJr00ho4TtzGgNaX6/s6vXGe2N4CdGdwvaOcCWGr8Nq6HpY0tFYRPN9b2/J8UsY0aP
vfMuWPKcQYZsAr3T3dbCm+Cu/k1QyT3N8xoImUma2y9QcUpDTidjAwFhw0nPpgKXr09yG7tOoX68
ZIE2HWXgHJCaKqKsSS4qsJ86HoAdIwGgK3z18qt/ME2ryN/XJ8aOfoLxxdFGNMZXg9XT9Wt4lvKm
PHN6eu1Zz10W1s2bqCUAVmlM78oRpVPj9j4AumjNCA1RMNjazrR6R6BJC3Mq3XKP5m9oQOEWtJtd
4Ar+om94/IjnfYgyGvb8VvvNuDzPe+JDbFFLHwi6kIA5ztPLlfu3QMEmAr7dcmVKNX5P3l+xtXWL
Sez3QupPiWEEoRATQPP1Pf/txufiawFqkDJMQ4og4FFOIgg53tFyfp9j8gE7m8QvM3ljjQ85UNs6
3opMpuDwt7WSXrMVo951G3mvQnNa6H8/d6hZ8WGFgRy3B9mbguDTP7Lg+GCo9t40rB/Z+Y0KpIsl
uD83tGF82LzJE808pOE40zggcIHQ0P2co1th4iko34TupPhbEH7m5zZSaUW5xZ2r3g53Z7Y81ND9
wSjuhECmsds2mIu7/rBzgEJUzv3QTvwIchfDIMGIY52kcY8gRSdF6WGfJ144QA0sEnDOR7k6ScH0
ZrSn6zxnLe3xOFBbjA5w5YyCxqR1bn3O8DJPY9e4lVtUdkzQJHmnZ5ISxzc6A6bbDPXi39ZLJ8F5
Hj2ZU9AIgYpW/lVLMI7FctoEGifhAictZGxkmq7KYxzmoQNPsijdn1ljTgZwIRibgSkgjX985rtM
8yDWO4FGP2Lf84aMpwABm8r7M+E2Ptf8GPfg3jaxesi3HwnNl1NrsendDHEYcEhXKAStfeGKrUy7
ngWYxzZ2O8vrf7hYYBsNBlu36D5JSYA+JWAson0vesw1m6MEZIwGC8ZYmjeKMAuU+ChIAOtTZOU5
tQHtTG7ByO4ChIVKB6Z1cnNQe3ggADFVY+61/GDqWULRQ7LlYsHi+BwzWT2IqGIxXv4x9JgeM4rg
p46FUm5odNlwVpaN0B5Bnc3449bd0dfWddN6+x1HEhneq+jDFyNzdgdZoNDwBOI/oW1M0xmpAYdw
JMsefyZkbokdC+n4OJAcMiXFoCixUy4h08VY9L5Vtm0bDoNRKJ94Y0o9qgbaKE7CGYUJ9imZN2Te
AI86A0CWNC+bAmBDMXnrK8oorEsJXIqs0acyn7CfLSv52rNFEnyBtnZVywQZ5aQS3lXaUzfDJqkG
NftQWz1iujsSsijLabf3UKEH65kBa0AxkzMvRvPRDHvHE6Tf3LSwURy0rpXxkpRuUBO73jx/L6l6
n0AvuqbcwkLW63ki96aI6h+0TxCfXocYcvDfQQnje3p7K3E6i0R6tsT65DauxsfLKxY+AN0lR14W
BCaDSwkYRT5zsCpYL5pu3/c1Y/SK6RiBWZpViFd5tmx1IALZv5nJ01wgEan5G451d0ESW7MsiMSE
fDbNLgNUUkofYraDfzIjb3DEgKle/uZjwMMNNHbreklS6ZXj0Io/gZPuKLutY1X+qXCr9lfMLkyD
E3FwvhuiN+rg8efYn+swzZwQKUNmn5nisO8B7Ohq3RRYZpd0OeAi04y2NhHV/Gw/PxX1p2a36co5
gB+4a+7UkRltgAblu/Uc5FzytY+vbnvbLsXbnBiJJKG24ro3DEXXd6NDvJL6+eUj6fGbUCZavTCr
ulQGsPG3wLU4HDtJ7PE2xpnAt40Zglyu5Dh7TBq46RlJTDD5dR0Dtt5cOwdm5MSxoMha7wKsK6WS
z8D3nFHLhGKZQRdJjSiw7fbZP9iGUjqpEF9+7MekALlS445Rq1iGFgeMyuhI710K84dc/7nK3D/i
HnaPG/YmQ0b0Di6auhkhoIHV+o9qmTm3ct7kvV8ykyUcfU0EvsLTwvAezZwbDF6pd3J3M/4R6ovr
9D/ymSimritiHeHr06i67R2O1rbuYMl1/20oYuaGBnmJrPiRywrbSlgXbzCjo3XoPJE9wndacNBM
IuY+g77K/RPHjKKdfpuAYCsUSo8yfm0WgR7dtYxaEgjTraCoEDgiGkbKyPFj01Ph/8su4frVlH29
PMIbPfkY65Zqqfm592Oz2uRnmsckE95UK06Tq6t97wUXZ19Bbz2tbBsH91DcBOt7x/EGWHGreRAG
LCeMggHETlj4juL12QRPKIWJcpLgBJxn1hNkDZ17MJxx1bLCLJr1Y+FiTNW9BMfo4WixGZsJDCjG
FSDO0AGpG2oPopFn+bguITDidFqMVK+7HQGX1ZkRsIpcqy24GVlJ1Y0Z1Sn2VpqCqFlhmlyA6rC3
Yc65IwuTDfmRXKUVBqZT0MVWkRSzIsdn12eYzNYzX2gLgQ46DB3YtHyHs89M4GqZ/NzDMAMkQh8+
ru/zWh1RTxpyG2fU3xfnVMQxDs6G7cnvK+tfx2W724rGQZISkTxC9ZAV5dvi/L1E0NDPfNjwwzAD
KJsKcdFbwgRmR4hbd23SaRhXyUkhfA0Mp1OskZFvvcS8lPGwdPEZZMz684SVmPQrnlbQEU3SsIB5
w+gQe0mYzZGUkwXq0KffeVxpScr1JfFE2SkbJ1wzJimSBioihydIZR1ZpHGhVPZqJskPCPKceycz
/wdxMEONQMNp1erUXzTGOavACjcKuU4Ywgu/xCxk9y4fu/66Ddy6xwRcDwwl0rxqPfV15qZRdGrR
Y0TdNhslvTtLW12N0F6fzRNOsfkt9mPnK/XAqfIkv+rTvS494A26gCGDDTtF73vWB7A28//jCIul
T5vljGyY25nKEbWM7m+LVbptoCiKHzauFYpvyRRjpf5ws1/l6JQweB0/sDghwAzkS2kRQ4xdwEGi
5UezoE6nWRb1bj+OelQtYPWMv+90jU1yEq0c+UdGaHj8KZf9fMZDi3okLSweV4xRoP9h6vQAjg8v
FpWqTYeyFw7kN/3GXq1gYnejjvxKiT+6P9bw4A3GFpWQjOcMDHA5mSehs2WSOjwYBdQ6GDF1Y9nb
meyt4nEjG+EG5KsBkoD0c8/oo4HCws8gsRCWBm1pCo0Fz3XLFcoOXsPRx4lIu6CtxE60CutFpy/U
HkB/ZL1hfRCr4JSOZLbh5e4czFd5jLnPT8sqe6DaGssZXkmpmHB8kuKdokFZdnzKL3YjqkXJ+3S1
DEUm+T+/HyvczqliXH4kRtf99BurNTlsVR8BU4wbuMTFmbYwLxpfdb2wDAnJiAXYVHxLYMPGRLhY
eED3/PgTBThWdb43ph50abYZ/YcdbAKT1/BT/MFHB5BX0dQG/RLi6YDv/QaO+mr/WArmZZDKmqwI
mkWuqumlbqjNzqB9lzYz9GXnmsROQuVZiycblVaCk7HyDcDsUxCeFxBFvJ9evCcnZSjOg4swe2Nq
phyC4HqOSXulFzO1cPu/kbaRWJ7NyJcMxmj3/JJmqdu8inAX9OwqW8B3vjHYSwLsDWDz0p6metIU
Tx+yExOoSNP671cegwx4M8oIH087Ynz2dhxxLwgI6Uwnj/DGVreqpuq54zc53EwUqQqCgBnbnKbf
NyGKN3mBiNoJeMVSspViUZMvCt4v35+excdr4PXPDizyyFtDZ2SmCe//BgpCOytcvA3zhLjI1CPV
NzgYz8eIfztDiIYoVrc6waAsjuuj6csgEkd49Q10zlSCv37AqV1SLiRyDl2CxaNyMLn7cbKCdSL6
T4g4Finbof5tOT/+EPN7bqvXUIpajSGiGMAfLFAkf13zTFl0kFFMlRNHD/Q0nDjDiD7X5tnwyHp2
Min0lNTwpqzmGlOoAsiuoQD+4ZX2/fv5jwSbW5i1gdRpwBBJm256hti/D1+No2OgaULQteDSkiro
VeqoLM3udkD8wjMfwPfzlme+2RlvnIQ8c3Aff1UlOVjUYcQJOdc4O2m28J4DIMqM8bo6HSk023S7
4MR94w8fdFGykvVW8zh3uxHbN3OZiJz86jOOluWKFnJn8mq5w3nVJoxZ/xhp50b4lv+2i1BO7VYy
8zS0naHPr/XJ2aeI7SeWaxHfOQVHHE0j5yH8JLT/aRHD6ILybeEuF+fxjh2wTNIp1kK8FjQ1i2/g
V84rLlP3EoZ7poYJVH9ieIHszPEmLI8bBdZ6C2LNuVazafsmb7DLRbN5vrL//slfo3Tdv4DMnAUy
2xGbynjmKQUK1r9W5NHM1JYCjvwuuLdkNs45y/fp+RTra4PsOPViIth7+gU8qS02+XumDW/+XHE/
Zy1+b/Y+dpS6bKu/K3brI+zKJAGHlBnyFLFzeX2E8d9jTfoYzAtb/IsZ/yylJq9P/JsQg6aJJ8Hi
F9UVDpQd9lfoDJwUEm7eNmE3uIQYngQJaMQl+lrRPGn8sCWqoysdRuMMf+orqCFOI+wLcHXHk2IK
7JH83+gROCUAnQ0jMpDQ+OndzhF21NJnOt8tOtP544eEotdq0Ov2DNIVeKpX1KjkWzOXp4SWux7t
Z1HBYXOao6bYJtRiekXIXKp0sElBkPcy5c+1MaEUaxONwW/G7kHKvGbzOSQafToW6OVnJmtbtGO8
bHpWVtWFSTnHYLm0XApvCc7z/l+ap35YZ3pdEo/Obk7C1y9sKQ/D933AXBYSOgUcdC8HFyrdLrnN
nDMlDrBHKTalRKQZZre+6+91lmE/gAMqzDUf1tF1/In/NqMxQu7c6czsr04OmxhoZRenQtnQNlO1
nuBNjJUH/wBSNwimUruRMs3EMjPwznOLZvp24UOP4U4T/so2MpD6hZtw3ceOq248Qs0YLOJCtyEQ
xReNCQZtHz2XMEXnHk9o6aqp0MgLT9CMeSSWeIP+LYFBRqJBJJEELt/QKiEqDIQe+UwkoksxThdB
7akomSrW94ZWrklJlEpe/aKrJVXISXu5+Jy9Xs81IeojW1nhSJxr6516s1uYoouk7InbJyjGGoiQ
NjMyLebPXe577dTZ9n4eLDKUvoYXNCbqj/4k7IY7B2M/4Jwx/45JlMJ0SFHc+MPIm+0E/Ux/B5g2
9+TTtbjPBvd1OXEi+lNH2g37xI/+trD+Cvro3Tv5rxSoB5C+sTQDGy2DhnfJXwyYkW0LaqlIK/Ks
AXFzn/sIhZgIW6fgBYwd0fgCYc3cf7Fg/ADSS6cQgd8zw5EnUauOciK6UMSw3FhWBLmmIvJ+O8/w
//63qYw7pWnszm9PTY6SZEsLRb/BRQB4NyT1UzS/nCPHwkx8BY42CIBfJOLIuJHvsl+UM0HgShCe
g9UTAWIndKWjEbT2XotEEceemgcx8SXr5JhtC+6bwUstdjAFOKCwqPTtsqy0vyl7O4C9mFgOBsj8
3g+5nzJcULyy3c5QS9HVuo5GArfOir04508FDzlOamo+AH3ix+OTYG3KqCfZ7tdl6tXcKxrNG97B
7UCUfsF0qzA7Rsxut9FiaXWPWJgrlhsRVHbFPI5a7UwqX0i3FAOOLfaTDEf0j1Q7hrnki7aAPYqn
5M7BVEbWaoz37UxOgCHkFQlpM8ZZ8FSB17JYZmZpX+XSIgKxWBpPjCLiACiSiRUBGBwAUlRqzH+y
IRbe82Ltl+3PrEJkUm248kpRMWourQYvn9aXXztQN+rDcvQR9L+EYnkF/1/rAOFjIQXYbEiZt8Mc
7jCes0OjfGHlaUzZ1aK9ElWnBYC0Qw5byh2RtXZkanhH2iiBotVXlB5DlVvX7ZIEBguqz40dIziq
WKQ1VAX9ArEQBT9JmD0IiBKGlPzqKK6tp3OS6RJomctCzAxmGcELs0rjS5bZeY3cpmrrIz9RCEkl
QCNLdVr+YjvK9hYxBA1Mg4z/sqVzUXd9r3UAkTbMJpVjuB5cRQBgakNVW6FEh6UGLIrBam1BzAlP
RxzILsG3ZNyaWFSu5KUS8UOHR0kWO2/HFqzaqwOWE5+Y7AjD027X1MJhoUFOxcLdT9ge0FnDZfPd
r1fCQihnacs/2PXJ1pCJBPF+O6Z3cY1uXgIK+twGEigpuW3FrGn2qGD2ana/mayqVcc7F7mvM9ZZ
AGhVh/Jka/bJmvtBnnJcoer3MWZuXJlpHpPtDjZzJ70BpC78zlVf8SGZp6iIs0b0GRFnQz4bcRPW
rhA24PnPOcnOFU6mJQWceqgP1MuM+Lg23ZfvRQBCxCzUx4yuOHKkPusqtIxGHV2tRJweN91XzQmW
ROtoiz0FLLlutlBhFGpI110FIp1skiUvYYu6uug6vFT7eFpr6CvG93CMo9Fub0NP5BjaAB92z7P5
ILg+7I233HlyeAHRyjubFc344x09+OSphiEpE7N66DxWBF4Ah0qs0DO623+HINXlMrhP9VeeQcH2
BGscpWAOopjDnuG0jUE5hSWRxVqOjtyu45PAp2L4VxTWDtP7+TQMhRJagwidHt7yaO3S+GUjJtrG
uGajjvFu2bqiW4OC/5wmjopOQHTj/qnoHjacFEkP1vAk+IahP/JaEoFhk/65PrwIUyd+dbfDEXzk
Y2HMnvuXx/rUYV7nkLigm0SYi2F7tIH+qj+2VlhoiNi97t+DRgDP87hUDaY3UlXIKRdIIvykyBCR
HAKbz9B909NDX4zkokkGGAufqjX/TGiYXieRysoBWgV4QVQRH4NgtvDkUuvbbSqEWIKKxbQNqN9w
Ab1RRRQRu+5LChGnbaeQrA2sCbFZz+AV++4xilpqjrHjAq/opZO5W6DIef5zAM4wmt0oMkJF14gD
fOVv6Y8TaKVzIoLkSbQaFdsQzOvjt7syZizpf8iL3pEqXTpLv8wIoiSKfkvvoU8vgatHYEfsEfbu
GVq2mpmc8lWCaTvDH1fzskb+chuvxZm6PzCgVd2S0z3cNuq+28M9zy85ytF0wuJdClgOMGNGau7k
zywLONLLBXcBePMh+v4TvQIsCfOjeb3SRCS/cUzqWzVMcL8jV6OpB0U4XQkAETjjP+yxi/HN4SfX
6/HJozFll+aWyqQykvnDFVL08EPItWLGkyd8wbGCT3CGcUuKm9VH2zn/Ikk9vOfRXeZv7bfZgpJN
Ep8YDLWoBhcvRNB+JGiFF3/oJUmHX5Sx7JWOoa77ztsjcunU41NDWvoleqPyFvZ31IiXPZPFuoJG
EOWTLKF0Uq3jewGU7sKbe+JjinUD4aNfmVH92G5oSrTcY+3RKUGFRSpqxhb60QFgfOGnBt5zbAEv
lBEnAm6XMAOHILFhrANU5KmnXZSioYvzgFodJjSiZGmXRQIF7OgTcYruHmt78Np2/QSEjyokoaOP
BuievOhyaF1M4NPpl0I7Pzk848pW4DicLiT/s84e9YV3X64898A3fyggOlLfwa4ghn33L/E8ujrQ
MeG53e/Ln0jE7ctFMxkY45v6A5P0kJJmHwFuPo6NuCqU22geK84JEhxWXke3D47YqEs+D1ENFDnR
6FCOe9beBAYcaSw5WoeeiSDkw20nBFdYmDF3DYPhxzyNW4c9i5o0ILAtNz6b3KVtcFBGu1SRahz/
mlPWkSsNR0OzRA+QlSRJvGuqZ1nypVL+GEoEFIWYzEDtkuw5gWr3REl6OHVxaoGvnhpH48XoUivn
dnhF2gDoZSkEUEG6I5QHs3nzYYMJ7Y0sIBV5ka0ICMmRs/+gJPgJ2pe2ar5ojhBRDd1poy5q7OBu
T2MospqBXmu7CGqXQ2EZKZOrqhCDTjA852RHc8RAIgvOAjmzSzyu8VNzfO/38gKVwE2vOPLDu+qb
k7ql0J5M9vBK7rt5oVNyseKRAZI2RBmxGFjIpftq+abn3xbvxPBlIW5kAEq4sVja1piZpOh7uKPU
EkWyuo2iODfeUrlst9Sa/AFmxsTl3LtBbbeGNszqo15paWqwUi2peEVXzNfQ490rmrOQJHgYIjQD
0rDmzqi89XXhVn+8UWnrkjCZ+EddfhB+L6QpqtrQeSOxXy2CZhVgSiEeA3DETrZ5loT+m0Ym/YWQ
PYSICH20PnqJJWeN04GDOfoWQXbaJ6fgaeCUm6CJLMGOOZtOYwrBIUTNqT4bjJLCOmu+TCYaLsIY
RHMEcoD3UP+g1cCKXOC0Gu8jb9U04MptnAPjQ8xhmTeeoqT/IlSJ5DkyUYp6xM1HYj3ZEVuaPRbU
tCfsayNGCx05P9Sc1ypTaDyhUQs2dCQu8OplUGSTYoCHOvJUgIhR/DTzKgzONM2GFL8A/AQIcONI
xJc8spbEt2RCufALQdS9oNaa1HyVJq9il/oWxvfVmQuxBQ4Utwfv4ZPG60Vfc0qMDrYLiqbpEGTG
XA7xLDc2m+rm38z6p+OD5ZKhYgROwIiGbjXW+dmv30Z8mAo996s2DFe0tAzvuQZgmca2tOgtGLEA
avOKPuZDVGPSzkgtBTC+3El8723Wqrg6I7f09ExaGZ+U0pTjh6HgZ9z+8a2s1R6ymqdD71sS3gV6
5/ieS08X32qe2fZyKgSDCYRGDeKM1CLpFVMdgnqotO+3fGNiDrtUEJWr/3//lSGo8YxeUhTAtNGc
h6lnK+d0QNxLCI/HvSP43QAeLZeZU0AtwfaJvXCBTvAL34+vP0ThtHiWoQQwpa/jeJmANjNPKIV8
oPpXa/1bouqDo+e2WRpxXPrja2xtP3Ke+P1Ziv9/MkkTonfh3UY2byS4++RymTMTIfdAWXgsX8VP
tC6xMWAX+GhG8QeBUis53XSrL+QCGfi4wXfqZkvI/LmBIwsSkw4ChlrjvKTDhfObqzHON+/3U9/4
nrv8vZT8lqr+JkkG6nSQowj66oFAT1sNR7DlHDM0q2YWSpPmluT8KFxYlwjgI1Id2Qi0wdG93lxq
2W7aeh7PypPRPWFh5ttmBJE8fioO2gUDlb8+KUXCmuWobKX+QcITozMsYp0CWBXQuxU9FWkHjz4M
S9mk81KFnoscRK8Z1kupMRS445kPG9RxSgoFQZvLVnknZ9tgQQNgkp4BdqcqhIdA2csxSln9NqJm
OGRUeXjlBH7cGT+cWDyOmObZ3iOfILBAUk77KSSgQ9BYE0so9t9SPm7FvObkHWz0KcMf4tdvY3Y5
ZFHUPRH5f67FFIqE6D/vGosTPFM8/0ZXqaxLKULNX/ADdHPOByXPoiRD+bOTAPp/+PrgqtLinmBc
dTR2DUYvNXC2tNS8rzNlFN6rWDpP+vkUGgsUaqGV1jzq5iI4GIstzfs8YD2rbgxRhg6MtpdvuK7p
4HSYwozsQV16bYy+eUyyJgSzgU7K7FmXIq+6LYfi1Os8lyEkozc8LBBXWoBGRCQIvvfjRqbzC9LM
GcyHRWuPpLfMJnR/DVZLf0Dpz6e/0WHR9mOHw0Gz6svEUmT74AvE2/GzLlespUEaVAe7AyiPUsWN
HBaKJkW1obV+yE8ON0NfuFHM3pEcgYDQ/AB1fTRp8Ia+ZvsBqxmV+ggaguw0Ge3A66HRT5yU1CeE
QfuqUsLtp6L/+3QjJak3i0Sl65/O9LJDj9lU98ehtv7ZftUrIZ8lR34yvjo2rXZW135KKQo0AX6x
c47AARXwcHKEwx0jHDTCpZI5r5Ax/xh1WtTPY1Nxh7A+M797UHN3DRDvQAzhYjlmMxCN23RI5WIP
WKL+fC7SzTdOsC4nOkTvwDabwP1BMmun1Kyxg2d0TmaheOUbiK35fjZy/dP9LZeR74GgMTrvxFl+
DCxPl4jy/7WP6bIr4HFtJyV/fx0YE80FeKKsx954gx3WizViOObFYrxvedXOjjGpAZyWHzbILWqA
SLo6BUQ/1GjcOoyU19nV7AHc+FsFkKJSS4Af2lrunUg6MrzR8UqFpf4WhdLLezFgPSCQru+LyB1F
EknXO1/uKfqjBWbgJrFZfBn+7XmL88H3xwOYZJ8Op2LQo0bXHMgh3eKkgRJGW3/TNxlhNA71q6gP
MThbnhvTOQktdgrFCT4p9y8Jz5J9QAbjxDFC2+a6AAlzq6SGXhfygQw+edWqIPiKHP9Z8empJ4gv
1isvOrNoTgcsJ4sdy34U7AZCffMR0d9/MbedkAn14PFLg+jCr9+06hxSUacgWMtNpHlNmsAWRO73
bcqwt3y+d1+L4tgdJoJhDuBdX4x8gTvQAz1GI5ze+zJmO5yy4NFQBsRP8JBUypjo8F/Vs0Nh45Ij
6Yav4tZFJs5xoRWMA5y+tuV2K+MroXkucwPP62F/YE1e8iaYKhY0L9djfVYZOWIdVN0rByQdbN82
8Q995bAaVpp/nc1RlApI1BrUwDmaa283bXod7rwUkgMug7EXas9g4K8ZPmFkbt0T23WPuMf8bsJx
869bGF6kDhSeKfW3d41wjj/qWm/5hFdz0juf56iLM2dRclXH/pY9aVXXSfS1zVr8LfhtOQgQbrh9
rDSJ4wfW/adsbpBiQhlcKfpYZAkbYEoVn/kLNexi2Um2TLRQLnZdNOB0UZciomdfpH0w75LwV0xp
9ordIB+/KafEWTXs6isPMys2AEvLBNXk3ETzmZbTsdnb1FvDvbtEptuN7sOAQrxqN/H8gWgXJl5E
+oThe96jaEioXyaz2Cy7uvT9zIl0XwArvDvPRXFnbxk0z7VTwHZya44X0jpdFplQnQtp96ijL+BK
uQ/u3bYSIsXVIkFBfifEMNgntSH+yldzJhwVuTKcThJzwgzWUa+x2c8mcei8PN9icMvzgg2AwaIO
gc7AJw1uS73zApaL+CeXSiwxSKwFTfK1Y08FNt7CJE74kC6lMJxUbNSAI9YBVGRlCwSA5TBQuVrS
FIwbHgGcqYSXEYqYxUh2HCuYItXLpDTBIKjET725pMAKkMusHnPCmhiA2Jdh04Go9z6HFHSbN/gX
UPIza3thNy/on/5Scoe8QgXWkLERFd+D0j2Fc/ikpu82mkfjugJZ4vNHPdBbMVemggidDTnrtNKI
hGIYXaiR/Q+JjcaIia/zpZ3YXGTAvYmdyyK5ibZBh5mhjEA3dgBYRot5XrQuWlU8Z0150StWGt38
oev5/hGnJe3mgC4OK0N3Pi6c6UEvtMdMnsQGssGEZUApShTX0ye3dE1q/mxkFtFc5mjbQ1t6ckQD
OTwseL3koiMWTYvMF9omeN4/JYANr8ylsZPs7hJjPL3MO/lK1DEKc4ZV5aDOmySpzoCzbxmHatSq
CObhNjOcuWJ7Xyv5eOJqxs7K+7+W1ciOG4CTT+FS33NxRLNUdzaFtgTNmc8++BAFeiqaxJ+AqRSq
LbgB+x2q0h8wDun5nTEYWsMm5tZKlcifcclnZrEjIoTvnOzE62dsdw4NkeWF1SiNw9qaLL0aYO7A
0zWyNJ7aqtedLTSfnUjB0whL5Dyo58zd3XnNmrsw7nxK50mSQFhXLf379udpKhRFT2RtTt98yZco
Q0PlamFY8JIC/ffXsEQE/Xkglin2hyC7vW7JSpY0i9r6v5NAjklNJgo6C5EJFarvu8S8MmDCS6Pd
PCBgIXCqqy9ro8DiUYA2Wwpzxf797D++6dZxNJ+pbbIBX3aL/r416J+r+/xLU0vHzzGnAcpv3PwM
NKbhE2lKCfg3yzKa3hkVdOPQ3stEGb514I6YnGHR7zxMglJAJvI3fLwiEfcph9/TDC7T+dYw2UHE
tR0gh1WGJc24wPlqo6PRZFsvTgr8FrSPybEniSuk1A2a4nlUm3R2+DNxPSiK6Ell1BkqFCTLGgMu
dhL4ZQe3PdpQmHPbkLU9qtRgtQaQBqdLBoBAzgjW5ZzmLsecRt1LYt1cZgXpuXugstMtPZSHWEg4
0jToTvJCNVtdcsAaotu0tMNFFbiDoPYknfwwQCXrUbi96w6hd2Y3ZcJ8DoPe8+Vs9B6FIPlr+Y4G
kSe4D+ZYFszu8OIWrthT0Jnx2FNXX3UW+w4jjkC5HjwS72YNALx52/As8eOO2sltsd1ULNTcsmie
RH1GKl9RiZ+glMu4wX9+qjLYtoYaAFMeDE66qbZiyAwvdsynB8dOqMQu4CCctgEuXELo+nU0yUHR
XvxH/p1YtK/3mVqDbF9hkF5VqIRB6+t1tyHioUeBiIXWp5H1Voo7hBc7pbbKXMvPmuoeJ4CcxFnb
gNVDUUpcq15kkOZ8QQP4hsBTeumkX91jw504hgoMlo7D78DbUTFDo6vNF0XNDVA0gUihft4Otdvt
vybHcSVCHG4Yu98CEqC6bXNzptNGF7G8kLiopwJz/zQhWWGCm24+rg7ekWZIAVYge9XQF3VnhGPa
Sd2Dg8LtKqKEMqXWTnctQP+K3fSjfu13upi9YnmmCxDvR1QRxAjmaGYIhHMd0TkKZcCdB7cgl3Fe
T9tpQepNYruwBLhPZefJ86WlFh2I/PuBUIpRAtS+Ag78lahxdsbB4gUeh5jdtYBVix8NmH/CZHDx
SE3LYf4cwd1bHcGXJw2RQBbKQbYMVznR0+hmgSe9UJwthJkETxcgteq6nCq5cU0aiWVHqOBmwYhc
TX84UUhHosrGZSkhzi3jURJl4mr6xnOTEuIGwV/rGeYlZndxMYc8moknpRsP15Fsdou8XFDEthT2
wiYExp0XSmyEL1sHfneacHnVi/A7RmuBd46oioYOLEUzPRDHvkEEC1/pRwlnTufElha5imkybuXN
/crua3mdl28V1wClYBru5Mc+uULgu/15WZe4XiyG+w8EW/kV93eTH+uiZYPLJimSo3cshN9uJ+u6
kfsC47oIg2PMRk7e62y3KqJwgfF7dHOxc+P+CX4dOdXNVdskl9efaRKX9kcCYFKCxMFLhXfgNquz
6tBFDhk+/42cTeHQ9R6RQjPGJFoFQ+6mNINk8xkrSY1fFYjwkpJwYstWM/I/a8XMGLuE1a+jboa1
TQ0B3RenFSp30aQEJuJ0SV+h4ofgt2E6UZBji8z4zEg3tlwGMk2v+S7ootfCfNAzzirytb7IPHqR
TKumEAEpGf3gtqtLKvMN9QCOLp6glc4zkhZFgctpYy/otlIOFcHspdhLCFNfMqeI/EaENfjrNNFX
+AQHKGQEnxfJu+kA6g4cVkpe8BOLcbb1bCBUJx4fzOa01/9h+ugrfMPREesV/Xwws4GCAG0NmqaP
UmZIKqOEznh9w3gOaHIhu72fgn8iJiKROr6Ks2ZmyqeKuPFwoyaqQHnCxuObk+X3TIMwgfVfBWBP
M6xHRCpFOBi/6nsi/vP+IIi0tYMm7d/VPqGW0d+0/pkg6t5QNjAtjanTtCoLwLmJsPIAA1BX8XFo
7nSJ6nomkmraHOdc5sdXtC0Uxai9kZ6dNv13IM/SbyR4NyX5EuOgMf90dnPsHxhRgA/Pd2zlMbMP
95806GvcoONWoxWBgNyFq8GtCWLcl7qyMiq1BEc/nwpFh+X8AHW+CIx90XaZyknhQDah2Afph+hi
iG0YToT6ik7gV9R4GR0yS7r8uEalS7W3Fi6D0iTcX/1ZwdkbRYxw2T1bcoRPfuvt9e9VoxJOiakr
NPrEFOqfGACdxiupPuM+HK4jJVIpG8SqQSv5Nssb3XeZZ35ggU+wWJrHKnvls1EebharTOnnrwiC
LPdkrzHw8S5dICSlI2aBdG08xiFiGBbQ0rFYfbAa2EKzXBxxRQipplI/JqJBmDFbYLhsTH8fahnv
f0I+EDWIvs6ZZBMz7oQbA4VfIfp6Z5IzZvdePvRFOzJ3RE5oQJNpI39pIFPBBamMoJvY9l/2HPDe
gxjZiLCHzD832Nc2lcewiOXASOMSXMlwzeYkJofseSqSROLAL2zqxF+QmDRVqYrNOntfuN3HZSED
QsU9oe5d1of7elA02QPGF8wm3Z1ZwkHw5VDtJuPBKzLb5sx3jzfXnzLxMzY2Dxq7aAbXCjv8KLfU
UndO3Gy5CR3us7igsaIKRMJHQxQah4s0JBlSY+TZ+17X4v1TMFIstwFrUUjrgeugngNXHjEnk4vX
UWA6FlxzRHNCa4fkB9SEsZUdSTpTRP0NDsAgGeilacF4SHhTceiPrZLmYFhMI648Y/VKCsZm5W3T
fS195ujq0Vikz9hMuJqxLO3ZHalucd8cQapLf2KjXZDYMwlB+VrRwvljSQilOUJwsoddkuFhGtNI
1HAXsEHM0AjjFs713m5jycBE7dTLDfGZm5YDti7CA0or8FN4Fz6smmkqIbIoNK1CT9BIw/WR7l80
ofWFeVBVSiYRXpzyH+1S6CFg4kByXlARb65g63fjQ06exr0I0G34cBmQARTGUBukaHeskFEgGzp8
yqB8nLJl4JLZiOq9i+oo2Bk1Y26v2OlYedVc9UdJZoXOFKsX1YgV4ldn07aTLiZc47Y1BfbfIVUa
9/htmGJuOd3U2TShFRitwVUyYLzDe86dQTnVwn3ooLWn/mmLocuWUb3u4Zm8sNgm4L8E/zqKaTn4
a6rr02s4bOK5nD8pIrt03nYaPAND60v1DxLQEtgFULkgnjze2oQsodrGGhVN7kSsgNCWeAeaPHOW
C+0TM9cO+DfXGmHNIjZNaSIOv6Q/o2IO5hrxF6rxN3SOtvvJ5TMwJtAijRS/vLvYwHDQkDQah3sf
Ut3JPK42TxZX7xmB+8aF7CDoatzhUXFVyXLZi/KWC2ZDyw3K4xz92kszBPqm4cjEn3p5o/JLJJZV
LRSY3nTqtsbbRPLZnZfOwknRE41DOCiptZ21o2vp0aAQnThptVrZ/Nc364IKvpTP2jVqJXi5wO8T
BUQ3oVugSbPiaSCovUoi8gqGxM1p385D1KowieZUQxK9GH/GXEVmwIZJ8hUK2AdT5iac9d9lt57v
htRfUDVrCMervIYbWJM1mdGEfpIUxOF3Ya6WnTXpcsZkyvve4BUU2gf5FmjOdbFdvDsiIkCtFjeU
PMsB8i0nET9g/eG1jY8GsrplqHwkJWk43UsCO6iAthXZ2DR/3apiMKmj0B00gwMmNm6xN+iPpFml
gTPvqYnCOVtO66ZCCAuvbF/qEqPg028aOr1Ji+47pW0PqWdsroJhKjkM0AnFt7nk18Tufrz4Qkmx
jb1BJwjV/EliKPBrqpdUKHrLCB72wKUWdNGIM3wjd543/9fC2JKSiHl0i1UXcofGZNTbzWImJR1o
C0SPvnLhWPbKcRDoJqFEpGkeC5hy8JTF8UQo14Yq45sdB5mJ4GyGMQlsNxBdmsT3e9Af7IuAsuFn
+i74xtsAQ2i/Rs32R74Wsd00r0pUoAgXXerw+HDBfFuhD1vVFtac3D0keav4PNYrkpDQ7fq8qy1o
6x3W8m0P1At41+eeCvLpcae5TRUk6gTKkG5sdBzoCm50wcJtL2F61YIZW2NzewS1B9CngwPNUSJw
ca6LsVCqlzlCaK9maTSLl68nud1gaoizLosY+u3WzhLHVHWfR2en31aXVFhYrYg0+AwXFVQIhB3V
2G7Gtn0mMjQRLEyN2FZVMJQupKyVvXGPG4D8WwClctUzL+4PDB4v/OEx4/N+Aaxt51wJEoC9DmZO
J+GK8p2og7cGcg7aNHfazCi5IqkWMPQddEhzGsC4Y3vh8gdnK0FPY/3A2ZIRGXkz55knsfzaeo8V
hIwd0G+c3l3uAOJ7c87dxsbpj7NWHtVRcx8eVwkNWG+6lsV//hqVE/Nm+oTsWF4dMHu3reC+66r0
ai4F+1koA9Zfx5ACBdq0/qfOnNciF9oxHX9qvCdyVGUqZ8cXFor7Suu+mBYDSGsMnS6lmqXwNMiv
C1BNApbS75kRTS/36rPCPp5n9dywlQpK3dQGCC2WfG/aqiezuwZxfSqKLPwgnKHOActoOS3/cl39
o2/pXms8x0kFBz6NBaGoSvf2ZcOgET4o6FzBRd6q/NVSdi23BzvntKoTc27R781d3HMSggcZ5Dh8
dHyvRfIKc6mG0C7d7YeD/0VleDuDEZKW7f7FxgRDHGPafS596f1vitq5dWJjew1xRR9SEgtA8w+c
zP3Kd2YAOEdvMwss+D26WwfrvbO/zhM2ODUL4PrWEexjENgeLM2eVrMXatwvSi5ZPJ2ETbwD5j42
1qsdC6alUMR+Za7JILExl3q6jAbPaWs8P9H3C1h/bZ5Btnvqaga5ljAgXmloJE6s24X00KLYubEB
eIFkHQaHFKXQLOD/a/wOXg5MO7cc3WJMColzSzzvvPg6M8zhPkAhTZfuB0vi9EhkY3Aq7u2aUjau
F0C9gqJZrjSkILT2V/leLOKK4c4cb12NFEVwScyzFkjn3tiqmySlSAH2fTlNlL3CKo6Ff/wdX1SM
9uaqcrNFJf1cRLjxfAMzTPpjBaH9Wlb2MHowKaAkOJF5nI3ylWPqwPcLHfeG+A2OyGsJVngpxcxC
tj/Oe1RPtkNU2NAsOWZ+6zAH1II/x754+RYE/5f/tUnbqjOGLxwYwHbhYP0JDf7GjA7ddg+TBXQt
YKmjQlwM5ZyKjtkmHpRB8AZwBtiics/il/LB/u9lYuQCWn3FHRFTIDJPrP/bgSqwChSriQTXqHt8
ElCRMMXZtee6++rCmrhgIuj6uTGFrqSXEj77rskVXaQRGVhOEEn3UM11r8w1Iz1smz/AbuymxGOD
K5rkLtyGTScXRQtve54NscLsx67pEXJO3tzToRYt4VydvWj32WQGDx66lo/nW8s6GxHBHKXcyBfR
IofZ3JCjFLgFw6zjRuygF8VrIpMlu94T72R47T2lgnAr8rlWfWU7Dh2SA5Uh9e38Y3yEM+Gu/TJu
pKyn2njwJTpoPPfpEEwoV27kweH0aKVLiKefCBHCtuYZ4YA8CcT6meLEzfmJOqbRHb/AMRoz7O/l
fjXF0WqeJw+/EucFW+sQy8dG1+sjOT4NrqMV7O7QZQ9mXRT94dQSGmazsnZIgUyAVCBNYpN8wsV7
kpWDxOHCMBUp/zZcTWUpbPmZS/iE/nEoLBTiiTJK86OssCi4fXPaol7G8eEoaCc2pEuz0msXnqpk
+Hajl5doahbOSR+fWo5x8xYB5M2Y0iUnsbyiivPZj1M4V8Jm/O0tnuXUU/RJrNNd+7GAxLFcKhgs
8NZjAtQpgyAWp9L55dkLNIUJxTN9tKxAu2TpWF3YjOCdO8pBXT1Q1TdTvLb/qaeMuslNryiOjA2k
fcotI8ahsEnqDhCutY4kHj5tv1aquh0K3GNt3KN35M/6/ITHG8HBwdxROnKf1giWUC6p2y/dwuEd
kL4K9ihCp8Ui0N1dJ0gg4oskcziMPxx16/+7iv5ScG1Lznwyyf21leKMDDLGt8xB+K0mTxXn5GH7
IvV+/BsXAFL4qBuRVJgOtDRkhBrytaujC28zvPnqKP6c+znz/uHNQqua2hof1ZWHJ+bIAHzYT9IW
KYbOVBLEJ456t4wznYqfb6KIpSXLC1xB5vhdHl9YyFcx+6OgOBZcLPWVOY1FmAk9BgIPhVbU4i8u
DZ/VmrZis/Fllm3pvvi7h9WbWheAxmjc649RcNGV1Po2w2acM3yigEW5GyLuwFQdQdjzg8a5SZ2i
8plN6VmIV0pZGs5kp1w5pD/ia0+Vnpqer0lB5Sj1FjEl9LfsEiasj5MyAzM1yIxLOxypBSb/Hc8S
UcCc5+ogInKFSGFQwmLaC3Eq4VjoQsy4jQdpjAERBo3FkYwWpodnZnl2P850dZyBCDFNsRIt2Xo4
LO+sqhNx7PCyZMixM/AxwBEDN9HrM0Q8ots5C8Ff1FV3qqfTpr2epQDq6lsGgiWGpw6if0XziAHu
QLp3fImytjZmJm2MOrIozDbT+yYpTLNa3CnInn1/yxT9WO9Zwiv1gqCaCL+y2mmnnXIt1AkhzaaW
l3+y+NQpyi2/ctqpt/dFI+JHDezsaH92CwqpFSAYKIC70+/w6lga/s6HCCEGI+QtquKiUVurC9M5
nfnmHKzMpC1SxJ2x1ZVADWHAVRrW4kDnk9YWCkV9A4SaomA+HXzfyQIgqBznfUEB2Cpuer5sgaQN
1y3MAs+OuoHWKD6UEIXJIUpCgHqpRaB0xaAmIBpH040CbVAqzeY3QdgWOtKJiX3oMheY8USU7myJ
a6meYhdY+H3dThLZYX7WfnycYV3la2xmIyZb2WKCwBbj5vskyGLh2t7IoUTj7wuoNNPZkVdmvToC
NOgZmJGX5rO5DWC0gCIwvfWIEnBtPRHnIKr4iqs4hDcZpkBy1qFfmRyxS6SlPqxORyOcBAadFgdc
brunbbzAL2cIPTxIOVn00yLKDc3I16oC7BFfIvQmYjrzZ5+TqtlzjLKLmt3xcUN+R8XYWX47Skpb
uRc510Azv9yt3T+U93LL4vvJMhpdmr8rBrqbiXvWSW0b0XSHi4G2+0JIiplIt2gW+FojtibUvujZ
BB2rC87Ov9sjFu0NuYgwD5/5bnGEK3vOl64mrhjNoTiBfS6MM1wkLBqXNvujKV/iRhskZCTvmJuW
K4qQSFnwdt+nEMEEMqPDUo+U9SxbEYgTT3ziyxAW/vV7d4X5G9RRjA7ehYJZHXhN+tIu4tU+S/IV
muUgQEOb4Hv0YkBg+IyN7emafEVXfBBYwIZUJySAEweJvHld0j3tW4Y3aR9eGC77DmxIiZcutBHj
MYnAqb8EbYZ4tn2jk41kPXEgxvbYytEnqJIQ11NagI3v3qWOgUvDe+OrpoCq9dZu5wVreN3i284g
HHr9MzPgyHyGLZG+0Y93LbFXjg8bi20mks/rS2WwqKkT7BAsP28c70oX5b9mrzFcxQ/dVW8bW+wh
NJlrqHhLusgdUuqkzRyauguAChJz+jZaLZtS/mC/P6lSdMGpxqmAb1++c9vH8MZ6x6pjhksXxShM
EK215nGtRsFCOf6yMURKCtOOtu5ERiZQ9avlW9kpMCOhtMYH14JFODE1ldEdyyZAAheyhvonYFbF
G66E6JlzCAGOpm80N35i4FVcQgakt7TetlycjcpOUmzJSsL4WpRAYmZ6PCq6arSA91cxmm8/amE+
Sjjss9wrxmqMYWIJCRd5GHTCjOPlukjhf8ZPLKBEPuSiZeeCMkv598jUWM31ypmHwxzbrJhRk/D/
mVEKWruEOyGIvY1FjL3FJeliZLZqHDRx7AbouHvQi+ra/C1hkK9zqtXoLSAD3ZKvzoaTzpQtPNyc
se+nnDFq1M5HwG8gy1m1RhsrGvpB40WFaG7nY3NmNLRPRjuODaOZYlCJXcOKKbYcfLLOAwBVtTdT
J88FB0Jfg0GSV42/QeCCHi4fkX/DjBz9lhiKKwkq33GWknoJjMnVTYBWlxNU6JSTs3W9xqDLtRjD
qxd4E4j4YiplVbdxMXEwzzKWgmmagZgQDC++Hh0Awmcx0nq4Tp3g6wcOyH5Y3S9HA+8my3/+9RhA
lztVLbUWlD+yHO0WD6p0WWHtt5lmlldXHkxCnOlKvlRaPEbRNfi6qRjbytzN0PfkKfdZPZNDp1PQ
x+UxbKBChByDz5HkcRlpNRG37EwRttz9T7CBeyhIgsATOpnwxNkKfG9jaF76jBiuyZt9/ln0dkPd
AT2qxaif6fAcfEj3mg3YqCFOysJ8Y275PizEkUEhgx7Ry/Wl27JjHz6RNvurx5/WT/2R37SrbvZD
ho5blZTtn2CIQXI8RWWnm44Jd3uBY+CQZUsyDpakrwe9cxFFMjHoZrH2ZPASVECRWdkwPjSvNyPN
2amiEKhtrAGYc+S7nJSdy7xD1JO67WyJ3If8NXugnF0jpj9KkdhRIX/kTTCX9CobuFxyi0qBnn+1
PKNdSF/SopHj4RIYtc5D9Rmwj9OSejXOFCzt1OKDGP4reIjEn4V/K0KiHlWQ4VusN7E9hpCLte2+
Cf22TKciZ1svE05dmyks3mf1H978Yva46rnNE0QIa5msJ7JG2XdCQoWVniMWQpluuALxvZjPRFP+
4B+eMjQKk11Jzbpb80Hl+4QXIG5x26ulHZBt3zOsisfQVMCrekisdFE0fW7hAbF+LNEOgN/IC8R8
WuLxMMEhUfRietqlZxwIlPEdwpD+0xqDJNqNHwkJj12xLJ73G9RLfH4R88Lx7whdimw56vTkwaSX
7DBUBLY63NS38eKzAWg0/tUPBBiqeWX/A/F7eLtdfJzrGqtH29BKU84jqqCC6LnaIlJiX5/kKkYe
31uRO+lVd4I+sqUT3koHKXGxlwQqHbLv6BJMBUOW+U026ZzNgw7x+tMXdAzsjrqF2G2shTsFMjYT
2Zoy9h6O1E5+7XRM9igHkU/OEiBLN4x5Buo+FMts28HmAyC7jM7jWpswGzZBLnGRyd3TYEIx3qoq
6SDzB3bSy23UKwbl7DQspeA196lemnBNKsUCjwALT3K9zQTg73s5AIQnKumUL+0amhewgC7chrRE
dQNWVTs/UBXlnJ3LVLAv2ZiQXutAD4zm47kRBAyRhbnmIdIoTcwVWVPw3gZgSLJz+FgLD7NyYwNe
KiB/hCUtdkiqQMU06TM8Vr4d3oHMAf3okk5BdVPnfHi1tCvrEh58bghs8BVdkZ28F5JP6j9CL4ZC
FdHb16hpG1TcD4RN156D2dfU7R5CtN1ZA0yzFehFqcmbUq1g2YCSKr6tH1TFXah86fHLiaF/60Rs
z+ssE9HiT4O6zREA7DJk/qZ8WlTgHwNS5lmN0+Q9fUzAruXlYInfaGV6+ZleA4xGN75WIh5eiZke
rZ6oQ1DxiNL9TiT/735rylgB6jwBmeDfjKV6zHRlbt1/7PYTBSO/d1yU4dp2VzMndH0+sDrr4STE
iQnEIhxkaoXITqUmQvBNhH7s3lDq6slRupY1nGblpa+kMQv+qpDkoqfmfhb2qJ0Xs8r7/4DWNhIE
Z31JErLCbxxi6gucw1Ubfmlk8Esf2koQakLIX7JsYYAxUmd330oGoc7OpEjHZx2Csco2dUyn4XRS
cgENFgrVPZej5pu4XFlv5EFOiOTwKixaVlRdd1kGtD59xFrruuabIha2HYyCC7iuvk/WZKkz0ryg
90GU69EzKbGzoLg9jc8iwkxUuJbvU4s69ADPoIBwbpLeP2+MIAGNRNBAIYfkLMw2lldURhQ0FBfW
UG2A2rZwPPz+7Pv+gKBOVSPPkCdcdyW0WEXIDLKiZsVx3okThlraWizM1Yhn8j7kSjf16rOveKnf
tcl5gyLcXw6/2W3BleZW+ijx6DkmECh+8sUGoB4wCOtAZ5O7+sApImb8iWB4OaxAEq0xW7UW7/Qn
pk+QolK5YjHY3tskkwhRUczo6Dy5EYenmZM2zTzjNmHNlrv75S6DLZix1KnWOXL4+Je3dYfArvtl
A6QISTv+dehbX1AGg4LBFlU2OX7DxiSgAlOi6gn5+RQODL6bN9fwfsESXldJSC/id9cnx21+Rm/g
eATIiA5h+fyc1jijMzmE6I3nQk/Bum/cSQOSzD70IJPdFCf7Cwfpv5EjkKZ4nSr0AYJyJdxyDeEi
7gLP6+F82GPpQWNx7Ure2viPvQ8TcJI1Q02pfEotogPOkAWcLgp2vaiCH4nlX1xzD4wACuF9aow2
5GxbtuPTmSU5Dcz4YcpKaLBzA1tj/Z7InSg5WgGYzdfwp6xKGbzQmD97ftR34lZHdQ9OtGCr5g6q
IcVLctvPlUk6McidfjoYF2dHnp28bSaZwfIpqqbxWRLzKfJjiQOXNx4Kz9JLsuM2VEZz+e4c+p9V
sdTfi9allfffFcYRZrAZkrCYAjkkp/aLzXb+3YpzhxeTS03BArt7BWLi/5foOHpz/wQw9ku2Y3X5
XxeANlf30tAmLjM6zQSNL9sfYPc0qgDoZuxla+97niXFupsAAH4z6f5xMJb81z5fq81ddpZDCmvb
zPUqgW8k5HakOgt8P2Y5QpZJ17mYZ4nFAPlIwin8MeiqFqrzNsSxMczYChvrkt8H6d4M8jdnQ/7D
t0ubMnMyJzRGvz3iErqEOsRJO5FzVMl8EgAto729z4uQFq5DV5HkoaT517bNi0awHccy+z4eRVEE
/czLZWtPPWaeMQ6uiHelvNlpqohXBzzKvFxn7UEp3DZuKEZ3InceoNoYtBA4z1ieGfrt+7CVu3YF
nVyI0DzND+1Dko/5KPfFLj2aLZahSj1yaVugWYiCZGubD8JUZtNJOhTlJwNDN9LxL9nwoDZyOwYg
k3egOR0DQdqwkz4ilvdiG8aCUXbErqdDi5qQlVfKv7j7fOyG3SLOQR/EV+hgJqJJA+YS+Vs/Sg0f
VhScynVQzrSXoND9BTXJycCr2UaCxXUeHYEXiKx2K6wgqpQBzV1zXyx8ZfqhJk7h13+4bDnzbBsR
6E8jrAwfcF1+lX3zGUtcJMzbzn5HrKcjsj5WRhC6UP7PW+PC2zyf3uxqrmehcfzomoWexAvyEZGi
PWRLQwf0iWFUVUcUfH3Yn9pqPw7d/rFev2dca8apKEyKMNwwLplEeJ9Jc1SusO1d6U0LmL1ICCIG
phm11ynfyUKnRlX9BQPLt8S5jVVPO/efR8yX+BY0gsiPH7iiPEnKR1nt8cMpLds/HGBCDrtz55jP
uWXwwZA4LZXL8omqS23wH1fzhK5WjP+BZtfjYUtr/C5Bm7AicQoJxht1uEu5XgS+faPA/IRMqq0i
R93qnY88260hl74tCr3l0Xvq/EPKLywQsmYWYaw8em2RgHiCyOKim3xcNli4IvoRMrlcEiAKj0+l
sgisZJBjTQCLtDsQb2dOs+T0yASaILIafJz0+cr4E0PpP0nK+1MJDNWW9bFVg9CsPzJvK4RXoUmC
fgDsYCjVlM52eBQ/Tzqm4pYv6lYyBW7TGij4czt0I8RgU+kD4mxX7hvgwX+29f/ZQ7e7vgFVDAre
Ho90W68zHUGD0qSD+vZ2MQHD+CjdGgv9HGAJ9fla6UC/r7wzy5j1DVcWUN3JWjB6S1UEeNFa0Rgu
ofo31AJXq507I1xNX/rew6rWBXhfy1rSFMcgUBfk6q/bwDcc7J/ahpub4bFYZb5yY2iYgG4SCpeg
Gf+jAcrQ4yJ3fz64F/Y0Yf+WDTKiUs7Fpi9VTzAaZdpCDy4mQXEfn1yNLP5QdyNpCuCyiAJVCXmQ
Y9T13meI0HnHF35CScBHoNqajwqDhJRVhCp+QyiNDsV2AnGUGMw+Nd15+orfg6obpmMVwYpL4Tom
iojLhvY5Ar++uGdEZhFh2HfQHw202DCK0NWPXgj9KZn2g18mnKu1Fgu6wzFxds8gPllb1ragpNlq
M+quYcSENg+OTGhkpBnxJZosjHuFanjkuGT6WYYuOzyzGQ2Y0bPcMLsDCDUV8X2gExINS4lsWo1W
DIOiIUy74YtwGSy3Bel7FStjtI9IOa8M6tyEqreGrMO0nLM58OoliExxPj3xbWrtgNHER4kN4Wvi
WeE8CzwvE+lv0wSxuLIQzxSr9FIQg8Ysja7l8/2D/SeE9NCz7S3NE5/OXcO+/az6rdvqlqkn/xzN
aYoB+i+i6PWrMkVj0z6RjPdPephnd6h7kyPvsyAE2mlvudTknc5NQ6c6tKdOWL1Epogv1VirWYJF
s0xSO646smLXhPnIn0FEJ1vKMjlFXPD8PfOCYPM1zVwSBU0Fgft0UWC/YfN36bfF+hIUm60UZ8vl
ICnpsHFrYkAhA2zkqppZUqyscgeZ2Nsh1gqj1ulB24UyiUFgbXbXNk7jkKGeJAu3JfKH/wgzVh/x
idIg0v+fJPnL6LzQ9ybo0z8dhPB8YgUW+W0KWy9c52FQakhClpFXXbT9qtSUxJ262a+mib4OnKxI
obuVmj92pUQJttmEBLP5i/9sBFt1ku6Cur26EPSJVqIgfTdcLcrEyI78dpx9fKeaAlPMmWPoEO5E
r4yaXCnk9A6HY9n8PKVNZxLxsJ2/lwktGvMnxcyai9MmSoXcAorNN7RUkPA7qMoNr0I1Yji/p49u
CZiTquTgu7U+cKW0qHy6hLORvLlyfHNTKVpaj7gZkP1WTZu7/BTl2OlnWNdJkkJeghRSWw+rIdts
4vvVbCS2rKWxzibihhkfSy3+NgeuVW0oTIbvENy1I7zi9iq9Z9K4t4rCfdIpOh2jNIoIvNfJ1Qsv
u65XAv2fIr15H3AV5YdofOuSXPN4UxFPSyWCXp3UKWHBMogLPdPf299tDfUi2C4KCipbsZ9sLxBp
hWD6aoDEDlu9XHV9Jx9eeIN4kAJsGwkLPwbSqXRgyU8QLq69Rjq+K9DcIx7o0OeCVXBNtAW16mFh
4lh+RjULvIcvooxGl42MHukBmLzEI/2TnoNcIvqm8JWPbPnMGtkjukUMm5c7XaKQdgY8VFCe3NQz
pLWlbUj+9hpjO++9aM5X3UpVDAyh/LT2tZM5hMQ9rwO7iBdg0mawgB64iZ4ZzewKh0d1cKIzWhgN
ixENv2Yu6JvYpfLFrbh0dnB/YaGFrVdlwlAqNoTxN0qwlD7api4FyQjjy2cgvfwV2Lp9DH1Tormc
aMxyQHq5bzNmKZtNvCvQN5Re41KEt0zyj5JE6xF2j3zNrOA9umiZKZLKNDwTChrceSVXBgunU+cM
X4UGfO7TcNxx1bHBhsxng64DacJjOlzAU7/IK1bUBN+ziBi3hugzD76sAxPePGQQ+KhowPVpoDOe
86Wr+RtuhURGfRmylcbCal1pRdyG502aSoCl1U5OBxwxib86FFn1RBKjCrR5TC5sGpTNM5I+nf8c
VXMHJvwQ1oxhmTPz/de8fmj/oyM5lEJm3qXmYPG24OcP1z1+5kR4S2CshDcVid2XMD1OJWF/KbHA
lGhSVEpuRFcwu8Ve8el+Ke/cMD39MuBe6hXLi01igoGsMZGuhXZtldMX7kfrBSVirwNc8jcQKsDQ
2funrJ0qOsz3iCpIzkR5pNmGZNZfkaHWP7l5mvJ1lFAZXKxfGBD4RyTdcXfJlw5cqUHmTUvHlhFD
jEVzUeUpbSDwU5ms1+eUsTHr6Uq0YOZnJ1sbZY8VgX34Xf9jgHM0lbsJV+vwkq5jHL6vF2oAuGkD
paZfpkIMKt/sqQudBdtguY3q8JrkqSBcWilSiXH+n/N3mK3xfEQkRkcUgZfribFk3qly7inwqGOZ
4XBwQSKoqqtqUIOTn1vEHY74qZ1SEmMYVG7rlW29zB6K1KnQhNeINvqMUrc3fGnRQe+ULDiAPoMF
2+u2aLx3eIoQvSr4x8kgu6SWoFPOhxu+nswi+gsTIS7OtBzsEW+IK735VCHO5H18ZqmkGa3HmbhA
ILrFPFSD5y71qx0kP+gJ8zz3vZSNvVspy8LbDPHhFnAoZmKg32U9C4FLEZiZA65nG2wL45bM4yrs
ZGZzNkU19vOkeZjlf1A4X+nJTUSlcNrMOcim2O+ASZMjWlmpexIYRrVPe5xW/FmEzH9LUug3KZsK
NUac65ldEN/T5kkDadLEj5IJAu2ho1+7hw/UEYPeip3TLNdRBPtAKYN11ePEdO3/pva15jzZuSXS
7syar6N9hB+9yxtqTipL2CtwdOWJ8q0X51D6J92QAMtA5yQFBmdCqAKDWzuugW6zVuUGLfraG4dZ
EU/1W8QyidIr5ogMlzSGNQpz9JXp/ImCapzkoRN3Yv29XhHlaJywycK5VHxWe8/r4Mhouxq/nALV
3Rx5ZWLAqx6VjgVbDbph/IZOZvZ8/D38bCJx+ATK6njX5fU+l7nFzRgcTnfj5zpDbeAlrhHzdD7I
ea1H+pwM8J93kQ/KCS1OjudZ2p6eUStHLeAoR6G9cMuedvn89qKo2EbooFV/JPDA20exEOcgUlGc
0bE6ea0ub1eTvqAFIT0ukFdWx6F4GjC5+jMBCHJ6zPcW1nrQPaCXdorMcNyp2c4lTkceR9rJWZbo
xWf99RPZ+qWmAp9rukKGaA9OyKN5snSVdIjq2xJ8pXLVhIqjeUZYZW+B8iyeUQ2lKRJwoaR4Czmf
sxiXbWDJ5P5VFGl1lBETQ04hhNm5vwlRfNjps5ch0QcyLnU11V8Akqu2BQb8N7TIYb2wf1X1Hz8Z
K0XYs/jOJwuAefMprOSXqAEEjfj1BI6okJAr3Vmj3FzLuMLyNgSQGI7BfJN3RqUaP/LnsNRvAo+j
QqZrQqnZ+2He+aoDtD9vbCSxIdzZ6kYBI17GBJw22wg8K39y0vws/uJ9UIfDWVguhKcAPtCPOIub
5PFdShouMaqRGOeSsJ3U8WFEKxsfIl9YBikxRzaquDMWrSo3vJUVbZaNRd5MSsvtMbOl3AipGCeA
3gAit9UKs+5BgGTmQRHP44vQsfiBXhDlzweica/HcbB/Pf/cVqeAgiDkODPSPK1lYRKXo714W+q/
iXLCH44Svnof40NJvjBOnFupifaktjvB0azoO9u47q0NGyoNvtSm3AmoQw7WYFPiEQFzpe4/OTZW
MDxoC73iQAKoyHlQr8cqDIA40p3r3gnpmBLli6cA0CxoyL+zK7wmM43oWBi0TLhClvti7f7o4PId
GPxpVFyW/VMxG3S4YyqUPPMGONn7MrUvJC1hTVGCPlNQ0kcLD4CVpyRtV9yXSgOcW7qbMcKud18a
5xTdkddLHoVxQV2NklYB143edV5U+27vLsXdcy7FPfG44eg9itQJrlGJif0GY3rX4SQQ2BqSK5zD
rNkPYTm1+zfEJBY+jCx4ve4MAtsUxawl2r1avx0fkBnxha/AYxKHA2De9pLvkbPnUAbzSqd0ZJ5o
3qZiYeuzIsFN3bQtVH69rE4AP/nMMaPZizo9FFU9SRmtNGEtYn8MktvCCxt8zFQo97HhPGEQ7CFt
hUl+e8basqDAYAxl49nv4CsuuaAr0hv3hjAz9A91W16+Hwd/WhxfxPzcneNPlbzMWYRRpaoAuvOd
ikCIuGfm5cXm5Tb5Far85F0mIIF4xfuPN5JenqUgO/WIlJWsjPZS9D/MVZYUqiyeNBLx0JT6FaOF
iudWYMyanwvZxwfiQqkQVj1C3KxUFMzzbAEZ96hxaa0jq2lOE2w8kmn8l0+uTw1+NMeJaoaZCZ9z
6CEHrScgi4Wi1S8ZxQYGAZQ4T9xUxXfLZaegsd3EyjTTpNYER1PjG/sFHWNXgL6NZViBi+ZzxanR
ZDvkJYSz1LDhb1EnZqjyMvL3smV1QPfzQXeIUtgoL8IqQ9e7igf2KLrp06qW2IR0sIxJqLszsHqA
smW/2+OIj8/pudSuQGaI3AeUsGs/BH0XFfJh0E93NtPF0POvsTqblzV/bEWyIGU8Xzu1ZqcSLfsC
JZnkAavG7hb552fKFiaospPwUygcleUUClTIssyfyC0nVnyxIc5k/C8jqov8gW6BoJEyDr7w61fN
LF1Q1et3pUy1ef1QiTj+gDZj7TJ8mYZRoiG1WcPDZtPRpEf8hsmEjar5WVnU3Jm9jWfCjF7fnd+J
0mKbxkFiIr2e29eXTtaXNDFK245HKFhHL5a0H3fL4TQ/WP7x5DMInzja/WH+UCHQscCIhKzNDBtM
9EwFISjUX/lK1vXOAGSytxIL2LF/G6BkoFyJ1HOFPJumnPs4vXh1BTdO1CBmzx+Oh+jAz8ib4yYX
c5hQs6ZJdhTLcqH99A7bHhbSIKCBoNEdRc+d0JsbeQMJ9oOkh+OMLvLxOVcaBdKd+SdhXfhHOyC6
0wFabaYAZZ1Zq08KiXbF04nWD4OGcFo//PW4WkU7EuzrShfACfnCvI2B7bbayO9qmKFuHC1q4R7p
m/I7UhYcrNdU9K5SUOkF0gsHWeHF+A7HcaNeyMa9/lAROzl4ULNs2D7UFwEpoxDc0oBGvJ1xK/Ig
wSpJ1EJfE+d4uK0VE5E2ZGPQCVfsVEgnXmJgIfUooYIZ8sqYm8dul2CZuMaBjgBW1U8IdIxs+sBp
3HlQpJEWfxa7t10YXEP5ddoYf+tpIQgo82g2t2pdhDQihHG3fMCjTie9OIppbBUTBfF/8JBWf3TC
VALjTdwNLmbd05N3DJwRJavpwNRWBuKqZtOrzfFJ6agaHLE6N6+x5XiloA97ryahUjxvATFNSboH
THH9l47XMGKrtxlpvm/cCrQLt2ErnR7ECryw2V57PxQmzPLoyveksTL9PmjYyiTsLmpBp06csNBq
TdwyvUhRW7zCAOSPwk+lrXfNb+TRtc+kxSglMlVWsS3hf22LqZSosFSclss1xVzZSy8PI8WwxK2A
HNjD7A+O77Fh8is0i0WlJOcR2dzpsWiZnMeu+v49UMpZO9rly6+Fr1lr/ZuZ36z1CDdYWa2eKMiO
vwdHLDv8AbGFvOtf0ej+G/R+3B5m7YxuUVZhHt/DPUa270TeVzIofS2I6uGRAc1QSD1JSCJUx8xM
BUzpDM7Bg9TbkfMbbXw4VHSgxTZOfJ/Z3kPXXi6ABmpDn6MlhRyNb7Oq28/yHjIz9KvD4jF+Nwis
7UtoTUejb/JPv3TV5yorCTT7mA99641kJ3dOZK0Uqh7n9Xda6QSre4tahsyB7nbn9rZiJzXMHuNv
MynqockDSJke33JHFjPYispMxiKfLFIPDPbxiFBKVlIt6Wkn8fVpVR4veGJKZAUPuirvaPUJYwTm
vbLVvTM7FYuTE21YAy+6+XxOJZ8UW2+fXQy4xgFgzXJXqUKtqjsayfKslYP8zl7hF8m0MoGuwhMG
1V8Z8acwlFWQcMO4qqw4fXq6bglje6JMwaLUQVmF/vjLAJNW8Yx/g4yJ7vKA6ZIncv0ihKcTLRC5
7O9RTnu2DvJ0kCY66LyLmNZ2sMgL63plCsbcHcKJBosFcz4OO5EhB+LX5dBnCuRuAWl42GmsK3t4
q9xnlxihoUsfbk8c0rdUGz5ulaotJ66ia/LrjkbqT8Y4PfwhPLGh1k7TIKnGZpbhXglYQKJEIrXd
XRGOZlnT5zpqUDnQzpiJPEAfTLQ3rM1M9aehrnNoAn3ooDCl0l8+LivdfzBnDTVhSWw28OMPJ5Qk
mOWTRVIllQzWPhjtx+JTy69acL8/jiRkW2RBIbXuODHVtIVxBl7+CczcWNVIlfLYpaK0iWXI/7NW
KBdS7HRcQUJeJnnRi8a7NTVeiiLvpOg/epJB8Djhrm49fkyiqhs6R+dxaISTX8VdVY/4LgpYWkEe
PE5be6Wp3neutadycOXC4BtHmOYUGwb7wG6lYhcXykrOH0Z/cZMTK7iIm53G7jq62iCGr0H9arSt
jdRX+440z9Fl3p6iNLydOts1ECWmryCgwnyEJjxnhDqhi3KbErCdmFHWQnLMbo9e5CKOE/K7dlsZ
9JFVfsoOQXq8szCTHh1SYiaCznXhbm8O/KF/NvdhB6c7+iMREiKXzmOKhrTlqmxVty04PhumXNBR
312GSe6H5PD7GJ8ZPOr4BCFDxr+QRCtY6OXwJApDHSrA+s1M93Iv7Q2ktCxz10DMQkjDRqgRPG0K
Whl3pQPkA2iLYwxLWp4Y/pgMzLigO2yHlnf3Q88T+4VH0YVVmUBhnPxHqfqGOIb9mCxLhsmCM1Ez
iFREQgxExR+pjk6KpzSaw22S3bTez6OXGqZ0ELogxdFys53wEBziueeRWBy472MhCcqbzHPlnrBR
ubOneVwfRk8TYaJDJWTjMVmzvMC7Gu7/ehrDEyYqcyeFefpciq/BOsPKZUw0OghZIMKww9ClXBEU
fDoAjt2ZWBRXd4MFSaMvcekMkvYA7yZXuaDSf30/+bnLigD5p7lUU4ZhTuI+ovPHn6nrnlYpCMmv
2W8fdMvecyAJbvT9zot5HmHxW2bFMYweGpz2xlSFowcgKcVKDU5YRz74+nFgdH0sY2uZbxZLNLvy
S9OSJgdjRpcwMMAd+2miJBY8IRMQH5mvPkBSEhQpgG8eEi4ka0vGE3trxE9ENB7ZIAJEI5v2+41N
7LKK5cs5C8VR1K3/BNG0a/4MC8M9GRV4TxRfn+TMeA4VlKCU1TOfCIkrDZAQnK3wIJYwJr3SCBol
d4HXM9jm2flyHjt9EPPntdUC4R4676GbHJLqCGKATqZB8gPt9o+bYt8C1BmZY0Jc9FbL33hlEs1l
omy/hKABFNKPblMQRJCD2/K69Mx7katgR0Q8SX0IJ5fANHLT+shtViVzwq8cu0EOo9LAyMd2fqOG
nOehING0mC6Q7b1kENkDQOgbENjRRo2xdb9pfYHSz1a+tjTi5VqllHWi4owL6VOwNfu9EwhdXtn+
5KOi+ZC16YC8PRQVSlBiwJrx2D3bNciD1DoIN7q/ZRGDnIFwE2LZ6U7qM2t+WC0gYR7Ym4q97qL8
nQ7sa2qpMzrMDr+cBRPijsOpIl8A7MARogVqQi8r+qdNXQ6nmOjb1MaENw79ttCAI52nKfdtbomI
biSnuYNZ4H51m8z9PGPWJCnpxGawna3/oqIgD2fQe7jEiblmX/1wptXO/0XE7ebUze4XSj9cgZyP
O3kLnC//ZyABNrl/HK1En4DBY65qj01leOu6aiCHSJbOdti/7bdMQPAmN1FlX2uuOBUrKf5rfTcn
Xfbtz0JLiI+/5PSxRleuTfdQ79fT3XNx4nZkiSQUs/wiQiFW5QAlYbwU4bjS1pwkIhOjReLFKHbZ
Q/8t/dDG0aHXNqG8telQcoDX0B8o1aHYwXu97broGoyjb+M8CZIn6ZHRAyIskp/OLuMwEVvpUxrE
c0uPXMWg8sY98djJuWvz7POzAV1VMzOmJqKj3OLcYl7qUysN3qIgGCr8YX7GfNnkOGCom61rKzkj
1qGdQl8U2B9WIOaE0Q8kQImLk4X9huDiW8qipeh+cxsH5eKxiHTinG8Fl1oZzT2dPDTD9ZzNu8Wj
5EAaQ4aEV8Bw+rWa6rcHpfsvwu69WfkHaEngE7sAjeIwk177foTVbEUXHdctxxiMbazCv9vuD2MA
v0nZ+RbKiimjMemxklnF/gNwvXWB949OmzYH9LeKtHiNa/hGSgUOUfd91fOo/gMUFI9z6OT/1qGl
5R+EPBDEHnBlRPIduPlUjht/FR5+xrY4w7gI9c8whsuwnJBIUwMrTRANgiow/HB5okxR9u5+2B4Q
qR1Jsk7uV7Tk9zTAHUh/spjzDbXLvbvMaa7CVKD3WJuyYR0bjWbUR5Z7BDYcf02AMYo2BRct5SgH
nwcucmRgqg1C25xvJaqC17jJC8uD2ZxnCN1i0nVt/tvYp3W2Kv5F/bg1xv60U3sH1lU6D/9TBeP4
b1mk/0PGjQQY562AwYGvKd5qzG6ak1xQD5Up5tpLcahdme7AS1FGzQgim9p52ooPqxaQc19awFs7
kuOqbVlgn+OyCG5uIs4ilQiQ+vf9kkJuBC2ZfYYSNBrTjnGBi3Mg/JIg/iQBQKEJyMaGnRan+vbR
OVtHRMOniXYv7+8NRoDg8G7m61ZLztvHKu7L/WAP50tVp5TIHa4c1zbEm6BOy7fMv8DMxFo/Bsk5
mACTUqvSa6za4ERg9VGjZkzGkYG5lL77FCsCeybLidv3HXcsaYVrQEPohvvZDxu8fe5i7TYh/Yq2
xAr3bK9qocEiSItksLGMOlLBoq3l9aSaRXZm5kdkXd40F6SfCxMN3Jrz4CLgPVefBZy5QhRfQA5I
PxaLAvdwVXck/ALov1vGkwDxMcL+/NNLzRrUbWUbk7Jq4XGLxQhxblPGKMCHIFMrbmeU9i99HZNx
ozbW0NPnruOKOQP4q9Uikxd9DMbFMGiuWFBPleWgYFsI8YxLhbp7QuaDu5QA2o9P2FByjgz2Iq/Z
YHbM+cvmaa1QGeDQ+7i4EHf2MdGyByXpAmsJYPWKBcWkAI5A0m8WZy4lhTy9qd5iWG/De7nk8vjT
F/fD/Fm8SkXm2pxxR5VBjOYGhQriHGdN5D9AIp3W29fbxgRQp2+R+6PL2tRcefFFUHodVW4U8dD6
QG5vFvD2tbJpVX2reZ4NYU/RzXSphM2SVzcEyQW01AuagNwT4q8bTD8YT/voOGLdkayTT0zwhpu9
+yquyJKZ58S82A1s8Tcp5LXIT80JTeyeR8JJHUlbVtaX3r+rrg+Jdn/1Sh09SteUyXgkCwXiKCXp
RQjzMTDD7I1NS/8OBImSldIX6xhL2jek7EAc9l5mK/Aq3r33N0ULy24cQlgEzCrrUawAkznOhqtm
3qmu3ONxNpWMTJGDBj62PNmAUvO8a//kmkL8Iahfe57YUsx/2bOc/W6Lp75QREfGJ6jEt91pgxu2
hmlRZNBP6FwdH/jd6UjIafU8yMa+dnGcTLio3eGJnbCPsxVaPKwbt2rY99TiqdBwFYdzkVMrmfZc
v2Dy4aGPxcAdmFaRz9kmU2nmyb/gNDWjufJXQykO/4ca8qxy6EHgfqFUOpfeTIo7zjRkLdECgkHE
rI8njocqnnrIsFMNaom1nkeB2lGmHZUhgbyXd76A3bHCDwcMk+kq83E6n0is+EcjGcQ/6MQTWTYL
E3l40qZIyMRAKeeGMQO5tTNv7/yAhC2CEDgLr0xkyS8tp+HNiLKKs/6sVfwef5ZLIeVwxFYp6S0y
WODCgkAJNOZbis6rF9nSHeirT4dVKIqJhOmidFmdx/I0tHY2C6PyMAg+6/enLdgnJmfS9gyhRq/h
0eu6nBUVfIcjNdtgIayXdsK9BA2rwtl3VwJak/dM7xOfEYJoVVxN19ckuKDLrfVwC22c/DD0YETl
Qxf2Ca/ywtQUW5xCah3CBwsePguS6VT5SHH7zjbPVxu3ZYBW154PwcwyAD31ALJPcYg5q6R9nksL
HsVXC2PO8uTyHEJ3H5OXGgp3RCSsZQMnFJvQuCj2UQPyODBIbX8DkF6ny6nX6sOaUynMYCXxKaF5
hSGL5x+rDDt0cWosejbPVJxnFbkECnlm9tnB8zQQkKlTtMT8Xgpv68kr4rEY4cX+sV88EtRjblia
7R5xQMYsQrBSXvek7UIml2ndgjOaaj8Pwp0TTRYZFcjUFGJw5hSoLUBZS2hy0S3BXBCCHAW5o33b
9u6oSvNay4rNAQ46qBA0OT+KJjM6VRYYKT+pYfJTl2jJ2Sf1YzZaOqmUe6lg+xihrQS+GS76Xqtt
90gBMH7uyIuXG4SfSGD0LiUizCSW7TqnvXf00GK7vHguKHlMg9YKJSNTxMkLvUrszUu2b1RAZX3E
2P1pFC124dwIgd8stfb9UrgseZx+xxEvCRIy8BtpKefLR9hfz16I3YwErTwmtzoJSp0zWePYhPIS
QNwBp6VHNcyUdiJrYRvJGhNcBNKVJYjuJSfFP4pJRFAnW0xMXNnojb1rK3vGpa22oPeTyzqYkCOn
eiDcYppCe90Apw8DM6oww4Tr8wUgTagBfF7jz0H+LEMzYg/PtamXFyN4q/ycVlBP3fPmc3jQNMoK
5YO3rH+938kRuikoJp85ujm2/uxO5ypfTDN++bGGApQCyxzl4RT/hJx08c8FFlKflUiaygKkOzXQ
atwRX2yjxCVtX5uvIT5yATo2CgjGKZq++J0h4z1ZMBxqwFGZbCaEx6f79hGvblmEGykIxfan9Opq
PfhOmmI5nPCLRRvtFW/J/ZBk9qlQqdnQ1sTIyz44OpstVrOPVU7S/viWEC874ZmEfnAFG1ksxQ0l
Mk1NL0QUIYxmr6Y/RdPuemoSgiTMkJT1uBatEM6toWTGOIc+ZYOsal5nxIbazoo3Zk6t/URUvsuJ
Kq6Yw5L6DLG8VYMUiroDrknjwcLM2ErKT9GltuN/x2c5MbpAvzsdMDhblbIPyiaw9XQ9y+9WbfZ9
PE9gaWk9eOxEMxGgBoLj6KKynLU6nehfIjpfQMKVtoo20D6W3IOiZl6dHnYCbhFhVzXYqFrprL7k
ubRXn62O6PrygadrFo0KV8bj+zAzqqZaFJyPXjilP5PyThCUR49Sb520Mf7fuOjc4kAFyrUwDT4B
S1EH7EjvIUP4HVzkK/s0aVaKvM2GWDfZVlk8L24MeTe7gDwtofYVOA00pZFAKs2hwpDhkJta9W+c
BUam83LRaY8SRqMwyaetgBPTxGn3fkRnL3ab33uMgvXznl7sCbqlcPGrBcSL86JQbBG0V6dsP1QI
jV6pPCoAU1+I+2FW1VLm8WawzR9SNoDAdO+2CcSRWbHA9EL0hyEP9nJS1qEr9pV84fJXMqIxkpBG
z/p5HlgKC2beiB0pOAocuNg08gIbgwkayf+RQKjq92u7Lh+cqV6tbcqE9IdhbrjgP1DM43Mbqe77
W+u0Yj9FSKgOH+HZxkeTfWp4/FBpPwaUOQRDIM8Dz3Rtj+VxpBt4YXNVSD7KZIu4Jdz1yIiPdB+D
mg/6at1bQDnFRnTM2NOJpJXG9PdBwDhLzp2XgfhppuFT7HHjSkb3xRnJNprQT0wcrlY/hyDViWrh
Yby2tpjXnWPIV/FcmCxI4rlyBOf3n7YJtPGrDIrO2Zn7W2N/kfrGQ4iONNG+We7d6/V4+5q8Nylm
nClwBsBcwZ3TIu10Cu4tzEfVNis9RScHnCYDwvImonyrYZZaGvjd92pcnWVXQWDCGNfCP/TROK8F
NTH725I0HQ6KU/waSn4BZGc3u45C/I6gICmLJHSyMmOg8bfpMCNlPfWJGw2yITqfhSBMaoCmZdVD
cGptV+7O5j3/RrnNjN+x/51mNKZwfnJEC/lfN4/K8SbJDCjSppZpOES+tTBb4y7mDU8yQmn6G0FO
XaG3YWsof3lDQhmJm4LfiIS3valv/IPipP9fxmCiqpyr3fQK03Sfe6yk+yIv/wcClm/jDF6FdKMB
5V31zS7usrEMZPSqS2YilAYIntCdqBjLuewcsrFzn4SBTfmQiTZ2Fk0PKAEQIi6zC3RmGR+axyCH
RG9ryFHl+6UevAxeGWoIUia9mTaimgttmApVIs7i7BTf9l8qb5yOPZDySehufFajPe1pfqHZwBj8
p1M5Jv92s9fGhVfqrXKUF5VzkcJW0j3rg7PQFCqZgs7JfdOWb0x6mzaWD+mBpWQdQXMU4ZZ2ISqn
kulDQU+7wILAuyolpDMwxOSJg4TrwaSrEfhb+XQuncGao5jsFgRLprO7F4tCnK9Jga36Z9Lbnd7J
iVp9164iwmENGLFJGP4kN4jqYHcqKnjEuCfGPk2QUfBBfqitMI45KGiNRpNycBBHhihbxR7jmrV+
l0seD9WrbXKRr0j5f09GY2pGeLDOjnuKGx0FGnb9u2i8whYa6NtL0qtPvas7DhZYxWrBDqxCmawY
E3uPz4FtoOD8Bwvcr8TGxaQzReu24qOJKBb/racoA61B2r/yrmblRiVE3Yx/amJBBDK+ML37bjKs
EAhmPWxPU2oX3w513l2uWlrJC+PYQh7GseKZIJsgrF5RJJLz9f2TJ98Glr8pVxDMBHiAWOlVFIr2
hNJt2hwITd67vM8clInMv7s5T5cSQsrpsAkQrTCoIh9p36yOE1PYepzet1ZYq7WuvHnTx28TwjdB
tzX+dLyL3b4qzXgJfN2WeGEwAQiJ3ighUd7UZI7U4qDXObfJfAHV9FD1IvnX+bKI+xuK5TcVA882
3gu3tvKIV8BAW7Id4pPFKF5xqUw7SnUHWGQj32fHDOX5sz5Hrbc9tDDZempSWSg9j+yYdCartLsi
jZV5pa5aKI0k6j0cMTv8sJHKHumzIbV9E/aAoCtOVZWFmREL2OHqEYHowc2IZCQVoA/wiLgKND2Y
5E2NmiBYwJniMtNSnP7aWNPllhGKVzDClEih70nbZnnLEcSJ7FU1DgOOwo6OWtkTLvJn7cRHzX9g
0r5vCG1eltReLoIYCIrGJVG9dHmscJs3vl1mVO1dOkt5lscdTLaNBbixL62mUeHsfDfqhaahlFmH
mxiDgWzOXOyUxYCrcUjFRBux7MpkOLWkD5M/XhXOua6e7jXghHE/7IbrFBS6V7JlTgegqLbINBGR
bfII0aOC/OQf5Cqt4ifuFceWASpd3Yt+MnLbkjVHCk5iQcooLIBRqUAgkiBOVdR7paGQ1OM5iLUU
X1bKgZUBhAXyC/csKmIORJQB2cfXyatzLDuzxRbigXSVqe+DIMeKXPlD3PBImKZ08g7TUJ+WmWcg
ZwO152xSq9mOG0Hh+l9dCiJtq2HM9yGkXjqEK3rqY//F/Y+GuveDdZlE3LNOHFbC82MrbeC+8FuE
R6Pniaz3jk7RPaqSvKlB2RzsO5tMLB8wYdY8douKAGF1U25n9uspATmPtEoYIHsCNb1BzXoPA4aP
AJfq8WGCka25p7AsGIUa/NDkjwb7vJpR4v3mivJ4kmmOh/K4ASGUdjq0efGMlkgiynBS1XiE2/NL
wUD02o6DIUX/qzO1GS5YST9z/m889kngdWNitnG0bgGn3j45tIK/OZ8Gp+jjvtt/47HXgHGC5WzG
NMW8Zvx8uHolWqAWyqdfTYXKBfVLha0NbZeP1Mqw0Xoh+yE16E82zCvyar1+wIkc7b8ksyWPGQ40
VOEHouk3n0rVWh0nrPZPL96Oo9lwrzHZeR23kKw380OFm80CjrRnpe9n0coFEu6x68i/j5+eEWxk
cOgAjf3dlxClZ/q1NnGXHWpEQkaemhqswJZZ8i7+SpHGeh0w5AEewK6X6ubnaWIW0kMhQihl/m94
h3b4RP6NgejASUulCLXNTBQqh+ezmQsD5Qj+21WejN0nhBaOLgqnKzI5xpecOZ5P/R6CI3Tx1J9N
CU0ychAYa7nY4JZ3QQDp4lqModhPAO3dq/gs5IVKm6fElhnC7SzfS9JsYzlffGC/zDJDyKF+4htk
C9iDN6irl+BajE45e2PCF9IC7X4cXAWR/+iTwPCz5FPfWrZNHx5l9Fdd16QSeItk1Yzsr8hjO739
HZYR4U3iBJpgFC9USA3BDpNYhoBYQ4txTk+YUEQvGAFIa/Hg8m9+eiJhMgLUyC643lMZqbQV6tME
kw4y6se3MmcNwEey5031Gs46oFrgWbczE4xr1P9K3sRiKrEx41RR6Dt99Nbn1YCUZ1+X8fQUtka9
vSs6jexqwD2yDEzzNHX26Y65LS2ce3DqIhaTmTs1fb18MKyaWv9LzHwMlNwSQkgvkXs0ZtVLiNR8
bZ75PY97j3Su3uaDUI+QqIDYOMtuuNs7V8j3P9cZ0rpyg4xj6uerNUnAtfQCn1QOyeOyiDoQPznc
D3vETxNdQkreh6FIiMDqmgLcSRu4qaYZry2H3OwjDmO/wIOaoHHAqriHftU+0aoOEkOktemlihZc
EaLaSx+DAZoi3nw4T8FczJRjs1Xe972RI4lAG7StwXOjZg+68toZeiGzZfx4FsT24KExyXMIFnio
+16Xnkth17MTinbL/8vZvxkpGLN/GcWIH3NYcieN3p21X3Aag8JJ3Ms8t7FIhG1edca6UJftv5gc
kCX6JZQpzvM2x/Y2lkwgE9y5OAt8yJ0sIxZl0e/25bqglQNgfaXwhtITXAEenkhyBBiA5QGkELhX
tHShwnHpXmK7YPPZmv6aVoeNIodllZdbicinJzAUobFpsCQpbb2isCh+YKdLmV8WxbN+T0knSfj/
IcpaNBapbctZRAUcQF4Z9oXiefVz6Sl/fdsiPvdCRV46Rd+Ww36P0QiEM4xwGwQOJCIEfkvZtypO
RXxCCvEkYpKvZr6rqtPp+mDjbxJmG+/4bDFohOvmRUWKjMR5lspwoyhed7BI3aleihKnBa0WTGtP
6u3wEeU5J2XEMNZ1diYIzLxWKXt3hk/+eHfClet4QzsyObvfSXUit+EftJu+AcBTGRRTUkp5rfP4
LehIu0iNnMzTSH22bEGI6GSGH8FpghQG/eicNk6Q4524MIozESNanFjzdXXPkip5VarAd7Un02RF
M3r8ENFlX99frufSurqaQB4Y/MCu5Opxxv5SNFyO9ZRc/G1JDLR78XkcBvyHDXD2rZOhICvOBBRQ
vrikxeRN5cGML76GxK5bPh/BczYbO93nCbZ5A/IrD6le9NbPSwtC/idHETuH5zgCSjuEiTVWWVHe
ooyuxlOCgi3vXLM7F8jLRD1Y5eetY67bRjqZsoTGcR6S9fL/A+uT1GbjJRPnlo7F75v2piojXpXL
eF+0EvFYZ2bxDaiQDi5fJPtbV8/jsJjyVXOrWCNpGeU40+haS6JihdC74in/q48A3rurhzMurBns
n3blK2gLtOqoEEbyJp1WNxTeKtaf7MaWm7QEuFzDoNCD0Mi+LCb0HIb3bne1JOIU0SbWh/VgzKqg
NSbniIAmgeRW+wYJw+hab3xxKQcdY7shT9X9Wcaq01kAdzBZsT3xLO0mAyDx1xqEqPFdrhL3eXU2
NR3Cg4UrYjoOA0kOdYtkMybjfDayQ66x+lSAPvbUZUB+4Q3xZdi91iNiEz//EuQyhXC919VzSJpr
9HVo6WZ1f4rj+u6t7MYZa0TEEj0nvCjtmp2xTpdpqSZ9dtq9/p7Vg2azjaEw74eW0jKXAyuyyjbG
u2BUXLOSNk42WrptXW6S+bxjL+ZiN86G6i8eMVmj63Iga51liMwzrgnHHPyA4ug7mVXnxVB1U1Ly
NvAPy82+8KfaJUVJhp8e0W4Kr5P14eQmp3DGO38l6sW71gj+pBnHk+d/liVhZsBiOzBuK8vxr/9r
D/TPxMTP3zChfgWqoJY/ubHLHN7PHZvoPLlGAz0JBraETHRs79zSwLqMOSv773m7NquF8GfbevaR
zfgabjpP4Bo0dJYRxQ0bs3quSw9UYwjE+BAfT6bNdugE4/9slyFjBWK+2DrDsil95sSwW4MzpV0x
P1OtxaaHI8ugFCvDCYV78QS9GczI6+LIQJgGkzpeAdJ8Lti3faRsWMFDFz3HHPlVmsxgls+uyZCW
pJsqk3NqUbp6DGyuVvmoCLF6pulJLcHpoGTCcxM4q3ZRoxObEHa6M+D0KYUlWJP6rOa203JU4RAU
/ggFpJtD32Wtt6gl/mi6Pob6sKBBxBuT9ZtSWoTBQKBIShjWoyZmGNdEn4pyKtlOEligkPbzq5dO
UeDGn2VYi3hDHiGLoIrRVflcGLkoQx7lt4f2mjUOAWlXf2i0Fnv8uyF8ifQC+1TdxWwhsa67HWBz
wrexOTi3RylYMTfotuM9/b1/YuQOJrwKBVKzqOQoKzGekMYa6kXsLdVI4qIPb/sg+4luvkSkILn8
tskbRiC5VZ8/42z/c35uIuGFQzibto3dK29gvpMQIKC0ppqLLPblKAEFT7Pt9+Fodsfrkfuhgcu8
aFuCZV7VpYeosX8hhIa57pIOV6CRypHA+cSI9rTOa7i/ut9DFRcoClFb6K52B5zk1KxW+Ym/XGu1
fBTtd1sJo7yIG2B4QgWg456UGEhJoFBkQy4bcfsRGnb3UCN+TySWUhjDvXnu/watP6o5scjh+o7c
IsGi/QjoA3pseXeCSXmeR6g6qPtYoqNAwvZvFMY0zLlpxYE4a2jfjX/VJxYBbq/hO1q0s+lEjwnd
VcvI9+y0taSozSkgSXQbq5chAK1B3HnUmV8hlHBs4iqYN5xD/5Ckj/5CN5zsb0+vUdiT7lqieRf3
m6Ux0UuSVspQ4xJCsAkyt9jVmVLBJ9T2aD6jOFKVJ7XG/NobW+Fu2ZlCWl8Uu0nQVCBeux3khlPF
JFNBpRCKuN7WxH6rMP3JYQ5Q8R8Igd/GeLJno5OqxN9kodm+OObSdKE+RKpz8VQGGNuYsF52bsKt
UJMdOWWASid97ihjrIg+5EH1LBOu89nGqayU7sZhg9Ii8gKhCZjlT+tK/F9aVZfR7cWo8ME2B/P5
NM2+Ll381hnrcc+MwnyMz02cjldy//ISH8BavsLYO6wKL05rkBM9UMxj7hA+YLzbbzPVe/H2s2tx
t+eyzgINUtKQfvXOEGqN2e6nyakgIZX/7CqjJuzx87XQ5P80osIrCy9mTf4B1GHsUOuGyU4nH0JZ
aXIJjyjKB4CldciEVgCfysd9rGXPVw/2MsnAB0nR1J+asWZOLJvkGoeINIjIm27Hy0Uy7A416QCg
RoD1eZnZgIX+xAnWV+IxM4KZ15P/eYhRkTP2dOG3mE5omsRrW5MumSL7bRYExH9jEvqh2F4WjKAc
gDniJjmbXJo+Aa+JycENC0RicIWne1DgKubeF8t9zdVMLJF6kVGh49ss0addI5im3fiYvW7ZV/Er
Tu0XpmsmpHxMTsXZy1SXfx3uiYFhP0sKT9usCJ1/Zp9W/oX47HmgOL9x1a76Ei2PlJmWvD4NEKg+
vMzmCoXioC9G7QiPeaOO/M1auNs602ChO8Hw5Egj5gzmdSF6tjT+5yOE+d2imAbt1uBWYBMLgIjT
R+QnRt3EBSBUHS82mrcUhTCkTJjN7yYHhpwYXArPwzMSgfFetRo00hULRrcdxJMLwRgtLXDQch5j
d/0OlaL2JXW4cFRxOckJrOno7+Qu6uFKjxzS7KvS1rF1+yd/YyUTUJZQv/U4fJXQQBbTwGvf0tCl
yCmdwFzNHk+1iYO14he4T8/kJ49UEy/gbXDW8Sc6v7qAcJHIJtUm6/PdPz7oTA+bHHf5TOqoqNAu
MgiRuKdUhPdf4amADu6bfpyG8Jdv7rPKDN9wRSQ7VmBFZu78ALDeznVnK8eRWKwRbGnEzY8Cahg/
2ks5meMN3rYwfpHHRpq7aRdRYd82yRqqdc6dUDQWPSyfEHNx9LMkonZYza4v+kT1Ez9rrGAT51DA
T2NltNZ2KApogfeyU/OS9SFa1Loop/FqBvKy+98VFYwaMR/oqN85N1Tad2q8zbfiM4GEv7mGuCOx
WZabPXNGgV7MzNvNDh5DrBBejufRnBklWj6WaWSEiZWkL//6AP7uicJGpuIY14Jn8s2wAtC60aAw
KkoyCa4wyxF9Q6IQDp5ramJW69captgPFxCYYjDEn9TCKHSYn8GhPlAj4GBX5imOKl6+VFI0Pr1j
+7epw+aozhprni6ceFyeLPAINrC0rjYkpsHWvK22+rZs0d5QEr6tlfqp98J+NXSE60e27Zlt/lt5
oZSmNfc1TPmiHaXJZnSGe8tp8Rah5EEjtdVPi6FBOFriNisztHEI30tg3VEDV7vY4UlVY5ghxnC+
mvaKJOuIdGEIXZwLkJPrFjga8t0XiUUA/zQ3pnbv2RQMu259Ion5w1pOoNfCs18qmh5qNqDXSheC
CBYjOjKp60W7BWNQrRsVC4R+PZMVcPh9zJB3Fx5vh/rZC11fn9BseLcR3cNPOjOr2D3J2Wuhfdzq
LfWN5wGOYvkX0Ro9ddfRdsZvu4/89Gv7LCoxhYYOOeadPqymX0vPE8V1kWQlLlInoiQn6QW1zulX
1yC9mhU25aMCQYp9mK+1WnkOlCV8Cq3191XBdfPgcNKoDen/4TvL6DPTCIwt0f7T6XlH3ONVpmjD
zprLk1jf9V1GO3ozXv82cYxWae75yudk8sUVB4JNArPh1yGZI/L0HaPI+CFNV6Zm3zS1jDJbdYbI
bfN3hxHyeFtVjzj5AiW/ZPaznDXejkszzdeu9+0IwRrz5X7qMMZYO1gzIMgs/uLo2KXJ9vcXVXcT
QXgUWtmesN0f+cUS1Y2iq0moLKnC+YQVgUr1vaHLAv0s2PeaMJKNSSDwJ3OSe2MzVJNg9tYYQAdX
wjRNcnGUpN3AFvTL5+rHBV0K0kFRPjNsGPCAl+MSRsIO9X62BWR8JZsQhHBZvBEu2a9nNThenbI7
o3JUAf9IkF8WeJMG+uSxelnwh5IpZUa2QR/Ng9HoSGjzayUc/n8V/Wcn5g8QlY5P1odKh0ER5gV3
Apeb1zwA1Q8QvbX9esUj40R9TqXSxJpVzpx2fRwYq3TAtkkR18dtMs5YXhwGeQMUxz40CH/t4SRf
zAmLrQKTnJQ1DiPGJEi+4R3k775fsvr//7vmSAUcv8jTrh4FLMHaDKVaVl0tieB9hTzxrUQBk85H
cmgaLe5+B6i18LAfcrz76Yq/CwG4IDeizpb5xk1RlvmoSI7hlCreE8iipUYURfeAQnzqQNUqJvsQ
xt+GhV2wZdHIdw5r7JiKPHOaQ6+tEd/zqqNJnIjBTAK/uEQshTqUAXh/0Z5Zm7e15g7sdtiKNu4w
RHCsiAG//iHhk+PdIsm70QpT04ESjCkQszCAtx6NGJRRLcOdhtsKvBao3gh24YbQbCB0MgAWHk0h
Hp1XfdH6zj5JmlAmSIMQQavxhq+2zu6iRHJF08dDNgVoJpONSzCkrl73GC7hHZ8JYsgiWc+Qf409
LbZmp/b2+7dP07zHIzWt1fZlNzkuyj7iMBOfUDjlFJtKt8/rgnI8ih5P5gjFWCu/QXMFjdN5bek2
cRe03xp/RPZdKLGonlRkuQqZ1ZMpxK/vMJmimmZZqs1U2+ufqUnxpbM7ACl4rYsNp667S+4N+paw
r1GNvHz6PCVy1wLPyqsPUpRg5/93v+VtQ9CT8fxObqgdOhY0doL1OpTRZtGYlYnBQY7qaDoGQ55b
eubGLo1lonQhQc01Xo5qYy9r/CSlxQvpy87N1NoFZ9zjvwnwUQlSoTLMTQ71wj2VCJ1FmvheapIN
4BDMhbThUKLEKuwgL5SZuQnIXhcFbyijPtgnJC/arHAqYCXYZtOg7TXFfa2+zuUse5uQBx47uNdH
MnWhPd7TvznNUYU+AAbKJgSrmBuuGe8poWoiLqxdwEfXh23xkET4dFzmlArqO8BiYwucSfoBc8+n
L8ZqtfavzAhopZV0w+D5qBlvbmaJxxa4yxMebg47YP23rUa+8T8lDlv0iLOulsAYUD4Tss7/s7gZ
pmZILCaQlU5+p++Yp3UW/xmc9E32DxDrUjCW8lthlds8aRCdGw/Uk0JbJ6rNRMm8DAzZboWu6mX3
r5V5EtyCkLdbLV5jnZjiBwYC4NBnbEbaHhzlk1mt/sB0PytaYp1ZZ089gE2+Ej6q18Nza4/muQDK
fJEKeeCUSulJKKN5FWvB1aXhmLJjRdtONtgXc5VOAg2CkYBDzaB2X+gtAZA42Urg47YhlJKIZmOG
1tGX+YGisJoYZiJWfbXVZq1u6xVxACaGs7WiBJRCIQUWMJshEdXglpTfgvfKjtXV4xGSHHrejNR3
M8/Wg0c2UQazuMOPFPywfo6JT6b4kV0LB+SsCTkqIYX8HjaegM36f94+ix74YI4B7SGT+vl6rw9V
RZeeoMtopfep2jN8KT/fV6ZyepWccrZmy7qtQgxkXpLZuAIQKBIkU2mNtxc4orzzZESLwXhqjSh6
lBYEpgQaMMCt9i4/9pubBnmqHHpkvlOgKLDnzL35DBJzGH9FOzKrmzGi9hTLcaWzjZb2+2Mf6OK4
InJiGOyyH1YB8gALEImy/c9CFQPht9IT/eGvyh+XSmfAB3QFrviwePTFhQhwxGDCmNeVF3HE7gkB
KwGdwLFOsVBFIFZZIZHULp/6rylti4bf5Ezx9B7VvWU2Wr5CrPdskJOv1TTdmB7Qekml4qQH/mb+
JMwup5/VEvGQZd9mVCols+NSVX+B/rUCrHWt7BawoJQkTgUFpxZAGpWrROIwudK7OH/BW8Ab7tzj
sZaMSc8rnszlzJTUHmyZlY9q7hGKNjkAeANIVC55PoIjAyWKWad6bh6Ejy+a0SSPy1B5Ohlm4hzA
JvuHC7ZseyoOjiE0EsbtiE/1cgW+ppYftxqoesPJ14K7dYEa84WNe75pDoieZg3vY71nrFqJTKSe
7YK+jrM+mFNtrc+3L+NA/cUvy5oInzUaHPKARDtTRottxy5CXzIK7bYDD5305OH0oVodauv3kcLx
Fd8jHGTK7Hl7j6fns4jpeNkWpKs0bJJXDon8FtVaIpHnmoBiXxddpk8UxoC5m+h8jVPbVRi35DM5
/1B8EhvMwzIgJgnJpv0mFCNpQo9Cr1BhFJebQgBDM7QwvXKrIwZLuyghiCkMH82/bM8nmQRtCNVJ
Kyyq07lxA+VoZUZ9Xt8ed+ZhK8h3O+W9XZjfVzqVRqrO5XmUrHYz03VOO3hbl8KE3JVQBoZTOTSX
IaLLWnF12cmu/+GJyCjqSPWwgcbE4LgtAFOt8ByqXzRoYvJ0TDvCf2WwWKpePDtpUCFnq7/+0LUY
25m4YETl7qPINzrwp/SN2VD0Sy5jyKh6TFzLXYy6bkhOoZcRly0JOhGh8khQdf21Ur8Zw0KfMHA7
Ys+XcFnqOk1tAX3CsZWLV5M1fdR099pJytcWV6udICuLV2V6lrKYgTbgfW1NnRZegDrtX4haK/0K
Ns6/DMiORpCC8Cg9nQ1RdfMw84pCFn7qxN2YynijBmq/aF5il+9a5aO4uvl/AjgY3S5WqMZ1Zz34
2jNA6liS9AZxy2vHmdXz8AjVJCnEX6lyy7re7pCVQy5HuNPKKTwAAI1CAZN18saT31d1TWHXh1cs
GCWaYKMPNAT6qD3diYz2TlzhvIX+hODDkzlGaYOSTMGmSduSOWkJ4XyegK4k5Y+8B9QD5QnyW4gb
/UFRlyidbc95yip1JhmzdYbDhaazKWSWjO/oKRegZ4euUm68hxUlAkVqMiz+yk3ChflwTTYRUjlH
aoeyYowgafpK82SsjBss2jl9j1fTp0oq5xeM6e6WLAkRwb+ZuqcMfaUhJV49VreAN3z8mHiBozPG
m+LsVLkUn9B8mOuq4svnH3ZhswKte3hk4rM7C4MUvsWtHsn3JxSkeuRekLIXt0YBSAdUgMnzY0Aw
CnZomv7DEfQjJMuoncbEg4JpnFobpmBUB4Zrbi+07++z5041npsWO/SNgRIFSexDtLvQXeQzJKvl
7s50qZqxvjcSkHGsAlOGPoBnQMeEkxMKkdGCn5BSfwJo44MFqYEbXHxiiKzasNJRBgiRd0zx9Zff
jPkTvv2w6GOQmuZcxizBQcaurF+qW3tCRveM39Ex1jEKKc2YfVZmlATyQB2W6HQcHDdEjZAyHHcs
9g2y6ytbQ9fDQ9P1vAOD9XssxvQHdRdAlX0oXcVwouQAx4b1cdwma0lee0h/jiWH+HZphl4Vhugk
2aNjyxtIvxOpyTTuxJz+q9D5HaVJJ73Rqta8U7DBHxp1a83/3sFKMlSRi07m8P3p0aiIy84x+0+o
+2/5C4AlN6tphNqHH0boeLIUT8vFbzRbc0EZZZfNmJCpw/UaP84NPECKbb0N31NDUQYA2IfE9gHz
lx5n93sbUymu6pH+7EUS0Ht+Mk9yCMP4nN7eZhpD3lSdNDe1knvHt2yS4FMzQp426h4HByWd9rSY
PzbRaG/3KhScWxIvyMum0UaLvELrD0yvFiXGMIZ8aTlSpvUF/8ydCY0SfBY71jTKZ3KMCR6UCQBM
YGi0TwDgYNbfcYlnyuH5IXTyN1z0sGCYBUA2y+wgG+PMsgpoHStmyKeNq6KwEtbfYgBRjbZIwbcB
a8dBXrbGqHhfFpa+C2KkuTZYVRdmqRnFKZuGVfMMcYhNendNEXLxFSCgxwVCjvSMACzyylcKzOR1
Hgnf3qMM1k5u5xAmQvcOIi+hTgCZW4P25VFaEBr4wnuFiO2Kaq4enQSWCOJMHjEnd0PaN34zv4Ws
M5l1kcmd1V95zz7Nzik2vSQn9wgxIo4XnEIdh7L+/hyh5cgVovRfVzIpp7rLS7QhAT+Xk7rQN42G
hBXQhsAFfE9J1L+z7+fPslwplxTMIyIFz7UeFk4+63d6JVq6pf4OzA4Kb1NCGsYsOBh/EqGkwHfu
KKtBCrsLeVh4dkWrwApDC0MNabsgKj1c0KVqjEFzC8WsS3RowWoUUDIFTTJk+I5IQBa35rYoY94s
vjvUWzaifXeZgbSZ0/dXNdrYTiutB5Wy9N9nB0VNiDU0G92Ya0vp1sJn7z2TOCCqz9o7tKwwgUt7
vAyQqoCb9V2GVVZic82o1SY0F1W5l2iTXpPWXC2tRTKEAuceaRqqsKcrRI2jg3DWhL4T3c4w1o55
63DWfwPJPllCNAwyip3+2+PVNL/qhLuihhVa4bYVQ7JcMdmnZTenRLqGvdn2tRMCMEOaLcFRZ2ce
eOKIzzLwQYQzzPEaxDn6eu2PF8//6i9MfTPi79MkoSm3fCR2YTvZB8/YEqIkbyvs0aRB6Gag2UuE
15FU5ReFEEHY+cCMpilNcvc6mU5j2w6dzgDx2bimC7dxkmgwaik23TmNT/SOnpbiShkd7+c3a2W/
PCAzV9PhWkAsyIKhnTIIcs6SiUsHRANCsXcQ7rMigWRSHOihC/ybLQI1YYGFw9HVZvujCjfmQGC/
UuZHfdm8vQJ0YDWiNz6x3n4rEOrr8DSmNKd0P0Z6T2JAYYKL2kRC6o8+0q5ZCNxetLrw6PBhKFvb
WyvBh4lcLEVb6m/vzXT9Geb3q7B2RkgP+KZraJtFQ4ISUaPQYuOanRSbtqKn4Vp79erAt0h4LXf2
aDZQ61p9U52KeU6dH+atlvVL6IXKnud+/rq/69RIv/WLpkyCVJJ1y47zhB70T4SCzzWe5JyQoq5o
VYCNItmNVNB9Fex8Q+YJa/3r7GsqWynHTKVRkQioUIb4rRDPXnETn8YobfNFg6REAajt48wWqCZ1
yq7l1+FjRvIEHB1en2NqpzSYM4cYlZJFp8xknEUTLccF0xj2PF8nMcLNokMHrz1fXY68zuH9gWVt
03pLYKJaqWONlNnacQEAcitwMew6h1Xkv2ejZkUoaxnpW6aywRbx+uwCrhDeCl65JTcds2WCQrgu
pzXXgWHlOPgTMK+bcrN2urk3f7VD0ocksci8UEp7qPxFNyg1ve6AfxFDdBxZNbM6UAwmgLnyNDr7
zVrKI0Svmwx3HOh/RBhbtC/PQLDrN66wJI15I0CboVQ20Rm+ROo2UzfnWiWWAOlqS52EcSvC9Xdj
MepjcP0p1Jg1rHGXHaZe9sxzSCqD+dFzmYO25RtI+2cqSFmfh3nDjLjoXy7yOpC4d8YOcSVX+dcE
QZ8kq5wF72yG+HSbyWmpuJSc69sZ1Ys5AUVBkBn/l8zgVdLc4o5kqeZtwW51az1dksEZ78FgBcYL
pWdvW/PoSXr98uknf6Z+SMrxIyBBOJ7fzLDfSenWtTuEP7TgcUpLOamUMOxUwNbOyqJMmOh8aYAD
iY5QgsFGPVrlMzRGJroGioVTjNXtP5zQjl1RFL+QOVAy14CmzImGO6wCjyD0zfHWKodyeb3hAFeE
Udq/bG5hvQ+yAysYAxj0ZaferatmB1Pdr3kwq4f/PeGleJrvkLCrIoicfqvrXUd69muSJi8XJCyb
N/DeLtbEOK7DZ7yVoltv1IrULdKznL2nozawF8WmlTcIJWdvjikmgM9CC5ougdEerw5MtH/FQuLi
+qNXp+sitcZ9lcBNFG86Xtew9wYoUgU8F6V85mMM57ElRlYbTuIARKnuWQhN0eD90gcpL0x0xUNf
dXyf5g0qhPbXQ0ULJS1xqN6Ze01hNyC8Lf+5zjVal7ZQkU0FHN+O5wL4zL9xU1z7rcw4tcHwS+6v
IiLTjj5fQyOG0/GQ7Xk+9mLastB+EhApWKWQcZQfrC8k1sUleOURTMD6S0mJCsJpHYNW/0CPlHaJ
D58eObjWwT1jtJEvKOa8g9T+vfvk6xcv8xWl4blIS/UHE3lfPEV8hl9zQVMrVThzc9s6FKEG7bKj
XtohfwdAxA7SDLKF4/rZtcnAFomXTdgCtuH8S6VZZGtzI5Q9ZhnwpThx+419yIB+yAoSFuS+7Qid
f3xxazKEni6ZxyFysj2UswBpylWyhncdSPfc4V/lV5RP9l9pYX41zY24eFTkTd8YJnCq5lAd1Cpd
IRMnS5GxACSwVkVlpmlkze0H4DvuJ+00vT89zZlWCvA72rSK+f25Gz5ij5Wsao+kogTX/GMVIMqb
gA4R80k3vrhI8f1J5vDqdrbWK/1CD6BLkO0S+xdz0rSEWRLTKMuEzSFZgKqQJ415/lSTPwLKuaWl
3U7PbfXpPij73j3s7czdWHrGFUpqlRTWRLAQR3qXuGO86+Lc+/infSrJc6ujgMYsqLOq8BI6/LHG
IRG7dxu5FKxwZfMsH4djQVt0ql0Bk53E7ei+YBNxQFDWyeL6d+FH0JHoqwgGDlpepRFfns+iQacg
wv8dcXHHD1Yz0muPYbNWMH1jSDgKsOkTiPk3qxlUMXkClamp5BJBwv1P3n9po2FZ7v5rOenMj6MM
goWB+LJtMOVum8XpOcT+JAAsQerImGHPGP2O78xVhGIPKD8c2CPaDOF0gMqN8Jl9CV5yiadjaAGD
ZvWMzcNldUAzbic1wKukjWZrW6DHIvGKTAt6cbWrOjKlKn6pKYwmQ2KOtweIkZUd9ieGKXZEInHF
e4uKKRoZslo4kK+wOdiVFcJO2IoKfNhjeRVrGlejLZtjpeGrLh5dSnJGYgJsfo0ukLpzBqLLXgzn
9RCkeHNZMTOIVeCPJNaM9xcVlgn2r8quT4L4kXENrybslBMEJnSMCvo/rpNieZX1cY+3DAYQRIkk
rrvLE4dRaB7X6vxWOt80k/WOHT6JzpGmM7gNKwIQAOZvIoymthWcG6XRs+ZnWFpgYTbAGCj0nL9E
zSQII07MqVdwvaUynjtDnZxQ46Ighwv9QjS52e7HJgH+Xk2G3ZSoLrP/ln1DnBnH+E4PWu/cx5Z6
WLY6/2AEvrLYrdlOAXHqZJ0MKyu2OnfB+MFEQ5oWULL7bjLSsAxERuCpGj1yXvXFFTGDZyTbAptQ
9SXv4M2dCYnbyZwYUyAFnXQOY5G8LiDWDP5tS6Q3WlW2oyOZdE3BotGPj3c5AxP8vXQ4agSE6tlD
SsJEydEPn60Kzuj28BPDDtL/XRzDV407cyXtDXVUdFpHigWXj/E2YF+Lw1V0awFaiY7lQOyBTYL7
/UjtWM0LUv8fwk5wzY5zO8dG8ksYDjyPwd4Bf9ta5sOmKnkJRQzXj8R3cqUBwfYKmQ97kukxFmNt
VSId2vIa1ObKjmgA4vlzr5Lku4BNJWTZpYgSVSNrI/bBmAC7jEkTjJ/4JHFAWsfiv+0vLA+inqel
T17XN5IaESH+AvPEfxH4Ej8GnIObcKgLzBqRRw6WnTsE56GrggJGdu3qQjrkec41znCMp1sUKn4+
/SfpD0/ng1cy294parWvYK7k/WuHZxWzPAop0HvysiFdWzGt27tuta2A3ZACw4OIh5x57a7IA8zO
daCqTvzLSyDrOx9Vn1zfd91Xgfehjn94Uxx23kdiL/WBtaWc8CIB78ESfwZSC786jwiM+JA4Saqd
cQWKO2wVNb4Gzr8CkmcDLqoRQeOBr97NPQK4Zh7JfylrynpuUZ47zx1mCThmO6bjjgQqxi/2rsSE
rDlXET0QtZf7/d4rTwPZhNOTvbLeuwqPTNcpuvdEyhQVGhuuIC7OcwPuev6IRtDGXrdi1+EgBIA8
sLaEL40rCu5teynoK9FYQhS05CY14F0hLwvoj1+/BRxJXWUm+TwLLVzlx7xBYzKvESDLOhHk4U1T
jUfmaZjbZg/gshhEpyI5ZU3PJEewnxAIQuu+AIQ5JVQUbuN1YX/ljTu9LdSA0r/pnU7MAit3DT0p
oWAcqA03prKTCY9SGh7CtJORwKYQhqE/+8H6rbx75KZL5HqdbSeeNMH1Ws/AteEAPVq9gXgf0YGk
iuhWLwycOtwfx1nj6DwGbONm4H/BlR2JJUX1dQ1r0j7MwYWvp01hGVF7rsJ3jd7nGEVmNFH+wis+
DZxPsZNHaOfRQ6+11K4yFiS/GvjkNXIf2Rt58wVIg3c4XD6Pg0G+ZkCNAZrGAEs83Js2Fg1CQKZ7
ZCvdDI15JqVv5WtdYX36fuannrlK9zjegPpzflP9DP7QPN3DGTTBSbOk+8L+pBe3JX7wIecosyVK
mkIjMRxg9D41e80KWI+pOaIvgpD0Bjz1fBpVJ0tJd9rQyr7L2YfbbVE7Wl3TEh0LYGuS/ulnD8kG
ME+/zN0KluEmusvQxxJ7cMsUjL7vLgdgzX7zpLrvidhIuCfFIUcQPqAAS6S2CvJ5NNi+DIc4RRCP
u17EjGGfIGZwsz/i/pAEDlVBGydzHzMoNUIWhgXkWsjE0mc3MGXxIAx1LlvjPoSMyhEZZGUp/bdu
0DkoDJAV4tgGY9lJV7/HExaHZ4hG+4R1OGxkgVpr16x14hc2lEXMdSg9VLzJtotHIfF6BFIbfGGj
OFf8eEVn2keaeBler3VFfyqsxZWD55/AhGtxhSGK4MdJK6idz8XeSI7IF9a0krZtQp7vi5t2FCRT
PJt5uZ2+Lc3o8t2n1CA7jezGRV8YCxVsvpxLK59qM/TpzCmMfTg3unVUQAk0GNhVTjT5hwEd09Jz
Ag6IsB/E/L08Y1jt30J8cjFuhscGrNF6oJD/ghtS/Xugre/p/mROX6R1Eyrg/Oevc78eF7fycbtc
0ugLvoOpY8tHvtWuc5yKSfSn1UdK3yvpwAHZOYg7EWKYeLd2qZvaoQ7xpQyaewD4b91AEcMfU7V0
BUdrGfgmf4EdM0AIFy1ziGduA+o1fY287RtrnrzY9A1LM14XquNs8gQkXgVGsT+3XNmu2KPvF7Ai
1nDnbGqgm+MJpNkYzRHD/o+0mDxy//T95vZqtR53A3XEBl39gzQXSbReDbpnEI5O26DdU+m4U+sq
SJKKBBilCp+q8J1zAyTZ6Oo4vSIXv7BG31gHjy2H98Fq3C+avhK7tZ38ClQfoeWyb1ifxbp6LsV5
0Zxpn11iC9ABsFESiEejSmrSL5RXKKdIdg6n5qyEcZSab7xmGO2FfH09csaZI55ejdoQTjmDHMce
tL9UfXV4udx93gi4lvklMtyrskkf7FYP/2qlHE0h10LWYcKNie5eUiFNmqZtMZgtC9HQ8LP95ejB
sP6TlaBe/KUQsY74BRvde86QEsu6y8lGNExgJgGd9TNvSrm3FqCdAFftPDvQ5+ryaoSM6N2kD9iT
KhsQ8X96rb3A0VU5Zw6ovo4a3uAONIFMzZCz+AV+kOBfha4q4TL8X/3sbR3BjdZL+Gh7kCdzpCAP
pj7xGXSPdoFNwPBJ5v7ApLAUnQVKWeMuPpXYSTnQ050ELRHT8zR6098wxlWtLgCfTdp7yR85lLUd
Ec4o4mRIFgXS/lDsm9zpsoXrS1gEAn0K9BLqpffB/SwqhZZNvD6wRdigrudOQh5ELEdOd6xVThUk
eYAWiPjNjnp2YGJ/6gD0BbZE1WAzCRYsi4rPcRROwxbnnfBAJT8RVQigz64X0n4lfTlFQSowCllx
RtUb6egDk6EXPDxoGaFIr1Xvz+peMddqIS+RVEufW8vIlmxcxBOlzbyA3C3N3sQk9TkLfb+46pMY
8V8IP4YZ3UbUeHL+JqawOnAhZB0ciZ32g0p/FW8F05JWkMFgQKfhCwgvp4iqL+kjUg1/wWwXUviB
n1NyOvR/D03QctgfjaFp5xAqHM6m5Hlyzk8JIcAVEPnYrZPmhIBZ9uHygMnhNHYD/4FyeLdTbH2Q
mTsUlIugiKeZiUxV/yvvYCVNpEVUH4RYvrQUdFPBYmwGDvRgqyEKk64lvBN1U9o4iTpMyGnft3M0
gvO3/tKwgG2nE4iQcSVGuguMpIsRum1otocLQfbKynboirha7pwLw74HIxI2wqFkeAvdkQ/gSkfe
hBptyAHu0mYEsZdx/mWPoqosMsL+uvZRM5tf1f83bIgd/7gOcsZeewUutQAeb4XEou2Mf/c592vz
01S4yQhzNZqpSxgu9b0309LVNpg5VleNZlhRSc70qlgG712ncF/BykGuqxXcbhSd34HOioyqOQ4H
5bhGkFVHp5pOUdJalXnN9/9G8IoSWcPaKkb1AHLFP5PMgoPVcJsrohlb5BKXcqjYnOPBPBTNmqg2
kRjN6NglpwlFg1bv6wKFXNR+x38hJjAe6k3WJlKKVoFtM+Y8hpdaJXW2dgdoYpoNG0kPCUJfkod9
NGKQi0JNpnR2wdOsBNcE5CLrEOfoYYJP7fZrLoTnuttK094xLG66Qg2GgwNgniIFXp20gdbGBODv
tgj3gBJyofFZuNFLsNiar3DtrXkijaTd9BUVZzBfqKZqmwWFMmnj0mlGlyqbbLUqmgFDpN7lnERA
w++zYFW1wfht93MieSIkGYid2kPqKOHWokO372WYqWJM8Iyuo0Tsri89SiZkajWZai1tFC+1NMeH
840ri3Tybk1wZXO7+0REe4MmKdC6gK8WmPEjrDksY4TSI2bDb14GZxPC+uxMnnJmmX6ZjPPRPsiK
N1EXHHNssyhqKtDDgkDJLPmILpD0dXth8VQAGIFKdcPAnCgR4Jr0RXpAAAIsiPpd9MOrgKSZhhPA
anmLkqcLv10rNCdU2WtubmrYxFXVqy2A+MAkEJzSOJOYQeyyLy1+q2MCNlFXgE2AkwQfRDjXzXlb
ZML4KpnsllTFL13D5CvLnKARHCVLcaHNzmFE/euU6wAQHFLb8oeWVsgQDVKjyKWVtfALeu7h13iD
ASzJC6thcG2gwrsDC2DPIBl55vLCPj6O0yelubnpq+vS0HsDfhbCx/U1Lk4FS6ixGKaBV8/TXl4O
FypmsjyKPWiyT8mUjlyyjNqF96eUUwAXFKPlqhig4A/S1CMxauZaXekKosKQ9RsgB5tX0thI0jpT
XtGYEp+6A5RKbrOUfhYDJ/U8aEK2GMQPWonQHwf0wjoq4MRrAHnoMNPFRedASkX+gK+QQENpGtWL
xavNVOjP58aTzYixtQPTzP955w3AGKAkyRwjVm9gPzXAqeaiZEuIL82/LVcQUZyF09uMCmWeAycc
sn46r+q+FVsnnLqyED9fCjxoCkjIQVKR5FJh0+/ljiwpyi4bUQE0fqXjyFtIH0y5tBLBoUpmZcLf
sprg7pccGGUkj3GjIsiiNn1GfND6P7h71JInA1uLJLqoLa6mwoMButPDZf607El5z46G514Aej4p
K4N4HuWIkM5o+AXrH0KDATrXPQdIYofyLd0WN7rYybMffI9mH4n+stEX2RTYTBLeiqdP40wE/1+S
IxXoUVCFcS47j3GsR08xzRV9BlvghRfY3G+J0CsPdy8IonhPEUYg6B+3+2Do2am1/Y8QEdOCv3LC
3I0gsZ5mhEkWu493CTgkR7GXIS1dyCcDU7pDq4lq6PrGY0+1P+xYPEZA8ACRUBHBYh8iGtyrkisH
pozo/+wwd8jzpW43B4u+qa1/C0mUDpOs7cQtdEPZZIL6Kw2H/T0XLiuAdvFRE0GOgFgiP/diWT14
rI6BPxk0HgZ60wXJAOuM94gg3OPi4jnzZ7TTyQtaJTo54OPZ2LaOcDSkAP/5FRxF4PaFfSrl4yGf
Xe88zNBY8CyIcsAK7h7ARVXdo6ku0dUdeUWvzfpXpodDYUR/qRwHYx4LqrqF1g3kPXcWaVkE+hpF
ZtEfYhzPlP+H4QRrkX6zCzMTD/3/F79JA+XoVw5esr0B5IIEwJ0YNmnhLqi9NchWXV0p/Oo+Wdjz
xSS0jftyLHIKQ07beiwYxiAjY4nacQWAnzmBWK+W4fs8JPzrpiDxkKlOX0n1mf2MZpt/WSSue+E3
fwQkBkfFf9Kyl0rBmurnkfe/tgzjJIXgGwy3xPqISn6g/lHMuSbRmqh5VptX0f38fWpYCtLzVDqd
296oKp5gDAzaUwFxk/+Iy2uiPKoV/OHpZrt9jeExFZgMkrTt/RBaMGcug+J0YuFjrKuMHtS7B9hA
dIE2GMCzSXJbEhMi1ZJJq33uMbnCC/XauquwdtmiiLVfHF4IJzgZH3tFItgmzDUf9d1CqC9+K4I1
gwfj3r4kS3DYunFOLNmeRCBZyHni8g2jKE0c0PrIIYThq9u/I60oG32k5SeZOG0aSf0vZz74Fp4q
BxiQ5FLT2FFUSI3yDuWN0dLeF3hoB+UhXYOpL9DwRLzWaB8XehfoI+r+Yp6zjfshRiuSOMNp+DXM
jlaFYOYzHUJTVDRYOejsVmV+EHxOV7Bew7x8YivWKDwTReWzCzYl7Dbsttv+16ym48zZn1V4n9DU
qhyNE17e91hj0nccKhu0LX4MRZxWMoyz7iTEtBUKnsdFYUX5ttlXb7KeF6zYBMqf0otCBiAyt4oQ
dp+7aTAHbGG72i2/iendhN26o/K5NG6dk5hokpuhf3jfefWBt9mAhdlSktHKCdWnCEbw72HawAxF
n70s/1O+zQIhDKMfvBi5meqYIiG85ixaj2zax1/I+93el5uijCZ4NQseTIOg+nGCgxVA7V14qQVj
VLR3S2ufDMUc31q/OpsJbEaTxXerQGdwolhFavDHDCuozicWkDh06zP0TPJT6xofgVGgF+8WCFiO
8pJGOKPdIzcaUKqFq0totUaeJE+6/q1t/o9zvb6k4TUU4Y9sxWeiLcuaNlLg6sBuNAd4VU9KYBrj
l+bxGEn0BVVx1CwviZv6NK1AtM8yUfhDZyf/q/jFbj4sJbjEFSZYNGQGv+udkrnTx8nbUVhVcqBC
ZoG5opYdstmY/4vUGCo6uj8eXRGDWYDhkjhT6J/dM65XT7uhdffiSdEpz//voeUKdfKuqnzBOGKd
vpFWHOstQUsxmgHcI+9Z47GXHcMtSu2+d/lae7yIz8XtSezoEbIUc3Uok++abpg327oMLOG0PiFl
AmDjk6WHkeTlE6qhAYteEMicn1QLv/G+kimd8+Yl6Voq7+R6REkNWjup4e2pz6no9wr1eAppc1PB
0JLM7ol72+MdHB7rGVqub1db5ghzrZZQTTShCYPdJ+kFs9wobr6DoJvSjaIn7299W5fTMQFJr40A
6P9B5IydskvCLR7yW94IEGtbrf+x1LKn0BCxE18zKY+PSUq5eoVvG9ZA/xCHjmt5BYkhIkfjmxss
jzNzTeigCJfIkqRwPNL6B2kd8BmCDW9EcU46ZzDlmKmifB5+cFa9Q67ZvG6bmvEvox3o/5Zn3phx
Il4veg2JJx8/JEXtiJ6hHeai2lmvu77bqGu81v6+h1UqA5MZrVM2+AXfEN+pSdn8lAxSKedMJK6Z
BIx2tD0LADzv6ToR9jpI02bEvVi71lkWIsYBO/JPu3rJBKxG1Ng5wtvBfJA1R1JlVzuf5tdC69KH
12iIBOitlA1+lRHVSqIPM7GkhYQJL5g1GeHJCzrnb9SndSIilBOjotxPuwaiCxKOQdoH8eu1Y0hA
qojWSn088HIZJ8KPRQbYSCMw39nqzKRMcZTSrs9XsZGjScYqja/N/04MWDgqpxguHovx5jgliiuk
Ayc3JbwUcDs7IOOzVZMYF2JL4xo9lHp+2EAEchWOWZH3f8SNTnDyIdup9w45iA70ogFmu7/C0UTB
zVkkWeNUx0FD7BE4RyD3HjdKK/AeaZSgO56uH7hEQFLCHcB0yIBaIuBzp5SimFH6xxflTcmyCzQX
64/bH4dKPIARHg+CTjECkYaXnsctDbN6ljtAZ6+NmfKoLffb8nBo9ab8krRQUL3w8JHK0w9H3N7P
BuNU5ovWI4fcmJ2fGnIGNAoyN/LP85XCkW033EXEw3UeNC/aMMW2rVbNO0HjHS1o+1h27AySf8+P
1D7jhEVWGbwvAWaoX1J/KE/O+4kAcr5Kf8Gzxy+Xqqht2jN8ANNxphfhY1VQE8+EKftaxlE19Tdv
qNB8559VV0HCeJg4G7CFS3RC9XuCW3v947LodGI/koSWDT/pCYfq5OZ8xvrEGwob1NB762x/+pJe
TujSeYUEOaRgeOmCM7n18w/qYB9LkSzgoVpT8VCDnaGCBOTA/I6TgQiUzjzuQR13m6V2OoEpJ8zK
/HpBEvlEPqxOEXxa2CUsaU8+KtpP7G1IW04c7f+irS3C9rxYDsl2LjtPt1FCz7Ajm+4yUt4kOQ9C
BmpUa13RLwHimJetfkD4N+HB7SDztACn26fJZz6sc9UlDl1NRLZFNfHVtlCtNcwMWVHbcT5U32Tr
jfLOi62EB8YBXcJuohmjzM+Y3FW2DJVP0Xvhn6sw6D7P3OBXGpyNeMVEBZNzeGMSWZQuvXGUPHPP
ImLnmmFTiUfPjoZQ9cX8XidFN9Lrm6DFMte9s4U9b209J3Ypw+qWVQJ5Rd09pB5zgJX37YUypw2n
YX8FkTBGb2akao2l3kPAOEFAdH+Pku2KJrvs6iKsGtn7sqQZhsosSScS3J2KhRv/NstiiqMUQKv9
YIu7dPmyLC9495s78eB5rMAwnorsKhiomLKkMwdvMGKGp2akjaRiOepjwsQnXyx/K1tzvVyKtDny
7GGmmHyIlYAvNRx5gzgypp6q9nnkbEmgPetI8eAtS34dQHuwjtDOHgdmAu9VVfPSGRADDSMITnN5
HoMANOIvjw91g9q/MYNs9geeQemgDTVIL4CVhe7ZErUTXdwzmn2AdH0omDmGvjMYQlFWbYghs2oJ
ixK6ADx7syByFATOs636In47GVJIcu8OCVxFQ0L01z5vB+0zKLScyz2nuFcuwEd6pjZMmDCNVIqN
YRAKAot+Gb5VTI5t83E0onmy8NBmMc3Fx0CV8fnraN03yUYdwDTkegPZ0OORSVaKohRN0QWR5xPk
vdN0BuVEBs36qs3EgczDAH5bvC5QUHazWETS4JFepD098Qn6emJdiCnB2bE2kx/WHwZZ4Uhb7unW
kTUbOw+tH8X5ASDKS4iRlLnbwXgsdUw2AogHGgA60p2c3K3CRraqvMoU4uEuuwWLAfUa0Hr451ob
+Ura8LqSb8VAFKDuxBp3x8vytShUSBN0fZoZeQzoNKWQrNjpb/Xb4ao63tfxya6b6a9qcNIgIuHL
fIDm4b23teJRJOsY2/tmK7n8EKJQlh+nSzOjw8yiF9Y+XX3sF+JZDURofqgn58182upm9Q20mxNd
n5hQ/KtgjigglRyG99reQTa72efM99YbRYHPS39OR/fvsHGdKyWsaAEElniMyMLCeyYlBd5tgVy5
y9D2fQxhGIKkLyaSZOiMBGoGLZ0D5/mFT18uGl92c1ZaiXcdgxUlsKTxsoQS+mc2JWGJ3llzPK0+
nMPUlKvao/atNfBM4MrJAG8TaI9oymcSK0a6wLARbuhFCB9ZwHWXRpoMp/QAZFbJktc4Rv6qE1Sc
qy3cNU5UIAWEBKwlk29tCNKL+xTpFxBhTajr4C+qjFUh7OZnVe1y7susdnwZfsjfnJCSxxMKgKEV
Sds2mGY8f/8u0k4L2xA9/dgq30nCNkGCwaIabpTNCYpJs71c+DoZ5j3OSrjCi6NS2K2x6aFypDT6
vscc4d4w84l5VZuH3DbzRg1LSmGifhvi9DAmnEy6GVgq08jg6jM4Z0ayDSgG9Tst9zzF2V/UCvkC
e4T2jsiEt0jjat/6pREHrdtesN9EbcwhmVJBYrC9fBz9jbXAB9BR4yA2aV2Amb1GQC7EXd0dg5vj
jIZVmypNhVzqr6HxzMNNozF/YNgLGKaoqTczVYcYiK1AaAhG9DzfswNdyg99MnNvoa/y/YHRGHBt
mqBPXvfwYT17is7e6zl2MggRpkWUPmTIXuRXE71f1tyujPQDva6wImLcsUD1Mm+MpDavKIJ5sDns
1v+chXqFqY24gGL5iS8V/whnPwlyhASuWrDf3fIaTMzXoYEqXwbbv9vR0Lq2o/eoi4kGHLhzsHoh
rlTIZuWLyVfk6J8l9N6g/WJT/xvaM7NesIiTc9HRRZai9jIRUcGPW+pvnzg9ihHn4aeQrDkhYNHt
9XhbpCEZ3iDhnZ+a9z4O5OCZ9w0pAiTdMxVkV8X3cFv4RSca31S2epyNpDHvQWECYxqpPL3VnKLU
g1G66amlHnvmGdbMq/FdkLlQUqolOZLx56oCKmLtt1tobo6YWuJfEaZJ+AI2OTGYFG3E+eGlsLIx
sOqqTAAi/So9IfVtGy5m8dTyk1wh0LKJeD9g3QQlNj5i9N9ABHX9xgHKqYLspLcXnVxZRVIJDJik
OBuy0lb3u4LpjrbHtAp/VmGfg1L0Hyd+XrJkqn7BmfstMhaHHHd0B4k5bNaE2Lfcye+NLT6hg8ZA
lA5nDGx1K5A/VtJOjVOeQWN0ASEhgYCIFpSEfY9ZJfleKnA84qe6B4ZLKhTCMLSgp2zbUSWhZJpE
2d6c8C1gQxqGKkEO4XiMsGte4UtODA8WBi58GwtByNr+fDifjBVbLklipr7GjfpFJaI03P8pj2GH
RuXNrlvk0kIXQcyayYsGCLvpP+UC+Oszhpi04MAUafloNGdx+NtU7zRrX9UHDhT8ugiLVUHT+8gy
oZpPbL8Fa1S5UgqwZB9o64bDf+9/ImrgBO6ZYNA16dogRh6Hpu392tzuh3Bt2Sy//Ddg+BEY0/CQ
OTXSRtrScvt6+qge43tQup0dMURhn+r+8Bu2x7dQPEKjZoI+M98aNyHz0D1Syk4b2OD61C2P2XqS
CQYey5sEu+teqSo7HOIQ2ktCb+LHVML3Zc9qBdO3el9ud7iTVtmsc7k2siCdNdOth3PUKJ3t2SMm
QZOpCM3BgFJzte+EGbU1vKH8lWltVI/Vx7izvF5tOaU1+Q8twddAjHq8sXnGHG+MlnpvA9E2B+ED
sejvSTG5gZz8N7JIoMftLcwQuk+KqfLgZaN72XZtR/zkmSi6aMG2dP1rhHfUaH9Y3QeILhfhz20k
DyZxvwrr2wR5Xt3zA06IFSQGHY9hc+0d4cjF4ukPe0G/FvvhflbDMfGmjG6xDYmUcQcVZ8pgS/Af
knlfxHqf+575znkHCL+ihcG9tsOIG5vdBAjdL8/bWKYohLAqrpBLgPj4ZXod5XJkIzRR0gV8pyQf
QG8BMFHsQR5agHs8WIJ4c87QNLEMW41Srb29WuyzR++eV/zxb/oLj9nV5LJHVXRf12bZ/J2lPpKq
Mp/X+YIC0f9LpH0Fqy7Z7zEO+nb0gT4IB2eVSOAB9EHHFbrMYaCCKorokhIODcx1rS1hs8OmCdYi
Lc52cHMgpT9T/DIBKB+wsPlpZRuf9I6dLV5/Mp+G3PgUFEBBO7UGRQYMAuLGbM85A0W2DPWrSeNM
LCu0WJCtQC54vv9Vzc7K5dkkTwG/KEI6oLv6n+8RIOmrmgW+o8tCid1BYRi2TqJgaNT9G1EPLhHG
nMFZwrwlaVyU7WYdJQtr4AlI937TlUiE3pSsqBCX8m14bnjfxzFWpgyTD3TtxaLpyrBKdPkl0zoi
kA0n42g8SNmVREvcKjpe7UqGGD6GBI1+CsuvX9xib5cBgko4ayZcW/YvuxryXOIVexeyT5f1xyFp
MdOhHLIGJ2ux75096Rnjs6XSQUosRxW/KySuXgde2x6iMitc7SrYqICbSdXckZ4LfhK5g9NAPV4B
/Cha3t3DzKxxhTnL4lLanNCw92kHFpXrYb24m6alhQs0dYB3tVHamU/4o5RRC7/Y4Gyi4cqym6rf
rmtNoX04thv7aIm4KvAD+yAz2OPnsRRp68ttMMZepeXl8KJZiozl8C4EEcPTuV9/Y/GAHEGO5pWX
py2eZk8j3al7uOsfCkDeBA61v/DntAzZs5wg7YlfSinmaJcOSJWB9bOKNd+RJnXOND5siCtm7iWv
DjrgfBi94VMucy5Jg7MWmkms6orgQ20cL0NBs7xMEm5cD+w5fhoNv4zey0YAYQTlhl9gxTCYxI1k
4DtwfQaFkHLcR9rKoQIkDpQHKUXut9LkNKF85/YAo51PE05qkJleARPvPdXYsaWMvC7llKtkK6G8
8WCoLoJguoHWh6P+yKdEj/ayWe6xHcUA2YrsD0IM5hGTD0iQJiYwECASvMAqgYX+ow3Bd2TjdgQL
C/893vttQcEv1R39FKTqUE7g88VTzlzEu8VUz4em3SweWyrIM2Nglgs4C/L2Bjf269Ira4J4Xu/A
p5fasHXS3gz6aUnMpaXJ0OCishXwF1HSkDGhu+L+BbdyGRpwLrkckLYwSYQ3N8vjdS8JEkyFPrKX
57jC9X6zQh0MW1e9CRXO2eJUI8ZTKIkas6sNqJ80iPyapRMR3gMbtMs4wTe1LACJaFlno3m2hOjl
ThUtFqeswaoJfnNAzGVx5ZDGXCzrdUmenwUvlAJp34wqerOBuH5sHZgu/6qh8UhJCmSvlvQTVyFU
sx6lfsO7X4TXyrEfTpZBfgDygaloDi66gFq+dFKYXgMMQxnbA9JogMtU5DSz8biSxrdFd8MH6411
zH/WFj6VaFrEj4qkSzk3ZZ9xoacBRLMf9N5aEE6uLKpbkebpjh5ea60Rp7v4b2Vcz2rAOs1Akoro
ciSKy68i1HtciMUgVVyu0qOuafOIwVttvQVBkg+8/uipO77CalWIf/Gab540ClFcv88kMX3aHlBO
79yVRe0R2IhnngNQ7MITHN+or0CKrZaqEPxCbjHxOnzTX99hadHqsqKACYI/AdhNDe9zBm/JG3LQ
6wVAEqp1cQuB1zfxNDJAjOf+xxLFqGaJ6grVASQhvOn6FSldbNZdN+xaIrTXxsx1D0h/Asn7BYfP
0Zx2NeFXSMVAThh3K+t4nnOZRKUduIlraTI5c7qrHFYBU7NR8AsKbVnYDoSXNXI2GoIgA9zd0TUr
6Hn4/WMl1lm8ezDnW8gLG4KmisSje+IOp7jUOuLJQ4jTmsa+RTSW8pbws/4j+h8VdQyj2Bfu4vA3
c5mYdCbJLKlTOtwfypsCA5yRoqNfBxUq5y/bb27KSnnddVYfoZsROXR2YowJ2EetWKhBVcQi6kW8
n4mAlMtZehsxVJ0O0IygnhPQGEoSzqK+xVUJtHc8zCXLl4PTeqSxwDteqlZJqwE5OJC1/p3i39RW
Rnl2vN3KZ4x2c0OJl2jIsyslMtvbpk0Y6UJfGoL3kk17H73JL/vntv/ILQktRWPszAM5P/Q0CUzY
CON1Tc9WHJpNWCkMg67QHkXZPwGq1Nk+5rKBmAfoc32RoLvJEJSDLK/iW3+Cc0C7BjjHFrzC6sUn
qpl0DVcXoQiOmX1n5/xdQRmkQi5cK5FD7CCTQB3XfTBguQsMjDVv3r438vzChdZZVo6cW7s9OC+z
5k9zlpQi6ubG3KuAvBU+AQk4Yvuppmi5XldjSv6pLT3fpp0jBIrPqzQXR0QKT+RlbCYji3+XuP6o
FMHmpjiExoFvfBP6cspnFTksGXrZxg2Qu8zquQmB+F/efEIELTvh3qwnmvADivqYUo4DD3nIHq3q
ni/ADF7TZJ+Oq8inC/+gEV25MFvnPd/h1givvkPApkw5X7R8G2L9eKVpdGhoSrMTKDkJPUrOpJk2
c9K4pAYs7SrcKUijXx+hIQ8HuNQ/j3Wag18/ZOWAbpmDvDBrPAzYUyxD5VTes/JhTls4q3USfZIa
PgHlNewA0LoA/79fu+bnywW044nLS5JxRu63wGPYmW3/06GHfQN9P0HvTlly5q7jocEl9gqJV6hj
/nokxqZdWZhOxVSPl5A3/4wjrxvaiJCT0UEj+wcEJbzPywgGxx14l0jqmHl2Hal4zgLAFIRPh2am
IeQCu50BSDdAPBhWmHh3RUHOLMCJ/wjLSxBqyn9MuKO2wLDiBGws/8xVF2Cso+XqXpSCYcC+OLI+
FzKXAi0pwYdBhMJhLEKVNzpPxdeoaSDSx6CyLmueguqA1KsZTar91HlH/fWPmSQfP8ggEmMpbEYs
sGgcqEbCqiQwghUH26lMb6Q/9aiSVO+bF8lX5JHdkFozkD0DeUUqLMwdUduWeEd8RnJgeEfWuShR
vNM2hvZVcWRji0I/IorzfK4HH5vm/6GtwMgDo3ZrB03FY7JijCOOh9C6VDB7ASKFfE2qaHJgTlR/
KcbAFnNO1FUh/4n0SbjYdI8afxe2CdwHSl0G7HWgRLwujiONx2i3H0J1q73j56TdPfbR3vWTlJDf
DSq1mdicnek58YJ6hh3kPQuBirqZWlFvYfFc9F7VvoozdvQU8sJrHK8YgLL7+lMYeVC/KFCNDhXg
sEw0TYxwMn4OLxVi0Xpo5l/78JXEwUWJpLz2XtoxogGg9pWNKfKqy76natZwLAd96zLwVIKRmBoc
b0DQqxeg/KgxG3rr+W5zmlc5+L2rPFdU97yQyz4r2mGMg0RcS2bFZdsTYpNGza3ezQGh7c2SZdPZ
Ks+rvSte8S49ecasozH7B0aM7jRxIZMShnNuCWIuzqCZT7UZza0iwZ2CyP46bEaCuCarfS2ltdJs
ODBMTKAcW6fn/SRYkaKtzMDlKUXgDvXnjjsemLouiJZJHAKzRnWrTY9alA1MZlPvYcGycAO6M49f
oX11pR/HcjXeGoU4r8bP9YSYSJ96bxgd9oLayC3N2/LGglETWYVdhya2MmEGLzH2rT/L5z1ovo/V
3iB1mlkkG66vvjrEEVuP+hlxoP2o2OyLWcItRvupB1rs67CaH+AC5Q4AIdBGw5xxd20+XMw/3lbS
paZo5UP6RGUIOh9yYeq0fjhj0fmWM6u/D7I2G6gTNr1Lfs+rzyWr/YxKdJyWs3I6zhZvSBgA85Hi
75f7f4hyMfJEKIjbGymRFLN/tQUSPI9gPAEI41ZyV+ULO01uex/MPJGR+65W8hPqvJ4fbWQGT5UX
jDPdCOCeXwZys45nZ6aOqwXA90nQ2Ua5Cq4FP7i+3NLRh9foBHSwXaBtypbnV90yv0a4pz1MH4MX
AqKlJeK8KnCybQACDoQn/Pg2uceVvx/CVJ5vCvdTUZgLGFQTyD1XAVrKxf2DAy9EP+dKysenlxRT
tuINeDTCF6lI6O2zlcbRnorwgUvN1CdAHsSt49eWKMxIxZ6pkzYV2wYwKhGhwvE0+EIB/Izqq323
fiYIK10Z6bPw9IKtyIkrezxlzRKHhf8dLq+py+XNiZsm98Y8HN9TVE9RQodvRsQDLiJkCZC1gZAV
4YCE3Izqh1DVGt9b8YoU+vF2bmuxJcDS/6Y5JpxczLYMvwzuZ+HGvX7Q8K1WvS5jn+rpncoJmFi9
Vekrt9frTCQTlvo0T2rHTFN8iiwpIX19NUFIpDaxpclBN6cveD2QRqKbnqsWDEYozTjrHcwTlFuL
KFfzBJx0dTyGwDCbLIqqC2xoFHOMT3YwkHrgfLhXtR04Uzdy7uX9H5WpXXK9eNWIf+01KqA7O4EJ
YMvjE8s+ofYdzHd1AlFxBqFUHd6DzIhD83Luu+Xyqm++QIsii3oJukdi9rU9/jeVfkP1SxPacRgl
OZ7iHM1v2g3OxDMqIBPDInEF1dKJ8YgmzaAVFkGPTwVU+JWPPHhMvR8JjAsIQCahFvVGGpbpABSr
BMVva73yOZeTjXUO7iWFTwIQF7tvnNCiDx1I7oNG6KWPocgQexGqNUsB9wisc+ufAC22syRXYfaH
RYa8F8stzqUdztNz/g9qro0IvgHCA1ZZPzHh8Q6FCnSh5UqFYcQXTV5MKvcYtOWv+89HwsB/ZPaP
pz8fyenBiF5CSgjOYfRogaCrRm5htpnUDM69Hv7FL79iDiEF1TH2CZ3LFOJbfqLzGi5TjP7OYAUi
HBzb1QfJScj6etePIxOGKyyYyfKg7BpteBadKQ/HONnMtBDuirYgmb+BKtUfZJ9T5YjdYxyhIV+I
perJTmoktgz1DbfMFq6ZG+Te9sb6F6t9Enpzbj+WWFBclSviIqk7dbrP8vyubJL8N+6LNygcLLXJ
8YcCEVKjG5GR7FTege0px8gmk+VEWUXhAIWtelI59gmr36zBWtgCLw5kGEXGbtzE1NZ4ot8n3l3E
ameQfHu1q1My9hT/2CBNpxFJ/dxO3Amv3EYGxDlAdvI/oSXtx3KgyiNc6CnDJICCUB9wMCporiFe
e4BFE6GVpTf4HprNqEGBq1iIcTLRtiyLSgcEEaF+B1DzJIJIarRO5bHBQS61hZr4UvKK2IP2FyfI
OTp/jsoZAyzfThtBrK+y5wtm+rs4lRa+R/ZVdUFM6E3kMY3HWRYK9Oeo1/hAIpRzD/uTynWSNfcN
1yGaiKeP7yKOcNVClOrPNkSpG5HDiYRZ9LrM+0zNf6I9oO3Gxg1znqLS+7pfA5r419MUPAzdAkut
RyXQongTifVfLyOTfJBGQJkQFtKTMRqAj3sky0l3vTZCSg2TLue1ncbb4DjlIlQhSfC6HIodaOSJ
lfvFTlYEfLQJ3lnw3Xs6X9yw5ikRU1Qj8bvIANif3C5rKB+U0G6XVV7akTq+OK5DBJz8HKtjWvme
GBkN89yUUB0qYlg492Lyi54qAiPyiZ9ugSLmYEn1HNdYtaWFZvgjzUyCSsuXuNB+gPjJ7zGtkQAY
9EQTZubO6pdnS0lYAwHRk4BUpv3qUPSIlXqF5CWdYCY3rb0LY81dI8ZeWi90X9vdzweStm6xBuNZ
ZrALnURaIE2FD/ZbYmpTTZeYnAAnlPgyhyMW7WK6xCjvqqy/mVBByFu0o8wOdUT8s+ZBqVmdmUV+
XAsvqRRcsRkZWGAagE5YM7ONQXcMEgxs1Lnk9MSmuEoP/aV2bE9TZJZwmc41EFhuLK7Q9/PvKO/Z
zfLpjivpB+vnnH9Uqukq8LxAd7kHi2xyIIgOk6d7ZXXciYLEYkGgINTfgtK88OrnF/i5WqzppOCR
+RsGEEYjLzQ0Ysfrid8oG7Z50/9Pf1TyPLEOtuJoi6RsWDkoJO1unpHpaqXwV89bSPhrT51tMvv6
qWgKHdFuUsJKQoKcGRb5J4eRy2H1wf49tCH1/2ME3mFYWUvMJcFHW5fVWo76DQBhb9t5dJ0Vb64C
BP5dxb1wxu0/oQKUqhpJBGBLGnzRhODUcFxqntD4+gmpoMWFRXpyyaKbSzqDWNk8w2DaeLstOUZk
29tINCkl18B6Vmu16DQsUpCBJGF0LZi0V/+tD4abt2PvnJbev+P0v9vuZFSJOv3JB17inaBSIQtW
1IZxLD3ZxSZErCCpRRKH5hVOvie7ApQIHPs9v5aFAI/iFw9L0iSTKw/gzvitK0RXu+oV/wVSqb6q
xXZuVplRZ+mgZMDnyH0oyVOSYvy/9t2rkPYnW7Vh0QzePTV/6o1Mc6qanNEVeV+SBq8U1FkxqGKm
ltOL5+yS6K0BPES6df9UfBwFuq4umvc/P9hOhfsjhxLEgqCdsGOIpaPk287g+3iJB8ihIJVoSimS
4MkthAh94nVnv/uyti6ljPftmNHIWUYzArArzpoPSOuH5bJkP9jzpHfB7q6BiDkl1amMcNL7UwUj
NtxSaP1byYWb8uHmLHTsBOKBUfTteDwjX/w0pvnLqbBE711B+ea0/ELHcsGiMWSRvIg4KH0DT+xB
wn9JHSL6VHoCQjnYmv1zOdRzAQwrLOzTs/BZTCQ76KmUy3JGptPyJ51vVX6bMl84rp24hJHd7X9V
4WsdYlELFjxeZrNqbLjwffpE+f+2fedAFncxo6iaXIERKvynSUjiFUeo+Qu8d2vJyIfztKGxxF9J
AR5o6gT4dNVtn8fMngWojMgy60FXEh21uoDjzGlyC+U11Km4PL8vYSQOlSu2LUho+u9MUA2nEcoB
JaPxilRQXsrDZtuaDPdPX5klSb7NtNm7NH9mnZCv72QCS+NlA+cQoBgJkkdd1/3M4duMJ2cZ0OVf
k6WiW/2zu/sbY8UWoC0ozsfTbivOK1y5KKDVsPM+VGuWdbs3bjDR+4QGxRfj9Ey2PSyC+HqOLt3e
F5rEpr0MJUmQjWzzMSMIFJuJuiptZzRET/tH2UXYN4iN+UZZ4HcI9ZZfGZhNPzPLvvo5SnTfUoZh
bWkliRdB2UfCtC/BDQrxKR6JgUe9Bs/aig2YINr+PnL+42Ko5dMsPlNHbVzYLlDOfgYOS/1CCI8d
RLfJfMeGyj68IlKVU3rJRWhaq1cCWc+cPKKqdYHvXZ8+666l7pqrDTDNb1GQxzpoxZ42sbgfKW+2
FboLLLIL7/KjwEKbD8bBI+shMk3zOe21Un/3lE+8LGRVC75Y52WpsPE5rn3hiq9qqMtKJ7Z12YIK
n6XePoUb3vuIGXKe0dH4/JBW92HoYLyiBOJ94mYeQdYFsJVl522bSdZTAXyIYWVJ9f4kzb6GgDiD
ww3wp3BEcgExv+pA5TLQXRsluFFM7XoEj3M8SNP4TRpvAyWUFBlyTqy0TS6mmqWvdNKIFJ5IBbGX
i3QfppmQ1MZnVw+z+LiM1e0VEjttcakP42Q32vDYtUat0efcJWnMzswXIs0kxGY0Efb1khk3hBN9
lxWqd3HE8KGDez1vMu2t9TqUTRFkGV3tfmLRAtmHHTmg8fMz4lLlIV8lWCDOivtEA6gEDeomVFiM
QDovf1343PBFx264UCr8dZa4bqOUkjT33vRWdPByWeKWdX1Seg+n15lbycYT8NbjRDpK7bCw8bzj
nP4STm2aE5n/ssnY4ue2JTRjaHhwRQnYmPgAraWFyb4xnF4X6K7GXAa5zDElNQ9WMGh4SlMsjGGa
2fv43qQdWFCXwo9fNgjKTVH+Q5TnvlMZKMv4sivpbtPbp3BUqYbObqClzau5gMgbUPLruEQfddyG
FBqiPzqLyOjp+h34jF9b7FFizO3DjT/zxvV9QlkDBa/LGcQbFIq2x150Hgz4IgZhExzWQ3PjEivW
WG4iE6l9/Fi+8PXdFBG9AKB7BXzaBZ7i/cjv1Ck5+LJe1eajfGgUTf/z3Im6glcY1cl1/M34I3LB
48YXoMsIgnl/yKVIgWmAeK87W1Lr85rF9Qx2kRtmxbkQK9o5SZglMkrPgVe9ytHlahdX0pzcB2se
yS7O2h5xygpxj/J6Lx6plpSYcz7jiqcW3SyCnzPN1q19ZR6e/9w2S0FOkLGC04gz/EqcgO/kS6lf
XxJuNvRHIWlMHFH+cgGdvpmhDjKFXeNepl9cMQjHr/wbP+kecAvCFa9zZVYYNmNsGISNqwNf8GfP
bPykZsPfiMRv+5xZ1SI2uHL66h9KeEKOiQU2Ts1APIyUKoLbPoAHMG6KGafPwxz/sr08NIa3Os43
BATs1XD78Zw3mAipKS5U3P9fBbaI59jcb5lQ5QxmZ3yb00moSRpXJ+YkS/tA5RTeUlOGVI/23JVF
5M8UlYGdhWopC0NmJI9V8nURMhV0xOSscOTPI4H89sP8jQjpd3NTQEjKNnVGcHv6MAt0gNxzB5n7
e6DMgVnvI3wB+QrVwW3JtmSb0HW54NtJZ76YZDJVpeIp7vW+edygToTlvRpjllOB8x1HryDPCG6y
GnH7wqg7TmnZy3Et94wAaHfACCo/3AFAkm6PmaHLFWC2Blvif/MIXmzQNUjiGXk+g2i8L1MrdehF
tRmu66wNJ/zE1b2XJkmTw5wFOTXo8IV7sgXIEHqWqoxk1yIchmyCrho6gfXA51aEZwdVffpXPhQh
5/o098oR4By0TbqHM6etXdgStk1FQw4pX6xwNoUBI+LaTO+03A6Mtgkx4tXPHkuB65OePUouAdjQ
HPzydkjd8k3ufQtQaaMfaOeGsYv9vqKQbCh5HN5fa5fnBQG9hlD1GFi1GxV2UR43ChHMNXVZLq4H
x6wDe5FpbwOBSGYGONC4weyRuxBs09OqSiwVS3xAg+ZXAUwUP6J5i+wbPIsrfcQrKAoqxRRTHB7X
OJANFWt4mMSpqyJPD0pR4DUQ3SDcs/iCIQIjAYTFA4YDD5Psbhu6SAD38zStOpFE2wDKfbnUAtl5
jOrMophtKQJ/0iM7q5AmPFoE/QX9P5kDoxW9dEc+p4IZDofz1w28Q5cTkL+x134yG8OjgRRAF+v0
b50nNRW0f7r+3uuJ6RjTnBytsK0wfQwivBrfr8NOsH+bnbXbI5qku935LUQz0+/IxZtEq5VgZvCJ
bqBRIENJBEqjlMNmS3zJm+fVsjekh5v22g0I6RK41EhbVsDzNnQhmuPFBaFixl+r/y1B6Qbbh5IE
F3qXdEkehbadqBtwQj6jxfRafNxuhDG/bdEuRBngJXFNoS5fX8OamW9m5mwPcbOCNd4HcRr9jhUf
7vrpPGvWBd8tExJvymF3HunHiD1Gs3nO2ats0TpK3o8aahE1cobghiH1QvbaLZPTc67pjommIb28
GwvpTp9JTYkeDRJHd5oMjzjo85GHjMo29PkJqNZ44cfV78h2sb8uyPA1G7IFGHC7FbmLbDhZlDQN
w8IApCcICg7kD1NPtm63YYhY3x7yC2QeJAXbp5qoeSPZFJIOIhTCoQnXCLCAC+iWq6CrDk1sS5Bn
cNxuaNo+mH6wfXgRv47KdJn0GK9O76rKI7Tal4A70KvHS2jpmPtjADRrs1nkVVYJZhn1yV3p3ZCO
pO9CVZ2kaS3eutuMLxfft7T4mogU0O+TqVsXPFtKApv/hg6lTxHaouGw48dsaodMQLhvACVtZmaC
65JmOHO0z8OlZdMl+Ah72OUbB5PIXyzdvkv/9LQph/xivgD0E3gdiB2f1vIsgPOR880Fd3zfXKpL
NffRUSV6ibXNqbQ7/c5jxpjRahWjAEonee0iP0y8xwBZR7FfhTUxkxelZyceee3SHXEOYK0eojp5
2LAaZMVWShHNLm0ID/oG2vY+DpxerRxE1pEs2qB3LN5h92EdUCp35pvRFGzdZ3iveyqWqWhZTBpQ
7qfdKZf2LRBhThX4p7wdcgWAPtYzoBBuuse3r9SR0HbM7+Zdg7skfbuKDQcNYvIaEXI9Wd3lI7na
6AAglrca1K46GvXsyV5+C9Rfa3/EBL4e45cp+Z4zSACLco8kn5+561gUk3WAEpeY6IZu+b9FaOKf
nkz4tlF2Bb7iiIMo5r7FodeeGNn5Ni9fput8p7uJeOlp8RLX+zV+YM/u2nc9GfLcL40R7SdrLGhi
SbxGbYSxJ/bSW5AELT3tgzswkpJhaHpTANx5zTDAWAX1fpIlCFWtGd55PsFK9bFV8nQuFpBjVDuD
YpzzunspX8gNNLHNtCYMiKHlL1Hz4s5i/56DOSdR13bYHkdGw4RQyjquJsb0Sk5a0LVHe4/Cqg3s
7X2kArBOyeFgwy/DOtmONB/AI94H+XgDygKH2RO9cOxFHz8IaO2qZ+0qng0bOGVUOfMJlvS1o0lR
ngc1BRl2H4c0KJSNC/G2ryygR11fj/IVcoFPiaanYvPMLjw0ueJlP1vCjXO5VovTKLfo3wevS96c
HTymQ4h93tT1mtpmj7AmaaFj7Fwr2Te7npprqr0q+ftOdhmTjCRd5n2bCOSDDU4yfB3eboab4PSZ
a2scLGETou5ZqF4ozmyB0RxEaY7eP/XhckiB5j8V9YBjZaPoGjbMCU/2aoT5GTvrcyJCd0oZXizx
KaQFaQiNyrjRtJYmxRAddBFeqftlrH9iDGXEyotme74MsM+t+rMMBLpfxg+7lNZQuwiIpEkVpm73
BB+ykHqJBeceXMQBeZijv6beazjPFYAB/MIsMZLVz92S3ug6wmrwqBr+KPkGj4kIpHkchvi2d4zf
uRQdR/2lnhpYyEyErE8LgOnBMyDmJgjTLCOI6oZXv3buHPdmm0j2OHSg52VqQduT2JlzrbEvnrPS
2/3NCQ7FPKpVZAe97XReXYJQJH3bOsA0eBFhsjyJ9FwTj7aIJA2kjADdWvY4YulwfV5xE37PQI8c
HvxGyAXKwZJcmBQ68Gw6wA1K7RGOyiVSKQd29cd6uC5sn45MrkgEw5EaMfhvJUZWp005TGAUChu/
HEQCeaE2cvnuDH13m1x0YVvpPBRgXRrG63hAZWVAsCGpnHnU7fc3f2DsD1xvA9qo8zKhxGiGA3cw
0ZA9TyFGRBYYGPAz/GyqL447OT3YDiPLd8uDjQriSxfJlkRZwuWP1Vjg/hn1mX7kq75WkfT76rUx
jgV12LIY6l2D312BeW2FZHMROuQW3ByL3Zg5R+xiia7aMQyDkuRzWQ1R1rb2+WblwGzosXUOZIHv
MqRS3xiF3jFc746wJ9VEisLM6Za3WvWOCTcWMmKxd0jsZrPTTYxGhaML1YeTVZU2Eg0jwJi18ZhY
ohZW6L7WX1hFpwl4yN66udb30nvefaAS3KzhAObntI4gQLPOAygAxGPvTCnZDgYZN1hSRo5WY2bO
Xw049w4M+NHj9quBvZQDvFAZ53zK8d+WnN9OiLxuX2BpzaJkRwil6+it1yJi9phl039Q+/mAsXqG
cULF35ge6ls5XK6tIqPkwgKvn2eUtFIXa1fkpo/h5ZFDEfc2NV9kYyxukD2DXbH9za9FTaqYt3d1
dMwhsSgzBfBlUwlmJ5bv0bSImEkIfhpfV1Mr4+q0eY9rFbesSJDeMcU1BwDImg3/2mEHAk4YiQAp
b2kh8ltPuytSUM5J0YcYgZgUZnii73AWpR7C3IYNFqwZ0BBikFvUeGXM/j2N8ijdNjDzaIETwOrL
xQQquAyc7lSe9i0ofLaSXMbHn+1KldGDN1Svur9ZQx885hC5kxn0wgKZN8fIbJqrcDv6xg0f9dpM
eYy6fn57f7v8a2lk5ZvupHBvClZODSh1R3FSCtayqtP2LlUGsFdkE9InOxiuZT4Y/IDu0KFjjCPG
cBr8c42Kv4AT00TQi1Fk6z++JZYHYe7YUKMNn18Z/MheQHQa4oPVwV8SxpeaODoLVngk3ZvPG8kv
T9fPId0l04hhzEbezFIhGNBDh8g1rovdYmTe2PmIRRbb3JJ+f8zhq66DPUCs/FRSSb8cxFfod2S9
Tgd8t6ArmFns2Kw30M8YOuwJYioCMgrrqMEUNbem2TfeB+l5Bkg2vPQp8WrJyUOYlLWBtYdFCjku
GdloZpDoyq2EcLA7JGMUzM8e/134lKJImjSQWFYgNvZgoVevoMHObz8axYncNtNaej1V1iVqvJFT
KEn4F5K5NJANt3lQxRC4ZMc4UZcbLJ9ZBLvT5ZLXFzx9nzzCHgusvVxJOOJKy9NRwfrrs1T9hqf2
7ZJ4GrUuH/zSOeWrzLhopM1HrBNYhNZtFt0DWD+dnZ7P5TPVMuMfA0T7CFT1+zQZbDB+V4N5yPYk
IV9EhKIpUyNyUlc3lXJFnDTPLHEMD6k/l7zFLUXnjyLs+CYnvqWs8kqgoVkvso5sm5bHN5ozhvSs
FPwKqkI4JauLSyglWawdA2qJFpjDr+6KMlojZ3MIMzIkrRtRrzeBno2asdd9QE5q9oOxolKYXe+Z
w1k6dmKKNFtTG2MmMjHtJsXCX49wA8Qz+u6lGyfWPHtMT/aQAzry0xwHZRN5ZKT5V/4gOusSmpLr
PMuHRlTurIv5MK2FjzEUT2GJiLm0w6XQLR1zmgcDSCYOad5wBKYcWJ7UIl6SUXdTiPruUlCkDJAV
4SP6NYlhhLQoKOAA+piLZICTuO9dv620mzDZCeuhCnCg+ftCBlDs0DvN2rBOXkC6KisPK21t1Vt/
o0SM7LupYX5aa5XM/WlndrO79rIDm2KuX681LrFRzNVq732/XC/FbIrsyI7D/akx2Njj/54AWaWC
PZZ4t801I4jVkl4/GhlvHVpw3DD1FyDVnk+Q1th6ficiIaw1VpqlwQuO+EAcSeps96k93hi3/IEY
lS0eOgcWcEP1PqmCXNDaqec261I4j0oJTL2m3IwZBKBoJWSNSbVTcljfrilWWrC5BrxatQFWQbID
EaE/1rk1RGlILfUipS0NiNRtj+F9gM96F7i4DQNXaFFFTB+hve59RAN29BTMg42UNYPAQw+6QdiV
XccyGtPRN9Q0qZusJp3sdaFy0rmakk8T00BhxSt5KlokAKn2URrih3xAVQ8PD6hvDibGjYGTXr4k
oYy002V0o404kghudY5chU7ShStb/9WthkuZaBfMI6silN6Aqcq0ahFO40BoN9M323hxIs15BDDs
c0nvlmSIPQwhEOIaJVOj4fy3YgBACFFsuvBrKscKrFpSM8ATHP7xq+70fywRf3SMKnHGs+KsSm6v
LlA5HGrpz1CaMh4X5NBCw+zg1xvhm2IqsWHdBoMNVcErKe6htleikjN7qrFZHV5KUHoaBOsaK50i
AqQZ91RdOvY2id75La5LoY6fRgr5gPsiM7bW50b+gcZZf6sOiGeBV9pPro4xqZ3uEXhaktRA3Q31
i2b64ODFW+A5DOik3ECUGOcP+gZbdgBOLU2Bx++9Wkc2Daioz5OkRBMgwDg1kdps2Iis2BsgqAT6
MHToX5nlRTnSIFI79IgCr0TLwuVffwNgJItTYiOlqHs+364rn5rI1q6qmFs+tTVAjO+1zGQ3DlCd
q6yav1NUE3cOczTE7/EqzLcna+NQhIGhXbhXqtjZQROHRwSiUL4Y4K2jdP0Kgwv80jOGHs04CD1j
vxBp4lLMGojWFdMzS29FdacDXg1fK9fiLxxMCzHNsh7bhTqqF7fKWUMqusU0k9ufqYOqLfy3i2HO
G8Rv3qPNl8uhdI4cydYMYH6YbC2nLhwi3Vp25pKUUO/yAVxwDmHo3XPg6HJx26PzSrRbKC25rte/
y7I1ADiiw7jmszsgCAdQLBOU23k8ywOzOyQSy+p1RAO+Fx2JrtdGcOsgzZYeOUqE+2DZrHOdM7Sc
CQd/H6oAp7N3SxfQ2EC/6mgXMxmh+QSVal766sowPyAQiaBTONTnpRhxLxMDRKN5UlPIZ89qRPMr
PxVKaU6AD83p3Ni/6GwPy+K22KU+FkmEwyKObIlUfD1j3ZRv/nGU9oYtpH/7Ma4VSz1Yz0uTNb+K
XXZJY4VDqe5oxmGSrBAUTf7q9y7mdxtSfAheUXdJPTbzbtK7c254DhhyRs+/69hrTj+LgCJvevsE
L4kfXFyKJ1AGqWji+mTZD4UuuVX5ttmRE9sE6O4w+ikeqOvcZmjuNXwwLCxfYo0hxG3cChXTttef
b7y70leFb/1LUCbqeBialCKHwwzE9qzN3X3mBthc399ugGFt62ZWv59k+vY+rkOEAeozlFpgz3Xk
pJNYKq1gaoq+2Gqwi2HA4yXzX2Y84oGYrxPofaE2hq923A1ue10cVfigVJqZwdVjC4rb8tdm6dno
AVB3safBsGVF1v9rwPS/01zbeVQ9hxrYSGxU6UeQrQLRsKsvBOWsJyl+MqWeShDxf6eqU5I/izkE
Qp1CuD6bNFzMoFxYN2we3FSev0x7cPYxRF77AkAXBGCh7Jk6HN/0LGAp/TeSl2iZ2MGnx9lfQGua
gX/6vn1S5o7IbgYsZpAuS8Ue68cItZMoTBc5Gs0mtcQFQPPoJi7TwE/QWBhXdga3NV+zyzcSnYxX
K5e4WsxyJZhb947lsWmlLrsJr9QiEY9DuMIyZxvdrVgGqI0sUI746G4Ejwz2Ss4E0xpNcgeSTSjr
pnwG1b7bjuF89PsSgbqCe3B1lWekDvWKQZ1i+bO0xDVRiew8PJFIZwdY4hBdQs+nhXnsafAzusJF
hmAS6jschYWdFhiDaPWtNma03kMm59BvdadGsdJgYy0MQOssvaoUBYLt+o1YLSVwaPpCYo8lNVOA
0h2LFBc4jyIOgsjH7KbGrH3cgT4D4TiqSgqVY7j0G1NzzKA7bkTvsm386TEbhBd86zFQC8DYK9/K
f0F6fPelgEd9I/iYJVZRqPl/+yjBpLKTVNgmtpphaczoTMwcinNbScFBCvF23kiRRdSn2y/7LwrT
FgY2KHnd7I/ZeFOqSCh+a6O5rKPU8PYjQpjh6nhm/5U7Ln58bhKN9AjJpGBUxqobY6VsrTv9lPR7
oYiVf+Bx5HAgsUF4YTCbp8tu0LMLiKL0ynT3Uk4VGqz1HdUlH9BiGgdep9O4VXy2WJmQ+/qmvcn0
eOudebMSHnR1QL9alV9iS8Piy6zri39vB64OCsLl0dddTYbK0aNrChVrUaBLRAS5clFjoBp3mlOm
g01FbnQCKSWQ1jV6nv2cnoHxbrfHSfqPlrTNs3Vn/f8P6p8gRAc1BNfq66OCpzTcyeIEG5EM2vUy
QOWH8OYiW6lHg2ck3LmXj4s8akzdSri9pKBC6mQXt+lcJrt2Nl3kANBJLONMQgfH0zjWn0qySZiL
hU6yKfN4YojN/IQG6kAAXfXhisGc6AbNRBeg+K7r/3HdSRXOETueyToeQNk2lZhdWpfhXePujSqg
S6ONoSMEH4e6r5UmABUmCXqrONrOpapY9zk3VSKhOF3G3bI2b9Iy2DFUrdfG33X2R/QgDdjcxxYt
d72eLsfMCiZAGwgkEZNvrqDZUP9F25zbpti6zenme1H5nY9+15LAThJ23rz+ou1D0U+9Bkl07q8o
ZiokxlPlCc0hHk4aVH+gXHASfTxDfAejQaRsgIJLlNGUEHPrMnNOR24t3HkPo3neRq+3waj7d/Fz
14PKMik+RDMNltmrrzoxBTM1LH+pBhCnHxBdOqL32S3uHGBuqkG0eQzP3AVseBRTlXttUeUj2lr1
NpmarT8jYSBH88BNso9b1teFkP+J7bZEN8sCCrIA37ncdIpmC5tA76ZEnlJJRiDB1gVDTqHQGEyJ
bwbrTAuVg6Dzy+Dn0nmOsdWx8DDuYKxKXrg/GvrhVz+BhldhyRSC1HEKyw+2rtsCX3umEP0WPjU4
4C4ElBZSvsr6O+qqFAncHTy/bBE9TyNpKWOlWbXhjydyQ1zwA2/Z0lyy0aJZ1biCmWH/9Lgvk4qk
MsN4TMcxIL7XfN1Trf+wfpcDrz9JlitNnSRRS8u2Zf5d3qljlw9treeATdwXVmL0YWXLwspVhxlT
qZB5ZmvDuSkfctVQEpURdSllmMtlA3KDoAr3LITspGrOGVfKZeX/sY33wWtSmzc5zCUEmyJBXc4r
uxJ9MSb++0Ox5mse/Tj//l5Sw1Rfm5z+8GS8UpJ7J5Ea5JidzZw6ARn4DH6hh6eFa634u6tp2+SU
LndFrUbp7Quhz35VCh0e2iGzfM04aKWFi9qFk6dKq+lIMahZ1aHF0kL4La6Tzcwrs1T7NqRBhK2/
iKilfJI0Lpu75Vb9cvJgUFZtBSl5DT60ct/zPkbaWol8APunyCi3as9tIUbEgfcHg22UOt1Kpoke
yYnB/FHcA0g4v0hTjACKXoY4DyJRr34Q+vTmKNtDmcJfGJAKNYD8xVSABJReehtWBDpgDYVqpkdP
eHcc2PyPF4+wrpgzVVg/UUVw1iAIqRs/Aj51ATV639U6OCfnUrM+3aoVwqTn8xpyDVUXP/UT4tva
rJwnV+UMQ/oXvmJOy4aLgeowlUAkSlXOyjCJqzC0w6Q+vFJeCWimN4ZlvmdodhvNplOGt/NtAWhu
OoqOqQqKD4AmQ2OkHAnQW8/13j8M54hyDpbognhWq1TRm5Bs+QghBNkSnFZhU1YJNVWbfD6P5ko5
K6mtEW9Hb8vfp82u6DNxvkd68+IzX36mAbF4s6aAluJBfnsQx8VmIZQktLnSldfK0AMo03qqfytZ
SLihJkwmyeQ8uSmcIYXg1vP6sVLF6SZMfwwwdMo/xE6rpJRXxo0s5h2thYoAXw5MgcjK978nIX3U
eDXoWui5mC6vxBbO0UGXjSIBKlxv/YoI6d06X9Z/3HyLnnPyr8lQ0BRQdmuURtN4J4KNHSE63NJ5
knFJr1nTZEjKdRh1+Btv1q2paTgxUnufEunoAyE8ad05CZIOj/Xy8XhNHXyBIXwr7nIF8pdk1djy
vqgQEYL0TeVBoeNkAItdYBZCFcw2TCVoAiYKHrH2zdlqMAGM6msRMwhwKioZEeXvYmzYdmlYHl+H
cDZiUYslGCqQH3lL6V7AS33ckExAhMnl4W7q/hjzr+CRNhsTUAwMd7cRPFzWK0nIsVTNReRv1h4d
YwtsxpYODFBu/JQvTB5VhqjpYA/8p0FlFukihHuRVVoBhF4ZyZPit1PJ1ESf7w1gyUfD1sAARtUH
y0haUz12HQ7cHYVsjkabV0YLDkILKJAKBdWziJloYsFYaEGSvsWisvpIrA7dI1X9by/pmCeBY+rJ
NckKXIrDyKDUXlGlbzFXr//uX5JlbKzj1HwdlXgqN1C+q3U+/AM/lvC1nkO2RBA02yOkVmMmihJd
883vE2x+d2ZJWcjIif2KVt+SkZmXQwUqV+xmTZKJJf1MMg+XX2DTFA8Bq8Hd3tWbVm7Cpr0lTAaS
OXHnDQtcJc6Abj/6fNS70LvaEz/rj4OFKMZS5dG+cJtDebVqtDgAh1la1jcLWSlNNr1E7NUfQOOf
Hd9mD6Mc22QLLQEFeYotAgBvgCnkjamnYiMU3/sMfXxraePhufcn/vHapxknxv80v1/ri4f0HZMP
qRuh+cTxq5WYsO3ZxYPSA7luVt1x4z2tmN2ONRotEKLYhfv72Sm1IMxe94XsRyu4RORnx9zJbPRk
2S4C3WdMog1/Jle4H6y5Rzy4835LdkMVed0YUhICY7tuV+tfry+vw9kDn3cE59fLeVneZX7KW8Oy
oSqayZqTJpbRoAqwJhZmi26nUCQ1j9sw8Tajd3ZCXU4GdkiyjZuT/X6mJyw/0y3sFBgqVQ07ZIGQ
m1oL2zuw6Ii+sEMtyh8+lpkVjRo/5JsFF+e4PleRv+PcTQNut0R7L8oJzmyPFEwDOE14xRBX5cnq
kz1ixfNHc4OUBk52L7MQoehEf0s0tHbMEmiyxGv6r6ljRgWb+C8SBhs+t9XX4XpEUgOahNvH6n2S
MnRcZl5PQVguygx1xm/0YctGbCibXYWhlxDJwYKsa2wh2Ln7OFwncJ095N55L3uLgfTpGTQW7Wzs
4KCQLPoCqiP7w3qGun2gH8xMSC6DlmAsm1dpR4vwD/6BDprbNO5EDaxLjVPy27YX1UZjKMCe3GEw
xUhG6p8RL/2s2AecJtHJjHP8ySEnGerUm8jlyuHVx1Tw+N7/qaFgMT54A/l3mvti5nWO+Qvr+igk
RQiNdxX+hu53DIZy0DOqPG99+sQr7j3N17OKg4Iu5ijsPl0bQb25L3EfHboEmSfj3YO+zyL3np7g
OeVdNazMXWTi+8arSP2Btf9BWf3MSU5Fg2/4XmC8sf71nQYca+61T4hGT+v8rYMJNUjtk8evOLQ8
WDRbIdJxAoQ1zTOk4DcLoRNo5Nd3Oc+fwSoo1ueKaQwbPDk3oiMknXVwqZ0aPXFONUn4qUn5yRdw
ESCOQqCw2xMo1So6FtW5I5JLjjOYb6oHiuhkVqaFJIFiu6NkW8l8gZ7P1jnjYWHvdgxFUJ6nJBVY
Hw7Z7m1uwJs9ZUmhMYR/y1MRDqFG2aCAqQuOrXxPWCNYmzGowkeuPVSQ9csNHlHtNeaJhGhdDJ5b
W5Qlugg2ylJldm+ROf4/Av9W+yvqu0SsHJs/GSCPLGS9keVPb+PjGwQRY7hykLrjNliZ26lf0XAC
xBZnpKOQn19R5cClqeUOKUvDnRATTNZF/ySf2iF2n3iatMxzEv1Qv/DZdmr0b4ieFmhkieTpcJ86
12YTCLt4KGyx1zOK9R4giWoKR58p6o64Yy9RSe+kGSkzFRBYCF2U2y8U23Dyohyalh1SeEtbHMvP
k1QGP4ys1/uviA9htoJPW61qUoDQdqdtotbcJbi7d859P57FaN0Ki2BjOZtKI2LLVSlrx9Z8rzqq
Wuk+kPF26O5a7r0YJpqVDQBfKavbA7ILqLRHuNn9SzeNRLBctBY3cIYfYRSY9bKzAJex2KotSo0v
0ZZ4BM+51NEjuIN3BxkQoMAxnn5a5VoEiDj0dK/LGzpyKdxIUwb8j0UhxYi4VNSnFT7fdf++/0M2
JbBZs6aFe4dxLIXdb2bQ/x5iY7gtsFhJznuQmT+6jJKLH7//31vfcK6Gbl9rtr6bZ5h2+LwbGWTW
CYr+9XFft6fwgQ8H+C3LgaRrkq+hNJi+sYu/ksKJOVkmXjnTGAeJ9SKxxHWQhXW2/YeBXlnBzz9p
ie7pa4wV2DFe1MA0YT7iCDGyJZ0czJPt5PNukoiCRE1vUheY5Me6HohTAzLFBwu6lM4GT8im6tNp
cddf/oc+0xs4Ur4ZJm5MhULaUVfJTT4aJjcnXrxYCJ+T79kXC4Bo60ux4cIq2p0UWF66cxjcl5nU
/GonzvZV2foCdWPGeDezoJdY2DaG22f1iuWFbkvt1PgE84MjPwstCXctlhYZuzRa8YzKXvaeJf7k
nri7RR8nPhfdldHaYVTBj1hS88BryFforkMtMkNyo4ULAo+UBzT+FaoNrrYmH8bvUpzmYEfLd2/v
WRilIbCEdzEBRNav74XEPkityoqzRR7ZyfntV1ZPRYGpvk6Bw2vYRzcvhBvboIuzqt2WVEz2aaaB
QVmoGZ32QNeZBngfFkj9QW/k0K8UKGZqARpyQtO3YvMHwNQbMoGprut/m8CtlYthiaDPv9i5+b4q
5CBNq3JbhtPaw6LQq4fDSfaGQy9Yj2hNAH3P172u6zWcHit6sf+U6g7GAFRvF2Y20GnWz/QMXaLW
kfELuaAw7ll6LYy6mNGRD9VEmzGXlHB4ZYfdW+86YLRNfu7CkG0k1c5znkiC/1yxda8BlxKRUeVK
AzuEI+BL7QcxGLQLfl5EfOMjywL8OID14Tszjgy57+ZPLl8jXhJ/A/sw1CJUtbyRZhb+HqMPRaFf
Pt2yhEJ3KjIv2oD9EMYW8etanU6hFZ3N81p1xQWasZIqfdpDLCj0KNp27/pjrUNkVMSCuev9TFh1
cav3dnmFqb0EQb9PJjLS58hWPwk+duZ4s+moBCNcTjgN4t05y9WJKKy08vVFfSHZcfIt5HcAdyUy
n8jDgYlqlFESgsjUe4U/uh/IqjWYqcb9HG4UX/IxT5feUHxeyR57XkZjjsQpCLMrSVJIB4t6lXYG
aRMq/0bcSj/Km0e2Y1bVwLS6kR6oWplpBXWOnrBlfHMo73EleI+f/fqfFyAMncIhzr6GSna195V0
55vXj5+7diQYLzAgEO/GiwGlw7S3iLRgreTVOffFzczzJN/6jX1DTj3a0KBiMelE0GacPY8UJRAg
ZQ49mCn9Z3DmD7OlQFSWmo3/PCwA1IIzHBLOrBY1kNceRIpKPCjImuO/hLYdWzawQDg2m4jH5O1L
agOgNWM96VWULNT+m6L/a4waZaSO1pPjaBlWFI0PpPziBWorZnJKS9LCu1WtWD1jiZYmb0w/wxi2
JDwCie8SWG+dX/DNfOjfIUjIjksHDQ4OHKYAqfpFEapSD3zShkthsk+gUkeV+0+Pj7msfsopSrX5
6CgUIE457qCyMG8PQw7GUUZNNcfJuJYR9Lg/MnSkxH5Piqaw8gsrcf0N1OkCEzJua84a3mpaxwhH
9ckjKumFZGAz3PJ9lieEPXFcI4vCXrLGmT6cjypgevVyzspR7SpHsOyXCdcHBHazSaBZ5u8W6klg
SJpSNTCKed1CLCbDHqTPvsUFFJtd6SzoSmzSdvftei1QFVyKJ68wvvCOIuJ7XmTWUPVdJOPu8tvK
QtSQ4u4STP8ARcBN1E4N0Xckc4VZNg5VlK6gRol9i0blKubug6UTJXMjm6HIMu/QSdGwGSJOn/JL
72cgHqMuiS70xY9PWURH50Ms9qzb8JzPoocghOTlFTalnjIwO114D5N0yTf0uN3cykBte4v7oAT6
a/Nc+lkBsVnlexMcyDsTKOzKWfrX2S2AzCl7hKURPdeHQ72+vlaudg4Q3BbOB1KWuwegj/+9Uioa
SmhanJXnk5yIW6Mw17msSUi00yC06uVD5p0Ij6CuHSDDildkMJEUB6hxoSs7y2/Y5sNbIpaL+DnK
doO0cT3UE5YRxWKoz5KTWpcYZc2+d1bbo4Shp2Sg2Hv7cc/dEmv6QEvwCgEZmXf+i62opZSgeIQ0
gxzcKaY/3H0Yk+4ouh2yXR+sPK06d/QhD1glPQ4I6cG8aTf+rPfKnIo6j+VwkzGdTBhDP9XqaunO
PH4bK0tz9hC5fIKRtbmVqZKl6DMZDGnt+oCw5VgPahyXWGE6vZAUXJ420JHNQsb5ClN/O1gxm1Ag
Qybl6dd6YYzhZovSpH4REHRqFLkbhTdrlUtzevtcL0na5eMwkd0UH0P/PWUSLHeOeDFvEHC6iBf+
Nw3GGzL6ZCswJk91qKRT8dqqZOneBtuWDiCA9L/WYHBxP3ta4PUTHKqygleegnTYr/su0keGojHR
OJ+UTKp/qK/Ly/69bbZRtMIAiCJ/0Cx3W/WyNa/27brbyRUUXCEtc1LTStGXk4RBN8dEeKUJ4bOG
A1S6iX04TTcdvvqn1OSp+96GTFYacHrXivoWFVnOHq95sf1k4tGrKOYwhZZUa3jEozefqAUHgZ6R
eyW1pbOrI4dC76zqN/lZCyR0R/gyR1oNQIT0Hrj5k1DWBModC+AwjcpDpooofqL0j3eB9v7RvDw/
0XxQx7QalyfhoQU/giJ6o5+Bs2X+DY25Du5xVVhrdmSZmhlOEuKF1qqnprZrsWL6Wofj61j87lJJ
THDL7uMxWMD3FpJDtn+0M+3LkXOGT1aAZYjlBt4+27NU4ds0znXp+e4LYD0OHk7AZzNH4sL/+VON
rqcGAWH1zh1WCAOrdjEgNWyblko4Ad0P95kGYpqko3V2aNn0ac2OlG8KMCv3SryYXQct46HYgOn5
Xi9quq8gciGRbIxHHt06i0ZM/+JyCu+uZ4tSRIiXORiVRfnSvQBfDSos6Ju1hcMHYT8874SSaDY1
416si6fp0TNU+ZwJpQSD7Ip9+E+QBQrSSZ9dmpxCsDkxV8fjX5V/PAYkLbL21UAaYvthK4zT7ruD
NAUKfaMKWkDg26/+0p7y4iyyPs3KveV2uZDmaORFQ2+0eLyrrbs9nQ70r3UsAlr3lHeg05psD+fG
T4EeCd3noFr1VY/rCM9S8iTbsc79m8xvmlYonS7wlbDKHJ6PwAw6Nh2CF6hijf/vuLnbAup6nKL6
31joNnFZIPlxx/J4z7zZku6cYHJTrMKfd6IJpScmZhrgIkXNfIC4s7zOfT0gdcj5/Te3TTvTspHB
YL4sYMdU49DVlz2q3VTnpj0tjtMSW2Hxv+iet4/crsS6JqEyURdKwcZa002RREDeaJO8ogf73yPv
o+TEf3VRuOc/iEndxd0GYgCyEvYySmVs/iPZc5zkMvX0PogZYj331h6dwzZ0l17A3GqRAZMbSPkc
uUZo+oa87Mo3Hxv7L/4yvQxcAuN0eORlxR4tV3CQ8DErALEQ285PTXdDVUpT+yPPNELp8rsUR2qN
uog51TrYrydIyrsi+5pmJIYZjhkCSA+k4wEdvATcWf3jDE3R9ULLOy1Wt6agrYHxG5uGW2VioOfj
cKTra0NPfJK/bye6ikt1G0B6u1jYgXG0xsTba8yLfPwJyXDK0VswGECLKTI6rc4leHYvlu/+dtaZ
cVP8OWjgXltJ2sHFVqEb5zNNIOXn6T4RxyjKLiia2BGK+m/k8/TpzBrlpVfTMfcuL0bY14LAYEaS
9zX17Pfdu2z6HTDQL10aWSgGflVUr0aXch0483WyLSqh1R1oIfrTga5GhEyu64SZRWP+OCKWipAP
pa5uCejkWS1mMrTT6I5D2Oo5KXGP7nCa8rsljDEvdfcNBg6qvlokl3GXEb2OyAaZo4eSkl12bDZx
OYpjjpwW8QtPUBLbF0qtxiMZuF6MwrTkbrOZsNw6DRi/phQ+3LHl0ne6vYsZpSW8Qhilx9ZEPs7Q
V1Nv7IdDf1Djb2MycxEJ8n9WTTNbMgu6iGkRRx479/irRS7Z0GuEsz2R1ITGkoDidixSknFncmP/
da1BZDsQwf9i+p8W8rz4zMnHpWy6INdGvNWv2X1ViPvlyU+iRErEah8VEAuOApKiRuiFR2hdtH5w
t1/D7Sw0UZ/kTYLK+ksO1aUtt1ZinNReda0nKovaUgvQwqJ/GIWAy5rCrQsiCCapno0ey5K6J2El
NmhNNT4Op1vcfolXCgbPCigblmoOZXmC3VP45yd9h7MRbD8UeYT8YejnExkgDiaxNigSGQZZ/rdk
Qcg212+nOEAnwwxRIZ7PMSvxSNVyXOKmHBj8RSsfuODxf5dqGlj1bmcobaZDmO/a0nLohWlA+m5C
HFxLS/EDFThrpCu54gSrQWOuw5dvgT79hh0bbbUVdXwDx0qSu/a4drUZ9ygd/bEaJqd/p1a+SbDa
FdvWVOZZZFQoHZvUs4DOitWuLSZZIRdO0jQonrERvGYfaWFLMBn3Pxih8meQ8cExhcNNyidVUJuj
anmfJFVMgR9lXdk/M4QsLUvxm6hfOBZoYZiibfvirc2kvvAtMFYjthGIFaTQxdPhzH9G8iXQK9vT
HcUTmG6eVJU7KZQOSSYpd0XXzdk17kUl93JvCVICFAZ0ohwbOdC+JCoSNdNnzN7zMJXv80rr5dtZ
qaH66HCCsomviJqqQ0HYBA3VdpUx/VfkkUOZ/PyZzM3lHgRul6ei2+FghjjBjkXNKLuFWg9tWaCS
5YCE/+viR/gz9x+7qKSheqUVsx5r09NUGXvEfu8LBJVbrfyskgQIsw/qEi1EGJoh/Jc2cqgXknWm
tZk2ye6Cw+7Y6105HGodSgO5mhMFb5f2sk/z5wsKvkJJ7cTS2DF84p6EeviBj1+FHDS3SgzXqxm7
NfZpCYE/2a9fm8dy9bpc3UQNXVsOpWfUYBmE2HCnSEm1h8BrmuPT5fmJ5u3J5I9daXwSiFiA1P2E
j1j9m+jaye29KW3uvNUgseq2u3Q0WfC9zxsqwSzeflV5eel1tBeOwiAALRwgavWW1JRm/9xM/cBl
AH09LTfmw7eihwZnX00me7ErTvohF6VZcyDg29SXmlCoY6B9K2pmYu44Z4aL6wUXxkExAMcENbT6
GNeAKw/Qfx/fhW4U2TDQXURshwqhQMqp9wWZpLsEA0xrXV4g0Xi+b8Lo+zmxa7kLrgKdbAhKmq0E
ZpB5Ne6AMEyC0mXp2N0tJiUkh8EnrM+dJJ8E5tvaw0EBe/VJCuRUGMPq6LdyR9r/P1mYiC7LLgC1
iioB48gCYrHWRXZrGS/dYdJ4JlWCUd6X0BdYK1R2eUmOBJEZqbqfYJjtuSlhxz99zUz+NjZxFbWF
PaM2WQGJ9scGW6v4CevT656vA2W94gpaAjiFlHWbpiLpzEhc2W08GKRGhWyHzfE4nM+I88ajfRgy
irK8uAtY2IkH44i2pt9lxDkG9l8+gsuK2+Axy9hijSoOPfjOiRsU5JUdXXmLefjdTS5WyOeB46Ll
YzOoNRTXvNeu3rjQPcl+ZqbK8tHJQk98kfLlchGmIMxC/nvlF2qMh/WFLvz/lUHBfs9mZH8VaelH
DAvLZ3adx6WvfbhWkAM/MA0PvO1FNKP7WlQNeorgPGAJRJ/R/y7DKFR/+STmLcvRAIvC/iODPTyM
MX9N0Ym//cEROAh8Cp4RHyp1dBdTRNe679VgSJh6RaUNADXxIQHMYsE1G+T649VIT5nChu7OJ2WB
5+u1qqFh7XxreXWtAkF0Q//GrC3gevxGOeavBLRmAYMlqM/LttlzWdveyY6Qn39WJEZjZwwLUFHP
hB7mm9PacuCvHO8PfmNAraa4tyCMm6EVfmBiaLsQSoBpZifNjL7HVKgYWsyNguht7O2UjK26o4oH
9aw4ULyxr95i4FwhWGRSA+ze7fUVZTovuUF2QdXbShOC461g46EdCbtFdilfRSuzn4IAHTm61yEK
gxEaGhXWTBBdgjBmAwmJ/U1VycEpGOaKnUaeGcUhvdwHpTvz6qSmsiJT+1iuTCBMet1eJ1X6ASk4
pww7iQsxOv3qNcONbfU47J0zYnocUDtH+G8pK5XmHQQItGZkxvICW95/NIaTRYaieu6hMVwAJCU/
q+RyV5DUzFot9E7JF1CVFYai10b17SFa512dyfxhcWdN0VmeAc9kzrt0fxmGJN9xH6BKMkyheHdM
0PUnehRX2TxfaKJAfxSEIRIaL2B882SFS0JXvCsGKipLHMm9nFxErChzCyyIWU430UBtHjxZFqsV
SDX0oTLmxLlZwcfV/FjodT3nPTtGMDgVVzf4nhJXD/AGT4ZVPz9sOc3kxUd9QfatKHoWqwEdYGKz
9rEwePjwxtZmvqaNHc1pIkT4mJAbSP4QOZ5QlEns0JijJR5ctXC7TEdVuM7xHH3DtNDgMbToWqfK
Jw0lx72iAXtdy0a2zS4E6zaxMjvqUJufjY3z1ZH+rlXlLfUBkqn5CxP5eueh6AoTSCY07KUowhzB
JnN3ucqqKmbuOqm8GXJkcTyVj98B/doTggpWVQJ4EF4cjxPULVAMmxqt7NQp+QbWkTIMPuAk28vh
j8enA51JwkM/AIGp3e0ykv6tF3cg6MEkTD6GqrX8QVwH8qOYzprJWLyfECuEBc29bqo1r/rX08PT
yD72ULEPTNnDXe5cm6wJlY8bFX6Z2ZGytCTdKE6kkUXK6X4wD4rkYbKnpAOryWkllt7hnmD5sC15
A/UGL2RUARPV5TT+4jFVa8bqi2vwMKxUxJig0vEaTPNMeSZW9gUtoasOG/sBEYIrAIJWM/F2hCNP
C/3puHdp+CubzvZ1JOqMgYGpZwJQWbWpWG01eyyj1KIE6CafUBgYR2tBPmQyClQljEyEcw8oxbwF
YeoVGJ7+4pVQjNcij9nzh/grzmRUyOzcNTRJ3QDvqaAERfoZzIz/vjJA1I4LW9lcjMh0L/ZPy6/H
tcPjmxdQoc5Zv4B5dEZf0zWv7ePvospniuVztd+dhRdN4KvG0DxgKa8tGhRi5aEat+ByfLsjtfWb
L8LdGITJGIjpEAkaNW5XLlAA7FGIwJ9JQSNcnD8ktqhecHENKLdR/fonmgXuPR4M6vde0as1Jicc
xsYbllCqIm8OArRjmjF91ijOhym1kP26bcTwdOVdU/JZne/fHHC+UuPLhxWGSgmt+gtda+7lhVx7
r6ogZMpxrLzGk2JxjderiyAGIw4nPr/ZGl6TTWDjTAaWQNvMz00m/Njf8/L+enh1wKRTksk0weaG
tGjzqYFgOemoXx/JnZJqHAoNDzWxZOnenKaPu+TU0a+86Oz+v9MOCdfAJ6TnurOSJFM2jtUZ7Bwo
i4YKyOJn5DBGuwsC1i00OKjqy23Az7t7MxK3uAS3UY7mK5RtufQC4QKhBFPuBmIW7AymKpZXPaux
GDdYfmHUW/hyA3v9Ln2zNoJ6RF4UR7LXuuh7aATegNPA+iBNr8kYWfzSAnMZacXYsb0jAjfPxHmF
iPmzbzsv9BBhdDEbtZJmHtjh5WwUFY8vslyjZKJhYBAZl7GlkOsjYdNow22/lTICMgw/+U/7erMH
uzvReFclqaQCwQv4ICdLDEZf6YpAunN6lGnM0UfZV7kW1KxwJ3k6KLbCSbvpunCGyzinLh6dP+OX
e9sRaxW+U5BKy1kYVs0CoWdhGQDyUGuWZ/ABuCyER0wX6cQDxwpdA30JYkLSmb8v38QXDSRfWe0h
kAkis0JIH1GSAcB50ZAWVOFYCQ5hiock+OZBrzpus64q2Fxroqy3q2HGCPRVFFrZ0HDylYgZjnv3
QdVQdKyiZVTIamVY9hA8hQrRt3DXaGVw0QXw2Z5B4lXYp+cuCW2o9tHgIEzFGId6O9D15ttCp4b7
qaB4FIdYLpUk7/boaDTdGCDETFdYedvN8zDsodVpoM5Xtthysvqvp2Ah5+daEkyNd5VAkc56/LWm
sQALZxG1D+thT9UDCArJMrfqCrq0X3IH22L2nARegCwQA2n28BWrP2mYEVROVf6Mzqs3pEGfXyoy
LdGyvIooxXkTaK2uTrvaQwP1NI1quiBoHjaA1gLYWVbXW7tnuRp9NJNxJOFNHO2B7VkgKPnvehut
UqhoEkGriP62I/gJibCdnbMbYWrMQ8B5tGMCUe73JIkRWx5D1xMk0CKZ3MoAriNgiMVFCdXYKbwA
BEQrSCqTfYvokoCu5YQz6JKTuhYeQDu6AKQD7yDP3Vn8yJGSl999Q0uiYWJJ/FNXr1x/V/cWkBd7
T/UQnOApnSTKMog1iDGIXFWVbRELzpFLrzPghSRr9Xlo0IXzTIi8qYSQsp51u8Ca8GPUmu0ZELO+
jxgY03pHkjq5t3/qHlcRWXITNhMYlik9brALuxStviZv6DZl/0J/2fUrdCRdLlPQlwlNs7977jt5
XGYI3ZpzTkJR/BeJXhbT7Va1DAe2x5nvNvqNPeaKsAVjbI+BDLsgvM7TS3zD4OOA+VFWrtShpnC+
y/tEoH4OVjKPA2NPmk1vQMclegf8E9jER502kWYZ2gnxozD6OXDTpTVhEeut+TKWLfWXqX9UKLSj
PAb8p4JeXnEmQG2aAowgiiMI1acWo+X7A8LXZXYdTbA8bdEQ9Hq5cL3Dulce/EHWTPWV47zorpoO
PkK7dbXv8oHyB653aiZB8VMIQOVmeuFkHk3bpSozAcHTz1RilHAV17vE4ovY9923XeWV3AmXWbx+
GJKmISvgmwLdQO6Xftj5/Wuoj4UimGOCPfJpRPw2/tVMaG3A+nakvuCfDQDeHR+wv00NnvKrMjD4
Qe0kovvc3ZJqVd5XK8N05b62v4Ll0ynH9k2R5Z2X32MsOjaaFfeitzsYlFKX5FBHFWz1bMyM4fpr
LiglN3Sphaggjxmf4ZouD7ypU6t0iHG0iwTkxnZuWRsWIVPnLR//EsOuN5Xguqj75LAGxiAI8LNV
GTwN+tGsGgfMFDa+3os2B7Gr1I9f6ieWxZnVJCPeKJcZpgTv+UBhp4arBNN91eWWBAQhg9VTXp5e
RBS9zKB2vGt3UDZ8Hbutwdv8Ealsbx8P8dILKNZsbGncoqQMBamFuD3obWn65U0jKUIQBWppj+1/
GqzPlpF5aa7aHNaUlm5O0yjNGtrMDFPCEO2ATXu1rJ/zUBlE+0irIilBvLrRtfXc8WX3RlGfYvln
WfMjFx0cTLnEIGWlykNbMNgrSoatJFMo5t/tpcJnZSkJK/d2s1w78hDjlbHA4B9is2TYkpZCti9L
EWEGrEkPikTT3SqDDM3pLycyz6YeWzfbkt/T5u+EGcIecFWrkPt3MlmhtzGRo+Ks+TkQkm9qmdQZ
/5dr0wf8q6sR/lmjsLV+DDan2C7idlTFISiE5Lyyvv9xZ1512dkkQr4u2azQ1UXcnhUQVpb0jNJX
i6finbtIE9lsZG8y3A7wns2UtXG80RRJRUwVIauq0+BGA5y5jlqEi9d81NykPpJht0TX6bZkCAkF
XM4a50ZdJHGgCtccqntLrSC5tlKLR0IarhW54bIgKWIfbeu+wMIhr8c6faTn7mL7rjq7xJXawb6j
xa1lfbFRVNAmrW1ystqDG0pp/HZSgC9wb93IIS0bmw8iXiqz5C9/IOxczE8z/xAhpgwrxHS/KZ4r
yiPgb3+pt/lDXXOeSd4Ne6UVeepwfY/1g+m2glmrRb0WHst5y0e1Gl125L3kZSNhDO3+495VdKa5
PZPD0hK3dilhQ+h4+KxigSVlJiuLj1JoMNUpUp+WISNhvifISa1yhR80O2CDe/yK98vmG3T3YzDt
h3+ymul/a9hMMlH7sJDtkGE6vilXKBZdiZE/FdlA9vxLY2FVEMLJQgg4XiZdpqb7MJ2Qz8lZVWT7
MuaxANYKoVVFo7co6UjiYa9jGqb+m/i+vmP11M/Rv6xm+zdoOAWAbij7fPwy/52r6+S/SkVywcFX
ELsTSBwwoDIiTbqO92QBU3CMWMQDairbaWqcXFbp4SOq8oiC19QlPunPZmqFGMaTtNKsZGljNFn8
XhbckMc4iPTJUXljoPDUU84yxh7kwHBB3AmAAVZ7RYV4mgppGelbVqUIpe3IAWg65RDxPPerMkO2
WzMaA3UB2Z5mFm7LqQ3l2a4pNWsDbhVCBiwKaclbpukCkOI+xhbyS9UXGLOTcoObE1Ww72dcNwY0
nxeqUDFMo5oOwvHFj1kR6i2lxqcbxfyMj8XE1R/4rxnfoTXxOxZw1rqEnjEwNJrPDM2pLFKUPFlo
6QAd6ltELeOO3kMRYkDXYqs1fkOJwVLdZ1PBFu7VsafjImZk0mblGguZcrqI+IVy4pC0u8NAinml
wxUMKojCl+PZIYl0QkGqTVtRFAkTXLW7BS6rsGHgZJFgoNskQsd5U5cAfALSrKz8yXiV5LHx4B1K
dCTPMH30yE9qD8ftE/xJUe3VgVZni1/Nwdx7OjdXY8gqtVPBnGNFm6oosEg+DFX9Q9AeJKAWyurl
xyb+4tx7M3H+cUlBSOHDGENT4FtQGYqp4cR4DTMAlAX7N1J8ETsj0+lO38v91ckLCNIX1Yr5b7X1
8x8t1SvdRWYC3ydHqzEhtTJxgHKkIhRmzl8JnKJubXt2MZwMkda0dCx3shY/quIG3vYUhc5gxVgZ
J99JBNGzQn0T7xvfc23zzLN/0BQYsYnYkuSE+jEIlJaqv/vRMfKq4HPQBIVYTYTqFZpnbHa8X4+s
VHJ38qnjS9mN0/R6zQT/yLjSvKQ3Vr40tJ0ItqjlDtXT8Mo73NiT+l01jRsJ3WuP3+aEw8p04Wue
E+LeO4NWNaT8Cnlv0Y4MWCUIJH5KPOOSoebDeYjmMn5jj9Aqh+f/yiBQ/5/+6IqFXIC+msQWynlP
Or2GHlr4tlq8i74Ja9kBaHVHbyzVwm0y9XqjERZjrt18+sRpWveWIhdTzH6wg7/OR35Fr/x7nWG0
mVh0Fx0T+utxtBFJITft+tUAooG47Wnf2vVYqlobgc4wz5lHIm/RDS4DxET4dIfqQG4ht8RbxS/9
o+jRe0jSMWsiKh2AsAjyVWCQm7D/rNbtczM0+mfafEzv119wfoNDitxQC79c8ojGq+sGSUYI4mhr
WMwF2dybwc72l4a50EM4VxleALedZHknvBP/MfK5LbHsDmKODB6RcxTlAGza4ICbC0mNwukRZxsD
2i6/4t/W8MnNEf5I64y0TXAHias3rKP3FgnVOkgGcGZxojpdwbBZFC+xax408wY+41jYCCq3TNr6
ve2y/oeJu0strKx4dJmKVL0tR6m+deJgpe+zYTB9nd7UsziA49rigJsWUuUEP0jpFp/XVue+pIhO
y+b6sjKb3fT5UkMssKNpUOwGeD3A4HRu6+lOEWZ+CpXjkQ89o8beb00tHe+9qa+Oo074S0BJlZcG
feKAm4b1JWakwIyUwOsk3Zof6p1wcscD0zzzmwmIJMI6xg9He8xsEc1mDnWuXC1d7eX5gW6iVxbH
7EPNAi2oB31CoI5Aq+D6JhMxZIRjYHZLMurIhNbPI6VrsUAp8w4M2/jP6bh8Qj3CzIvNmt0tQDPL
cOQPbSrKgY3G/cdxYWK+iTzFXwwIBGe2mOkGbuUnEm39Xc03oJ01ibr8AAIMXaH5H0SeHLbnritY
MVUPgEY1B3h7uagTtUin9vO2Aw/V/8Yz6hHXxoXUuw+9qGIbuk16MuGyhQdaAvO6yJEFha0t0vm5
OxqY8CD10l8SDRIaZfn1HrneCMlBmGqBtTSHFzCTopCJ4oGIovFB68kvoTo+9ao/d13toW/2grNi
oHuI3JsnYwrd7+8VBCtSWEWyhMylwc8RTDxrT0kjhQBafRjiDeTQMafWpFujuj4B4JBVOCGsNiJP
+cTqgMd2AV5pXigx/9XzAzbiPww3KFGE4ashw+52TxwZCY54gAFesOgeUw+fzMsRHRukLj2poY6G
RKuIX0CNBncFdOgjuPeZ+RDHMiT083aA57bB+0JDRJaQ3X/IerXpjw34FrqfRmLWv8YLWT8Zpt49
nZHJ487B3b8NBwpv6u6CmGXIK606YgfyQJSBTjPskd9igQPobSTzNZ8vAaz3f6Iyop87n6Nbh4um
uP6/SgFBgWWnUYuifVjn7lJv9U9DK9RCluZHN6kHK63TUajjV/JTbL5ocS2rTMtg05hNsdwAxAW7
2UfKoUN3diKED/5oHahNz5zXtMGu9yn98Z37KzmEz4oIYkVA8/7lxsQO7UhcgyT1/srYONrnU0h2
ZIKzA0FNnhzVvSrKBFkou1gAWU8hKGwM919YzUHPjbtz4fpFX/qxTwvn4f5PUAy18fJTyDeMqrjr
s/eo2lCKWKUsafIGWBDe6wj2EpspQLLkXB7il4jN1YoJpUzDICtP7kByxeuLWZuaVPDOP3V1RK32
KHMmCJLk0/txY/aEQlZgEpyjD71ZVO9IbfWKIzJysmPrNub2+Zi0eYCon+dv2ebk/dyhNoztCbqT
QpgM/hXOIACEUGfysfjqfvnD51iW3C6Va0N7Fq8yclXoSqy7iCtxiVgwU3VhnTd5wx9OkzSmyG/Q
0+yqvfNk8m8JN1B7ctk8Y60RGJPcKY7TuGBW53Tbg917Byvtlai9TrhC2DWXPzlFqQ5W4liMeuDL
dPAPMzws3HzgQCsR+KWvx1F0MDuJ3tPJZhT52S+1b+GnaiYv22Ig/wwZ+xMT8S3ejPJKld201MFf
zzwlcGbuo9NI5dsJzG01H5KL18jvF1y6zGoiZV+80eMwGKc9aSQTOMaY6FBTqfu+bOgav3NR8p0D
isXd3z92neUZF71e1tE6JZRBra/U4FFJE0rNbIgn5w3YSI03ZfMDLB5OMi6HHn1abnaGLETMkTKj
EK5O4NnOVUf7H07zTaoXlUvQ2B683RFaHS0SnHif0oOJJZQivS/iSUwO+dFAWblAFZ04iB/I0Pk1
sJkAhixPRbf7BtzHqhaX8uBW9SaN5vbdTMLCgaLJnSh0pEBUl1F8Mkh3nGFE0pu/AtH7tKWMdKwf
A6NX47k0dfaqxy15FophGnkJi8h0zFCECaJXu9U6ACwKbzMP2tX6y80sXLwh5q52XWYHrhZemRyf
q31v9iCCANIju7b6kCoCkcAD2rDSf73M6yJKCdB+TDQQwYkWlyeZ5CIrqilH5IqMG1YZMebfpML1
rzKoJd3QAWfnEx4CF1XE5QIa2Y3iSpqSlubgNq1mj8rYI6o2jR0C53zH7MyZJft3e0hXnBjlTgvv
UQGsffmc2YHYC9+8o/XXjBGsG/B14ngAe/0pMbIPYOiheyXzPMdipNaMlw+wAOe45JRE6kKfy4D0
MXOrFPAJ9YCmcGg/ghFHW0VnTzslzjtWSFI3ukRe6GN33CDRPyNRyOoaowXuBi2O7zn5I7dZIlyC
1VrTZ0D2yO1XjdVst08EPXqvUtOIRYUu7dGyqNIIQhHBUxLexQDSPF2eYtCFnLalB4jWX8vlCdCT
7XUS1evYtVSOq31tCmPOkdTN4kk7V+bUWrrp/rFkGrHK9btu8/19LPocR8nVGMR6bahzHNcLXwud
i9RYXYHxIlP2eFfrnF/Bs4J23kkRl6cZhzlRV8Scx39lr08ZPBMZ8PHzuvk4Bw+KD7G1Zb3lC4AT
8VBR0RSBa28ObBp2M9zX1FQXKTXKxfduxbwYDq09sbR2lnzWHXGVcpf6IvIQST/jD93frcQVwWli
RyNc+cJm9xYu4W7HwV99wihCwa0PrplA2jI4vvhI1ItOV5vQHiWE2PolAc/947yPJvX8mNwjA5wN
83WaLLKMLtmKEtM86lfIm7JmlKE4tg3qOmC2GGeOmsXaYr1AUAuq3Lk6i5BuunTyRXKyT0Y9lp+V
MenvE2MyPLICTTR/5pWkelv4PvW/RhCAoRvL5UQcMgFVzY+rMOeSNxtDkwCmap3PlvBwDFmJzz09
jSfBwbbJm1Vc6c4jkPMgvKyzH2d/HKZiDE/+pG8Hew9LgQZv3Y++sDKK86tsbDuQDJFpzUa8IxyI
KcaTYcHWG2JlGVZgMlHSaGpjVEqkeh3DZ7U6mhTqNGitWEif2CquYFPHUWxA1e7eYJ0ub6iflJbp
y82iD47dGGhyQUq+RDu8lB8S6+DXhxoKzWCa+JH5NcVo0ilzaDht0I9ABVDKEPkWOWilcdulBsYB
k40WhRjBbE2qycYm7Zk2u0Wr/Jy5zd3+KETOd/nOmfmh9kMjHnDt17moqo31wJwGHn88TAiD9p+i
XKA6xxjqlmIzN7CLsErLO+w9js8d/725hpCR/e90U6jNC7TS1/hpqlayNzZ303FL/ctT5VTphXRz
sE1DfHSuc8DYVYAiCz2KTCEmzmdSyLHt1TWZN1EKnmIGMjvWyArerszd7vmx6F1kH6B68YDhqqPb
MHw2N0Md7mCAZas9juRLBhBUyFR5ds2EL2DaZHLuF7v+DZ8wReYlodfla3TyGKhCbs4jVF39ctoZ
VjSsoaM3fGmMlQIbLH1L11XHH7kIX6Gqxpbm54w2fFDajxRaPnRVcYr70EgKFTu8v48DRJvf0+Fp
ggDkU3ao5mBE4pOcuckBvvgJPURxKlqsjV2p58YYmTwu76HJ4hwr/5mULhwDr/kPIZRLRbYyVt00
ja2IfK2Dc+qoNbbv14ojtKdD/6Z5gjeUvCogJTsjOxc+FXZ8Gq375B3BaAvOp6PuyXrTUcQ+y6vW
PHZKnVIK12S8jhjpKeg7KDZ1dU8knRL2P3Dk5EVbM0hRMkUiyYjorU05S3/gQsKI34B2sexe2XOl
VGonNOF+qJr5eQ/brto5JdMoPzJvrulLoYEoS4fir1EZl6pFIB8cZUgFnkXTKW/miHQxExXvJE3u
4Jf5WOA8p5KLXoS8UP6uMoJfYEW0i3jVT9rUGyqT3iMoZXay4Mq3/RFZDyrl/vczNpD+cBPk/R4A
CGhE1nGaZOemdxbSWPW97faE6/81HLzZudsdlRG2t1ZrC9TINFsq+sIz3nHeJYRq+YlPXfQZPVYD
mGL/Y93HJgv8G0WO5UNUkVQikCTY92AlTGV+s52/EEBslRAwGr6BOf69oflFy5XKmqg4vc70fobY
Ac3V6D6mFbZA+g78eNL9wpTlGgfL/6h5JdYRquUHbF0bYt2RL75+oncjzB9f/Uld+4m+gp0osLhu
cp4VfEF4V3hCrd4ShnkHaWHQ5mzmPgMzisInFYQunNe2oWp25lQAu98l5ZGoXltE1KPJu3hllYe3
I5HmDttIsVhbaGiIQv/gZvizLjoCZQ1HHy5wt5abhKcXij8aneBd3PhLKnvB2v7YKfQHQzP2ZbIS
fdE2lB6UMi3BL73OqeMNT3AGDT2+lbUgFdP3063bHP09X+rFRME3NudiPwSAt2VRvwCjvVK6EDIY
gI/k3YoZlJmu4BDKuTwUI/XnBvZxqeuUj2hCMPy4ez51DdTcWvonR761rFE37gYKcqFZYOPwU6Tg
InYwyg7Is8HJZsPXJPoMhctsf12jDXrezSh8D04zdAIqqYb6jc8Q09Ylq494OsRrolzRLNRgjIkq
3sxU/HstFbUjOlIwqoo2XiyaiS/WRIrqeLnqfQCCdSHHjYDAneimnnU3mZo1okGcd48H4NgFOQdw
3QSYEXuWYJSjDzh1vlSTDbLw+aPdT93SOyJ0T/OsmV5NWf8hcWRTk2ogorcLNHIO8rdWbN09QzTg
IQhe8/PbcB9VQax50kYD61ouxGntkv9aJUlyTkNw2KQ9iS02gtFHAdg7OrMYxY7w7ZiJMjTmD3wu
VsdJjC1puHzvv1bsZvef1sApbxDSG9CVkPO3AuqDckAfgr84/xoqI/L6tgKZq+2WMx33LF5GCx43
UJZ0tusrXSJrLdCKkzmz6fAfBSelknFXvYG63U+gpXof6OoQ/ltrSdXHI98A4jWtv+jNc3239ZLM
dFzi1a8xitn9r0L7z/X7MR9giC7BNi6zLPZst4NkonNcXG3rix85edmL97LY6d3abmo0VBT0Eowp
nZlMKGRM/SxIf7WXA2sUChF1pQlk0/Mji9PIWw6SidtEhcgJnKjwlAWKBz3eqRKBaygxI0QRek/Y
J+sCDsWDkwRcQ6XioWkSNyXLiGGi6ry/vYTasKC0TDLH/I1UfLhJhi1KODkUnfKdujfwbB6/8x2p
GtT8ldnILP6QzlFLL9XFxhwmudOUZH8j0zF953gtlPre+SPRx7tYY7frqhdfMYtr5WLhU42dDXMd
u4ZCqkC3UJDa+fxQUxWl65G2mMlH3Cak7zuuKKfmyQP/OFR3h6mQXoAVIqv6ELyM+Lho9dseJrqm
7vtnC0jOoPqglEuh9AOTO8ehtWwe8Qwd8SuFheh4xk9F1ssCEJRYUoxq1ir8xNAc3iOP5uU/yMXo
Gw4MK5rPoPtKjJDI1V1XVJir6BRrC6BdbHcpBhjolSAQmGiFyhm9er9AVm+nsjsJzaIE3SquDruv
mrBckss4f40XYq5e2kHpUbIiUfhsRQAFjj1rdaiZ54U9gE3PZIQQ2e5XYd6ocZXXPs6CkKWt+1ab
5uQiSG13kNwa660sziu7Ue72Yv+zTuJO/6IfrM83MQiZE0e9H0zj/BoGgpSNj5RpJxXq2bxxm/5U
mD4xA1PhBavU6+BiKKIes84bNmVnYtHvkcDBMYtUCPhstCcuMU+XO0CUUU+AT4eV9ESuUVjHTMXE
+PawI09ykZ9ZvBJO24jskJGjQ9iVc2iC16pQ6pfb9qaoDqf3qqlSuXXpkaPwqrPbbMu/C0UpUtMJ
l5EYp1gHabbkwmG4GyHt+WRp0WsDuVpG0HZYuyvdENyga7jP8aK6P+uIZClKvYbFmzzwMQU13Tg0
DKNodltLR9VTIoYARkhk/ZOJ+AX0CTgkEqqBLceDv8c3sxBda4Kx2yMG5rnLVRMjR6QhatK6N+b4
ibKqr/kIIpKMxW7sUQSAXT/6L4zrlNLUD2+0eB1M2VsovtQXC7XYpaYoDZa45Sj8mNzF1LXb1VPb
3IzkSOFF4zvbBz32fLw7LI21a16PCp007+hknW0H5j5x9tC6jDRUUOYPjMbITfJSpi10I7q3QfDi
3uKxHHqeGoI6y4YlsNe5GRQPDJRzD2Q7HEhh42GS6GFTewNTABWdvltQzUTVC+dQ7EB3QeXpX580
ORhR78pAjb3wq4Np4pieVNr1hTkQWui3YMwrw49CtI5ZShhuYP7OKKGtm78TMY6LfIn6CGPY2n5G
uR53FafFYXxM6FcVvkFcUoonpCUDPcbV1FutoBHx5GhDUTLZ/d1/49K3Rjtq3pVDfiLPLnmhoqV+
T3clBODryFuZ6JlaR81sVpU21ob34DGGy3RaYebXtlFMFhxHrVTIs6Sq3C6IbZ5BilX4UPLD6GVU
MnYYdH9VFQ5UvwOXVLngcUooGAMZi+XZPsEvj3kAPDck0SUA70aDXMmTX8HATrUi8PkNa8yL9wDg
8YCPmFE7oX92HIeXaykCN9Vp7zbsH898oWrkJ0LB/AC/m0z5dR7xCeRzX/Aob0FVQHI9ro3oksFb
0BpvGEFYA23/KXAsAObCHvWOm8XBWkP7ywem/r5to9/0Tkq7Yqv90ekM3fFdhK1Fi4sT9hwChk5G
ZRSilbp/Ais0+AjqGYcchorR77gK7zSNXUMbVHxzhZe3I+ewfI839uB7CfSKSG/r9c1yag+cDNnW
7oWdRpbHwN9eGBYOKeaBq7cDDpgtcgJiGwO/Bf0rQiW+YxeJhvD32iEnLJrViZIWs7Ewky9cvfY0
cvvnpWFenE0HQThGWnwRNk6fVcID37zrvg9/f+SrH19kxr07d+TcWrAHaBBQXRHO0f4VuoLpnX/C
JTaI1s6gArz49afOTc/ZtphRU3rPdcrqThEvfqC2+RxSPvco/VOgVuB+IZK5+5EL/qzi6FuY8QKI
0o1IWwlTZrdkWVWzhCd7LqnYJy0Z3NfpZFioPqPApHCuhZdZLwnd6RzhiHfyTEpu6D606sQIVpsJ
fZmDm3IMjOubU/dws4vlzAsJqPhGMVEp8ujoI9HRNLB9kEzGet+kwHc32i/z7mmjNzH/RirYLdYq
Nvqm8NzJGZOh0sv+SYXuYXWQ0tOYqK6jXFj59YH5as3kjya3vTb1gTk6yBHWl+7B5BdLee5caaqd
Af4Jx5IpOrePyVSIsfit4Ib5ZWGeH6get7SHka62ds3PntQkOhJ49dXqC9XVngCddRSL8UApVv0k
syjsH0GhQWSed8geIqfdAft4Rlse2hPXnZg3X/CsVLU3Z2jMdm3LDp/+Fd2Z3nXymrJmUPargFoX
MTrPKqgFTeXmWjVxIzrDZMl8qYrn4JVnhI5jMe+Mf+fuqmaSkyVXV7kbdnsrvFqPFw/4cFFvLWlD
vnz6Tax+pWigMfTBigyD7/9KyHG5XfLeTuL66HiqCysbcRg2GvU1uD5dP0v5a3iayf+CwSV6RIOT
XamZriVC/Ws4qxIBMeBMY0Q0ic7RHH1So7jZSc22a/GdR2FtxJeP327LsPe82FDq5Pdq55VbONIn
R3G7xbzcr2OlQH7EnChRV61IHhCqOkAEAkyED89X20ELx+fhMKSG7HDaAKoT99oJ5HTO2LSnFXaZ
4ShhiQ5lR2eU06ZWgWr0qt5LOc4QwMFVQyH466hXDMcBRKheGdR5Jjfw61kq5Ku/zv6PRXjrT3tC
3/o2X5O1hy5DybzElyawp189oss93YSVxuNuK7dstPMdW7RfH5rOuI2H0mdB9OPtJ1ojHRSZ6xmQ
CULjHvmfS31/crtk9iV9a0c8WfOB9CWOqavlp8hot/dgPEGCpZma2d0t9Ll473z6ZuTdP1MFu1N2
ZUOhnqA5GcJoFbr/UZ0TU6lQHKuy6FCpWqEOcpM3wIgd9DIvPbkJYv531N5i3QZK6l/VeMhretHG
G1igFZ9ye3/oMRr6LriRuR1Tr0I2CCoojpGpnIq4nxVlZ4tqJa4CaabIpEzUMbAnCR+8KB3yreth
4kxSth5LjOHgGB/94jbmOc7j3H44P/FfdhfV/HR5DN8IR/rWDTOrZDYgPPDPwFgC+Kct74hcs/1f
YTWy1vo9n0Ybaib0LaR2Z/izxLkiNV8BiUHyrQu1DXx629xDr3IZY6jKnKwk4iX55PZWpIQKkyi1
tqnohP3KDn9Mw7uD/yBBiUI/tzRkhRFZQPtQxhzXtQCTi+Uya/uLy224HwyM9GRfTgppOqV2RPZV
b8QLq/WQY5eE2b4txv8EI7BC7xBO5Rqj5BO4RZrJBNu9bEPjUf9Pedk6/LVCdQz0CARcN2qMZG/D
0PtGBH6PDp+sfhJHw4TIcQtmKx6t17/vCOCiVVSVNvadeDBjhpgZhfZDdKENLt7o7nh6LxKSx8AH
raCAgV7HS52k6T0Kus3b0UC9b1wmmDVYyawKqZuYAZ3MonryIDGyLPZpz9H/IhACLZKXtCDcbRy7
qkhVJ5pL6nkCMQLpZbswNzLQ/jYEh8OCo1geygsuqTTBEBCVPqa0PkQAG7Skr6H6oD0AW83yl0xT
N5/36JuEegf0b+rDag5B2oYsOdUFVw6IYcjTHJB5zOM4TiP+O9uxC47d4qlRxRh4iFj9zmkTMFwu
xjFmXIkYRSBPKbYZcCGmYP2maDytqBWqPfBWNm1cdyEECwkytIhKdEogBnqJMwkG6ywtzSn9gtbJ
NN9GLz5w496ZUKQpz6uUriXxknuLk9M/pHgwwi+T1EkUfHBc+iWy9uL89VZCMJI2I1ZerjzR9yVL
t94Lx7YHfc9Q+8Ilp6nqRBGlNGCj96xrNDbGE2wRQU+TDngUGs/Hl8hTakqQF1Pk8cJj193aw9vV
3LB1OFf7Wv8EO/EeF1Z7OW7k26zULZUOczopxF+EC7+iNgjIdMl4rsFXue8m8q8Btl8URowGeKzF
isbLELWIuCh0EBnv7jR65yQeIJx/YQoScbBHWWvsOpUSpDP2rglAvjWSH725WYLY+cOuc4zsWn/z
VDvBjfAdbrAKc32NrJQZRmE5HtZfZT7CJ2N4IKQEEs9/OL6YP8Pur1/oawY72ky4qYffbvRTYLF+
vmUQy4lj0XIhvfyybWXWJkrwlJ2rvavCLgSmwbyrJVwf6lQDu6nUAj9LjGy4MetzoXuvb5atIpVK
82xVM9o4onlfCiwIzdkBg2AOg0FnPeYuYDQwQqtyL0Hs2J2lZnjYwVhMeBv0RactWrNTffJH7Z4O
kiueQE8pAebdHzl+qLhjMzErM+o7q9RLhP4NO//755ZeLTemftgwJqdYQTTT+E83vHaHWbXseO9+
NfplSTsqqwfTkH5vtNCbn63y1hICFkMVMOwaLCp9Wqr415Ory+13f7bF+Yesn7uOcOKtzGTpqrFM
vZRbN2igH6kLXM1YWbx4lVxknfLsDX/Azy096XvN5oZOlAhGYuV+1pvV48IwWdAmjPjn6YPieTdk
lIINSWGPxK52NA+sdx2joybKO91Y447Beg7/ATl2mBy+1TJcZTvTZfZJ1R/+a+4NBd0wSKq61Y2s
VuGJnSBbU+P3fb4DnyySEYduO8a6OD5pPaPD2gti5jxWEb6A8SZB3TiL5M00BUpZxMpARFvQDrVA
6dOLSZLlWOTf9wkHhb5DFe8LeLfpUHenA+qNzxS1TvMhDFPqzCpOjqDQ4BFw/CHU9mYQQbtZxJQi
pt8HcfzkNC1z0bJ0c1igq/hCYKt2JCayLJzIE+V1LFpU7MO4qFGH8ZDId5XJH12phxiS67m21m35
TutnNsx5j8v6UNZfQDosnoBdyY1oZkMAeI1xx+ne/8/0bUhWSnSRik6cGk/3Hu2HjyV8k1++ZloW
UyCwwAs7yNeUwi1yNZeLihGDs+31w5ihPsCOf5qgyiRDRdGuWyngtQIttDzYuYjY/EdgeQwXJuzm
NQ4PCVaBl+U0RwCLbqyRfLnsHZa6LAaQIRmQymzNcHHXoCwaEjPgLVFU2JRVmxJlg9Tq8kkXfbYy
2k7RVhNbRl/1gPd7I04+1FkMHniFJfI1gKEiQpjJ9GgP9tS6d5J3wBbUuIYrc3n+q8q2siapTlGd
Kcn7D35+dHIV5xhEVBNcVwld1LwRxQMj6/AoTFqyDfaUbE7RB+aa3axhCa+NzW6h25wDsxbyZiIm
sGQyD2QGU/LHGKWxCUTyhl9jDgTjIUd9phpOuWcpEBn+FWPYwYYvZpfvT5k9p5SKNeAggCC+W8Mx
tYN3mB1Sw3i2vbLmZzZbj5Ty3BiU058WIM/u6Capt4L0KtiF6qBgO5F/e7vkfzkLuR+MQaRx+ivB
UB2Z7TaBc5dfz2sBiSAZQEzkGz+mXGIYqVl3eMM15bNcOxcb6b02reB9FIzDlEVcmuVkrcJsObAg
w6hHjL83USMMs+dG9bcXfFYsqa8yYDnUpppp3Nl2ih/0ISMACL3jlVBZzthOt97xBCkXw3BaTxA2
iKaGlLlHpjenRfF16uYMgqHDQ28+SIPqtJ3CfxOoQdGQ4Pr6RsG/fnE3U79cj7ZCuUyLT9AR9oai
FRmnfoLunYhNCO3SAvUvmBaS9q1vy+KNPHVGwmW03zs9ftBVWCFkLCGZ33OlAMSbCD1kuJ+dsugT
MVpHOp6wU25UiCnT9CwHKkV9lssfXpv3Y9DGe/kalloLMG2t+tgPpee6rFUIKj73On1EkwLCe3PQ
cT+gd78O3qu2UbmYzRYJgHCwPeiNyLmw21BZAvHYp7nlHhmU/0kTSyzTaWzYQBnLKK51PZVwSWJ8
Cl2OBHYqQ7x6jCBH3HcHqa5beJCJkB0e3ewh+fG8Foy8E1rZUGzOgr1BBGEGq43GvS4o1Jl0dhem
xNhwJWOadl4T+LysudOyN+6PS2LIbN2MxvH9MKjHHA3jnTmr4/wqlqQXsfgaHyAzjMLhod6AhuKG
F+H41oibd8CCqGMa084MfcRm27jrmJg3ioVXjZNOvJI7K/ejj0zbnO+OQOv0lAPqgnofgeAwXbEO
jRsG1kyU5xNlUt6f3ErQisFEx9NdYfLwmBWOg7xD6sF1aRK6qzZlCIaBQD4WiWLQMfNJ+qdWJUGk
gCFT4VcR2ucYXan1A/eJKZUYXp7rcvYi8GFkGe85GktBCQeKmgyrmDx0TOAL4fNIDa/BTfFYlaOM
yukKlzeAjhahtJl17V89fSXm2rSunCoMg/DpIQzpYEZ1zoDeVV+wRJuZ/EaX1IgeqP/mcbxBOvvI
4poJmcQ/AajqIYgFZHm4O/Fa+QMQGB8ngvosMcTL1w6YPH/mTEVd/t8rCds9aNOerTRMLmyegkNy
ZP8CnUgobi9D6PCjXETkvnkmcVe255yXg0zQu9oQt+H4ipkFCgF5K9zVjlV/XHd8Lu50gQPZjuOX
1SNu//XcyHSArM8khjXj3ipCh2EPsjRZT7sVNseDrbV5rB1LCdT8d6ewSOZVaALO2FbJMz0bPwOE
K8AcCK4ghC6LBsHJ3ap8CjqoBVkVgsLBojP+4/8lF0rABG3jIFiBsYza6sbNualFyaRBUT/9SdpE
xmXWE3q6O0jJhoQPrZD+tErsVddpNzbEiiSAyJf2IKaz9n+q6tHdUO5kLjY/wbpVpyqXQkomLLmn
eYFdEdmg5+cfEFVTr/WorOCeJiE0TYj2AheK1i+A5MqdKPPNXM9xndp7JS1vvGekX/6wzyBfRmSt
yeB48LKVqwZLTxnkxprllObgInbP/dsPdD9hvD0C8gbyp2we3ueE7sHWHccQHsNixZZjdyx+yZeK
QWfM/hef7+qXLZVwxiRSX+fNwHHGCv4TZtauqyFHiMRiwtf1aXtOm/8s4/wJWjchtN5u+5hSr4UV
7l+A6/7fgp+/WW/m13ffjHRJ/Lnp3H6MAgLJDaEtS2ZE41Ba/faHmRZAFnRS9pIgyYy0FqlADmNF
eQrNTCgrNNuZQq9v+76bzhFVnkkQJMpiU3RR7qnXufe/LppxE4my6t9TJySBfhBx1IRC9P6PYd5e
+OtW6MAZCTHDUct7ODC9ZrFhMOe/9QO1VEr/lEHfseqaS49qgQP9EVbr0WO+ZFO+FS63hxepOWtz
7s+lw0pyjCRE+LcTEAtHZoRIERuC75UAsvhLh4WE1tE0uZm6/647dmsYLpDnnJyVdILLoZIFoMvQ
/W6+TtS8EbzzjjNCsMya6DDfNhBsJmBwfS59zFP61kIWOvGVAsjz3MYuDLX5Lg8okykL8bQpoTth
0/xTK70g0RybZtdarNH8CkVUTad/33xhXEFHWE/6KiUly0h0EIPw5f3QmgeYDKK1Xo6WYDDd+BDr
dCmYyg2Y9dVBiOypls1oqXr3TumaUY4+TD9YLO6f3hPqpgL+OQ52MJPFyNsO7OoRw+ktIOhDnulo
fzTixteNP/stuilREw3NFFR+0v5LQnIRXxqLktmKI/aVGrTpIvndVydi3hhkVaexPcVLccsLU29+
nLoUu9oR/5/0aQ5WE6iCJVTKpXIX0QLBuO372kRcHEEZk7CCuFU4jkrEpAt89Y/rshNYzf5g/2yW
hIv3CH1GIFXqgwDVJeqA7JyuJ6JCoDNizKfN/HzPrgWFJ7zP7orwCZYkuSPYibTND74FsB/gAaAC
luafbJy9vDo5gkfusCbn0l/H0O5alSzFQoiyxn+LDSrFzrYgsc9xXLLeFTsYwBXh3ZNnscBihCB5
lbwCiyQoT46O38ghYGHczJMzz4UxrGgdzJ+ixI5+kXP9/lqSURAdIqYpUji8FhxpS8/6sV5LM49V
JsNLJA+YZ6NVWOlGqIDzf6Bhxp4v/6uWVsoR5V5IDuMulcpn1kQLBmHdH9RQga1OOT+8ZvLGO9ZM
4WbLMM+nbcsRyoVLw6T96++9WCdP9JQiRQJUiCXN42SyNsg/jYmyDeaX7t+IECIxHqLM8NatJBOh
u9ezcJv1kgVyDGQJqoDksNnTHqrE/1vXAnbt00DpdFBoVJ7YmfNy+PYpI1WMnYD9iP31pZ7bZswv
ccaBuGy6nMDljoqTD2c1U/Tjvo8i3Cxy4CC+ENxpHMv4oKdrEJ6i9M2RFCeipa3NErlHvMyaI25e
c+HnDDAryR8mLz5eW8323JYBE1DW//yiFkIMqeDuUFwC++Sz5RHjAfkWhpPo6D1siTkDBZzyJwIP
U8nFS3e5u9vE+RV8ODB+Xn5bbc0fr7RAJ8lVCa6gmq9bpxglE5Qr4RObhy+00GgqCnjozUFunaKa
0FzrEPE4uF0RYI1Tftqxfw7gpvcZGIRgPX0Y8Y+pjlZG6uNf2+16cnYl1V3fKml+9WrISRiwIIlD
Y2JsrDaJ7s41uRvQb+HGTUpfDey2PjfntLeW6/jfduQxsMTWpPvMwtwdP4IUZcKi9cj/3/jSNjQS
XXbCb3PmKN4YwiEpwDtQVulXdaCHkN1q8zJZ4lneTSAQ558vtE2Z/2loPG1AYpN5gVhOLHQtD9BY
C14+cAJ/QxftUFm6fxEghRTt0IR/+HiKb8q6/3XRuXjeKKt7U7+vbqfGCvq24Mj9Ho1Kn0PmD02/
VTnZR5GNa4ttxUc04/5DLwSwKe9b7zUGlFPU/sYfsYmOl40a8OdIetIwnttdgDXWqD8odpvlfWwc
HO9QVuVvaHJ3iXkAH8AHlLLwDoeWnKRwLgH9bEvZPNftRWDi1H6QDYP59If2qrgMuA7PFnZPI/wg
yD+5w93Yued6wGdlhl+5TpCGxt16mkul8Z1Q+TBt2KsOGTVZVXYpaLEvhM03Qj+L9+Od/OM7doIs
nepiRh1tuZvGcYB1mjjYu6aV/wKBU5CWrrAw+TNjXTETMMBf0xgXJzZ289Ln54TEguZQRb53wFTE
4gX0khqCGXIL/VLi5BfA7TAnLLvJ0Tb+eesDeLslVlzqMOUstCryADIsC40eR8wiDrSshEmz7n/M
j3bq+O58TzfeSg4DJ3L6AL2eNRDqQ87prUnej0SB8LQZkO8HqrIMYhkSD+0eiekSFeAcGWsr3h2T
ipkngZ4CfTF67xpLEiNoTEFDxCKfQ2m/zVsbfZx5RjhzU2oF/Kub27Fi7MthrM98U9ZFD+8Lr/vz
BVt+R+mtfx6WWeRjwJuYn4vUQ8Q0/fjrR9ChlVUwUyEqcGQC7cjQZMtgs4Pp2FOf5Zu3BPbIaF+0
6VReUG1PN44EB0YX+aqEjPt9IM3MdG8R3HSEQ6njCbU/eGzMw+eYzi/ST/Ur8HCd83FcBzSjPKhd
uJC3fZvdsRSrM8e3qXZ3a+UtIbG/lrV3rMWqeCUW8U6Tlk49NTXYGBccXn3b3+ejP7VnKKdWdZue
0K4SqLT83ldwU9WUdWcWgZIxkfWmU4vrW7z2m7lyByd8KmU44Ixv8we4uANYdgCIOY9ELLxiWecg
zHnOi7WLbAvZBgNf9sFm7EuBcGHauDgtRPmoj+FM2L+SDxiL7tMZE7iehTCKg0sR1eGNpoJPrdM0
3D0WCuFavUHK96Hj6CT8SQeOZX087TTFC8lW0LRdGhZoyUdmwNkvO7xsqXabejyN2uZO03NLk9eR
62mp3FxE62YuGfMXj27xN/Rsl65IvfHDABhE50oA0kVD28ZEDtRWvFggDcfMDI2tTGSF3VVbe4Wh
Ofupe4VUBvcCFcxcdIF1q9T9N2099nslyJnVnzUyffE2GFiIUFnvkWXASvPCJDbeySTIWoN6gvTN
nV/ot4A/XFTjXmYyXrl9aMs+2Qo4AkvPIT2NHgDwvVOUsCV81iSubq6e7oSgIpmcCGYhSD+TtKVN
9fr/ICdZiI0P3hoSMecUQlIj7leN+xyL22m+0bQH1wr+6BpMbg3Ze93+SbWbLVK342/LZhO6NqLI
EMtGA65XdvN9xU14Qp9Uoe8hMpOBC3oh65Sy7nxahDS4lrJHyIt0cuXO42tmW464iCp+IiIXet7m
Bd+I/PFR7qZMtBgq5+cc1atVt0+Qfrwwy97X9koSvJf5NmyLSdBuOfoNQNLmDfc1/ImdrcwhIY1+
FPVltyZiv04dlLoiQ/zyvCP8/Ap17eAfKS8n1WhOz8RPp3j5gewjcNyBxWrHmBV3sdlFvnkabOkt
Pq308yqRGPfSONr9kWez4LDTnuWFjw0akb2zFI5u/SWwr9p+SmrXBMqreMcFJ+Dt5DtcD1Z1PYZ/
ZlOQyQ0hMdY0/nlZ0EH0jO59qq2oeAP2CDOPT/CK8KNceHUHprcWYixTL65A7bthrtPoD6aX6wWG
Vuipr87kEkdEF1rv0xnUbcivrkFLWXFm9/voShsPatFuxaiiapGTh9ghHCrk9fsrkxrRJG/m1M87
lPUJ5iLW6+c+nMj1i5NW2cGyYoDRFTx3LbRG8UrQo75t2smGLwfPxIlTJEtQHoy/p03TNmzRDW69
QkJ0iLsJFEYy/Ur2/j08d1ZhPS+iWHt8yJaehNsLYoihHaVaZgQIUuB3tRo5N/rl4d06jhscn33h
K6rH6T2QDe4kgo6Wo6r94hD8yb6d3vhehBdFIhDz71kwijwmdvV2y2Y1hJ1Nl7nihZGugr0us6nZ
AIfmt2KR8BQndYCen3RCCZDYHjPDdsdjKUABbCZPkp2cWLS/a8Rj7PJg1IYna1RO1gYzkhJVRlUX
wuTcHXIUGgbIXUAOI1qpZ5qKvDfEek+iWPd/9ch6/MjE4CVio33ZufR6mWRNVlcEZm9QwSZP2wJ8
UFUqD8TIVUCNcRmLJ1fccLPiRRHE4kCcD1wRNVimCjG1euU4nX9+nvF0oRNgAotefBsB8qR7pi5+
F2fyOJhEhWSoK+h9wElaVvQG5ujLIIUD3HhAwtAHTARIn6R1yrXimpczeMKLyEwmmbAoJicBI8s2
TNBnw7tHgFl4JH+cDYVQmJkHDcgnO7PvL/u6kdbIjSZmCxj02u4td9l7vFVB11ThAVOFf81MKp9p
imDa/HGfNQ9KyiU0RUvI5cRo/FPlm9gD46r1ER48FNAjM5eaPctmoOdgM/+TGrbgV26RDLxEH1pR
yydCG2KD+iLxVnzMVV3Ex9ZOzRzIlwzrEew/XcpgZjbUncBNbWpfCtezf0rdp1s3pVx8sIwTUNg8
YdKLjdIvn5Ht0G7x3Bvn6KyRuhfYZnBoA9OaK0r7gzkJ0II/J+lWB6EBANli7BCvIYnxVeVHm8Ig
uy799PU6TVin1nBtecymD/srwcxV8rR8DSQDzUJV9vx04uoctYQYMR8vfjBmgdju2RgLoJXuIiBL
B8EOoecAHgql58W/dP4Pdmy0H6remIRp7uNvXiuCcs8cQY6MP4/aKTzr+WIeDtz5WJT3UMDBXE8W
nXQHhCgFDwV5WxB0P8RE2/yY8gY9q4ITJG9JIPnT4NGkdMsFHQcW2A8aky5OBHK9VCinrjetZQKJ
c/konjsGy97KcOMdW8b93pz4d34gH9vlKsGlaHfRVK1CEWsn+d3CqwCQ7K/CzTSUvoYtnLra1kbo
458kOXbKpPKCJ3gu8xzT/1JxRoflghHlf0Wx5ZUCT9MWQYHQH0pap1A3I5VRKaIFOsTuKa+XRnSp
i1mqjk7vaQE3N51b4SXUPQ4LRyokNBg2GoItLyyrILMMAQdYM1rF0RoLQIfoDPRUB9ODQBB/wOXF
FYn9h078wnThMA31XQ23+wOsEeOHRL24s+SBhM/1gK/0Bs5TZDBIPlskkLTzMpGFlhOdCPweOJ7B
eH2WeIUyJoKI3NyqrfsW6cqOfva+rRvryWTRW9KXX1AKnxecnlGYKOewCsP/JYmNtJmZtifQhOsF
zsYl6Z3t/y5vGmyBy4yMhbI2YOjKiDL0VRWTqIB4qHCpU+sCiQ0bkt0FhWvMgonAKcKOSCavOZbG
fCK29f0otsIU8ATXYq0scFuuTRV4oaI7fLBQ7Qao3mqv7YEaxfDle1zZI/DUCokdTNNrEO8RaA4u
0YfmlzJ+o4HAWFFwQKslOxd8r6v3XxexxePE8cviH0xbcRLQWGYjV69RzcmpWdNQiecwL1rhQLCM
sNyQqu/CpG4tYtuGO8C7jTQFMXIxiX8iO9kdooXoSoAOpFqGqXkzUOb4Fhc/v/3nueQ6XbYUtq8M
bfFteph8tBT9JGaRU16JAf6xHmZM39UsUmRpvmVzDUMkV8UUdHrXUKz1z5eckmM2S5F0roDalABG
94bzEHOEZF2kuGySAaeoG9k7y/zZAlOLBy+VgH377a0C1tcCnYs9Xt/p0XDD5PxeJoVcnF4Gn9JH
t9w77Gnb6KH+L40REmqAeZ+c28HDkEudOsxRAB7nD9lXTpPuaD8DFjIYEfbWxBRUDwTSqc0famO/
spoVTMVTT6hI+o13IYa8q4A7qsLyEQSLeTRkOXFvwee86BjHEvJtAjqtQztkcVOXP4LXhyqUUV5H
jqhHasJK4SRYP6HFLHz/mMa0Y24Ex9vTEmyIYpuT3Q7dUiRH5V1krGO1pGHedASB9K4plsHrh85/
FqDbCVGsleldO3pCgZCSGuVGQ8X55sjNB42j4sMhjYlYTL5tiON8p910EfqV9My8dMhNRc0MYvNg
BKXakBNXwWj69uO4AoWXmcuHz5OLVThckdlqLxTucTYIXC+1/Xg4/MiFVOQQkjglbbXdeYsbFxir
DktybDa3IaeZFyKr2rGPvKZLnNF6h3wdZpK1xl7NAQfQD3vuQMPppIYS+I8ZvbTIIDe8DuBy4Q9s
aPMsAJafxrGDJPFIj6fzTsnVBHDKBO6TTUb8Ved1bJBS5F8ItIVjPgPkuUY/QR/2+8GXBg5TFuWQ
4lbYpkI/K9yb3T+MfOzecg7w1FwfV+N/be4ncWfWPNLmnJ9epYUVzBJOv6BmHfi01FaEiOSKxpLE
F3uMd3lfYh7uVS4bJX6LDeuZwsS4J5WP+lEulyIDC+AzBCVBHRtN6hCCOVSTvELSDDeMR+7vzCNc
S2KfxinlFHKshoK2kBv2M4VY4gOJa5QEtp2Vvf/eYKaFoU2rsghwdCVtle7kBZcDAaWdSo3i9CA3
f9FvcJdpv+40GfqcKOLaBBzor5Qx1Ne8TdR5ErxqNfaipyVvX2bP08XXoFCh4Y+v8WepfakjXwV+
numin7qdubbZZxmx4ElEakZ/Q0EFNv6P2WalM1MSXK5uxfkrYyBbVHe1BJ1qKz0EbmILM6iE5SdZ
BlxnUUlRLhyIs5AJ0ady/HD22exyxs9yEOQmCxtPyi+vmko5a3wxIvgiQVgehlY5Jes/HSQkqst7
iQlDiX3+GK2WHjBBvz+YsX7h/5p77YPYQaWkCMxiC/JyGaZHrPOwHv4FjJGbuFbDnjQ3QQaGlbZV
X9ZvRRuh0f8Z142Fa+aUWwhWu3wVg1YdDE/lXcEJW3V+NNfoh9I6jkpcEciGNBFecfr3qwG3igX2
WrsVpKWj8Z+PEdJUP0f0c9/adXHf/gCnB6RGk3wTCdmCVOmC72qbHeqvbslLOGJem3zut7arrg0t
PtY1KGWrjaQrPte9tczSYkvKXfmN4745NjUOfa0wfFvK2V1N/hEQOM3qd08Nb1K481nDd4CFZyMw
Nd1U90/iFNLAYfcXM1jjhZv0GN2WtNDfX3G6dGwqixID51sSjtWQXH8r6FL1PPcAWkWqcs+VQRMi
2kuVJ+WeLEkJP/ni0PrRtDdsLp/mfZoyND20MU2B9hY/cVqH1IStWjHlKDcdBa/OVTAGXvzAvV1a
9EJFW5cM6fKvwhQJFDt8Ikz3YORZ/MG3Br46VOzXfRR6rUQOJy8mq5UwGD57es3wty8V5riGmG0Q
/iJpekEmUUpHyjJnkzyAO4X7T5r1/rjtCBLeO0tC2lvCu/xd2+nR1B8hI3eHn4LtW8JLVAfqUr16
ProAT+5V1U3aLHXO7GfE08TBXazZIshTONDoMB07s803O+4czYoBF0T8ZMwQlDuimc9CnNCgR8eW
61VNQjIFYHv7y2LbBr/KBWjz2y5phGA+U3FBTsiPcEhd8CuuUaI6zhwQFym1COUJlZX+CJHozHts
LjfTX27NW0HKfkHTAQ7WTizVNVub5XSLVzNN5QpDoba0Sgm53C1+k/MAw8MhewfbNYKOCDwyuPr9
WzZHkrs1hyjRBF7dHMguQsOjbkYLIyhISPtamHPZ3g7FRk3811IktdWaCswUKwdtKbfHVuRq0o6q
KCeJCSmg3njo1UpITqdvY0GRheh9u3R/TwXXsPKrQvxDY7v2xZomWsUBjltpaIluHfXftqELPDl2
GeFKtaZz+kXMEliao6Px8wP7XuZKzqoiXvA+25Ey33V+/7yerow7CahdazxGLw0IBaTj5x5fLpad
NR8Uul1YYRP5WxgO2h4pKDCI3vFYRrQBE4AfpO+AzV9Vgfjn6sUb+8hvVJMY1ZhYCs6y7whalmNF
6jAKt8l1DE8h0szcJeL62PsyWyPf8S/grP6pqAysTcngcXm90Qou7ldE67Y7wkKkXAfqz+gL+5IK
jsv3HTCrPkcQkYIzRCssyUJCcKwUfTiMAPhhtHTGi8t7acOaDlH8pwKs/doRguY/T7sW21+oKXMQ
JixGVOQWn+fRq8t4OYtMz48LLtc8PTUVEBrA9QWSefsO2yTbZJzKFfMTCD416Zgrn59YIcSFN4Se
HQxmNQ1MnAevPMxnczQuacRphDDJeb1c0aglTVvQCjll8J9Axuub6YsGwVHqnz3d5QHUFWZ9pAqr
5iiY2qTRw6rwb/VsCWPERMh6WDqmKnW186AMwHDBoQSCuDjdOvhxpvWJyUYiT4718pGX6jt2Fg/5
LdeylBWUJnFaUGQjze93MVn+1hE6An0Pzi0X9kzU/tiD+Bnup3ED1YRTYgV4o1ntqK2dxUBjRKsl
OKsndNPVzleJ8RJiXaOL9W1ASHzPd6Xm+GPkLQsRhIfvcxEegzt1m6nqoIwO84z0Rfu8ndyrpaaV
qz9PogiyYk+EMRdF9/QIIxOrMr+Op7kkf4EFsBhT5okGWXIJfmFo0d5G7Bh5w50BtABjAsLoW6Eh
MhqRebWkp25B2VDM7F2S2AQGaEVJln7/iwcuUO84s/l3EViBUmZNUB72RlVcGDGymvHcGr1czGSE
HKUdX2nffutBUNMb+B4foLxwltYFMSy6ZSqNRdbhzvCRFWoUp+DnkEsaTnyPl7tJNcEsvEVBkfxQ
chvYwmnARsXAnNIIAbpDWOFn/uX9dOdi66ub4xNWJxdwsH0tVQI9CTLvLYC2Z4d7oX3bxbCgnnuz
9is6BR2sLwxLbEOYoV2lOi3S7ZoDldtbyEttDEpjOjrrzJbmllYHD3SbH11ZKokFQMqIBTYA2jV6
gZlmVX9M/uqaqUDlgLUPu6+4+r7PkGmryRrlbefCzmdNRTWfw7tVBxrLH2oCla3JTKBDupwwegur
Vu3uyBVcIJ7zCsJ+hwa+dhuotpiqnKv1DTY+VMGzKzK3btkln68xSTAKe0TV8rBGrB9Skxhvjf5s
+GUXxTFOeY7cKehKWpeTIDFXWDhYMLbhXln0LNn3PxXkuUTuc4IMVXEQV0dOJIIZxFR3WZN+X2fJ
oAuiFm7zFg2ML66tgUx6jTmynqF6v5LVW0BJsNoXmsfa7byzycVZGSp3VBDPpC9ojlhtBPxczWWU
Mi0xGLKqyMlrM18BOjOr++On5ek37GI+k1JUZO3h8wQfyW2FM5KLjt6qSbpyEZmQmngvKYTatSgc
3RZVYf1zahv5VCRedR+QSiNrPT+CSlXuG0fMOrSq6c6pRTnyFwS03Id4bwc71ihiEIwD3ayfiAUC
FkoHExuBWWCdU2hTT36osvYfX8HncU2mUyp4i/wrZ8pTRNGK1ccl2fm4RMQADAOoXUVCefIdT72b
NN5up2jQyhVkgywwnfaM28gyysZTsVYKDjpFy1MDMJ2nHdIfQy0fOLlgcgPweW7eZDwdrvQ6kADa
PkPikn5vmJ3+xiiTpeZL29wK9zYOKWgRXC1Ao/vo3g1w8WNXuLxZV6HWnu6ZMY7ZVac/wg0inarr
4Qmd4c15iCN/o0PvR/WCyF0Slt51PiRxLOuooAF3/I1Fz/oJzsw5cQLlP6syEfBFgGmggqaJnAxK
kxl/jEXvHV8BVmwSymym4I0xCJ+i3m5q+ahBfdseUxIKYN4L7iYjHGMa8ZtqsCWlm5S/IZy5Rypa
rcBrYmnFHJcJKMxWGbz+xwueQURaYkp8MQDlrW/G/kLLkEzgMkhT81VZuwA1gLcE3yyOkERSkZ56
1qkz4eqiiXN4FkKunDudJYARZbjwPtxwTQkmk/Xlu4kHBc30XIjMgl/rS8kPN0PLOH6mTEZagN+B
FoQUJP2YA0GDM51oSlTBxdvuNAQBbkH4F0RKlYJzTNB3JWoPyI3or1VzdNSQlidUn0nQ20isUuIl
d+cVSoJefNrnVB1Vyoq9iAXYrDnA4QdxsZ0b50cKnoiMRsszJQLWaPuSZbg3zgCzdvCzTGA4C5Mv
yibwH0EcHNdCPVnlCsAZzQDs+qVPEUhidDSJMMN0N0JVnE6CkeCH3yjzaAgusrjfa2VdOQZkwBGt
ZwU1P03Yg80rKeDPo16ERg1Sk0m8g4TK9fI9S7AxQ6dNKRmzalB8YdjSJHaDykAGKl424YWvbaBR
8PdwfdNrbXxS8tjXJJmz2EG7e3QHeKdPJGmi33tKtiGuyWfTYRjl618rIExudtaNotcZhgWMNiII
Bt0S3f7jcS8PCUD88CKwSaZVSpqGMtC++e2h+iODkqxxt9i/LmVaj4iuRIwz7LDE/GMRIpYUY34l
FevC1tcUBhQSMMzUguGwAxibPfdHdS1Im+eRpIMgwylXJGlulJ/NyKKFTXAjCwblyik7omKcSwco
chgfvoBLV+rHSfscxBBOuLF9T/TS+CLWfJ6ifEL5vnN037LsjmJgOj0fna/Hzax+nbSepGZ5SCfU
3L5cUFPN74oSGaWqQQ7rCu6JZIRJU9C8CpX844aeJecBsZSN29z1Br9aKRl6k2sWnd96Sg/qQtgq
w3XuTOEhYH3pNc7NWOd6Hmj7kyVjpQBN9rGC3QtndzmfgGR4070z14F3hlsnu5OCtckybsQoi2vS
G1rqRWuWgmU+/A1/XSehexrcihOv+pyuH36D3QggE+SAGN+1derw/5wS2QFTUTvIRU3H2lpF//jx
qBjwWQax1SA55AcHFrluSMBBDRD0VUmabJwXYVii97m9SrcRaX4/9jGUAbJELtxkh/W6UucQbTWZ
WyboWEXD36ML67GYeQxo0F/ETmk8Df9WjX/+4q+30fE524KbjrfH8bru4rhFF0Y0ddmnSjmkjR8Q
rmALFL2gWOFTaT/mSRG4Zbc3XqPSsD33XIpgrXrkBcyM2tlWE937etMT1V9zKMx67czEu5VZCqO0
a6wpCP2sySOw1InNpwK4Tf6RLrb4ZszxxlLj1ShAGD2ahKQCiZ7Vzrz44piKcFI9mZMKnnfNQhXN
aC50Wd7RyrJTOYgY1wbQ47do28ywMbpo2NpgPPONMR7zlQmAQxDsELcn5Vg+40AnegvR0sKmqj3C
+h3eiLDrUjTlLeLAdpXpWZW8l2eV+Geynv1KCi8B3AaAllOZO5XpuF81HODyOUqGWn8mqYbnbzKP
quykajP2ZL4MQQWVuElxThf7hxc0YWUmPJMlXvVNNFJSYkjeKKdHC8xvW1v3VL0DOuWukyAx/e7d
apswA5W8SWyJHjsy7n1etjk6q4esjCo2IDVhqMIY9NkBT6sUbMaNVReJmCUjrr4b8NKsoQUUbonp
ePjahd7T6UdZZ7mEk57YtcHXKzeDU9Yr7u5gVM3RYCTIdr1+RZUZqER8SI/zVOEM18Ovy6OjPuf4
CRklQvBpC8GgTTNUJDRrMxtxZ5cOHfIW93obH4GuUTxAqJMZZfIpxrugEpxbtaX5vJ3kP7ieqop3
I9cxaeNGXQdqW11lcmuivK+Nl/1iteUgHM8c+vDjhIyZlvbd40XTR5CUUfQfT5FAJrIyc4yP1INF
lYkKxlXiQ7kGlfC3LXKKM/LzVH5C780Bmkt0azBrUVK+icrBnchA2sgcxMV9DG6ZpF0qmNvRIx94
qh0wpyMiIxPvQ2TTNOy7khb01Zp5iL+DZr1OFUnmaOHrbENFOBx0TLcy1zM0mut8K9Q+GKyflpqD
FAuOvxCOKnkA/R0LxmmOulAtDWTgW32Q9ZHaPDsCt8wHT5AA9sOBRWf4LGfqnDYMQmK+/J7EutL0
0Obg4bx3KX7FDdu6J5ylMXRa+WthwDUAmsp/EwVbWLtMUhPl1MkXLdi1QfpEIxHA//2RcKOXhpqN
NoD7u0SWz6rsgCK2hGpL0El+ZWZP1OGu0sp6tROEMzDv9ZG6HHDRkF5+cv59KeFTtG+QNItWHIse
MggQETYSQ3iIcvKC5rrPOoU/ovrM/76kRPg9EttT52I624Co3nEheudn4dxCC2a8sMp1tgCX1eaN
Wapnj45K+zcQ5un/ygiKZc/GEeVhaXEwJN9o2kF61yw7h/EOE8yKgsqyYMdMCe7Aw0Cy146jDOAb
8W+CltBEdRijraVdz8yiILoIOWdzSRxX2bsb1wuqCLviWr/3TgflDXjJnZAHKkoH4ju80lAlHJex
9UgEfWgS2LLGtYZwz+CvP7m6IfGfXb9IOJ1HKqk+LY2mLlF13kMBMuTcPKpBMi02WKEbAQI/Cx1c
5SnHiIzOe5ZX770nncjR1/NgYB29FYcfBdUZgry8XRqmDCZRz1+FZeABZXKtkOSrKwQLPoaXgZYv
bQDoIbGIk4CVbqirQH19zoA3N76kEP43yaxJDmZ2PGgaJd9wVVOkzGjSFTYSpQQU9q7bGKpAEC6p
jDtea6R7VToiBQORZ03s+1fVhymIkfAsVvwRJRR8jqiaPqH/dLwuzmYJ0qlRjUgfii6UjM2oiIbX
mJxUn7AHKO75hduayU6F2gBPM1jYyGoiLTS0+XQK2XSz3GmDI5yKVJqc66VzOOot7sF859gGgWAX
DvN6aIfZ12fy7bK7MJXC6DZGrpv+YIDlvvHbCLqNrJGFmrFy6G5CeE2gOPsFxXU6F3n6Mqt3jNJK
ROkBGP+j4Fkw/eBmL+nZTNRPLp3W43hR596TyXFFV49nxHzom8YiJnAXR6IQEbnHhcyaHNd52O+y
4NsulEQmEhFVDoa6SWoMLapwBFt2mTh8kCzsZuVy3icRuTzOeBXDvtZm3d2KhCm9VAXbGiD88g5B
+n4ojplp1ovYyfGzmRk23AfV5K1ggIUbCtnhvs+Ox5O4WN5KZpM+FV/OFL1Q8r/k7fiueIPLX5Zl
H2X9+6D/DW5mR6GD3em4xq18WA9LnZmKlDKqw7vgxgHTQf9T3w5YE52J2DlQkPoELdVcUVdj9GgK
8r8yw1HrkJB6kXf4gJx9/Ssw7qOtSKIlEUIgGuZRa/AWny9JYy8EZZRSOHGydtE+0U+rAWNI7+xk
FtcuD9JigFZ9DHP/9Uuo51ZqAXufzXGkHp/+Oj6cvJmGJGShtO5ux9JOoPg2DJ1FZO0PbJ10p5wF
0VeEo4/qQScbtitbH+aaC+NsqQRqPgkJOwrqUQ4DeEG3r2jIH3+dq+BKB4ibgiCgjLV1R49TR5BK
5iQF9xm1OG6p8oX9q6WUwbFIg1C6LaiAxKQ0jiduDTWw8ecKwe74oGCuP29SK5oL8qcKFe3H5jac
x6E65nwXpxIM5mCEL5iGuHivghEQfxON+5AgigAZGJ3I/fOkrh1oJd2TXK/NogLcUdbcfgvyX5Bt
PYw96SGacCUuy4fb/srdv0GfmISlqr1gnHvdjR5M2t4vae6HmeClfzoC3nqz1vNqMnsegzzt0ESs
PTkRIyyGM8pbXBExMQGZ7/cAuUbf38z86jpxK0ePAMbjeZ12TLZq8ExhBDmG0K/5HUA4rsLbKSQ0
/3s3oJmr15OUalb2rsxPHLpT99de/H/y5Z8JVMJrN1rB7Vn8cajYj2K1ky/BIejyySxNxZ/A7erl
iwD9JmPj+HM4XAFYMxFm5iiov3Hotf2yoLESyoeS6J+aSpleBz+0TEnJi0LX028Aj3sSV+ealv1B
MbCppb9HkIAlgm9C3Jf/CaPmx4yHK0G4ory8/678WPswUzJze3xy4jGDVoF0X6lfSgEuE9a34ZTF
OAwiB7i6//hCdR4rZq8W7GhI9RgPvqTl5sFwkut3w41FcyPy6IkH2Ee4kz7U9Gz0qMvLAF6LqIp3
6sHDuxWX32YBu5M4gMwOQYtjDtNnnmbf29SNpFWvXTw2tmqKQyfWY4rsXi2ZKvrsqgj2wItx6D9o
XozexZ45yn0GUs9zKstx4WNPWRK/nZvWyYGaqjYxHHJ3h6b1TzhALEsmr4oDL/pRwka1Od+J4XP4
bcWB9D+0wYujzTvpKAif0bqEiR1bctgivW+OBG4XOfV11wuKddWR1lExT/1BsgM51u3VnWd0XxQ2
vcBqHSZPWriYhhV1Hf/mGDOmu4Fen+4FJQo5FmHRs6y8wL6iOR0D0r6T5HEkwq0lkSQyzxRktajS
L+3tW3RDwhG006Z2bW38P1ylSoNPDGWY/zyNtFGBHpjJ6kIDT7vEtid1UGh1Vo1qFFrnuHkTMnVQ
3mlbdRlsyTyJFDT6/t+kQ7oI40IDhQVEEzOhYutMC9NwHHzVpru3NYDlP1FqVl4zKe6sYl8OXbXz
IhXcR0mq6kWHZ0ge0340ss572NmsvwUOP0u4K/d2mGVhCP63iUowuBt+p+GPCl88M8dAloGtXpBo
Qy3xoI2IVXoU9tE1v23KK14nVD+3RY9jVQcAZOIbAZfs0nPmg+naAa2enUz8q57JXy8ipWf8uyIG
HNWA1nBNilwINZIDXzshtHHd9sjEfMhyJE0jfWUTpuqqXWx+p+iHv74yyAYqk4/ME29oKAIOjYGC
gWV/Qus804d63UJLNdKb3sczpDabw/VhrpvCNgHsNh4yiAYAlNFgBKcBsYjw//mlvYILM995rQ0y
4fmaY65RLExsNLb9B2ic4EL+85p06OOBiTkvMMjtR2t/tQjLF6npzgabnNCgiMJkNzT51SiEBw4N
bXE8BFkdOUS0ksCdCYPLF5pJix4j5y+Ayiy9qnWK0zNTPKuimoT5iciZcPTF618MNm+yMOmcMMs5
87HGFZiEnlx9SDSFqciRWFZZafh5BFB5lfC0It0G6xfdYpf8Z4uMhXms/6+wSuPBaaqGM99VIy6G
WSgiYLiUTO2wktu+BaFUfhVgbJNYytnkoVIPO2snNu5zOUdZ9dc+MVUwVXUxFxG8lQfC50oLCXoA
BTtOQ/ZcBwPbf8AMUNWomAY9Sw1plzPb0YXxHmco90YVD3TQWAKP9lMnZKxmjSa7kNpiEVgGCWfy
4kc0AoR65cjOgwLcFZqBoEydv9GjKcCNtJsSZInwfxwG73e5UEvgq3VKfqCEib91jJ8/eZrYFa6m
tEz9QfVI6YqotdLI0oszM/VH3AF7Yzkc3NXSv+6d7bw4nXH3M931P8mJ87+iwFqBWAzizmwiG/Zn
s18DnrDtS1GDqXDfrtVdj3lQEP6ArHVeUf3UrDEdgipLxfraGRxHiPbbXdTN2NVzz3RVCduNfn8g
kaY1OAjtnffLar++O53/ITdaDrT+HmjCKHX4071IGfczQD9oxcEhbCtcs7XWrb9QscqxniRL81kA
dK+MH742J1/SHOxTf/g6qded1NGep//t1ZaSEeFOONmd/6DyD8RrjLdrNK2zchKBp25c1va5AN4K
2Sm+ZrM7lPZjQ1VQ2RBSdPHhmM/IPHTQ1k6svZ1HhD9PCyQJp1dMHKh1I9I7geDVjO1WHyFcD27+
ZBltxGYWITeB+6bL4c/C9/spXMHCXGBi4U2k6OzHX9q8AKMR7cTeWu0JD61q7egg85BpH+31tt5T
kVjZ2TrtYB/jkRWdTKgej0Psv9O5hxQA27x72H5gQhQ0G3OXd1OMNybRekGaoMbqa2XKL7yi2DdB
7mWZjtztwRqTUBVxZqNDerP4axLQ1FSYlzrzjmfoVGNtfFoJJ015Nw2iVERw54+dbMpi0juKN8QX
BpElYrH/WiL5ORGmXqa3wGfmXYhCbwjnf2Id+vrtn1Py0uZEWOSUILXBYzKPnlH/IBjezIt5SG6k
0n5JSakUfRDuDX2sf4VWWrbfqSQbtXujOiJRPRYi9x08wjXiI0KSZ/A8d9tqIZN1D/1Qdca4ZemU
vvxWbdksqp3uLEoBbQKqKPcJUUxemjzta83K7p/5lDOvR3BSZo7t4EtCXltgUcaMa03G3ELzsN0G
hAiPIi6fZsjWdxKm56/gEMe0X8aSLn5P55mnvl2Pl6WXUq8Gk/UVtNd5yfrW0hq9qx8RfXadzdnP
b05HsdeRvSqzHZgRITrc1v0C/iWeLPdX5SnUrrKZgTJfgYEA3mc3J+1WdmCc/+XJsxR1RV3d0MfI
aph9ooiSt/dnp13/b0fx6yLH640tWw31J9H83Zbu3K78Jt+jQU/rpjyp7vd4p3RPhjN5yF/XreFt
wCE1ZwQgKojg8VR1fiEDu1t0TqkW0I0eZsqyPDbY4DwWzcftrTlPNbEzqyao8GgsFOVd+zhc7jpL
uGtp+MfQC6U2YW1jh/B4sVB5Uyl7wicfqCYVpOei4kaBuyZk/1pZkfoG+La9rMkht+PQ9VnYWIFF
na5IWbPDeDHJit0DHLPorjpw0rq9PSYtPhY+JZQvMjWQZXjkKoEnN6TkeLSleDdc+Y2OiWeuHW9n
LDXf+Xn9rgnHb3bTuxY2jUx6aACerTh55hxK9ljwbOIg5xyi8ZqghTlnoSd4ADaRBtbp2KVjTfKu
1MJEFL49Jax+dmw6jEz1L8gluuzhR43NlXn01vsvR5AQYln0peT4ZMJvliA8I0Au3E2rV5m+a7Ca
J+fv3KI7F9QuBXijr0LBu5ufMSloTNiRZ6TdespI3E+/WZ3vBpjslCoo050NcsbscSWaE+BNd/jX
Z/iYeC/dSCI05ozGekw51M3p74/vq1Qzum2GYY0MEfp6pn2GgTgrKG1RgzB6kiXV6Z0Xu8Y/J3C0
02gltUXfd3FfeoK/lr9ctHMBe/8wsKwFEKDG7ueSJ9FlCKjoWVufFc7n6NnFgNkdAfpctEPFJh9B
wxGtydDCXunvcNlMvtap3pYDmyIo4JRupsp6Li5+pj3YW8ZFfHFJ1Ht2ozB6PCPLOWvrpzAyRUOL
/0aIebA7+AtqKGXw1ElfYbo5t5apa9T7oiakpVaL/8b/3qYN26EjRA0LehMQ28EE7WKtnFfKAIeA
m31SUFpboAjV/BahzHmyGdqrDUI+si+cwnbZLYQY3nQaleQoRG/rqixvG1GBxHknXlXKn98T7K9s
9h36vVJQ7wSSOjI86x3TBjZ9zXVQ6gc9AG9KEsNBpSNrGfkBSjYxRCC/RexqvyNi3SMRiFj+9l9w
jYt5siI/ceQtdAIYAEClgTfB2F70f19fBKTAz/GJCCjWjaNba4uHS4TtZPLxdfcQrcQI79CTNJMf
ZCxqPoX6rw6tlpQjIzpRlmm26qlkV8mDuk+2h/Rt40xRMKv4ClgstC8v4cgwycI0kxsHZd5g4Jwq
3vFF6f1tDGsfr3Lld5s/UcJf9f/2azXOHhIgGRQdGQk+4XHpK1TPCvnf9YQkRp4E18yUGMshhm91
ruNV+TSiUz5VTpAyPDEziuQV6puCK6HnjmwB1kIjG2cvDhuEytUTTDIA46Hwfi0rbOmnkT/3UWYb
DIpnXOTvI9nUS+rLkMBA4DlujUMtNfr/6QFqr7RKx+DoOqzs1wCvPfhwbbV6AgLXG6ySjr1suUvS
7l9RopcCqLkVvgcenff8A/5OxZ4X2k9rCx3XJFXTxd6ErsbpTgcLYXvqHYIyYQ16KqOioQNEDZiG
jreqXIq+HD/PliTM9ndfrq8FQmH5MGPAK1DgD8mtVfLPDHlbWp8BAFKMfbsfaT7nE24b46pFHwHW
iSbCEfWvp7pNAqHdwG/7YG2sWt18BLjZEI5oF9L/H98NNnOxWLPLOZb71lnDBjNnraaWjjIjcCg+
ulUJkrqlJiQfrt3HoRdvrMjxz3YmxXLuNlGM5YEyMQHArvYn9+nctRFtoyVFCf9l/Wk+A8Z+Qpaq
VxCd/YGeNWry+Wp8xbqwJwjPKcdq3WFw0eJfZZS0dMxEsKFN/RxrCfty1kjnocVvNtc9Nc2CP3QX
vc2WcgO9aJK03O1Cq25wQ8Eh7AjmWh/CdrNTAGJW36zf9S783U6tgR+eWH9cMRnRf1hsYratTqaq
rItgrpbHiReZrxFo+ca4kJZjIQYe3k4BwXpdEHbq6v1arqvB8lUd+Zr0BAcLDHNwqLzW2b7QrTd/
QGN3Ppq/fxf7XktMw97krvsuLmdOeVwyWJAmefHFnpIGpZtIT4rCzTZ2eW8LfF/y2ZcWW5/7WAV7
Hx8sxu7pY37t/QtieDJEg2wUNXNZ2b+fA6AlGWu5RhnQdcpY9XgtPWQdGPelNJpBV8eiK+KliyYH
AFHQILqAwmSriePjRCO0xFtadAPD0JpRSuN/bdh60E0JNtGai8YumGTQcqZ5079gt8KorxamsxY5
v6+6edbyjgeQVXKrEy0toen1144Mdfuhi2WFpS14GE5l9A5i1C1otlux9Ie74zrvFXMv+CjRL1/b
yH4ygk/BqPPAZqKjNv6gad3HZpZ3m6BEtd2qr03m4sXzOzJugIBPqBev7pcotd4ibhKstc3ThaM1
2zD+NkNTpx1rFEZFntppQ9vCWyLhmJhYDZ9BItxzynbXmF5u+/CsZRNTPGE0KH1PCdvSPK6YjAtu
+hY+1lFrbvd1XCWgNh5wMmY6g3qEbSDmVVnd2hlJhDdYFv2lA83hECwGWBal+YXM68MUNWLoEaw0
qajab/kNDqKFyPSiFV+Fu0+whbn/bLXGj6F79lHPfA+iiZVuKfTr5KSLMCJXktANKInr2Xx/7qkr
18BtK922XdaVBQEOBtK8nnGYIS13PSqDExvPvg424Yn1EjczZW/rUlbkQkvn7uRC8R7CsVu9eMHz
ujTtB+YE8raB+Qn26B/qzQAgC/JV1sipwy9LGAzxkgyW6r4EXXqHAurv3GgECg6xO23Tu9Tzv60K
nWKdk53kcac3Sl/3dUvD7YK4xMrHxjBcU1w+r7ZsL9zk31ddWWAkxbWHwTox1Q7YjMinMxUMQca0
odaIurjI8rVXSPYsdmL6TMP5/LToRT/WPeR5g+5UBt5zbvYliYgEDCGU2brDNwcK5ju/TxBghqPj
Z//paA0FPx2GKSKdJNeYNIQzSPk7GcD2+6YTqtEplYNLO1o05oarqfV0FnOtmgSJzDfFL2nWl3zv
MtPteC2vmz7mBCcEOoAb2Q/lJ+WdVSujr6hEMmppCZRyMz89sj7PCpSwo66Wlcd+imXpyJwm9Afe
1sn05GVqABYOl5qPpzprMf3XIoD9iok1nDVZCPPSd5sdFnS/69xwkJWA+iKvT634cPs37znXRj/l
nEZFuEjueloc/212zZoIrzHDHt7I+5SsRWKPgvbK5/tgqi2JBZIH9FQnsjlMr9QaywNQZKudZOrx
mRRJEkiY4N7OVFYi24B1PzUAMTBHvtIalHKO9beXqpyjHx/hKljuitFBwJJ3EhFkPjTKl1CSnAcx
jl3Rjj968qwVxkhdiY+qmwrlfvSryf43hUB4aWDgcozTFMUgEx1w9H12Gdo7N7K/2Da71qKbUot1
GaliKWjb64iB3qwsOoIDvpu/kVBW5Vr5gc6BG9gS6gO3HJWBfqcW6NXYB6Dg3x0YLbij2zdAWhm2
V8/1G0UxDvDpd0ZCzU+fEM3joRKWn9bmBK+/rxBGRyZp/8nOTpBaxgIF+Qbd6tLKmBdXopODku7j
7N6Pf6MuwXfKFb+WFPyRxgIalYRxF9yjBIz19o9tPFo+b90vpYvrK23IoZo4Qet/8ggC+oXweekr
pZmdobpQ6OwoZSiFLgump93XMngU3BixR4G2Cx2kN1a0W0S9aabXXz5REDxzHLkbpIhI6fAZF2JF
Aw/GUF6AhZkWTvb0xK5g1o0teAevnl/gZOGOcNo4qyweFux/oC0gJP7OwNeU3R2JR1EfoSCU68Gk
q21fSyMTz75N6KJQ2LZhWVY7qebO3e0o2FUXr/z+nRVed22MGGbBbZ3CKaxGxIwaB6tT/2pmk9vi
TwqzMGNsCbYyPn6/IFCRihsm6Zs9CJBSKRsSU+6KzJ4to7GENR3KFZg7MwLSo1LE23KHCni5ECtC
lRNGBYigvC9YZhb3JauTDJcS4riqH3gwKb7A3ILJ30dWZTC/IuyCv8CqdrTlWYDlun6vWYrX9m+i
G27qm6LClgfnMw2+bA+ecqd5bZmdyxFrff1r3fLBacEvMi6848DWEzLlHvN2BWSCyRZuzmn/1wCJ
pO3lgIQyDGJ8/sIcJfoG36gi7SlSBKYmOyw9FsY+5Zqe9iFPG03Hj2m2yHedJq47I9eb6mK+AVzR
2HCIFbcZXdD/SNr7e+ohn8ixkrWikSMm+nSe1TqM85pvcQAphvtOtrf39IhZB7K0bnFE2AagFLE7
BD+RviBK0BVJH0Kh1nUawe5aUSph7sqHf9MXCaMf+pN+vkYoW2pHck0Qc8syv7Ba7q1/QvITq9vB
viVdKs3plUoYlHWwICdvnTlON5PalSRnK/VmOybMILe9U+o6CXdVsQ4fTPqbCvOl8v7vD4tTnrfy
kgrA1u7qCCbaz/jTpW2H2szQ59fN0X5tX7JjhuqzgZyCehxORu/R/2K64qFMqZZw/bqQ3x0a6i9P
+0ST/hJHAXUASORnJc5Z4lBQxUGc0KZr846kihsHviCB+PzIl1BqpD2rb/+blC7LGBGjjW1UlD5H
f6ibty5VkfrkSyEMpsB/c93nB+XxYb2Q/UBFyw8RJbkAG+Cq26xPhX/xxgBfQnfYxZHSePC+fLRk
1NTcelfNXIHiyqen/UPVEGU3IVPMoXt5wzY/J33da1UBOTmSmNJ98ajWJZCE3RKRkq2WQsUwfvPL
tsNmecsFzUFfOKjbRWfxBBc4MNSrTKU4MRZLdTYniVj+cweOe7vyyo5u49jkeoT8jrn2c6yffyT5
65FiOj1+mPD4tbdkcr7+gYUrjq17vE6LwNnOoRF4H1qw6wzD0SITk+pr0SiGHiTUOEwC2DI2JL0i
9DoAbkAI+lFsDUx/NXpleaQrVCGxhibJgG03VRxSENpeA3WtuW3feJ+Y4VcW5DfEWC5NNfF+lW+o
IoJrqduCendEQwLPy9DTtofPTMPFcpMIh/H9fSgIx38bGVhb1Q9/nynXhz0Dq8fD9O5k5Lj6SJ9a
z61+Mkzp2ueGMBzjxyteeMH7uOh5qP0GG81HfGDAynsLzEDcrfBJZNzIJrUwPwE8jn5pnZtLWx/n
b1nwX7fY+FJFwINqpi/7yUC8EMn2tTT8N3gSUOMYxkTIs02a+KQoh6sFk8W0i4ocwsC40TdIkZq0
kDDN/Wez0dovlQK9ffy4ZxL/g5Ib49yWFCZYNx7ckch0mtI/4LFym1bpDrpShCcYjlD/Xirt9+J0
I7AnqwSSXdrzbTJHi7uwlCkSBfVymFXY2uKitKWajsCM3x/VSsPWU5Lrkp8hqOGvQt31aVAqsNhH
ipk2K3e/eLUtW7vWkmGuBHwOwoHyVOxFWzxWqzDwhtLzsQ3iq0PeTkm+0Y/usg8lRfwkK41z83fx
GWX8lRo8ODkPl6Pg139CrHEgjhZ+bKFndNi/o1PtjFfvO09c5nVPfrH/WY5Y3zdbJabXGj1Ko6gJ
IkWvyOvYKMjg3okXvn1b1Js5tIcTooiDQyGxgmk+hT/yQvERiCQGTRsjUyG10XJ3Pfiw9wwK3Gkx
9jXCG1vI1OcAO+Q/Vn7uYABKIlw5MjZAcsQqOz/+cTAk90+9JnGiAe5T202SclP8EsdtwSmDgmQx
Irotcd3AKTEw1KxHYLpJ14amsWTWOeUVOSpiePFrhiO9LrGDz/sFJ3WmKVDoPhmDblkU8M81f933
7QPZuE1JRphNnH63KShCYEERpGgbiN4EIs02c45HcAcWtOGRK5t3Cp5owZzBiESUmuE99lYj6sTq
jzjPmkLb0tnAim85romnByfV4J+EeLoEODOoyoE++GqZ0V78aNQ9mAyEr2AQhQdikrbErJW4wyL8
ZZX8aqeiprmXIXJ/FOIb+i+plFZVba+mkYRhAGdV2TdWbTEuU3FyZ3Wn6ORACEdohIEXnMLRtgYM
xDQl2LVSHeqlTRgFsYDD5YB6HOniUlw1kJaIZzFEBWVfJcArL4AgEwS/N4P1TgGPdHCLdJJOFOd4
qPAtXdQldqAPv7wdnoSW38YUk6TEmzPeeAvTP+0JFPIWnGJaEaI+Uach3zFOtWKpid/e55UzzvtL
vaTfeU535I9gCMHKhVHh2fqPUJPy1N1Qyf99vHjAa/EpQEPUpiSgcXTckyKKbz5RqzkZszMJqpb3
Mex4H+zz/0ZXnBjLxbthTTycrdXxg+KF1/zhOEp0iisNOhUdISAmYvmHMNlwmoRkPxvn8ON9Qe9q
QMr+yGBoWNkkG0KoL9qporDcmFpKTBVh1JQmuG2Avnu9Gl8L+RkYQTNhFmeY98CZhtQXgxHYf2t9
7gL2mCUOJpfvx2MivunyI+bMNMjNyJfhVDLWPlHi51qyR3hE4mRse0ifq/7Mpr1XcNiLaP0XOG/I
dGcWluC1g7sbrlr+yvTBgF2SBLUc0HTlKZH7t0rReRFO9TRd3GmrEyOl6VHrMZeypUnBrfcCzXs7
jwCICrvGilTk9LpauAjfoPmU4KuZcloPoacb79uTogYchE3aayYb+Kj00iYaHxGI7CfCWMAxX7gl
yLLcuAA5XQsBydXQr5tZIxP2CYXaa8AxCz9HnL2IR2Vi43SLv2eePbe3oj+jsCEve/dWecPUAjdU
PveD0IxbP1IpoiCs2juUtZTV6T16Mehn6VWuRSrYCBi5pxykl87/th3ZrHrPySlIpVWCoHkJDfYv
fG+bZuSK87BLuQECO4cTKG0onamaLL8oz8Kqw0mwojMMfJK2SJxBMytYzgg27iyJV6KUf1Uj0UcJ
THb2MfdQsoRbdRzYi33ZoIUmHzIeR8UrdJ+BMqfZEyX7cc+AV3+v+opfKO6gElqracXjwuQB9BXz
/O/bjVyDhz1SeyVFxA6EekZS0mBaEsWh7El5MHGi00KzJNftSLLZKun1PEDHUVujmEMvTMa5oONo
tonjfPPkqI7YtwzoFQUksE1p0dl8FfRHTWBuyW4vkaHX1QCH4e2DMChPJ2UZZk+H9rxgOt3YKex0
imxmOqHjp1XN4VrgsFtVRLp9QmiHTF1DTpX33Lx8mc2YcKzShF/KAutLpaUA1qv9eq3SUiobZwhe
O9pthFiu4VCR5f3nU0B2zGZ1Y1XgGE66DKsyR3ArCS9yUac2uffGG+APt6Lc77SeJn7Zu8ZkCVuB
6O/IuTOTeJEpvHWgAyXf/odDWipihhuN8pk4uSEo85SMsZgaRUiSgNnlQM5o/Xq469+lgz2d8V1X
jEt/NpNIC2fZrEQlHxfFkCX70SiQn2dnWxCcBWc27YZL0Q9o2stlnkYnFcd8HfDyyOU9rClKw6F7
DdXOQWRSw5MxeRIINGx41KwLQNpWAhSSSf8Dhq3uaQSJJOFlczQw0QN7mU3ar8f5tB+LrkNAPJzb
IYYtbVXenbByip+qyyEqz+59qotcw7nnO7bUviQjaLkZY383z+X9B+eFG7/AFP5pvFmAs4onP1Gu
XQ0XsEpvpJe0peBUmxGdKAnH8daPqnbYAi0zSqibcxymQCLkxoM9gdHmGkU0Yxe83LgwbXIL6K2m
qK2PER3Pi7Wbm1WJwj5ThPlrXoNgmogd1Eeul++JGpaMcNs7cgD5R8l5Gsm3et3mYPAhmrodWEmX
Zc/zvHMhuFaxPMRWLjkXdHlUA9lbDSv+/L7Pimm2yZ2RUNplNhOBQvcjpAaQCTQao5p5asBrxkjJ
t7g7tuT1CCDUFJhn2OYX3y1Rd3b6ahdTbDQqry+1YmPrnn/J48rK0aBS99wwTW2nokmncg86K5kF
QsmbZR1BkudP21zPQHFpXD332/kxQ3Lc3110c3IDGU2ygy8tcFgqd20GYrn3dpbAvqMr0AvhACOD
iIEXBkqnXBAru5ZnGFWB4an/4RckYmXEExwifEcguEkO+oFuxYzXBBwmnufkj5B4Upuc/pE1NUfa
/FGkyRkD0npZ6ptUvAu5KpDKd9AWKcFdtbUFCRCFCyWzNTzZuIh5ukrIkwGzbIcyDu/g7Y3xyqJ2
+DksjpHFC8CBmSHubpOI3TdR4O21pG2eiJXguw/2JHJG8R1KFj/yM2Pf6+2Qh6e7DrZWIF4PeKwN
fbwDlOeg81L22kbDQCxrzOVU+lNCpkXQkRXtaVrwWR8Utj4Rk7vRTgHFmZGdHj15uoXb30G/rjh8
BqJJoiCAopAe4XZZ5jYxTtR1p2zqT60lDkK3WFiPxvWv2qd1FNAUH2y+R9z23rkbvE0LiaOYEw8J
3lUBT5FMHcINKKVsbFzTUT/7JqyVEimxaicRPhnBIPXHse2cwRyLb5Duh/8UMxRXtqI5lqRELHGU
FMRG/BhRmmsBvGgEet8Q0VRv1s/rEA1GJhqgD1ow/5Fzhr1FBRH75UH03eAbHirjtW8/4eUUaFEQ
8uyR7i8ofSG00iQlusftqWKn/FxasQdnh6frg/ei8QRs3wvr0sL693n1urLu1aTg0fCRYUczSv/3
bhk6y75YOWIfYWAtDVMW0nqOfB9fmfFZAYAXuGVnK7e/0HpLASJJgxCRUahTD3anla2W44FufsEX
PXn2mmfxfanJ8hfIEJd1jYqs57W0NNZHlygxEoMFdJ1SKYwP8uShtEICsjKQ7O4uSt08ZmdAyVp6
9xAsA2zmmibHImp7ApO335WFIoA2PSPIluc7Y/3dAWNcmxM/noBwwJq0IFr1jOYr3cRZOgjZTg7p
ozC1y9gtJ4ZD0IOpzEzrr94/U45FO9wqdxnjYGVwOWWckfrY2PoGyZzjF1WPGnrpGP+LCZTrVBWe
bHmNZcI6IEq2VRwGZlW9C0CBoHJSvmoLDywljz5l09sXv8Ji6MP1IQNw6ZTYHgfZNOb/xZyMsZtA
APmFG6/DN+unVlV4gLXFQhm2mLQA9OuSfzkrDi30Ov0OlP8CFnzSQSn6cjBU2UL1wkPCE+O7UHcb
Sbf24dN87HV/WqatEGKq30F5yyEsd6uNiM6lPrfh/SotlJWh7hlzHBosJxeQ+6c7nk2+3asy00BW
aFjgRZ+6SmiLzXwe5JmeXeZgS5iB4mORDRNoYywQq/4dX8n+S4svDs6DWI/8U+N+rarWk5uwI352
LvSY6EZuylJb31cQcKRiTro8BEXwYAknzPLt6qFZjD+a8mq8pVqZDfoIAMHLs9VossVc3wQaD5lV
p3bQw4QeAMR5/lqaGR/j3olgZ9FmkMwPwuV4gqNGsP9bJYbaW+e/fgejNPEBEz7sk+Bmej2MfB1v
+V6/O5qVaBBAEsV7dfe5YPqLqWThLUrhMI8nwNJ1OUu9QbA19HlhT0nJG09GL/szrr+VCcqRmKDH
31M0EDUkSFQ4G3uLqqGpsroIdC+ji7DRv5jI+xDlHvbFsbk9kAIahKHFCOkaTkberrPFFq9NnyZ1
iEhR3ivjcU+dtnEoprDypkpYP7BVgipDVpkDqLwrQBPqPHZGs5gnuSv0sbSz3HuDafi4pv7A798R
R6o3SZiYfXEfVRMAzWIB7kkpXbF8DvtINNQLQfm42z9IdymQzsWXKnuMktTM8gyR3e6FKnsmg1ce
br1mOO/X/8dCuVrqaN+SbJsiip08qDNwAun95jKvw+1KiQySB6dtjL2TWtY/R2ioqm/sZrxOlzSj
BqmM70OtVc9QTFoLxOwu0KolPXGdQvNtfVYAa4EB8ch9PF3/akfmTcScx4QIySXgmMGbrciusE7/
w3VbuRfNeXNYk1TwoBMXYV1iutCxUI9/AhKlHOR+SpCbz47rndZXVsmga+ktWWAXcPL9aPp44EHq
gs9FuWd2Y3kG+dN8XN0hwPEBk4lmMqGBHAL7Ou/8yvs+pUJfA9S6pY0jrwLvrOVXuMYaI/M/FOlq
MUw4FdcbMjQYPygsBTQibb5TCxg7IQ9LAtc97FDTpb8RQdYYoJyOjKR8bp3PVs5s1wWoGnxl261X
gx+dBfDEeYlGi4CnBGLTqRtiKW/uCxquLTaEjjAsAH9RGCiPhoC+xtoSmeG8s4EKaJWz/Jbk/UQ3
Y6gGl+F2r2wU5mnuzs0L/mBDIc9v3wUobxgaVeDMxGSGBGifzrgB7NXusJvaDnMXfMkYq44hKEtt
H0PCctd3TBZbL9v892YpnOLwc1kaSXmOEHg5Mk7rC9pfaCWkrrLRw0aNwQ4fXbMMmh92gm4jemgl
f5w5+SRxOEjxVR/IUNErBSe7UxuL0YPpBNZ33rwNfK+h/5EJnqlgSACRgUN3q3I99NO3DdCoYxTZ
BIjptd04TeSzxS1eSa/88n5A9fbdCzYzfROFVArTPosylqmdnT40X3sbmGf1VUVnPigBxjc6vZWs
yaWtJPZWVbv0nmjcajhyO2ShU+564aaJebXrsqZH74vY+Cx4ID0Q/8etXmjyxld3i+cribmHNR+B
oGxe+kctUmc3r345e8Iv+EjADYgfSrAxULybUwSb8M5SW+2qKNxgSBwx44IJ4NCM1bus7Kq0fz+l
uYJrEtDPKFXViz0a5+9yf2ea3QN4D34I3NijPqBzIYuX3EXCmnaazK39JOixIm3PI1odNCYZv+pV
q78/xQwao6gdvYxX4oDmDbzDCiIEPFgE+AgsoZsdRCrK6dzkuQzIf4XrjI67SgASBrhsgHa5ksvS
910/u1AzFCFU98MWr+a+qA9NjyaBSTMWWun5gFKV9oyWtG7/sX18wPEBSa+UUQhg/f0vd11FA6ZM
JMUz+JNemSCBpq57b5vVX2VCP27ernCaEoTphRlIcHJjyMyy2ao76/rQOKHE/81z3KB3h+EXq6Lh
QCzOZF9SFyRb6EXgUlIfI0b2ef+mFPWoSHBAphDSAbhtmyBaO4L9C0/kpmIHDLUIBow/0vHGBY5u
HPO07u0XjXIEiHfAJ7AoUzDylbxVlg7V2y5+mVGcRdQg77QWOhpzFF7INevoiQyg2KnoudDDAL3H
fZM+3vCCt1soCOm5OMF8bFqkI+HmKlXA0neEPrSz5J9/IsKs0Yc0VkRXgxPF6+7tW+S8uVEOSqFR
1TQb8TuS+rGNRvQd+UuiuLyXUGO5YnVdoyFyuf0Fi1vsgFU47H+8RmIRnyWzp8AsCpTaL98ccThe
yYMafIm8bfxxa9kbSSqLYmy1Eza8FCqN9Qbej8ALv0nPwXV8R6QIdX/xuXrbqNNi0FX7cSeg0drR
z5zY4OJQ5Pfi5GlwsNuVqrxkZXFV0ro+zqsHf/2dlhFOLX7N39H49v3FIrDeMDmepiYxT2Gcm6U9
iOnP94d2q0mR1jlo5Mgi+XvePXjiWwzNw+2eL35z06yRYEN1pYGm/v492lISxxi/qnyZUD7o74q6
d4A+OcSTy0WXg2xsj1xj8oPqd+SgSGbTvy5eafE0dlh8uT5dDzcOsMTNDA35w8WgFYwA+ni/8gfv
+ydWt9sQ3LaCPJ+iF1Tz2mJble0NKOquAYAOdhftkKsNIv+0n2UTb2LCVBXT/FQlL9tc5mWfDk3s
D/KWniOswVgYs9egmTgQDo+kcrGel1tG+j2W0vSAYOk7ICKg13mceYCv7regBLat+RHalGdeS8Ou
I2mh8SqQ/wcR7gv00P5wdwk4tnH41QOyFzFrF2isfW42QwM+BBgw5E2qD2xAvwk/cuzq69PybgBP
UaPYNkBYGqjEcOXj4OlBFshzBEf3uk8mcwGG5+oLbMiS+Mi1FNT8bCGMkP2udjU0vq7H5bSf55J5
Ihj6Dkh8RBGvYyMItJALajKqYqagKaBCbxxxEUUnheu180k2XSX7FkgQEztcD4QgTRYQQtWqiVi7
dbY+KRpBphqu8GCRATGQU6nHgxmyV3vgzrF3YhiQrecGcAm9tkv9fadO/UhCfxERxxQZuP5y6fVN
XgUzksW26Spyi9FYX9Qkg+D5GUvm4vxquOQU+8Tl5ajRFca/eoSWgxzs/aCWXbU+ruv4MxbRisGQ
qGSOVrgxv3CbKo/gkVyliYGphUQOiDj51vo2Ao8nU3UPR5X7PjG+RBZMo47Jp31UKnvFW/f0sajA
utcNALJ2We7RY8k2zxbdBFK6tihuT401fAlcankMfE+yg/oQb/qRKqqfpTrOZbM6W3xcSDrdIQgU
6KZeMUotTziafBGGQUlgNAjN6W47ntVbWeezFND/xPqtvgnIpgYvZ9QvCdSrsYrOTNUmWaTvLGvY
0VSAX+ZsLT6AKPp19IsxRk2KCWm2nrlSdIoHlzvkEdx4qH7a3ocf7a8D92TCetW8TfeBvUK+eBpI
gSyBPhlaFJJ0cnDfkRR3hgX01V/LlQy6noB/ifubKbohVxl0p/0VTr1H0UaLnKEC3hXL5Hvkk/FB
SyZlKV0i0yGcnINLHZtjd+CDzBk0lxv16oZKgA6+9w76doGxfuPY7GKAQQ9IW3Bc3S733wx1Zn2/
3QgBfS5keQNjpzYTcN/+UZ2ygh3u/gZpZJtnoI+Yt75T+jlgXZso6is9+vBwA6TVk39BCZXlsPaW
PRzxKmAu6H2FHrdQZOA8SgRdBcPPpgERiezvSZAcL5PgJDwZQyBHKF7xqomM0icLIcesCLiAdppa
rP7wfHBR5JBrrbsnxTCEMhnaM0qz6l7UZEdl1stkpU+a5+I99tCHZDn4Q0hwK1fmqpWBJwkP/Vnj
n316RWkXMEe47dE2MWFxQMzfaPNytSUgqaI3TZWgvZO+cjp7vXh9JTyXj7g5A5IcjM3X+TMpzIJl
4hotjR7oIPCFZ28iHTxHv8o5A/fjoV5Ie9PkBFz0tRHu2ep6FzEsf7Ck92vvYFLqv9Wny5ZbllaA
K+n0WKdRQlsOM+zNXa5wAKDWd8gHf3e42OnmdempBxtem5mRbI6LxIKbwgC9jaYHp6X9G2NG7Zkh
9zyxH7eJ1zuxip71Au30ldupDF2HU9g9vWDspCeXElRUi0zJR4jiVscRz2EoeAmyNgCb8iX8bwbB
0k4x4fMqAJ5z7pb56GO7F0twK9ylTpyQZqvWZFTNo0U9n+sf6VWCbIN9nrkhLvjBOVYrSBHTeFXu
8tnSn+Kj4uAH1SbYanXSVDmCogi5ZIWrW/WUEjlmOvwv5pq0VUcFASj1bq5fZ4BwNnhisOWuV6kj
3L2eSP9UXPf4RSkd+rI+7xri1HbTBj8tB6IspNrzE0RFmpPoJLuLDc2Ok4AqNKcaMPQ8qrPeuYHS
DJtfG+wwaZ2VJq3BcESnr5McVTEo9lP8HSe+p4mjI5XiY/wKIj5g276IN+Gybc80/N7YALzG0yCa
mDIgoaR8DnPoRlJa+wo55ZYehP7Z013S5DOgR7J9cNXT+47ABPv2WlK33TPqT//fryIE96skS9p2
iKhVRsWoGTfHXRtCA2OB7VjplQgoQDIJVKhOMNSfBBW094OiCjD77GWCve+QfH/Yz0jlKrkjl6SB
mnCSarHi961VatY/bLPFkY3wUhQq1/NZCSM/pzqKClLKzheRDYf7A8qvBFdSG274+8B124fnEd93
mIAt8Xzlb79htvw24K4Q8syAlc3NYa+aU5OZt72lgvbYVt9B4+rxG2ywUDQ+TPofPAsimQOgGw4u
2EpC+CYHanvQWqEMrvtXq3Tdv2Ze90TexxvkLubNXJa7ABRJjfDImZ+SXejYABITsQU0eBe4lf21
2Kh5iCqh1tOjFhnyzULzYEnykpKS3s8lfxOgdQAjfxS81+PD+jJD2lxKU60d+bxcOjGffwz9IsPB
esXnCmsVqVoXJvwi92R1SjLAScFAsR6yR4GFsTMA4bNeByDoAuNQUuiZRXh2Jh/DFpHjPYhEcTCG
QIEtGX083F+whfvvHDzwpJaneguy6Kae1PqfLX0zphIMp6PK6iSFF+T0T6pu3s0d/iUzSPn+RSig
IAOT/Wi6/MtJjDu5wnj80dt5K9rk8B9Eq95X5yXPxkN2xJmOfGYLa7eJ7T3IRHM8bkrmkcsUoxOc
m+JlX8m5gxPd3xT0S4kcvDgVBqmoLN8jmHGfWLq28x+ynaxBDy1S2E48E4YKQvP43GfYeG4YToM5
/Jf48q8BR6wQAMNE/qikgPeyt+rFL0dTyiFd5r7XqPta4HZuftByoYBVaOvXZOIoi9TWQ0ZkN7DR
Gf9rSPHNK8156R0gNCjtPmeCTgVqOus3eLMPRBmTFPbz0PoDRWr62/EsatiJky9BLUXRI+ynrVr4
jYVrR4FjvpQAQ6WHwso/uifcD7KmSE2ObXrrXnbdF2J3gQhHCDWuPutVax5llpLS/SX34l2YbU9R
nyvz26RRlAkRTa/shgQ1lMbqXmTyMnfq5i4/FKs9dxlazg/UpiKgpDBhL2gUXIm9d1Q3Ryr1F/BE
4+exQBP/ZDSLKZEtxFkHq8e9t07ATOgQdCnd/GPnM84N7KYCDAYBUm/h4XD6qism8FrpS4/rk9Da
2LBFt3liQK2YGY3TTw9i+bVxdMw7gsVEQtprCwV3Y96Z25zeIo3SA+OQ+8L42GXnhf2QN8fcdMUS
eSXzED74EQe5zZeV1ADLx5T57Igs9NmAQ+vVb/g+kHPqXtel1hvtYqXNlqRjC+pYHQa33+7R2A4c
9JLIlAosoNGV4XbSrkfoXQWuCc2Ka8yvpsIGnRz0B5pKEGUVlVCDpkECRkb0NnVBGNMeJDiIp1IW
lYnBrzFLNuuAbaY8dOj9ORyLqSSJnpqPM6PEHR9aVlXC9OksdOwDaYN0OY9BGzjUxcPVlHAVP+M4
UqFaoUHUaCPypuwvSCv0CuelRNbGYSbg0lAsirVPhVSNJTo5+h7GGLOtcPWntU2MDUuHRe7Ptv2S
AmYcQO7nuctVRwfxHHf2TuFjYyQ3cySNvbbDJqkqbutYkUhcVbptAp+FooVMpv11aHXfGav8XCud
qi9qUb/6uLG4CO7k/gz732zdFLvi+BI9UHP5geoVqQ+5LR01OzSPWCdBL8AW/4rq8FcyXzun5ehx
jygPcGqXER1Cf/Xf8WxeuD6PbpE+gcqDijjz20eTZVfYjBE4wTiXCu2HVgvK75hBtvRw9R5sLPhV
VL76oexoMNSsMiREPX4sFIgGE6D1tOWTpf00FVfvPTopUlmQLgBuH/V0X9dWEBGc+xsLieZ36CXP
O9IGBBeIGTdICwwNEQ/dQ6441I8vFxxgLeAnnC01ipDS+U7P03sgFStyzvVV867cp+mVvYU/85qx
s3VRjXJS5AkQy/rNWdnvGEuVxXndmK0OuX/NKPpv+A8bNisImIXhO54JdfqnIHKuXuhV/nqgZAiz
h5UrNgzmlf3ZoPuStZg6xhRyO8//vGmsw1YyRx8wNOPa8V+1VAFHDBwLJwLNonZLrU4doD83oGxp
9+pAK5WdNIvKH2jZC4JbSMs7yTx2tDGGgKQjfdec9zU9kxyPu5Z/bwXs2Ht90Ryc2zGTsaqzN23n
xgYhCuRt5txzxED/lswgSbr8TiUcKJTThYwnXOQUE1mD9Y9e9W+nXIXIHldO/ZJRZGEL8FUMx9Db
fRfFYivtgIGjdl54Wz4PwPpQ8Qw7bO6nO3QUXQdOvv/Rd64fH6SQ7ikIs00LmticVCCXTiOLaTN0
rt4G2AE4TsZU1VQlqdh4Xuhi3jH/0VV+C196cxlF0yMjHHFkBF7+foARE+aOkfx6DfAqSaMwLyTF
5Zxk8HuZvnJcWCTjniXGE0fgJeyFnFgrFktrApYvCoTD4Y68JrLc6DJns7zrgToOxu375NfFp2WL
YQZOqryJlyp84u2Xoc7jawhl67tnIG1j3k/h1V2nOPZHtO3vu4jw1s59YhRkBx3XGLKb8aDl89yK
B3CAlkLpK10WPKhfofRlqXy4JOZ/Ss/vYpN341NcrLhXzlyiRfZ4nht5249s42Lhd7zfw7jSAmmQ
N2zhZMOBtno3m9u1ll65UpnJ4b9lt8eP6ceGdVJkWfV/MqhKMPys149ipKMqgU9ITM1m0JhNS56p
IHukrJkPa0KVrBs32ZNKDgj/1/7nLMHpSIXFC4YIyX7dRlraIRbb8WQjGubPqYSjbA8HbeW1tdAr
gg4cQk9bKpdZaNtCdWNnXJF+XpTn2Vg/K0jzA75Y+in9HvH+JzlOebeQJjR3fBuRc6ijYlC2Hoi4
+bh5i122riwR+dCa07OhROwuS+PFrRPomelWqTBZxW4nK9EIWc59Y3BggHGzVksrnf1t7n/ovDFH
o665EvqDffda75c4EW+AntPzc5Uerd3NDE9EOw10PSJBR5KX7/UN+TQotovFBwusw6ZtQ6uPxUFN
4PVkBYUddj9halZh3xi1R8AXM0fHMEQWKTOzTDU1iJD20XGojN//HqHIX55cF1Y/f3iG4MH/7m/B
exkbuJjeBKxCVYL2Mhm60dq6lQO9yVulXTp6zP/jevmliRw2+2cq0VXOyB/Njj95vK5QqIj21ed8
jKxnjtEIUpMmwA9Gk0g32RueuuwXj4t/N3xOssqz+41KBFh90CjNN+3kyloOOEVu2ClMUkpbgXbl
I6p9/kci7R+oNA8Gi3+mcUxWWmk/tvS7lOSX4meEKfvm/HaxoBsWM4JZgNMLH0OwlhcN9IgZcmY2
Vh/+ti2ZhjrBLkhGwSGrlqTYai7Sw4uiwbPBnVJSFipA3Tz2nYNk/lFF/2yhf9j58m0DGbbUFucq
1ZjUTSWQDIhT2LopCSNnwH42yO08u6wvPLCXrouDRWZQBpnho9/ERoJ4R36uRn1e3MbBhPvmmjwn
jM22wYVfeXVN2qjPMOY9hfOd2nJ4Kg03UKlXiIH6EfoMERFkyP5234muGf/8Ywcn2lbovRkdnntc
Moj3MkiB9y7clJUNhYWAJlFTQDU78WPLnjRNIFodA6Kl/nH7PVlXB9liHpge/GkqCXEpvC/EV3EG
srsLi/MWSQIpEXtyZ23raZT5Fin6NR7Gi2IosPPdpr8Pwa0l99Fqlaf0ulp3k0hvMEMcFCVKo/PE
udq3PQoUPoVQBgu8c/bNZ07jk3TdtswO3z9TvWzTZ7kgnmkkdivp0sUHIO3kc4oIOogPxF2Jdf8C
EGK2sKFQLsyYdjdfLxdHJBwb+faDx6tlbmBVSu0NmKWdUjkWsgX08uTEa23GBoXaLrYwrKLA64Sh
V5ZKRriM17/doPPh/wYFMx+JRQaOKp0rbgPQYtfuVnQGzn1gd3cGS/2ovcUj6bv8jRjsLzWr3BsO
9wr6Y/ZO5e+ttEb/TaONGnY8et3HAsXEBbrAHWu2wG1nHL69TrSpWH7xrqn2ZFABemOyyMAbrPVM
z97MXnQ+M5bZQtYHHcCFGzT7gJ+ZU1+J/isU/HUKzoXKooh0+ReWf3Pa/lgSQVa//d6lJnsCmWZh
TD+5v1eww0tMB+o9PZ0vR6weHYWGCc0/ydFtbE7heLq/wJNQ1oCCk1Q0KublvLyy994aS0JCq33h
J2zCxrsdkoAxucNWjoJCs/oXbsHcV0oi9Dcnz370ho1Qedxx77//ka0Mr6ParK+p9+5le8wSNKhQ
o3sgKWA9fv7b7CjWWi45ksRpTPmHur2FOhToGl6LBwCthsdun31sk8+h+H2zDy0Xuz9koXTP5yty
IcSEYIo3MR326jsvf7rMkkSNEsbVj3xoGNwwmIRJsNE5N8/inovyEwj+nMu6NkO5c3dl1kvaMkx4
IMzOdlNpeOaMoVkKfX2y6SzWm27VT7ds24eFUGlHd9RkdF6R7ccLaA5fj01ezJAx4FidZFlYi4hU
/W9NNIQW2ImNs75/xy9208mUagvkryCevOf4JOhV/+G3pqtK0iOlkxJyYsREVqGIb76EqKTfVltN
Hed0Uy6WwV2RPiLDAUMO0P/+1e6gZ5AgL1FMARlyiyZLnkC98mbXTPj6bYx4hzxpZefwB40bbU+6
Nf2f2o96wl22iNNZgWqsS8LMBmbEzpIQO9T265P5ptTRFNPlx/9ieSjqvdzhwkDctl50XukqQzOv
0Vl9WUe0ogbnxoXnPFI7KeBSyOANvZuCmbWWIxE1M8c8sK5Pw6/McIX3CfvZg32qH+piM+aqaltw
ePgQ+v1C0Lm27YHRDPx1XydVYtBQ0pb2kSCenpnGeA8Qnb1f3414AdX1hHG/1emylWSzKyX8a28F
owEFpkr9tXUQ6KAf/A4eoZHzdH8nzLBGg3rgYfkULgL1XsackoIsoHnrQiE45qh693aZJKv267kE
VA9Gjzo7Nyz8Q0Zdw9FWEXx6rme1oPbIySD3+TRb0SA0kg0YVuvBKqzP91IE31/+RfU8itqcVI4n
0uO8WmImgmEDqcAgzuLHWjuW66fki0N++GXlLmCoVHHMwciz86Wjzy4Q2AoaazB+lp9Hph9Xj+Jt
JMHyHrLLivNutKOQBBeSJS7WfLyJT0WKYFhnbqjcPZ8B7ZoB9E5nKMs07pl6CG4IpGfz+corIhst
oMWn2M+iIGoJ1p7kVXIRwhNl23BP39BRW/v0jbi+M8Btw5peu/H65CHp4JPVRGZC6GVOPrOKrHIC
8zkuWyVRZLrzZsAmzvdp0b5mXXPabTNZeGNUijm32yILY0IJMu4xZW9eQKTNAn4t11KnQju6tWGZ
U54XenLcOQ7gz00gkJk5cZTOlJRNEt23LhXQKQX6QvfVGTkxdRGp7tjQ0Fpn6xcY+uYI/dEMm+UC
DBqm8gaUkEvAAxR2S9eYWH4AHCWsky8poFhUx0+IxGWJhxbfAS0REVnazeDXaXxrDbcZN9a+3DPl
r97Ekd68KnuJ6DG7uMc4eur34acqxqHU36FqXIkf1ASvlS6/wA5hepHU3EQPe+FqYadHk0sCmG4D
xzY+GwKgdoScd6g8lQFwzGefznouPhXjVpdAPx3zRIpA8iulaaXMKPTdAms/bohBFkxwwvaiD9PN
AHdCA/+Eg1bSKH3uK/ulnGZS/5PkijkE9lXPjvb1uKwOMMQ9geK7Z5ZN3wyyybrVk9NnYUxHNnD2
C1iiVMSUGbtrv8PwlTEE3yeZqan6UY+OOpPvW3Jq915pAjIQJ3qcRIUF9Mc1qlNHcWdtk6pgGMHJ
MngU2yiIVJzQc/k94esE7kzt3TsZRqt4R5gauev/KTbFmYd5rOwRxDt5fZNvqYSp8DKV9y0BXhUv
ko1pM9PrDL0B0Wp0tVD1Pzs7j7Lj2Oq+14D31j5tAOP3S10iRzD6wVsFzD9MKKq9jcopQqAFMz3e
Vr5ARwly9zJkLuyujWFG6Ud+52idja1IesyxpkoVudBq1U+pbE/MwQ/34B4S3q+Fdmuh33pzq8X2
WA17hWp/eqXjHNGxSCLddUPRoPrM5GK6I6HcNFxgOqdliDaobdHmiP0dNp37WMYnBU0AyswydajM
Eszm4RNMusPa1VKYztaoWA6ZI/XeY4N0OtTR4kujMOPjmT8vIyfTa5k6wmbA+kjA0AmyCgVs7vuz
QeTO93NGpbE+fEaZZxQ3Us9FlAVXtkbKU/cwV9ZfkI4eg8mbSL5EiamMHytvxj+m8aDCbmYF47c8
l1yHFb2BuKjj5tQ9mC9Wt5BT4JfSuI/lvpgb6q4t+2VqhfVlBaF73HFc5TrgZOLDtw17IVQqAy8k
c9XJGKO67qZgFo+ba17Uc9PtDVcSD43vJr629i4DDANbAfFLH+kshWl9A1NpEi4aQ3eqWMHLMHK/
GLnwelPA5e60apjbcPfQWyjC8cHxZlqbg4KUwkO/nNIV3FSHqcaN8Y8Cfcu0tB/7cSCvTg8P14Qg
xeS//fM+dMHUCU2aljRicv2wjR7dSt7kvniNknCNg5+DA82lvzlpnWN9OmO3jLgB46cXtPO8xahO
FqZFSo5AwC42LE4ZFV2hqDS4i0qSaXTj6hgmL++Z13twcyxAu12vVkSi2AtnvETY822QNvPoihM1
UsmHSFRg3N3jlxVD/BEXo5Xt4a+T/3V7/yhJ47FOIrXjZ6wrL/F47cmWYovXD7X0OOOD/QpRu+t2
qnyqJDERET5Hm0guORXlnw0rWzxTuesiag3SgCZgTxRo+HaJm728Inr0IJOD+rwXp1aeeQPDwk9g
rpg2z/mROOurnMrnItYS5XQHI3IclxBD5Xy8oD2HRHJVwwmXERqhKP3FbQbv7EKvrvllXXUsdOlG
MTRG1qCYL0UJ9qWolsaSTTos/Lcf3tJ3mZi3dQQxClSmazZmWoeIcdW2uLUMgYlSptk0ysfm5Gt+
F6ax11QnUR7ueFjRxxyzgJHM56LsT2KhaTadoDh5YS7rlop5Z2Y8aPZjYzAa8r9UsqOKx22DhbY4
ulVleqqRdvUiChCN9iJ67djdG3Wfd5Vtss0Nc2ToVhKbSqYIvS3/v8sw/dN5weqM+yRg07DFH1sy
OzH+PEQVDfimcOv010KGxPqXJXRCYapGHQ38tpPKa9m2lwagsXHXGrESn57+jAi3wa95XTfSZfbc
yzuZtMNhLSjPSh7R9H2PrPgwQmJ6dYvyqozazAIME43R3zaYEAvY8YvO9yFhxhEXbLcxBCg57UjM
5dfvlspVuDfTc3CfBAe68kfgKFmV+oW2NsoWAA8ELz7TlLamUKugKyEJW49FONQaSyy5FW9hB4l5
iWZy7VEYrTJHHdz2aHtBNgwoPGwlrrxSe4S64UjDp90t7lj41Dt5fVkNzDLBaMLMhai950vTGffk
uy6RV3noYyetxfV1R/8UKlMb9DCh7Cw14J7H244gEVin9oJdGLG71HBAoR7znQZtH+k1JyJ91ORf
2gsWWghODDZ8kTURCihcEaEI0JdtOJ0DDkRjhvM1cQx5HaczRQGyJyEd4ONoMUJkI0Wl3i79eLLh
U2WUiGmZajFUkwimu6MSvhvdjwCc5ZzFMDvKaM/NntHE15Lpsck6FIR6Bfwzr4xAvrTa2oLHFFUY
PkHY3GwBXt6RRA7XxnR6G05roxS0sW4kLH1PTDa6j1QNgpIQXYAh8PrvnFBTs8oqbOFemZzRW+QN
twECUKGOCHgCo4NRiri7HhCzaBrvKgZTFs35sjnvSLE6/2OdVfTmSPyEYGetmXk8zPlJewIDmdOi
BGg8Q40Mwle0fJ+Y+zCeUJ0tH3hXxZA6EUYkHCvkfpXiIXGR6evkGKPzc4k0mTiOLWKsJ2hgCg3p
b266gYgPqVlcY1CL52oHTs96QHkFjW0L3F/4wjbUurjp2KuePfbuzXfllpZnVzmgJz27OcRLrWCO
ySNa/H3gj2630i0XYfy+55HwF2wuJmXAPFDIrUwd7gYcnPUVCosZP7b2Mz75I9hqRUsCwxF8GSjY
b0VyMoHT4z0YbyBBRjBTPaZ1ePDzBdf+PFASuhGYkObVfkYTkiYFdWiH8Ox+xgX6BLettUVnOEz4
NowDeqP+K84f4zdnxAMBFkRp58nbWgj+SvZ4cvObzl2gDT/jbc12D311zitj2J1qWLpKjsmGBgXa
8Mee7GKo8sAYoXgX1sKl4Qqp3F08NguYHbI2Y330G952lNJndudM6iYOAfJBFoICgJCjcZfn+ML3
VmZnumtRexhrTFX29ddJCX2KaKkTJwgnVlUNcXH46DgCKlX0t+P80I5xulEKgLCbMzoN2PA+rbyJ
ESGv0liWGn3V+CjG7Lj7gOiYuixduzlf8wV7Q0nJuUFs1tB7F6yRs6Id3CQ57PeKOw8M4rBvtvMv
RInAmztvdJHuddYK3avCsxtbqNdzviZWknVCQFDnsh8BYli3iePFFw2lvfLxRviSbn2eiW6AB08y
ilYu1W/3aRXmyc0heMPTsUCziV84c3+p6invBfuLACmU3Y+EJt7vbbE/3+TkBpJzDRS5kHh0khfw
4dmSsWSl0aTK4DmZcWe7euoNRLVmbK0ahJWyQSernKHCrCLDYYpbs27Lt+YENP8pvAMV0YC4Iqy2
yjvX8CEJEQadac68qBYCP3ubGN5wnQ/eutwG/HGqgoq2NMDR6TjQKUWeKuaAgQZAusvEB+0CU7Lu
ejWcnkuheR0X4h0xNmtCkYds8L7dDCsJR8T3CAEFGYzNTVwWrotDv0MeQQ71D2UDH1GtHk/QG/s2
wHcbi2Im723+c6Xcs3C9kNoaU22YXovwPg51m0j5ESZOeNrtmLAYqCRjVpLMBkdqCZu1KNba06iy
cTF4oCUE3u07qjh0w03I/S9y2F/XtGq9ppqZi9I/sh8rlm01Imui3QWcalPfwFfwEAiLMNzLWSek
zK6B6RIHHy26vj39jf4wAmDQqXAbf9azAwux8COk93SbkEyHry0y6ss7jiXJixY/5q+ZQFsTL3uL
YuY+MBm8bjaMhaniIoNt12gR9L23w5PwAPIv/RS7piUcskTUHmdsbKtWxdKgz5IYvU1pQxo9ASF3
wbtbO6gjOGNNY//x5FfK1+zQFP4vDKEju9RJiKyaN0DwTZQmVzv7h36YgEZXdkLRFhizm7Sqfe79
cLYDHDbgVG4cd3VLVgsIo1crK4HXL3L+5QGhRr+Eg1vylPk0YI8DSjg8DAZdQGzd/6I4BdkN0lI1
X1Fc74a1ZNBTkafY3kC6Wo7qzAKDKR7TURFgpKNI48I9oH8lgZEOJ3czv9Q+6YjNlV+ni40jGXNd
dP6uRT3d56pwPaLInHRZsS62fjRHMFDjzQYGjEDS145dll9sVMO4mH7crbaeA1zm4ivxDo/xY+4I
/ot7OntGfrPr7WIKbYQBgI6k1uKaFL6sxI481eomFvHWhZ9idKoMMs9Zcd7HxfRct4maTeOdIimQ
DKE/r9vripbbwBeQ1wxfNKzBp6EEGTwRSXeOc9eyb5IzV/UcTlP1oMecD6u8A7FXmaFYvAzFs03a
jzvQPloX3pr/gGPGJSeDL17Ezn7eZC/ML8+ikV3Yrm9vfW+XTJBKoQMSpvFCWG2lkJBi/FSVsdUd
jZtuvXZrhg2tLhbMcxPuKwbrM0a+gAYC6OSWsYu+0QQqS2fj2qAegI8DbK5ylzwF0nN0r2yKzo/k
d/qz5miZp+xcAfn5mzUFQUITDXvbO+z6jyXI9DaKP37YTKDyDM5dywqDciMc8ns38P3RJWL2PvCY
Z2wRbOXs6F7jj9lZfLtaUGqjzRl1GWEoi0i93A5v9KNYV4oL3/VRbaQ6lLkXrT9oDyOEV9UGXTBD
xmF6llqkwQozpQnKqPCSfPaanKEOvxvy/hPFreqDnPbrwRua59qioun/N+pikJIeSU5YTybrJohX
AxXHRqaf/EEQ/tf+94UIYDqOBmaCpOwjA70U/XlQeAR14BT6MiIJtE0ziRSYA0IBQZ96vgiUDV/c
B3aTiJfPSsmPaIuo9fihuB61b/yJ0K+5RCxdQtz1SqmvfIGZLUUUTfkiEWcMBvCqF7PTKVTnNi8r
5JISY+xQYkpcUPGAQ37fdv7RvJzNTMlJj6KaKE0kRg1vKFwmpF6UHDOrOLA3nf/1YI/Sl1EMR/LM
rnXWtwFR683UFVw8js96+DiWkETELXeHgl3WdOWTPdGML2edjqSAXQ5YyKBm0QXZW01gHH/+/M7N
zSaftGnT/59OyuCs6HDPV/+KKLPQfHfWta53DYmJPnVinf7vH7l+DV8apyV18JyEUaY0h04mT93K
Koep6x/+ANqjPLw7KwhqlqUYY/8fZvsjkI/JgZ/E40w0DSYS1PS9nv/BiFJQIRJrQW4yGIF/naYd
QXv9Mpns4aKAIbZu23+8qoRhZeh/+FWkEM8c55rD2pgg0GpEOCvCwNSnuW0SbZDt1zr7qZUsxSBB
LXOPYqGT80WyJC/ipNIDWBFRpwzO0wMMxEABovjZT4mL0lYNY0y6iJ7evYNg7Ci8SLb56cEOIU/w
7Qh9qg7G3jRwppQYVXxtIQBr8GgT8MOXsIt3fMjrGZBPyOFauu0RpeYrmMnYikG4xPSU9h5U8nIH
EBWi70CyzYuzyHfNg02Qz/7YnDaiY6VZZy7ymAelcuCC+9CDgz7UsgmCWx2pbBEYpzugjKsEUScA
tjXqLE5v2akXA35eabINALTi+TlVp680ulVi46oHv8j6gKbg5+jwdQe3WP3nIRsWjtKGMTJgmWQF
UNZL5o9y49Zgbnu7KiwKq+9UeNtXrPsP83yaxcs6DnL0lgTcVO2CzE4Y0CSwM3Tg++Zy4R9ut7v1
yDaj0IRId8rSw+ByPSP8Dsqp0T1SxyHK2SuX/YZ2IqKxuTG4YbWNDqrKy/QtNKdAiHqZ22T9Ivc8
AtQIkcj5yBekIXXw2C7HE509Gwe/YlzPuECUH3aLw47W4qEYrDS7yScao7Oc/TJ0/kA5lip7B0qd
zlQ1caNe05AcKG9GQIaQlQmVBqqvlMYQgG4dBYKF2TN8+EXA/jyq5VHYBYRo/THj7s4ewuD6VO8Q
TQ3DuuhO5YMp35DuOpOmjxSQ3jXq64WPmFce+C8Wkzc3LzMWUuE3CmHfyeD2cVemsev//0UMtGdN
CMNI+2Wcyb98jrb3RtJiBOanQ8617/DoTFsr5XqJPtkVkj1CN8Oi1uHQ0pZfqmEuVagcDdiGhBgO
2k9F/zyV93GZX6TgahgDS0Un1scz5Rh5Yz5CqoiMMEOYqpyrrEoDkjRjVVOBj8phHQe2Ef/86tqQ
S5gcbUkr42Y8f9EZeltorvjAFgjd2q6PxceQxcumxyNnsvD0ejwwOqsAyDWfrA2qKJm0tw/lhmS4
7Su5kDgSwjyLLKmR9zctHEO27Go3solgXYPdO1lTS7mC3DQCTBQKLGeSXmS9szcbkWBTJkw/TR0y
4BMjV4mrGpuZ4pu9rYmCZGiXtnwdv16PJtaqwJI2e5W+1JpvAOMX0X8NBAf2I5REyXtuCM+EXVSa
8jB5S3kULVrnkEa0LqAdVgdzbxb5py7LjCHDYNiFFF0cKJL0XX1m/vp++PAJmc8TOrzV3RxqlSqy
4kkjzzVBzybkXvBsy5hEa+QaDzdgyZ7KuEULq5MamII0fwRz7Obj1f9JIDkfHnfedI3kXUIFA3Pb
PfxWv3cBsGrFjgQPCq/9fT8BlYpQUsUylzbNzeNejRFP02KPkawiHs4LzGsbXWnHmAmsqfj0ahpX
1avWHmCkHgEuO7rZH2BKWXBnSQNdM9wXPON/FH2otGJaMnP/rfTWktg9NaXzc4xkiUEU1cTznzHW
yzzGm+5jiiSa581r6T0Fs+s0TG7M/5KwTAvyf/R7ln7ZZBU3TSOll2ZrS35ifq/LVonJSOC/9fZ5
zhCpWCXImJKJGifhbjXkZy/25AV7+DWrS02gZBrQ8zXJjotpfBT4GXl+QVt39S5FQ19QTS2DXWDc
6pEQk50KdJTk4w5uAITkig3DxlHk70eHcpMKRy3GhX5vUD1G3AUVXiXi2gZonCyQxbSZJ8jvC3sb
loCQUXaqCzufYrTboiuueh8SQluUAjkF8nuqEB/vmZ4s5EbP/g2tUXjW3mUCbvy4CSDTX3RPZtCy
444gm/eV/3MMRHUsQ4GVgxQye99g/rA/6F+5Si+YoPwJvhtqxKfZbZCHYxN85DmZcyD/jdi6A+pJ
I0T2uuQhEghef8nZK4jBC1HbmSKKvVn8JUkCMttT48baG2ogAq+jO3N8fAeGBCnz34277wLS2Rdb
CIoMAKgyiyK15S4fxv8dkZGGratybELNF6MUO5zuPCIRxX4q6f3n9bP68X0CUTrXNbexcqwZb5cB
2gxeWFysW31qIyK7M6BrgW84tn2y46LGO19sMZzin1+G4RZHIE8HwlbzOjppKiPHNG0GKPaZcnn/
ZM/t9cTtFBM0hPZQxPxSUZNcvs6ZoF4cYqVzYuqW3OYSR9Fpl3b1wNExJz1Dj8EL13PXtHUy0yPq
TCLCX/Yvd1FQ/LVVtRvuRTI2EZc2ecnDHJ1pp/bpoubEhHx1Sun3QCjSr/IwMJhF6gY1V/+tbJIV
5nKzpowtYnw9k/PAp3N7cyftlGWk7sAiMKzF+LOCRpj2pwDtu+WFBSHcY1GKsKMr8bsGPyK4deMS
NKwcX1QM1HQIw9nqq2aTiiLfywiizKQbot4rfWd07xFcBxPZeGaIpuhmAvuYK8H6WpYwV22Ad9uU
JlA7bkncu3eu17Jf+F9JgmJaOyA10M+vJ2nqoDhC0y7l4F06I1yCrQWM9hReF6r+AjmbnJZzSMT/
DLQzrE7ox4u+SOeWoey6PTkQbF7scHqKreeTAYiNT9zjZGbGY6CV5wDj4eDxUczrarj7q+yewabd
oTxKCTvMSOKOIlTWSBtx3dvu+OvyXYTXsP+QWvgIlinRF/xKuk1Je8HTHhcTz+bmEVOPodhv30Md
8cCWOW0CnWyf3PNUWOGCzN/4oZAGWtECkoUZ+IViYfij96+0s7e80YAFaiwQdjO61Adwxyj4NnFX
jD9xb39LM9rGF82RoX4oSVcaBJgx7CZ/5wa6rUecDT37CgsHOtEqRWHBqP2iq/KG/UUUaT2x4HeO
j0FEm65PqyvJJKXyD+AGmiw4pnr4sVuHEuWRg5/DALCvLyDND6EDyVMINJYLYm0mD8vjD54UKgnS
JpexqJxI5znudFEX87F1j8Ul6cyOv5ciCadEevWIMH5U1QmUQ6nbLsgcDyQvHeaNOM10V5Wcg8gg
Ygy7u7kzENSRz/rbtrlb2PyaLYcW9XlCkuTN0Ds0s9ee7h6KKq3kS2wjV6xt9enX2YJOJkqipmpZ
vfPOiYcTwZpN0B+YLB3SPZC1Rpk39g7UhgHjeYncR4JnD3hwYtdkKG107y5rDz8eoe0qT7DT2hgq
QpemIh8zGSepqMHybwLlyWDOYapxO3C4FOMSccwVjA+g4phlpxumT/+mKPYkPzbEIKSbpH4uU7MU
r7oJ6QaGEpMHIUi5P16hKgzWm8pT0IKEZwNsVMgQAV5XtXmyHjalcxiVQjFQVKfRMf3ux7XBDrhG
kEYW5COM9xH/KDCKf0CViaO4+7xeBhMybiDXqTk3/JWFBsp7I+Ql2EqqUoPyzaQjBa58GYJR6rtL
xtzac5U332ZSKx4zS1Bjkti8KDLXyr2+mDR76v4iC83JWaIEvNxhYMV5sXHjk2TmxbXlBCBWISDB
njUYisr4C12s5ZoTDAS7qcLiAmcGmFyKZjOj2iKfMuCEagKJvALQbujnH/F6+aAhJfaKMiqUFEoT
MJ2qgzR/pXIQV2dqoYAAXr7hiqbjqF18cFpHu3JmOAjgrW5ISCh9GeOHwN20jUgkDroxzhxNh9wS
fcm7zX8WH8I4lc3jxKvzU9fSdj8ni83GYp1Kpt9P1YCoSlFRCRLT6IZ+O2m9fckDtSks8THfTkYl
AtS2LfYUjPaFcIr1wTAeBEcvMQuI7mIi2WC1bc9zZBWMcK1fwrEgcUA1stylxZST1Zf+9pT3ATH9
d6pLS0UG6S26W/YRg8IDDCFvKQQCfBFwknO24O6exXvr7p0guwmBJu+NLaf0+NDflSrkwVcAsHYA
NF1s76+F+xsngwUGVPHyLYKxT70UCtOAh87YLRdiVuAhp/FP4zsflWDZoCTdHki2ZGJGghhi7Rqa
0YNJ72z7xiQa8eynoG1NrlIB9Kk1r3v7dsaFCM/gMrJU0zuL3MX1OtYJ5xPcvzRCwH5HxgK/6dcd
hTTU7w8vttmhEJ2Y//BktFFuxCQUZgT/DRkAT1563vZVfNMUMe1HPyhN/ZIWxKWzYF5XcI19OzbG
BFJ6BoMzs0l8W+PjrjYIO4ldYm3Bt7IwCAo8L38YNmIvbekbY2NC3CR1p/2SO7nE0xMdWl6jx2VY
TdUKQHYd+rQyzsBpGOrtd06HFp+ZiZ6qtRTKha0DOZmMBmfo96rL4efUVgYbuUhW7zKV/ollljy+
9XChqzawGPFEu4TUoOmNyI7aS7Ozc2W1NzaZLcR7a5ysfPrelGgwTRmSgpXCg9Edot4uFwmIimSq
0p2PadC5nwW+ED93r1hwMGmX70Uveb1DA7F8YDirUW5NWWgo1bLoLP+r+R91CzU7uugAxca/ASMh
qEwvo1jy9kerc+JfS70mGlzz7mKW1etSeA90T7BPUy19qZc+WOpJ/9CXw1G9e+dbUb4JTbKhiarf
MAjKPaRitumEusiOUep+6rC3Hg6i4RiZHYW34J2/oy6y7M7nhi0aujvlrW27b/FRyp+HinOL84ih
cSPoB5zu7J3hkT+N+Ixspo9RT5o+UrvwL0KQnOCJC1i8Zmbl7rybRb+pwZvZrdf4TgknUItzuigL
kUdCKVqHnrz/Q0ourqYrj6cmv5D5eowIsnUbtJZM9Tnr1rXg9UPZUiHQjJH60pGDGfUx37ozwK+T
J7F2zeGDpZhxuPrX3SnzfhHqI9ZEKY7N82aSjadVwig2lflcO+f0GcAJCVMtX8UAJVCOGTiuc6O/
NvPfgumV2rRtsQ2kojRCJxXa7bpphJaUnCMPss3+bdNWxmo0z3C6ZgaPQG6XPexJj8YecZsnt+YA
hBnPhn9Lp4xgb+kuWYSFxTmCs8rIR/J6AXZMk5dIvgUotnlXQ/5XAded6pD1eQMblBbx59S0wHlX
2gf6IW++/unhMXH1M1wYuoVNdAvmgiUdEIp66Nokm6uXHy8QgpusWT/hHCYqo+OsMLFnDrFrEAoQ
nnk3o9pWYfbl634Sw5EyO5Q8aZFFsT0TwxFNZv/1ckfifxziSmAr9APISx1gqYprYex+z8iqZc7Q
wa84sRqsCvhZcmQsxW+mg1vpxDj043WFhfBEwlKXMPi7UHvjdZoVNU8hA9ccXO/KXpT+OBsztLsd
hKwR5iVwHqWgSoombTXlGSTgA6cH6/d5Y/IFBqPoDU8thDOAOdZ9017Jn3eWEywj4mSPCeUs/+OV
unknjTxIJQXEk9eA28GGjpHaMRXlU+xFOmHB4q+REHT7NThzSk7NpIGSCGEEgxDht/+C0ns2yC1m
w4RPGphqCA0D8H112Y+qkzkl7ZnGGgMArSXltyA9GYcrzMxF5b4oBqCM6Nk6RzLuYNwPJ+lPe8Iv
EeM2syPgG7bh3yS26cNfTQl7Octf6nwdTIdwLJx1M2Aj1GnRgWm9gYmL+GC9wmJz4OpCrkcWjyXB
xcyBxd/eCoJWDGbwtBOvOrD5NlPKs6ocfvpCHYjBmHrrdwCI4vgFScZYEmbQaa//WHC/+WtwUQHi
SoLb10ORM/c91RFx/hmoPoMasHwE/fC65Rgm55Ltx3hNuGMX1FJUStZO6ZGdScxDHhfIo84L/K8J
NTe/GeBePT4Dowaum1002hYehDRNHoiTyK41Nrw99LZE26HXZoCR9cmEse5UxDelHjtNAs501nkl
7mRtMH6XVnhgzJNG5yw6RyD0f/mUvSY9DmQ7GIlCsAjgQeiBRbmN+sH/crf7aZvNcTWVbkYYZQUA
I2xj0ic/7spxTShBm8N8YhK7AtorqcxG9WeMSj7KzcBxaceOts7Ou7/6ZLYpGwJnJQ6oed4lHG8N
FyNcZHyNG4vJsLWhSODZ4a9Ls0PPwG6kKnwCR70T0EaCRdy4+6q61yJIl8NfpO8VBu9aYBkCzAyB
/WIP6AJQzFBUL6iXGeLG3NafvI8n0fTApTY0CtclvIBvILcR7Gb2G+onSpJ5qJMfO//hTyeaxVOt
VDluQ9FAx85Z3MTwqrED5rIU3HwcoUeVNSz8+F8HIo9jmrtIvHfgfau2IK1BMYADcdEEL7qDvLHM
xYR4dpQGRM1JIW+xUaqUioRiF1Fs8Yb7s7AjsICNsYKqdFJISPnDPkkEMr4PGGxqhod3Rz2d6lW+
zaKY9XHrsBm7uoM4U1oU7547jwgzHiOMuz2EyFM+zoArsJCOjI2RDOcY1pqm95sm0cAMaAfBHpu7
zBK1aLc1ue67VJW5xMDbxT4kQ4Vs7Uad3bmBKQNDGd/6QXm41hOXKfcuRhxeGnRYFzCp2BkYhGTy
ZCdc/Cw73RHX9ZrIJ0Gb2VMlksFuFzSlgqZPhFQQiKz/D5SaqK53UGrJTsDNDSLEnscHZhz6MmIq
pxjnVptDMKPhTON2RTbOYpdCbA7gAbpVIxn/jpBCjyh/YYIJYU6bIuNaz4AdnmcX2hYIqy71XuVQ
DcYXiB+HTtI35H/vZbZ8IpS6QqCKpg5pVy8EbzqTjlGlYsgQOIdSY5ucH9YUOi9E7GSXVFhHQSzD
QObsgEG7h1svpRnL6TLf/MarpyK3fleQeomsCl5f0gkWxs+emUL4JZi9+8pr5X7GFllK3/AmLjv/
bw68syveoAtCa19Jn05bX/c5aL2jEBoSLf8cI6dP0MB6DgDEj0b8kaUIqsb8HIf+EZvxUeRkq2AH
ywBIXlKWvpmOzwAwvtXYTttQ7e8B0783jF6Zf660e7ZXqqCJ+F9/Qnmyov1XfMB+bjFwVSWe2kxQ
5JktGUg7DNkeQ3sKaVVg3akrA8bdGViPwf6NQgEhEwQUwQsm7KoLBdERO51gAKl0iWlXCTCz3ljj
2Y5aNmFHMhG24TDpl/6+Xcne5xznKWgL4pJyqAxMBC5Hscx7sDn0LT3bmxunUMRlvdsSfScEwNWt
wDKEPl1I9qrzPMjzZd4yAJVxwNtCqGWCxf0ZXREuq1ZciLvOvhZsH5XDg290VObcIMh5CBnhdYbl
20XO6XJDqw7y1Gr665Uy3HTkm2ZL4ZItZlBrLLXL/cqfCyHgTcOYMPRp+Rwbg1+yS4vQtoF0O4WG
GhaouJvDSDSu35FBQvkeY2ScvDLbBOBB1jbz6Ao6XeS6NsbIVAnc3r5ZrRS4uR41PF/Irq4c3DR1
5+Lm/UOsuZSWK87blYnazylT5/JoCQRMZGUykRNcq33L9S8SL35vbymgQx9RvE8Zd9vAcMXa7UlS
0sEFmF4wnuMbagxOn28o8Y1GSdmPC75BCFkXhsvC6BhYkjOFZ8Ut4c/Fu+5zhOrA4fI+rcfNEqX8
FdjwiBbYs5qaqbwK8xb/DzYmx7EHGs1gchtdScUx4aH9Z20NIcC8Wek3dHSwpyQbm6pQ88CdACvD
jAIdu3Vr2kEApL+oadx6E+XUB2vIj5ZvXATgs/MzLTupRR4iOCXJkmPL5vmErNtAWAWManm745kE
hQu1aqWvputh9uh1KUb6+JvibffH4rsTRUSb2I1K2+tE5HQIwOqQanSvmyAxfokooVuOpBbiEVNL
YltzeazAtVq6jpiN9ugKyXRNbx+EYKpJaujmlUtADeTz83sQiSMxoljhKPKNGVnUcu5W5XI9FQTp
SwRIdtfDpHAj9Y2NhA1Yj++FcdeLfIMAnuoaN4e2EieODxm89vdQn9UC5dJKHKBftAJZu++TvR6c
FeXruhZtyLk6zxRZKb3xUTjWbV0XMNWFowxSgXVtXpwBG4YNMbVUvQvTrIcBne82jNOU+tduiUkm
d5FoHk0dP4XNyqM1E1hsuDO6sElQzbPkl02OggQy47laLGJIrpN0zo/jfYLIlM/8IMjCzDZuRDi4
BuAaimtzsnGoMHaT3PiwxRjaiDAUansL/Q/ONwJwTmowoluzs688tee69kXaA8f8NaSKN3ma/U48
FWNxNupKG/uhyNFwDBLAyuehe8vyOvFJdvNMYSbnLb0unvbrJFKZH69K92zLZhvszJqalzx4l7V2
0Wzc6pCdSvBd2GEiNkRZ3hynpkF0OBAtE1LRBFdQQFXW/OjT2YngK6p8gqtljJLYrJpF5W5oYeKa
1wDpniTD/OQD5HReiWjAnOKbuhcfSb1daAjsLqeOulUobPJyvL43Dtq7w43+7XKHg48La1VDE5oo
LemlffbNgD4vHStw8a9GxdOBKp8jSwMkEnR6I5/35aAnDsXFdRq6imfIMvC9xvnXfhzV1SrIiSow
ozlJH2SZAxJbJJhcHe5PN4uZs6aWgf/sTqzbkpQNve4qGEVwqYomjjcI6Q7FyrjfpTVEFqlI0uk3
RrweKRpQdtFTN1j428GE14rvF+EK4uVwsk5WQUqL+irPdXmUxBlF7TL2/bygSRmKIgnMqGRSmarN
O0/gK7hFJAIxCzhk2vx0KvOWamPR3CANFElh3dtBftw4+1JNQKC90wVzVrwnsFKU2l/qDxtfgJlN
iFzZiFNW0g7mhQ4MBv8hNapKHFz2yjrtuVGqJyV77jr3yS9+TkItzGj1ykmmSaHxk6Tm+M1KXx4p
hoEXDIX165HYbraNkbaOos4/ais9X/3Gcjvqluy4C3HK0WSeXre3Wm7/sLKj/VJmz5LFq2iYXZqA
dwiQ15gwWEZEjhZ09B949RmvssEImjc5uCduadT0rEhoMg20JC6RHAtGqu9jzqdLKAMYQlbW3OTS
0mrR98Oj6si2CTr0bQRnNmVxOZ+6wvzHjmwflCZRJmNZEe1IlrN6UQblYpVM3VN0SVKZlvOfjqVP
JdJBtpNHxR+6JBdxJXY+gtiLkrj6etrZDsHs+kfMxb2ACkOwmq4CCKpA9HXU1jsRXjGea90pwZDI
qSioGXd3IiiDkZnggUCJX/mAOFdrGbldsHkdq4AUDmjv/f/WOBuPIr3Jql/ZHhX/CfZT/dsxxJm7
h/zT32+H1s2WRedlpJaBeND6gpzVorTh5Hj5opmSaNl5WtXLM1znLKViBbHpx7PyVuZvrAoMqsZN
9dDpBbrTaA3E+Th2t3OxAINFTcgA6buLekyfZKJD+Nhje6hIs8IL8SwBcDFt9o6iV1tTEijyYwi9
HHDv1bf3awkmmCyu40OX6brzxWhe+asqpzFfEb6TX2NwnnjkbU8WdMdtd7yIxMZdaQbQk2mWyhhI
UfD/duikyJ8R2xAMMjsMSNz8Erf2/j4COlxLgZLDvQ0W4EqYSb4tEf1ShjmZYkX4dW398CI2x+1/
haJLf0MHKZNUfosT+1pZWLq5n2gY7k6MsAM9A+4kE9M06wMIdaybJB6BidaXnAZm0CKefPfdnT9p
+7Lh66Fare4y6jLQBSpwO7+h+aA2QPCAtRqtNy1OTw+RxrgsP1gIDoCVMbWC0Roteb6HTkZ+ELFx
p4AiEOP8QueUGkcTih12zXgfg5D01gMkowvAMXIUVr5rr+8x2WWvs1Wad8iUk6VUG7h9D9KBunMz
BJ6kxa5fvBHgcWhHqyBpR/g2c1BTztJCqqTvqwnKqA15S8TRbNuwos1Mk794VbqnPD8r7UDN7n6T
dN7WsOwm+ezmmxX3ND4QGqMFGBpdnrp/fULhSB5FWuANzyFSqU1gVhW1iyHmsB9yo9cXhnGSuHzc
KMEYQDOuhMNyo5VqWCdupyzI75qbuWyYG0kt1klEPO8G4e4dISI1Dfvzy+uRy36kE3Z62GndaN0Y
KpXoX315Q5mt0fY1KZjVXutoSQpIed+wwSq+xxQGbFKclox7qb49eekMDVXUQGu8hJNJE6WxlIu4
0JPUcNHeWKrU3gW+aBdBTyvzu8qTliEVkyCY+YAc9bka9Ephbd+QHOe2ve4dtf+Jdhkvd4rLQEyS
pfPdr4Ufxtx8dKCJnyyVNsvQsWljoXooiQAsn14UpsnyZAHHYtS0zez9UoSpasQeaF/0Q8XJWT4F
72kkRsdvs+meEaO8P3q3FuSs6uVqlzZRxEKKI0oyn8/AM+1H8Abz3ASpoa2DeT83JyLpGaot7Igc
U0mQ2HCqzgPWy+NoCJ+eBri9DBDnz28C8ferqKU90yMtpWVTPDLdG4V6uXp0WriA1q+9K/FPh4mN
tdOG9wsSem9AcbpqocIPTZI6PPSFXdObVMhI/vyvqu9tpTjvJfgb9gBQFpTEXfC8kIMQOR6X4Aur
8ZdSvKAAsa8eXydvWFC87rpHMQdE9Ba5rc6FIx+lfGASbdCn+kZ4+YS631aamslSSiGaJicJ7O3k
bCV4zgBtFrdK5euwLoGqY9Pt6Nu4821qZGtEmgWt4AtR0uJwlfGWVQx+cnGqe5wW+dHfSYKuUUG+
R7lUpbYqvPLOt/+5ZndiPW83ZDQxuiqUR5y/tCIR3fQCbMP/rKP/+bIHCBeaV1LPMeI7Xbsjb1y0
1wjUh+u2hTt7VtRwXiBdxOsbVWTKpqJTM31TsnSBO/ZANQ7e/4QplSnXZt43crIMsA4k+rTv55P/
r2Fq1dZUZdcH7p0NB64EgZNGEhJWD/IQCxhMIrqBTqOb6ju6IEwH7xcpYR0/TsZf4uCAQFR7tiVC
QT28Mu2GHEBW2r9S+2C6kmpcpzCPINrfF4WPuCNJGQpLYO1XWZXx2KdWRsY/A6NFuhjxWjBj4xEn
od8zvrn/dfYMyMK5sVkOvsa76uXoE84LadaohnfOJ/iWg/ZyXuX6DY+C7S529iFKncTO2Qt3mZfy
DmtUoZEKeRGrGYPimaS9QhKl6yEkF/R10ANMp60fPYet1WLkrMFEgcw6P88djXQ1SEyyiwTdAjZJ
QJA+Esgcnsc85hgxmjOiLrJS1hoZK9u9E7hfW4f6GJlM54kZus8UutFAzUtN78DTPQtrzbPl+ZgR
4fADrpbVwsbyclZNRi/TPmr8E6bSvv2psztDWvTrfOD8AgRsdGF0nrWOYcegaJ2SwLeIR1N+oEhS
GkXNeqatVg/yA5dx2GotC1nBFql6syEI8LciwC2UJM8km99zMdi9UodG2fJk8ONfFhJe7TQQk1lD
7y89IcrGZFLkgQNvIBRKEVggddKdd+vowAAHI+KddJPe8iZ+3R3M1sTF7S23h1ABBVQ8uw58QwuX
E7ke9UgfaQerlFbWx4rx/KpDzyOcs00kpDjddyeR/uHXckZ39mWEl+BohAGLHlS0J48q92PDSGXz
S7uQZWR4fZD2Xnvi5SDwbia7Q+FdziRDrOAr3qDkUQKrwK/IZCdxzSZUi7J0XIGuFH/2nSiKretg
jnxXlyzUEB+JdijcfGn2DprPi2xs64Jwc841j/I9ELn7MNBDSa/cfBd2ztOJs/ggTHfSK7LDrJbc
lD5zUc8JTxqS1kjFQljaka+a++9ygu8J7hTmmk+S7PsKwb6wzfNNDBmS7sLLq4jOpjM9M3KGx7Rj
wPrXi0j3WL3RbUgsA41mTtAoQjtKttqcBlNIzJpHQM8wdTVTqtNt8E6bMcBkHYgq2+VQvWoX9zWY
CBRx5+egrKp9xqEE9zL5MyNGJxvqx1m9JxaepB23niGaduS1AKqEJ1iSQOwzn8xuDdk2T+B1yh0J
wva7YyOYVuWyFz9pWV32hrEWIJqkgkRiBDJsS+mt68qH4l/xMQmo/A7OhlTNx3CE3nobzSTu7ogE
8hCPJ71+EmtnDGN75volmy/rdcDM0WIJNNjDzJ9LcO7Tn4hLRODmtO2DAjue1+U6uogaFymgTzzf
wEnH3HttHZM1itS5+J/8uVTs4J9WqcRtGB0k++qL5E3Kj1LqYD4ws8wTaFAT91s15+cAru8tnOvK
a7VsmXQso21RyXpwzJknXUJcjCILLgr+hofxG6/u20jbmiBmrlZzOJhwco4j3vgWPC0sVyJM9j5A
u6zOlOR8k7T8a6cfIIO5uHo7ipfstiCruK6Tz84D302A+SNDB+57V2537oXNQZoBuhNAk46fDvRn
NuRMddFXcysVyNISub3hEtccco3fyesAkUudy/FjkbRZJ93UcDQOYdNtExg5kWSML80LRQfYDzDr
gcC9EY4ei+DmtV+2b6XR5USxOcdO7Z4xMYK2EZwL7QQ7H7njclKKgk9beRvUCaAGrcj0HBFb31v1
4SvRLVROBmEJgJ0UVZ+wMsURVty8OTD7KyNWzbZmWYq6mirbRBs6vQKYc6AOsGg63sQDwo/N/djR
9eQh4bGEKYrsORJJeqwNFuWi7K/rDxEEQZMBRW2s67qi1zaTKB8qfGMpKzW5+nnPuL7BkggRPjIH
awhqwWLhrJ5F1IiqNJQNXh5fNqqGqtMX6PeeyfSy4bcosYiPZYm4/yc/8WxYschgU2eZxFoN46m2
gVtjIiZeIc8h0pGEUf9/JV5Si9d+204ungvu/zplo4oo2+iYIpU7+X+eGmNQMMNfpi6jTv87JgJ+
hqWcC/1e9bCBdFyZdTaWt+1oqspv+UHizbL4lBgAX2g1qoHtpBZ/qtkjnZAMSj4qxycweCcv1m+m
XGEH4tzvbkoEfs2e8PWfOoXM4mIS+scqO6Wk0JscgqqYDLh24LqhJWwj7KML6fep++TMImMIAorv
++yx3T2A9egOEKW2SH9xfVJOm1V+ANEHtz6Df3DPFI2D58ZXbD38f++4jLkVDcOJidyDwJIVB45P
hnPEfVNpjSjLz7ETgZxdQEB4Ug0mxiMPKZvgWmw2x2Ggr3EZexBFV6Tfct+k+LgNbk2tzseWJ/mG
QGOdkAPDHrOGaYt/xpf2j+x4YDX04PgY2C1hjV5BK6bpYVj3gqawGLCAjzbA6fG0wYMAb2bGNwC4
SpHDyH4LzBqoaC28s4hOwQ2oBg7pT94XEwKsjBZ0p69w1uuE0jWRI9V/j/0NVPNJiuCPulwIztY0
YEzkBkskQy/HUdNf6w/EoxVsIYxGkoYqnoidZKKLPdKC9OK7R022Z+DADj7yoDqt21yrNcWe5UTm
smPkRCyoXRf84onhq1m9cf2igRbrjVNOf2hmD/YQj0T/XweH2nFgKeHAL7nzCX9fr/CqB4B4DHLG
/bl+oia6os4e1SfiwcRi9p29FP3RaL44Lqk16/tVLX0fOuydYs8168TxSYoTQ1c3JBCtyK9fl+Kp
XvGI0tYgvtYmSC5w2NUC3DrQuxVuAVg/uxbHuSdBoOzhi6RS4UILeKg0vtiLCepL0pEJawPPBbN2
FlJJdWtUfSS6hp7XgcMgnXHT0rCxpEtVOq1eOo1caK+Z/7zhso6UMWwbpL9s70qH406n1wmzxrwG
SoolCWAdcD9mOj4EodLoGIUoqMEbn3RnTDlvkssoB0/dSnfBl3/iBfb5XtdYwFij5N6j0QROFdpf
VdYK0VZCc0gnLldgJQPl2dNFnwt1UxBrhxsVd85TgVfuO6+R7MKJpqKupZ7BNUy4lr1cXzkwGany
4knZoGcw01TdwXOmvUs4o4QbwmL0X/AHt8SzAj/INhPzcoUAA6BPBmEl4w90Qi8+YqpimiFJ0fik
8ZWBgqcTHVE6CJfeYUccAop3I81qm+8uj/39/eJ5bh0yNN10yri3X9+9vpoWtDhsLad79cBA+ohT
bpp0FAcjlE6AdChv3eQZh+RMORDM+381NbA+57cUCNcMey0wj0hWdEkws9Zs1golXxnzPY34kSCP
ANHsVwKlY4LXwb/gYrf8UqTweyRntlDHje+moT5pm0yJcDkBfXKqEYtzaRqZk4e3Al+eakJkbe+D
Z/tde7qpu8Lkcsdbo3kC09lOrDr89cMxx8uRUzKAaXGlrYuJhKt3Bu+9zxcYYg0JhsbBIvcxJeSk
+DzFcq8Xt6n05WuPE/LLSS65vxkcW8Qvdr8AnLVyG/dEkUz84M79eWkkgUCKDIigFEWd3tZI4tQN
0p/oaVJ3i7IYuvgLQO2XYd7SW+vuKNCbDwV5Tv4+1ElPvBVUv/wJOqvJ1OT8SvhYXQLMMSS1YE7T
bVVSOOvMr6dfzpR1WP+EdHgYfgMhBBkCj3J5uTi0m8nlOdUH7UOQAyShlvbZmto7P5dvqgNZ2XjB
zff8Fqc6xyM8tAlXCh7ZKUMDaPSrtl6wV8fCT9mrNsA2lPqJaV0vu0K4iBlVJ0CNoS8c5BVsxy7C
XWT5HsCfi/6xsr9Lmgn4PUj5GaIbSGWN1tDkYev7EEZ1LnhheVIszLfzce9rrLlcf9eBE7NcUz+T
+ID5yMAH4MiB+M1chwsTmnwfrvfjMaZEbZO6yrA91n84MLz9iXEZZntAVQehwp/DhhyqxqSQi59Q
JuMpigwI0TVvjguXKLuoYrcVOMNFijDJBbKui6eSc1NQaqUzPKcBS00ltwWT2Kl3d2mEnP9QCWEo
j9KTlnHZBkUQ+DrYefXQWqLAQ5UX8ggUNNgc/llglqjsn9yAKbLPpXv2iwKCcEs30Y/RNaK77qBN
gAkpAk7h6+tcOcE0wbDGgXRPb3WJ4ZKjtSuW8NZiq4+iMJ0k8ziY9Tt+pjQU5kSr7E/ahnVzXY6D
pcMGYgy5G7gXkgAsfPyjY0CAQ4qrkTRiPg8Q1/bKwdrV6sxt+alKkg9S8MDD1QLBUsf6tg8+UKD7
QTy0f9sFfFGpf9uXj5iOGDEX7etBG8jqPwae7jWC1g+Kr6hEX48EWk7X4Vks+ztpcpdrKuAQPbZ+
tidz3JOhFH4W80E9rGmITtUOBNrdlCvfjV1J8VfEsqPyMoDnYIlA6zpf5XECYsfttVwcMp7q2sAC
yFAVs6bbWGWoymh7bjTU0aPf8TKo0RsLNeNR7W6HGkcuaW5FCesKphn2Q2mYUGsl8Hv70ae3TiTD
24+e9pwE8eJsrzDVrwy171Cqpt+folwTM01CAmye0Zv5PfDuWgFz+Ob+ADCa850LPcy5hZQUflWr
HVimntgXb+eir1b72aYKd+9Q2vHiNJfFq9K6tGkrlLWeOulltDx7cMv1doigLgev217GaxpZbaF7
pmPNVcHnNgTxmPgzXRm4VFFISJ+G2KpeU0KjAu6nYhpqsIf+TE5IBC8IS6Pc8qOr+PtvgjgG/uX/
YVf3z7sOS2+JYvvs7pWijuLjxadah5juKYcJXHkfAOIyj6C3vG9VciMYZSfPOgJ5lSRGpTN+lzqZ
F8KpgWefjc9GktmoqY6slaqg+S7QBTeFrp7tHIFQjFMrc9NAzkmtAZXCtr9crPtRXMwOgdul7MoA
lICK4Or74n17dPQbDJ6MGNk78EeehZ0tGQHt1kDC6zKMxHIDZhm/AGoKMVcGo9rttN9G9LvYzQSz
1uRDrq981+GSwKvUoADFrKk9B8dOj3Mi6K67vNXPB4l3x4wIKHIoL3T1U/y0o1g2MG+DZ6Gv07gb
SA6QtB+b5yNwro11O4jVH6z5yxLs8u3GI6+uUOKHoyGryRC4ZB+utfAGcAqeR/+bC65uiVb6affM
Q5XnHTAKcKdgpE/iOdhPf8N9voh3zKCNz/tkKqb2zLJxx3/HPuziamg9gRYgAbTB/Q0sXE4uiBIy
58lSzlMVQbx+SRRSTE7g3pMU+Yjg/aOQSZ0CQOCF21PpXlKoHD1ehU+nJQM0xW0AllL3VbU3q8A+
69YYOjqqKhGVCNF2syrqYB/tH8cqzdCZkhaA/yy3kF9hyb7mfTA0L02rpNCF0DO4ZTGKEVw/zazD
nxFj5d0mzNrT+PMWdj+ANKcSV/scannJpZCjiMhZCBn6nKDWJMcaa3LbgMHKldFjjePrxULsr3fv
0ndvObe0RfkjNRWxPcjIa1jZWhwV6vEKPjqpODukib6uS87znDXKgax2Dtgq8HXbaBcCd1UmUt3U
ZXA0UBwfBD41303oUjQFvaduP9wUo5SfaQsjEArzJ0OHjS4m3/7vepIRGvRPnliqsIfuME/ZuphE
Z12vyqDFLA4iEgNuXe1+K9M6mpADN/ErZUDAPoO1rFWGgLQo6sscfq18aCzHYx9YF7ItpxKUf8Kg
l1lM840e0jGUG52E6zOhG4F79Lt0VgHnuC8NsywBXFLxmQgMGgl0jLL3D5TR3gZcayGL9eMKELCt
WkRLNf6BFox0saLye2/pQV+5xlyA6xT3TcZ2CO6eRzKBQ9uZum5unXxBFkntRfl4xowso0Rop5me
QZTEmAp/ikcoQFgzcmTAw88nEINiOKerO7wDF03ZXWYnYltiqnEsTBNP+hN1AQjxJD16oXZA7dEd
6D187JG6alEVeiyw3EgfUhRie9fOwYbzGx+IL1XkPV3SFqJoKLFX4HGJWKgeaAekawA7+7vzmVeV
1he4QmOsr9pFxdzOaLVdnf9faD0ogK59QVB2QLAh6ChzcjcGNXLzQgqFYdS5K/mn0A4DziQdE4NN
3o+OB8h+KoienzK0+mYh8bF5vO6qppNde/O2BL34OMF4W1tiLEBaEYenHv5NCNY4LMurpWaP1Awc
bvhKG5yuD8R/AuhemOVB0EoSoKCHxF/0s1kkMDXpakRqn5L3ag8l3SwuZJHlElgM6GrQXYivr8UI
0CpaDnailwo8VWo49i8DuUrSlsC17ldOdSaGEzPpLBOzchYYBw4XHB5wc0F6Yebgh8asR0vRncJc
bszJ0LxU7Doo8y5LV95bFacHYXcGaZC+OkRBCgqzE/bg2mhc1WDIPM1QAjvsSyYkmumD8WmtUk/C
3r0DmMTEiCPJ5AOi9cassqmAmE3cLUbfy7NPXdHurS4jvZd9NcFRsuHdPUNRUugRAzza/rU4Wfq+
huewqr+ep0TIAEFEt2hDBRjaemFzP3dTs+2raliXFyU6j/j6DkSNWN0Q/Ppo1Cs+iddBB8SB0hkR
TznCKtdKIVLBOPsYlY6GxIBoHnY/cmm1mYaBTmc90KUAJ9F9nPwGXyMuZtHPOrfHwtQ+NYyrKNgB
A+PIW+86KND3F3+B9pvgr7B9rq1G6avO6uTPemOm3BOBo0MC7WoztommJRcSkdvGGCS4wbnOcRBB
wTkXlgwRjm+q9b0xfbeSIcHJ+MO8nu5yPrkVfEg1/Pe646S8mIE5KrgjwFSw4z6QwgBQtlh7Z1YC
R6ECHRdf02q5tWVR7u+vxvx7euScVT9JkaZKJIyA4T11B7w67hBySxVlHV/YnYJzFrka3zKWpr8Z
HQ+cePb5z90HB+vEG59XqsnluokNlMO/IhvAJ8U/iFkazuNXc9ryh5BH1OWwiRbfZ4q2QrA+EVUh
7jXFski3H/aFmzV/xIs3UmOBIZm6FlBjh7yaE/tDv3xL6P+G0RZ3R9PmfU45eqFwieMYq3+hL9Fj
6yf1kSzHyYuBusG07dzeUMtYBB+tNQzEQT+YnYbIvsqZ87t5WzOPrvdlLwRw1C2kPaOaYUW3pcEO
qE3Z93CW9k4Jna6MEfbaeY9Lm8yU+iXzldTarQxy1IKyS66+ZgEdNZqIHfnkZxufgG9J4YJtTvcV
Emuv60D2OQoXLWGH+yHJZTFAudpR/U40RMbLbkPVQibpoPTkgzXr7KWLDgb/8ib+IzFsLieHvygR
UINQmvKQX0RaNOjvgSRg4WvC3+ZHTqClCp3cK68NhJ0AW2q8N6eHiTCIHIutpGI0+Uo55A4VCz8P
cBhear7ldnLMbpaFgGg8bCpdNops1aCvjkh3JAXryZ5tZbp7nTMjwggnFi5YdeKpRNi2tCqMc7Z8
FzJdFFp2nW/QsgVRYcNzrXpjaDNdCGuBYk0O+w9XHceKdHQ94dJBqWTgwzV2jas+j0hDpa99C2S0
tgTJmFqh4mwEiPxATWgEuTxRs28Y21xjpafybJLEYNBNuZHrfL6doIufIriT4ypFWgmGmTwPnRdR
UU9FKHuCpilY0jaNDu1qIsvbiZbrys8EGUztQbTsfHPFkik36hXWeRMI7iLRxrPtI8f/S1BZ60Q0
0eG5I+rBXq/rx4XXtRI5edOgqLur+B/G/PDcrcfz//dh4eCuGBnyocgUJTAVEsCAJA19Nn11v1gp
ek8EFPPh127qr22TOyKzaUPmX8Dtck8ocYARCP9YKgxfIJ54rQax2k3FRWw1kWuqokXHdlp0KJF6
1xRRIo1Tv0zX1IQ/MR78wwca9f+3YBQv19mDCjQAEBHlRFtf4HyD+OqxPfWq/8qJ21CUZPjTEnPq
YWrN1oZqXy7xYrBRUymPvxW6EbBJSSzdHSMI9X7IcEuaJYXPahw99nphDP7Fa9auE9/jcnuew3Fi
N82y+Oc92E/4/OmgxstekmuOSxCZuXp0oeJwUA2I9OHR+ErLkJzRBdZhLz/I3MCF/rT+QVg1SssF
tatc+a4mtzdR2F32wFphh6SrLNnbojDq61ijN1kQybhgl5WmSGDBPGafyvqP58KzwvdgmWNz1OKR
9KBg7bsGyoMxh4De62xRj/elIW6bQekgiGUN68WMoCz3j1DaR+t+xv9c9I9Ca0oXCV9J19MfktX9
6jDyIL4/IGxMb3FdWTYy+mawKamr2ZB0xYV16+zK+nZsYxzLgnlC5KkuxeR7mjDimILKRdUT1AgT
O8Lvmsu7Eucr9hgnFljNmwTNgZk2VUralqtt0FowmZXRWPkMx3VwK6PYVAhatp3W01SQOSxlxK3w
ic78EqECehPwSOHKdUPMaehp2E3/1+Mqx8k0gt1mrqlhdhDYIEcYTRIbHLZtlGaHMjnK91T4MILF
8eO0BHyqN0Uhfu/RNOzgpxr6U3gw8qoWY123Xo+RYsdAwRi5ZheiJ0MWLwdPuG4R0ElXADI7VDqh
eBrGSD9ZPThg3rgpnSfT5//zmjCoVWapDDZ7lCq6m/a81iGdzcDY48saqxAplA/5ILDt+orD8brY
hywE60E1aQ/UG8dKMseYiyCoNrzXklMJxxeqoO+YRw6kjwkvQCkDoX2TFamBDLbtLLVMhWbCba9Y
8Iv+ZBHzOwnyGsejdbDBKg1XeTdSrpczMgYV5AJxyNxFDnEdtP0NjksB/ylHEUDzyGsq/GvP5bWN
TRnjXkhb4RqaH88Q1Qunt+PdGAB8Uftv7b8lvTFM+PmJinhXX8jZIfn8R1zwgDPhUCI9/RAQFrDT
Pj6eDM2Yjomf/MTQL3zIclAua7Ia3H4sIV5/F78SObDkJzjr99vmPe3gggKbEEO1J0FKQEPheG3h
Kp+/beVSYpzAhBJ6jjn4IE6db9yt5RLnXyX52vakaCfpse+3G6/ZtzlAPFUwMRBbNfGfWvYIXl8X
jtG+C5xlD8VdAkh+Tx8J4toKTZ910NztNhNGn3N1J/5s9TVT3ZA/Q8gc8pLpMPtxbA0CqnZ4gYBI
HgwdcECWaRSC3G5tN8vAh7TruPY1+CfSBBObW++xhKdzzeNNHMZQwKjrQCmTLfbUzneNtsw1JV6u
K0wN7WvTl+5VGxkG7vYStyYcFU/rZC7tDN6lCpce4AROVX146R0uWLkHnGGCcpgJpX48YdFOwMPG
MtcZQ3n6RXVx8/gG6UNJcNV36F/0uiti0J5u753KVnFWJETcf1UbVvSjVniE9oMiqKmL62Dp5vXF
WkiPOFktIAPWlqn3VOVk283cg9+7mzQPmHUB0BPRGij3xcv53mN/8Gt+LqlPRcsUA2IkgcXNkbd3
Uwz8h4h8OgWwcd9TljZkwWBrmE0H7iQVzrogctdzOtyWHsYZHsrery0VsxF1sYgAB4MSDAgQxHhm
U+EZSRlbITIVIYr0IyJxHB+fI7iQk9JTXimSirhME8wJbWp+ZnxTMqp9zkgzPNsi9WcR5bBZGOJz
DaCfkhgKEYJwGHR2Jit6Rlt1Q8H+lzp6x+YHD4p8rJvh4n9Vb2rr6wq0xXh11uZL5NVROKIJsrFa
Nn+m+WHQPCUSvWdcmB7Zwfy/kR4XDXRIw3x2SNyXXiGwGJwHHGClAZB3eqyGK+c+P9yNNTFDSCsb
MTdR6Y+7xEuUdcFpPWMvAOXDb54eE7POYEn/DwJ8GxXVQve4Q4B15SrL3LLDvWrRUH03ObMDfFRx
x7WnUm8lFiG/LM8RziMTsj7AYF/PIeRx783FVQw94sMYUcU5lPFBEOjVPu0ZWMpzS5TkB1o3lvRq
83Mu8C9w35pIXad78w/To+5q0i2QqwIv46jmeVp5u7j8xX6Cw/MbnucApEm2p50Mtr+3qFG4G9gE
VAi7m30AleyKZByOHDwvcXtPGTdd25hOqP9mtXMuz8JDw9hMx9mf9nkHLdQGdXqujcCR+ZfdKrio
e2QoTru7egwkVSr1YWCXIVeOTK2hid5gE+wvJiYioiTYzfSSOKS3LePjs4ntZG+1KJMD5BG2JL7W
TdRJ06YpBSPeeOVxphO9ngiD1zfWxWNlO+86QaoLsN4iD/GLMIzG77NvhPEmnZM1ZHfhayha/pEi
1DLEOUWT9BnM811IEhHe2f4n2YcFYnJRWcuYI0hwYMsGt6nUmGwjEPTSs0cVnhlYpZmArMAFYNyt
tuauIoKvX7IVKY4y5WBvAI9JL4tfCU2rmk9w/O4yhBHoXlsljLmGw/fvX6JZ/HOw+ieavOhZAHan
jlRYdP76qyanwvyKCPDscSZP+uyDEFmuRP33fXQKgAp1NXdOlaeGQ5lS3k6RLXoHgNs+TKh6p83K
89q8DwEXXoTb4H15WrIn0FqnXN/ELTebh3UEMulgxGtDj8Ofhdb3HrGAJeKjFJJh9hzmkHaZfi8J
Vuqq8+AVc4JLXIzH1NOQMaH6e1l1W3uEU4mGsJ17Nv4+B0/uWhSZT8utUIj0OBLoCYzW5XC2WESj
XvvsRaWQ1TL/PwbHAIo5wbUcjIyI5AcDgAUL4LJflXCB6/zPzid06PrxsCT2SA4/xpZQzT6qtgwL
/YIAPw7N34W1Ywp5lAg3YqT346b2DQdiBozpMPfriFldByLONBDDv8+JGNWSNxIt62KbVDR7TfCr
cAk4sk0xxkQAuuuZuFHD4RVUWAhTfnLNA7U2U70joB4U+jpkAYAnBhKiPsmk4SlJ6qbI2mp2rGUr
U+kzy1G2UG2LgU2UeMq8ZwtV+NfxUkVtExRlVyP1q+BX9N4rGpBspo3L4YKOKgG1GbTwc5Q0Hp5i
Z0QB6h073qbzJIwZpHZ3QBrpovKO/j/izMQOn+lhtvJp+IRSAKt/Az1ojzGhRlG46cgiQUtgGdum
2+GhDTUAYaaKq0llVBjULkaUAFzxv6Fkn88iX7o/pKaK4h/daHv9irQ8n7y76T3y69glcnkVTD73
sc7uZUFGEglZ9ImMlcktPsJfPaer7NSZKzxFLy2CLblcqh/2bLwUak4vrKf5UHzX8T+OvnLAd/Cl
VBHUzbwTC62AhSk5KTFQjyNIKE+QKl/fAoUhUZ0WNxqhOitHb2X6THOVLY62/+qft5sUvFO5aVOL
Xx6Z8d6o2lm/1AZZKdbjHjsX0R96DL4tW/tqjfyUe+8sQ9HW0e+M97EwXfJY06a7VXLIGjZ6Cr6u
ZOi2fUyY1LFu984lk5ivyHa8hDtnmvCwKPzLibp6a6uB/Pzj/qtTx2IOPJ+ZjXSZb6nd7bp3AqbP
VjJb90yx3R2sF0LU+dvC0SSxuBhvrciAzwJX+zdPdqm2OSif0SuZLhUvxs+yzmbpXW8O5rjVa0wn
tqxa4Ecyw2qKXER6FkcJEHJCRyFukVvDRVSQ0lTuCShkvQ9sjJB2rlEpR5Aff3LmeqdVaFRndOxG
iKXobuWNKxjwhVPdxhsnqTwE4WclrsJX/bet2/RWPyWK0XjLgcVeuzcCZzq3eMkObeNVvKLBwF2s
CprIhWYQDCGy4/pzZ2dATGINqEVfEuqfnLeSCXx2vV4KNp1DR6Amv6aJcUWnNWUaRwdnDasgvrPJ
wxxdWCmVtICmjUghLLux+oB5tAW0z1kyqQjpyiDqBxeDD8VTFwrvqn6qXJxQYAqC5iVikWGbEzHZ
QIYJaZwEUCCVrq1Fop6qvo7bwLC0s27ja5Itx/BK3I+jgfSim/91sI8/RjySiDRLyZ//b9vx0e/2
poEI/TsIDMjt3vLoeB5V9oDP79X5CcwQg0U7rej6kn8v3LBdczpNtKmv34K7TNtdJ0mZITRGgjuL
pbQXqYKtDB1U0Ryj7M6IGi4VmoTt70c6kipEHIPEyIjmhueT+HVPGczpZ44v8BPndlWZbdcGneXd
VQcLIuMfi83rMTLVuTnbK1D6yuhxr44Cdsa0Kfhrl42Og+nlvBN+bPloQBB2AkhVI45Jfjgg7pMK
/jVunjIYyUIWu7zcAfQmLJgBBuORx5hL7GZ/5rrIQBpc6sVrxWjRuZYk42TwwILal2XbZbiEUMGa
xofcPfekzeaczp2SK3DTgP680QHlciPBCbT5oj0C5SwGJVFCn4K46QK7iO7aIqWUWdSzqdN5LvF+
hrXYn17yH65RzYMvAnAwG1gXAEEUjwCbIRetr4zsFpAbPJJaBiNE0bqcp4hkjl8Rn/7haFCpzK7n
yeE6dFHI/jEiwegO4PgG0/jAdjD6hOV7OThSBmnsiuX3Z1cCzwM1LbIa0pqoQUR9MOkJ0dScz7RT
geRGNOdZHPQXK8k4DODjhH/FgWhGuuQMZhEzlZr2IuvnmotwuBkhu2W1iHs4ml0SwgR0DXa2XKUG
rRS9Ec6P45E36V1Z0XfFXdRU0sLryGJYlChIojTKhk0yF1S1kjQBgH3rs7N3te9WQ6KrrMvOcOTO
OOGBH3LLiqFBfWIEg9BucZHUP/1krAvTME5Mq9FXz3/u24Ry+gLTFuHMX0ptfCfYLF2mwgamHma1
NIm/aqK+UbCkmysJDXCkLB23urWc+S5PEw8GhXcVvAOf+IHhV+DQf14h2FFcW4/RSbe52leu6sPo
glPxddHKWOab3KvGjANywYSV0VDAEV+k2v8zA84umls6WasGznMrFiErPEybeTnZZV5uJx00glwT
TS0U4kLjZ7RBxXaX4Y2dlKbehw3pgI/udCWShclWijw9BFGm03i27SVaSNYMe7FZmscyU8JEbwBp
JvD3auVa/+vPRwlBjB9zBrei2o+e8V5+Y5B3LmpvmIKbibVcDnffQ394cioe2MDioddudSIehoha
Fpp57mEHPbmeQ/oU181c8eijLyOsyxpVB+/eTSYNpBOmz0D71IMLuHHKcWtIJ2ASPBN2q4/0mpXh
/9CNGoc7t6YRM9m/P852sYSf+CVikQAmM3Gpc4DxMPKHklk88YEgO1oPd6ujmI5PD7zeNvGxStm6
ajtZ4evADhyaC/nQn75k4HwqEhv32a10wuQEM7YOd5kj5yBa8ear6/4aE5sudnpEcLO5KZjm3+8h
HeXryvLqnBz4IFLQDWofqVp1joQ041OfIj9RHA3vyr5EUBkejQLwJAe5N17/oFgED7vhYEPSrt64
4jdtS1z1eujzj6w03UaBzu8NNE7ACFEDixQ+fCWQifwzue0oNmYBoWVrprvfMqWKDSpX6r+S07Uf
w7DIZCmtoLtdgDewX7D3Zz6QnLEeaxmIa4g2FzowayzoaLP9T2zko4WM6+iIHv7hw22OYdn85GpD
+6Z629U7RPowlUWf6PiOlCaPKgBiDFhBTtUWk9/M4NJ7owawDmjd6CJE+TaiB4Pg8f3Dvv8QSJ2K
VANISXa3qz61P9VqUUKR/U469+GaJAUyt7dFXRBAPVATbSGskx1o+rvJIUnqf6xdzTpWHbiI6AUo
zons2kfFm4I+EVFD5s0YE+fAqOreSP79SmFtlYY8u4LzOYuvay/sG2pEODp+Ku/Y7/FB/8r2bY05
nXk3QmhziBakkqYNm21EaAnvR+3evejMG92QPsTQXN6PNMdefcIX+oNBBJYmyuCxLxi6EgH0VBc6
g+9w6htd5RnfNWz1TLEZJ7gvqNFzgUVkOkMet5XmYgDO2FC0YQGK73BuubpbOdE/Hhu+wo7MB4vl
8y7f0oK4X8vnrFbZH/X6jnbM6v/rNu6zkgOI6u+9PcArAO/5p29RKnas60EMHIV+wtRjoLRfoH1p
2D+1qgNgVhXQNmEMOKoyO0LOgIt332nWCEZaMlvu0o/Vxq0FzMNVdoiXq2QdJJ45nbvhRCWRU6D8
5JGHNitxJgNvYWquXgr9W4XUhxTDpcNv9EQESpNan8BvKIa3Bm8wggzQtcsx4o9x+94b3YWcM93b
Lu1PLaAfeeQ8U1mRGVAzrNhTdbaigx9626rOk2QTEB0Md1dinsNvX+0Azkc3ZYSU+ILXFGk8Lo1K
+vQqzxHbvkyOSSoYIWp7sAtKed7DxUIgHIH9+Mo4S9a13R9SJMvSsb1jnbo3XH8Hz6jcd7xlB+Jn
wAiPblO6YdCBbJ/UCRfCDlJQ0aJJpFkVPxlPtP/0gyYKcI9Gc+bdj8FV5+oL0Zo2LGm1uRwhmA23
LArsJ2Ha14uPmrlNgYJHlK2dkniNpOuw0sXY5dn1AlS0bOnorO7SmAiKL6aWh+HtahWD4l+AOJDm
3wOD5xX+XmttyvTRDRb7BYUH6zz1p13VGg1vF6u7Pl453H4EsS7T107R12oX7MC19ub0cMQAVKSk
wIymKDk7bsnKLcprHNewkJ2X8A+GpcHCBpWviwz6GTH9kYHvVJDeTF7cUsELvDUtYApAlFp0dT03
oW5+96vU0W/FhEOuHxaVACu+mstUJub+ZWX5kEXtAlldy1b8IO8EzPBrHr9K5O9bWk+VVzhfwaKe
S5LQtHwuJR2dDAm8v4eW0dCl2bAfDAQ+5BCvKcizZoMld4O+5jDVBvsyzyA4fR5zCsoLfBMuQ1oA
yOIN4GZnmNBfN5xG6uDpYxUd54Zsag1qT7n7lQDRuXy24jINhq8nzqH2zIlKoyTDTLDqXf0c54Nw
zVh+C0sf8Ir21TLC9r/1/BiZYx6F4HBAkvqYiBh18O0T6sQr23nd4ddJM0jAJPUPQqp1CVRzj+jT
/iQFEfD/xcSqCixtlpbCoihjYRox6jwIQeSfCnmyw43z5TrChxwH58d2kvKa0JOgwS0L+BAKmuu8
Dc+Z8wnZ0/SrsycoMSHASCWeKVV9txJg6o1SU1qyTtwDGj6HhCBJyLdZquAPl2/7bWxzOpj3am9f
Jvq3xinBE8yE+gcAFn9fuFH/0IqzzausU9PymcVRh6AAV7tS1NilLLvD8SZJtOqsturzSI3AsTY7
Wt5ctygOCwTWzD/CT5sAtK75y/cVkUGp5147sjEKNxdcOg6OeP81ewAsKQIyLtGGI25nHNMXdM4H
ComeeWrg/YYq2STvbBgyNmH4KtSzoK64aAHpSRFuMQTAcOZcsnyN5sfUV6FqH8YsL3fpojlX8XN8
NBXpDvkhxFG//N3F+2rNU5rF5HhzO31h1hWYvCw7AvdMMyljvuTbokxTri0Nqd1o3Zcl5mk9Bm8b
IQcv03hrhDOWTspG4LN3fG+dDd8QYbTXm6uWn3kEURIvK6gsM+s8R8LlA9EVDcO0OXwTeU+yjebC
GkGP7lyAn1Ic/ZiDW0C+ZdJUB2i7XAE6QDiAJ+5+HsNyJyuSdkATKDn8MMQT7FWq/F2iWPp+rdZg
Ge/u0JtR0A7FisAeSQqcpXyTtW8lrqBNcKfrFwh7v5LBiUq2G5acOgs9eKPHcgei67HnaN2TF3zn
1BLchkjVml0Q/8LraI8+GUgqhoTCFrycCxNcqjbfzU0CiadI2ToKIg3xmi3mNKeDVuVMitQ++gsn
kghNFl8sRopoj/AwXzgkS9UEXKTxe6rj4oVqxa5zJShjMRiq4gpfXP9VbLuGIh4ZKlvK0BzR2JIv
kourx7AOg8aoZmkuCNmg9GxZb288qS79ofgdk8hfGNWop+P+myIFdc1J5aMHT7jpgUhL2XpBZHEO
MlZoUFqC3TpPn+6vuOi5wYYsOaZLE0YDTUUQGe8Z6TAKUpWAkwYvV9pgMmcaYFGOb0d+8v+Mij2W
QRFp997Qgc/hWx/9yYafqwqnZe6OdA4Y9pE3SXASJOAfjaxVHEPYKshCevqic2/eCTIyRQvQsJAp
EcAMDgXN/ryo90hbR5Jdv21iJoQo7rcgu4Magg0jetMKaIvpGkvwC9kXRKAW8v6dHk/OCAx13/yT
4oIIdE0hllXguf1djTvhUq4JppsSmUeUT+Lx9xxmzgSH7pIk45m0F0hmxSeSHvGFvwJeRnIw/vHV
I8wLHm72Rukezqm4ODuZJg/d+HU3J2aXiKMsAQiBvN4e5eHM/HTM2yxdsF3Fb7+Ai3e0uCgsRL+J
gPIH809KNIa0gHuB3os0/D/lSOwJtaPfW66mU52xzX2/oQD1mADzfMUIr+E6QzPfvtBMxC5HxAgj
Bzg/Hk+jEB/RQh01YxKmvcdkJDPUnq1ljQtZ0YGpFVpPs/9YQIXwlLuUO5VZ6YY97GAYdmmoKHtF
gOyChNCIFD0qkfONydi//HY2uMarjmOzapRTKi73g8rgwJRmmOCw8A5Xn0QB/TSmzo4bfDaIyT7+
4Mg/LiFYx5CqSoNOZjJedj94qUJ9oTvthurpK0JcOJQNwUQsJ7xB1nZsjeeR0y9Dywxm/nA2s7z0
uOZ/hIGIcVAimC4BbAon2hUtxfdQtPbp/LGohxDhkt0xgnqxRWq0OLvh5u2wTk7e1sWSVbEH4pjp
pkP6c3Af6+9n4js6WFYUCpJ7mDplpVOo3xYX6OXCVmvkVtDXSPXh0TM3At9oR3u3OHIIdz5GN4b4
TLY9lwfw9gOr2m1+2Y1mfYnr+lRBhpT3AsLiO0NqaoWvozMCroJUIQYf2jHBHUFd3oBxehIPzl+B
7hlst3085TaTNh3jb/aknjoboeUh+X8+eLEX69i9L+RCxN8L0duNbfk9LlUQVGRZGgrKZEQGN36y
ka46b8Rk8Og5ahbN0Ll4fHCAEUbM5uzK7cDbrJ6+m0bwrip7SpGhKqMmQZ1llaJZnhdlCkFM2EaN
IxF7YX0j5ML5bSsqAh5eZy+zpU8IPYv5w7VRkHbx4IHue6y+t6q9U+/oYMY1w7uTf927+6n0jDGO
kAiZsqkPii0iUBbhuD+45Wd5GFjKOsZJks4Hrx5ZnflFl79Dq2i26a+LKVrErgS76Lqt9NTPBFFF
dgqEfnelCRGlM01TLEt/M8HuGxSJSUPVCy0+N4HiKbySYJCUMC1Md0KIsIZA/CHd4ZsX87o2Qgat
h1cICH6+yFgD5IHRDpWcRW7o5hB4qaBIf6aWs9iK+FRRYd+DzPwuC6btJ0H6yj/GsD4SmTz89xfZ
CjpGljPykbIlhSgddnl2YLKh7rRcyE/Yjk7yXT+hxoDw9p1C9y17HtrsZwTSzCiV0hXt63WAMH3U
2mB1GUMM8lXAzHSuqmE+1zV0luZTLq4UQ6wTL9nMiduWuwuABklgtkJlzdF5mEaHsXv0tw/93Jst
hJOTj9H6fpl4Gcib8v1JK+hfaKztPn75clShIP4YwwvtTfjMOphte4xg/xc0Ld3PxqYelPoGbWWs
ApE9LijVFv9Zsc//diY1lB6fI+Nu9WUEOeT4Q7Q6GS3nPgKc/DtJUVSuT9MYPxuINoK7cPfkmY6/
nTkyJaSlCZGCqAV8fusqb/fWEiCCgOCCOOWN6opx9AM2XV2e73Z5nyVb1Lww3iGiXt6qef99KYOb
YpWHpn2vYn0XqL7PmG9jAVMz5Ri3WE2jJ316Yfg40CgzoCBN7peokhlfGzTLqEfjDvutr5Ew7Y/A
tpjsNRHb98rBraYpXwZVO9RaqSMdcHfBp/HuEQVscG35U9Xyp/hmV+Jx9MU6CK7eTq11CooJc9yj
UhazrXtFFPkWEMpO9h3PktR4nASFLt1bVIRcHXRnJqFrVJS7gqCccAKkJIrGrSvaTwwp23tDFyK3
e6C6mB73va25qd6SD6AwnMX7IvolahQNZKCS/j/2JHnHSkKf8UNLvn7kQ8MDoZlUl76pYag1RRt9
pcyzy+ecYzp1CpqJx3ux1Seybk+8nGKUySZaqUyWL7iBD00nMAblm71Etb3BPEb40nEHoNhZVehj
i03VwZx0nJys0N250y/sGFHESI1RvxPjFnIXkalwvXqk2r//+bRkrMkFzyP18UHvH6tt+y9LjUYP
m3+Npsj4/UHWj/4qHQaIaOlgWSFxXQHEEMNtFCooWIwWXYnXYBCXNLhas/rTBifs9QpWUQO0qpy9
ss9gturmG4ZB6r2cJGQlNc3ulPYjvhwr2qM9EnO2/xwgg8T1A4qeKu1TydVWfLBS3GTlkVqTYMXj
VKoLAg3BjbTVnvPJvs/es7cU2gImI567FarzZSsrZw4Da/WfFDEvLn5ZUHpCz28qDtxw6Y0GmgfZ
xNOXfBMOO98tK8oTSuvb5ejtX+BtWXJtqR2sJ8Pijkl25cdqn1hSPGgae/xx0JxEcPqfdeuDVzwi
cLDt3qEtEKs2MRW4nCp9ceO6Ks299LWmwkbjgY/nxMyIfmY199fupPWOHgU4V9sgBTqBX+4hvqMw
6Yl0F5gJVO0AjBemx25fBhAlH6fZSGgBXbC0l/Yo7RN9/Zk2C7IpMKZZNQ3rcF00hxb64NFG4Gfw
BuJ9r3Wi53812KQrOpJaiJGi42y5A8qWhAciHGKdyt1ta7HT96QbupkYV5fw+Y3KUsW4b26GEnUK
5lxf9pp237D/iKwlXr58ShQMrd5PyNpSmFIStCIXp7iBgnOf+SS/vkFAvHRlLGAh5qvJjM2znuFv
lcPjuy1gWYqnHrmpxVT+MmMyiZqqY8CArO4Hzbg19/IwabDbe5Tyr41DLYKT2o2L9ML0h1cW4Uba
T3qVs9HWrORl4h6nRQeqFf6xnU1vf74VLMEY6lYwerVeuRLtGSt7jacbSoaIPpcjhRvIk3h8oCDm
dkBXNBl8N2oDmcdt1cIAXjzR8jkE3R5llREXxMmnDFJ5jT1SZ+Cfo9i5jS1Z6KoZ5Dvk0GNx/4DH
rtakO2BXsy/aolS5n7pHswYDgbgH5P0vBedMhqB6e1aVQJBKKgylsn4I1jBE21d31m9uLN4KDDKp
sGJ30usRPnyHmLlYVL6VjkT00ypS9CcH38/LOd989hB9n+P/70SkrpxaWc3dUwp+IXcxchvd5dPV
FlAHGqVR4Y1yLb02hoVegAV5JqOlLUtPrOGfaC6s44W+eIUUObns0MjdfakVIh45iUuKPtIo2MX0
Uo8aiCZA15cmW/wB4kSzylgeoSg3ZFUQUaK7UVXYVX9yZsUT+7UunVG6GRZ1W7e1d9Z71UzymbBA
cZruu5qCZDqI1LeDz4lgyidP85pOO1xjw+WTk4qtD2KimaBlC9Kb4q0YA/llG6NNj/JsVQ7EgjDS
8xNt9NW18adID67sZJ65xEMRI21u+e3JMeNCaCpSRl4Umre34EirhYZgnClg3GDWq+AbvL5Kohen
DkaDM1FbXlCqIn/kxZBsDtJJ0VjridH2ZIWGFnJhyIYrfZ4eVbQhDEJ8XXafRvOFXFpDozUEM4j1
jWvhl0W0Pz8uef2ZreD5o7rSAeXGxYOSOpMCFPbUk9RA96no7vdDmRzA+xQggtNiGnwgv5FT75D2
lkLyvB4MXnjWgQ+cz74phKiyyVCQcFcCbpajPEX6uXoN3OfAgqfqul4oRlYA4Mbil+Bh/Gp2hVFi
glJe4S7pTLCHK23eWKbZSuMdC3AAF4xzrYb01RMwXuJ9ZA3bLO0fSgJ5ps6cJs82WG/xOkABvwkk
854Au4MklE7BTDLQMvmwz5YLEG5q+FOvCGc9MVXret8JxBglnyBD02UihJQ/wj0il4SI8aTAlryI
oI4wgHiJBzl+b6hC/G3FLKo4l8FG4aQ519nbF2Y1H8mloDPzkjgpXIJ0KGUgnoRSOEx15TOdemJS
gxwKe93sTD/1beUGqpHMlK6uj7KUfzeU843NUsyEJk7kkF1c6nllJNtzWDowQxW+9vYNGj+Pevho
nHtuyWMFIGL2m/pjMD8Wf66uviUIiMRVYeAK4SiOZ0/DVg1wgxcYdrQHsHQBcAV/3CYybu4v89lj
CcRTHxHbpchzX5PbXiMlHLJopLc1GI4lZ0HfUwaPpDbMVEqYDCYLHDv0I0StxDLpAt5oSJIUgx9l
RVIrudcIJUfkAnnCbjptqPCzCaux+Tdo46UxHJ+jYoxX1HlgXMs9FHd11R39NnzppCSW2NpD/GjD
KAyqKoX4K2fjvglCUDUNq+0oTTATJM/KWCxZkBGJ7+fKnTtyayuHaKiXFPs0ktDxAHQfqoaLo53K
ouGBiP41AG61se2dawagBXFNPGGNg5q2kTA/eB/ix6BzuSeeBqkD3wOOA2TOdAjyxACYbcHPzhzy
GjPEIPoTgKRLuzQiN4ydELMnaFJpT0hV4jvTVRo49OdSsism3eVRdK1BPs1bFeKPLpXgxcIYI5dg
JLAS8NBVeryV32QsUf5FHR0wCNi6wJ4n9ncbYY7ZQECP+rxRSwQXUciGQWqf6RZhTNdZtRUaKibO
6dcr8vlikcCJW3GPJ/A8cjQd5xcEZy8OwWEFas0aVx7A6tX/u4xf5oUo2y2EsLAv73ZzQxDC50/r
oSXTUcEr3Bh83ZYBtPI+Ch4BXqkb5A+auFBBWCy19vUGPM57UL8q/bEFSpz7voQx5fA9zb92Yz3B
DGfc6boxdBhnpV5rW2WXOlZSQArcxfRvpZA7lw79q2C7qjV+pzfu+QzM0g6zQ6ElHc3oAPk/9Q0j
PX1Hioqb7/yHTfVJkY3xnfFiGT9AGLZaO/O2XDsm60WlzqSiAVN5f14D7R68m4lzk2Hkz8j9b9Pi
W4zUm4rA87AQiSpjrxTQnxd1dCdzjz+wfDsW4fRj3gazCnCyr9i+L4+LBY0/vR4aeYkN0tQChZqI
rOyNuEv3zR12Q+zqAZTS0RXS5VRlh56IkP5QvIYCDjBUnSW+Q4RwQ61unDeDtdz16W9zUfBeBpRE
7L7Ic1arTtQdc9VsZCPDws9eFTSBKw60yIMzLEhcypZMN/woQo7s1y5/e8IuJBnft/DzwSkFWiHU
lpWNKt4fHg4PABUwTn694v3/Lz4sMsLjV2yf6IaYbe69Vzw/FzO/Cx/TD0Kt417uCjiTWfP1FMV2
CvSgTTZtxpv5APD9MoJxahhbHfoF5ZlhjKfCWiRtdzTVnSZCy+93giDn86MW8qU/a7c5/wlUlAjf
kzNSgYuxMYwUNyZ/e15drqmm091LjP/yzAj1RhEFE810CX5tGg6mGGgG+Pgyp56UB/bJ4iI4x7Th
4B4Zna4BzhpD+UA2eYSeXYP2lLvevAbwAs5STsKC08qLdlq0UfBPx2aLerAZfnXoO6P81h/v84Cp
B65XE9DUQOTZDWraBe2T2UCrzeQ9H+l6lkSto/2h82OtLDz/E54SC9JGBR6jNpQbzMQfOlW0bagr
aQMWE6/1Xgb0MdW93B66AmIH15rXwPAnlESdcgiV+1/MsBCld77/daBWa0Y3/6pUa/16dJnwkVQ+
LslFo2N60PNxHi1bxVaX9DtrT+Qiq0/DxQleaBVpN/C5wlRaevDhOqeQKT7HXmtrQP7/D1S4ienq
k7gYoE1IaoCbWXXCqo6WXTrf6zzZ8qwhXMPwARJjS7ITuRt3sthP3gtir2TvmmFw+lhuTiHlA5gC
ydj+a5YjZ+LKOf9ADZeGgfjhTge6ZofoqzHJT88Rimy5Jt28sa6ahysBJ/ANzPotIjmqtx5cqQO4
npq5D/iKcbPYMq39OFz71ySCXjFVOWNj/gnuF662Jqm8RY6LU3tfHbObCgVIKyvvKqnYGSYFCnhv
KK2w/18xcjgdMS3URZ5QXk8Evr7s1dQ8e2ORtOeEc6t5oJrNBsFsuO4XwPg5y/uWqOKJDmTQ3MNq
VWhI4LVQWs55D4RxQUn3xi9ZRoN7sLyAeakNcu+rkgpWVmyxw/0oCVkpW180iglkNDYxaSYSfRaM
0ekBSaweQgqhdqIT2rYs6Y1pzOuDhP5cCDP94mIp0eAqXNVmXtOj/dObdoqs3Lg2zb2uTvTnMPeH
e0dEnumVoqvzNlY2Y7qdcDS78y2YAcMIkYxAKDjYxXuquws2hm78rJAN2A3oEsTCsPf1SBjOfg5t
tU0dNYLqIuUxrQ/yQxDwE3trAJ0GNVeDJKO6NF13eAIPSZ/65riBNZZW41bjny80I3LQFmdrkbIF
swm8qG4zwz8Umo1mkl+vc4iMMTwhiq8JRc2HNGH+xl569dOhlO18m9gsPSA35kq+qyUvlwvY+MQX
Vz3pqIU9Y3k3TNwUynaL0SY4iTry7x0x2hBh1LVTMpqSTO9ZNnJ1prG69SyR3BAm3I1wZn0ph7EW
Gru+LdvWXKTdXuqPSx5H0lxqm/SnFId1nytVNdT6dDaQo+sX76eiUbjbHGy7l3lvqRQdhvJTgs1m
/1fZ8ntFVVCMlhF7g3aYurGmpTcg5U5m7pboNdmMJFL3ev7ZYHngqlvVcu6UlhjRAmNVgoyTU6qa
yVX7NZPAF2DKwJxO4wIxz4js2wBJeK2vcfAivLbXsXYoz9WrARDHYiXt3/O/LA60bl6RGAfUttwT
4b1rbZ2ZT+I09YzKBjmEjUBtw4BvWQuIcRlVI93pI1MuO2j2CEtxtoF+6lcM8OZJD4TbmiA1Rw3B
zqFpLUKavSvkYHHd3RO7Wh2i0nVDzdHIyrT295RqD+RH1ucAsE7Cd+g9BZHFXgrCbErQrYY6vkHj
svQJGW0yrII6jcMH2Jqjjo5Er6AZPLjVOWE6ooKwKFeaj3xIUQNHFXwJS4JtIXJkCz0RV4BH/cFl
hENNG9/hVNULPiLn9nFqDBJ9KcH2WLNuuDjAsOUpevFfme6RZ/N60XrVu5pfeVSBi4WoolkZpRj0
K5+27vVSVcA++CXoI4oGfc554ZdqHVqVeDn4NPpJyTYxCGT/7mRvIOUDlaerQApOnIvlM31pODrJ
4vwzYxCMLrnm+aNMmzqeZ7qI+gHp6izS+22hcrRCibZOUeAeFqNaUI1xs2E/qPJtPwCJncl6sX2c
8P/S19l9/xl6eeNwxFZyS683+Yr2BANt9WulmiNKgcBjpBiQX4t4qxSRoiMYSViB03Zmh+gUqMlY
efuthwE+FUQVEdp/SVi3HfJM7Z5a7zxnZjvNoruPpFDDluooMm5AvHsBx0oi1Q2B7MD84z3l5h6l
RmUq4aGcHIs7RrFNfeAUMQ4qlx8Pp7cyq6EziMspC8Bi9UVxCDwUNKigzy1SotkXiDyfNBe0Yn+c
rMd4xgfqnX7GYCqgWVKV8ZI2dO0CFvbfmpc5xKjM4W8XEFNgkOVI8ogvCOcWj4dC4Z+hUAuzAGoj
NPvC/ZaLGudQ5xxaWb7XUjJhhljpllyL/RmzZFcHkv+TNV04zV1ATx2+e/KnjJnTSvKmTgZD4rRg
qoEa3ViSDXfbVFEiLixX/y6/lmOqZ59tks5J3QE3AVoXJ5tE8kYAOgn2Rkr0S4WcLhvooY6+YzFf
4DVJOqlumNtx4ene8JhtVrvq1oap/cCXmqU4BOhqJ210tVtbeRNriXW0KFmHx+kdiV6dAStwu3ax
InBY+DqdW6J9rUAbmN/A4ntph8R4DhNDv67jEjrbhV7QlxtcPjtiF42oM/3hB3lFyBTN/lcI+t0Q
svnBlyaIchBx9LE8R7rwV3KFm4rVI7BPzP00t9YgQlirc8A/43h0f+OlWb5ZrRAtsVMo3D+s8emL
7urKpX/wihpc5O6cpijflZOIe0Eub+AWqeY25nuo8BB/8oILjnqVpHG6N05u6eD8AJ650f2Eh4H1
P03/T3BnEPBhBfEck1srmQfTnScHDq6WJYfK8BASHFbUPYPxBRA//2J9vrz2+M8zBexkMyG3s5OB
5fpKyQWrEJQsrVmz14zNAGY4x7LJBdH21aSuo9GMNnmAy1R/Iv5v19tOD77zlQiVIYgjEe/R6vjJ
/JvkI2AAWEe/0m3RKlciN3Jj+gzYlfPeODKp8hBo3TRhaXWce1TGafChSI7nUA02XoO6K1dGlRfS
c5649Li/7QgDg1tgHb3TssSid7m9qeowj3AnngcT8qhvGE01fwWemADfUk4PBDjJ31UkX+2IEJje
sCyIv2IT7uXfx8qi0v0uSU44THtz+a50M8VvXyaAd9y9Vf3veG/Yialxc9aU6K5+DzXRhgx7DRir
Mm8Xda11FQir6AZ23aST5nmDTsiOx/u/5pxa8LSzIA4JDetZbnyJ2WSvnJ+9jUl1bdiCfcuFVTQ4
Km5FWDm+Afk+Fb8jpUtgV8T+0HPgPLX1jb4t8oYCLokTAF6EvMfWkmw39RXBbWPIV9M3NPdICojn
6TG7OA4vX/bJGv5y85S96i+ZRaS5pXNeCC0PrZEvlMTZnkhzfK5fvOPhCVbDZPBZhbOVpPkf+1At
LCYHa4dtdf6j7mWCbwXhSQ55ZkLtOUxSTtfWa9jGd4Dpy+gsXfy9T+u+i2UIzTMCu2WUaAM0CZbd
hfp28fd6zh+VAsdgmHQ0aW/BS4d50F4N6IRd9+IEQhPXgCpZpU0xyfXLRC++0JMyRTAh7Sab+MLx
Ia798g2SaGCwDk34e4hwqLTBYvOlQNsu+t1bWhGYh57rBtrSDhxbUYOFHwVZkKKojlIt3hMOgISt
koEaNbmKTWwFVMgBijPcwECOVN6GLTlZwLEN/o9JjYKO0K+KTfnmT5UL6/CQAxoIquumiotRcetJ
EaOpCcpeb6D3KrMiRU+YRjT87S4+WjaHPFN0tNm/yVjjzwrKsxBbSx2PVPsddT9ZSIbLGGd397Bl
AWPGnHaTF1ysQh9lsS0n7c61Rm3PMhatfVWHvgjnp4s0fVExi368dL3SfdEJqF5dXtaL44lhhtse
1sZBWqVURO6CQZd0hnqo2ghOCIiAn+wSM7nr8CzuswDz4stCdcQ30IkyoK2Qec7x+nKw27kaNyUv
a+p8gkQVAOeptjAe0KwcLqQ2eqla+kpt3X28uudAfHQzFECyO76ysHyGBoAu8tApxnyGADvC7Ju5
6jhxC3mCf9ZZg/bqu4JQopywndKt1kXL+59Ad0/rtzTPUFb1XBPwhzm5EnezBsQpD5IIdYIPeq5A
tf+M5V2cCXmQHYtqd0ZFtfuDkvphyuzf0jR60l/XxZ66DNkLu7JQ1jUSqfb2y3z6Q25zQm3vivp1
PoIpSvJes8Wu7ryN9h36Y1aiNlxi6cQ9STLjwN3F+4mfbPJSyXt91tu2OQyoBPrks4jqoqFApeZI
EgzA2SyfrtpBD0R/L+vq0CsYmw0aLgvRgv+DETDTKEVDUryNYyNTthFZVvBZVXtLPJmNxikT7wgw
9Idb4zTdVraSlwu+3sViOd+qeGycgDXYPU74OzkXM3Y/w/cL+YPQu66PNGKJ/FPb6oaZznrAEjR6
1x80wImTCHy8KbtvczyFckHnJSV9lK7GmWE76GHEteBd7JbwIRQmqm/K38OfLr6UfjON46PgYKJ4
ihpdUBl8JrLzoxkOd17uQ/tASuJJA6238ej3W5/YVwF8zz44tEVUoObwxx2C7D/Cz8Yc0XDl5IEO
8XlI5Li7wzgs+97R/QJCisYoBIp4J8d1yvEgzUoU8l/mOw3FJZMgkEx9FxZFEMIyt33h2VOkVbkJ
ti3zL17YZZHQYgYEjPdn5DQO8XUK2ynRla51FvZFbWg0wj1Ny1R/97pjArCozKEoOCOeSRGc3auV
O6Ng9goGy/6B4xDCtW0VE7Xo8O60MNhiR4NcWI+Nm2PRzhob+Wvkg49/4vajoGy1WpnzEli2WGx1
Fh4rCbUIsUP8dZmVGGBL2NciS0HzzCPW4Lcy/RXFkSVgHdpFlGozFOOLHRgSy96SvdIEQs6+E5Ow
f2ThelwzUEjmnDcsG3SWXtXO7YxmcJqhlAdg4mUmIJGTcOjUUIQTvqAxYAyCRh7gcjf4GuV7XvVk
6Yz49gyP84EBIFG2V/Rk2Tb1Y/bC2s60Fa7wTfMfXovfo34CqwpmfKUqEFbnkIKUp00117S5kxE6
U4ngi2RYQRylzZRw3HWOO07rAL7m1P8AmL11flKb60G0BCW5CELio3WEeOFQiDWIkLVRwsCipEDK
gV0tCACeCqMFH2L1YS293a8aDg1QKgJpiE+sbrSeNAQFB9ifD/xA+kr2iNvzfmddVGRXejOZ0mfv
Z7LlJGvxMcGj6hhfr9s/HpocQTPLPSsvphpSMC6QqnkLl6qZd60x9XYSUtNli1gh90gezzAKWg9J
JHAK++baQfRV2HQkDRFd4MKJnsKXu3Ap3pQJeuFfrP8ksJoIopX/s3sTHrMltjjZ8ez/nLFW5coQ
e9B4PHEXUWHW2FoBcLPV+wxmeZjacoz6DpR6vSqrY4v+1oIC6d/oJgCehWAAe+GFQTVQiTaeVdAF
rZj+xws37k5nFY9ynXTesEYUOWe3mVHiD8HlUjH8p6iCsqQMsfRES3eJxXClLLchw2j3Ws6Nl3n0
ZEPTfi8psItVDhGmUqpHRS2k5F5lXXDSDlwr+7qNox1uubLUUjdrVOLh0bRwqxq7q3PqGUBTqJRb
WaZgOYYPXUoRfIM+nlURxnmRi4Jn/yHte7i661EnGSjVK2vMD03PSERe544IOuVzBXdpTU5cUvis
juMUc26Bl+obqL3/gOrG5fY3WkYJe0h/r9sufZKDaEC1tNHYo6vcqoGH5eIZZazv2gQ0hUMbNN87
tocmKEEv2ofThcDQJGTUvrKEGCTloQbycDjK0RBzCB8ew3I1LophPJzX4zesjW5WkQJSMEuw64IJ
1D6Iah7pS1FvWXeXVLQTHZdVGxwo+jlHXJtBNvMuTZDlio+E+1ond3WuZBqScY/T5yq9Al5HGaFq
uCEG8ZMEpvO638sL4ju6LrSP4APIp0j348ZmEsUCIBvFqO0+d7fyEKxcFzRSv5F12RfKZYIPtYP7
Q0vIOHMdnLKfaPnM1yWfXZVJGE2ZZ9/RkmNplK3AqSlcv5BfUqc3TDXqA9hv4UCdqxZl9MmKUS5x
eKBWyRxfjFlXlve3OX90JBSMgXBB0xhzW+bwBwwW4zUILs3X6Jb0/AWcuw07oW0kzAW6OVBaN0/F
qk7X4KkgNBO+fXkEsdn/OedkdsixEb55Jn+eXGa25r+E2npI2ayRkLJfMz91hWzerhJR64S+EIih
5jihCSbSFZsWeyoCnd4BVSPVvrkJHX3xWxInOLCmsuZPGpDvOyd8kBaHjqjAt5+GEDVhFSYP4fO/
EhTLYac02xrfNlyY2KSaUdOYUyM9I2Qkv/zVAzUk4P2aDhTtWLYGyo6xW+ex99nh2Q05A2yJsawN
8z2Cd+cNAUx4nwzu7PZHhbPsvwNElJEgdK700SCEvlr/EmhBO/JX1JuOgZxfY2ub8jsIdeMWMZrZ
s3NN7gUEJ58O2R0Vw3Qx/0v51wf2FYo3O86p3r9Lt9GHSc+PBM0lerr0loFFtIVm3JP4OHm9/Uf3
tmH6W0lHphkegaOHLf60elsQ9hBqEbgp1jAG5kZI2ZHVGM8ahINtSrwOhfEcO2J7F6V5QzaQRoZ5
hSWU+FhFNQH1LCE3d7QDL3fd5D4ddnVS/eMw5Q9WIK8C6kqjbfIQwqMSuUIRGYRz+uxAoi1HKrXv
194n6BJ1/Ye+mkuKgXtuXB7C1UjPypxUui274W5jhaYPJdUyostKswrrNYsUjdU0P8mOO0hgZm/9
IP6BsGsPnsEDfjrw3gcASlKmktTWex/X3WprcgKz/RqocJxY+LgijSCcbhfqywU6frEkcuN+Ioiz
vHJmBzbfox0y44C7XZqNJgcf8+v0tCsAzPUef5l9S3UC0f2bVV0sRPuLQiX4doO2VftZl3t5kyxt
R70JX8KAnYEYtIUm3eyzfmDIjxvsKzcf4YH/LPLVwlVKFfXVxpqs7B6HLoNaJqpwzXhHOp30gVCD
PZMbVSqcQ7r7tuxgw51vYEKFlxGIlR3MEeA6PDwSFcbnmivQh2tGF+mmL6EX7dBe9jsW+ZNEKl0A
ndvZcLNsaDRG9qTJU/EMpq0J/9hRYEPsauV35ZXehfApJtmHcLbZ7839qE1+65Kz+8U1Gy1+V64Q
u2T2DJONdWtSU8bHQ+EWsNmNCkSDPDRL44spyahNl7VfoVdN8CdEQ7iCHammkFCRkf3uIeMxcqQp
E/+/Cl8T5LwgU0Bjmw+Y7Z3LKIpMWaquFteyVYe8P5TkQAVn4+BJTPVoc2N1C6cMtoIGW/5zt4c6
O7OMA/9LaI5Pq3esf0Qy3AEuynCB6KTrz1h4Q2xols9TE4mHVroJ1+FXhUx4/QUdfX78F7Ey7zcA
BzcNC4deD6QmiZxe+g8jMSHIaNk0XMRYH11rZl2sXT3oqKydLV+mFA+IIthsD4rwxlgzJpwNYSkU
z4Uv+BVEbFFfpdnoJ/1QCfLGXbbOsZg0JoB1JopqP7xA6fp7wY6z1WJGfRJ9q4gPWVUfnB5ANpoJ
u6yPHr2nzJUgfS13geTosSOE5ZJxxksJ1Fx2jv1ronLGhK/R5ks61RKiqpQiNQNY0PlZVqXv1FtP
habn98+TflfE2FcrSIRhzH1tIiKx8v0IKt8O8X1jPm/BzMqvsoDk/bS8irDWTQIdY+Av6uK+/l6W
bKsE9hiv5IUNVSfWFWIzpDqsu03jHsk+a0pwAzuhRa/tG3byaPNWipCtJ71pPNDOl6yp3vmajKv6
2YynHvPOllD2Bvsmcwib4hkCOarcULSGiFbQKrJ55AiO3sP5imUFrXU7L1hHwgeOO60MKPZeLyWM
R2Ul0K39oGoIgfkSlF03oo7/5y+ErETfXhk3TmhY6s3MDDzggQ5TwRotepps+6261DV1U341qfhi
4vZxBVEw23cIUR3DVIR6EbCiOy6lbfXVmYAWoBVLVzkx4AqgMTQXvlI52n1hXYNdcz0PzZEOgGm0
wAtDeEqQT8izf1cJSugfuala1pbEdaVzG97QQxyCD62rOwiPDDCUJ2QPd7N6H2TyGIuSzw6O5tds
OUjMULJuZlCG2scLLhafBRzgx9dQ17ShtBMOm3E4aoE0hWfP0uuORFIkKTZ8kZXyOevtAs6jJNWm
LvpWoESVttSUwxs4OqiTgFgyKnpjKODDqK/9+QwPHVVvLq3OqtJXq9ciz18qxupL2HJrlIKixV0K
lFMOIQqba5Kq9/ddfcpaKl9wA5mMBqVRN4hQJyeMxEWv2OFvQRTbOf0OUjNJyFJg9Ns2VvUGAmZ5
rDosK7niT2aCuZbQrYphRkZt6oZVBKGbIFnnf6ouXkr44syIKY8h7i9BJXIr8lJiBsEB1EzsiWYU
MKDQpjC1GbjN1IZlGIU0vpgXrTapt8MnMeVFXD5iklADayoK228zbZVJTYn0RlcKdTsheTwG7qux
MVTmeISExvIECdHzUBNerfuck3XidB8+VliJkSfmR/PDdzMlip2lXpH2Bccm8FS4xCRIJDcR8XiZ
+3c6iZPLBeATxynY9QbVamTnGcgbDKC1UFLMp9HzCSrm5d1nt0Yj8RF264IXTwcDjj6V0JUOTjHT
aj5KC9d2hQGNh5i+mNacCYV86hH8C9H3ftQn6IHx1fbD3WACFHIBea2HlAQU8JqArJ5qcmO3DydL
r9oKRty9qvlMzNLG0SVG+YH4LIV5LsLzmwAP8tm+AdR1AzqLs+N4ygz8ChgCU7w4OmnD+1MP3MlW
44LCkecyk57PmsmDwbWjShqd/Ads3FPWyQR9NAB5cLuEX0ydAFX50BB9sfzBhawjhM2l20TEbx5M
328XEX12WHbOVDtIp+lXEgr2fBEBCZi4TcyyGnvokWKq3V4UOhUnWfqGesN1IICGASGkpHUps8bA
30T7/Vgwdi/twg7+s/B7d8/TLTKn80e6E+fao4lcFH7KxdLVr3zY5Pn2oiwBGThWKMYXLGb4V1cW
6MxVvEnGOYTBsY4Lc/AbYA5hUfGShDEVXNT0L1XGZS4pertyl15LpSHKvvsbiWHFiZsngQZ5JoRs
kjbXUMuFomjVpZWFeZ/9JuHBBje7z/LWlBfbe2YMaZriNw5R7mw2Bcv9SA6TPerfFjJ0AuSicLiq
tQ0EeEc/t9+mqYq6APyaX+1f/GU5P8WR23vp3AAiWwTawU5/4kR4Xm4VxT0FXjJ+n/4i2f6PJjuI
JwGrKfO184ZyL+O6cXNJE01oSFOEClnvSavEQIz9hQexstPHDeD1r90FfGd9QRFzYGSswR+Z3L+6
UyajmBj8YrpmXrFXBAyL6vkZtZRXaKPObK0UzuvYpEM495HRCQrCURbfPJctE1yyjnK5B0qehX84
aOaV3l3cFd2UjpOb2jCyOlRCa4b5kGGDLq4whHdtwdg8w+bCEWiPfxyEcwdqLCdBvwKr+arIGsLV
8RZJrahxkI4m1QiHs/GS7IUyvz6lBb9vf3bpiyNeg/OXgRtFArXz6wrvB+ZtC7VLXg+RVxOgSurq
IdWQ9D5kUWsyJqMqpD1uNrGsFFsNVfGlUrNH1gRLu7VT4J45DLhbe5aDhb5on6NQyXBcB6VWPn/9
5frXXG7L9advuCbdO+KfXKOJ6iFSRBLOBuVeOyqlV5EGXisjJ9pTSi9g1ClVxaCw74zDNa/c6BXY
TWxZ2ZH+JAPhyRW7VjiqwnsV9KYFsDIkebC7Hn41KfEZqdbcMMGyS6KsZwyXKivPq26Y9MHwBk0J
Sm4bEfV9oMGbRFNUKFWVBKQI30u6xRJKbKpKJAG4kFILsjKa4xyovLqeLGsGLgneX/5mEsK2vz23
5GAhnB7J3rT4pVmzWRbJipJTGszEfoy6HSq4SA2Uv/c8ZNkkhJcKuQNtGta3zacigpxv88SZOhur
Lubve/biTYAmoJ3H8aj+f5LK++Tub6uuBtjvHaQpuntv7Mo+ZP98zg3rVDa+AXEVQO21y8u+g+DR
ExwNNmg5ACWlxGHQrQoNfypMroOTbKDiGtAuUNY2dxzBoS6LlskotOIVPm3U+KWxAdCo87sdWIVS
ZPAXhjdkXuu1FqOqAn7gdEFAgzqsj2jgECLRTzPdgDcHbwZ+uWoA2K8wabVCj6uwh76LrKIV6JRq
HH2XRKM+lVfpNdK2jHl5qAgN1QuVgM0BbEPnmRq0HArwe5VxXiwZmKXo0EVP65J549j/GEGXzsZW
t3I2XjMlfnLUdnJ28aeKTLu+jZUl4Ql1Ly1hZWO5Cgk7tKKzj5yUHnqgRhk1hVAxnnpRd8TqJhMb
h+vVnLbISTXorXIBfAF8/OSrFDK9RWxkiFQF1MkcpCYq0Gme7GZ0XlA6eiuQJgVEJj1NbAQBGpnO
V3dH3ykjIm0io7ERRPNjXgoBSZm3kYnNMfK9t5LKz+9qy6iD7T5JFfc8tsEnFykMwYLcBtgh4wrS
+/a8KI1wOt4L1dwWTSiLNC2cDsXjy1/SYcFP8imaEgIz+lXtcB0E6VDzUH02Hv8sOXQhXDG26TSs
IAPC6uOZXcnZlalNEUVgLKIALOPGCJJrJDXEZfoOUwvd1tl3Vu0RwFErL+qCNmP8g567ElrNlhyX
i120VnPmQG/AUJCbtU57L2N4Y0Rjxc/TFij7tcEIxqCQxxZIBRm4XPcqREIXFFqm1E8h3U+tEIw5
bgaAOiFzem5WntDJ3g9bHlprmQBwPXu8FSbQ0LbuzqgBYzagmkBBJeNwNn6kBpdAVuwPI8yTO6nk
KqVpNrOu+vHvwvLUAr1c+LpJrPpRnfnCOVUOs5Z491sDOWZDjWrT4k7JyjvNXUObMdjZnF2os4Zp
A/CgVjDIRbeVzN2qERrJzB06pHnrzeqfq9EXurjlypWrLRUdaWEl1iR3M6k/1OSsxRfH1uQdwSq6
6ACHyRujX5IgvkW2WOvYy9bARfVG0r8bMzQ9l8xXBlNbby8+uxpElp+4la6jLbN04yny2S+lGo+z
2Q4AMgAzcxd/J91oR8fbeVGbBKX8aa4nDODclqMRI0ZWHasH3+H7R2IL5dVPaFwQWy+bDBB9/647
RigtGbypNm3a820dj3G/5nG+D1CWes6eCTRfkgFVs4XotnrUlimq0uHrt4tnygVPUmmVCE0b4NIj
3OeslJD0fOsKfpFFVNVoW3jChj95OsncDJiyGCigTRO/SGFhEkdARcLbv7I+ZSawvGUQ7X0W1Tp4
zqg2rVhsxPhUnjGTPSBcx+gmrzFNJxYVaeuzItIAVLmrF+fRthS1hfNinib6uuc/juhOYkm54FVO
VwmFn36pxOtTltcCmV+/Q1qHg8wovlHF3Hg8XZ756BMViSsXq1313wPj0slewAuLWR464R920OCl
QCfW7kAjGBa/+YKdn8GMiQMoubYRH6m7KyYdHzGBDIadUgF/y97TkLsDroDe4GHYdJtzT29h5s0Y
ZYGJrc6/3vTHOicQSxYIZmcuEQP5QfihoCY0rrophBAhgCtyaFXYazpg6UXQsRDX/IYrCgnGFxAq
ZC3TM9k5WjmBLw64jhv+fSo0wxo/kg4gyYpZRxH0Y6Y7V2jWaYzOshn661EdagYEVy3IuZ1WaVdn
oLzIvlis4atfatLMnsvkwed8BjkXxDUMkYaRuhd5r/0MkCZ2bWSNRcx5XveHA2Oee1FnzDOF4IzM
qisvlzPihG506g5yDkVqbnyFMPFlQR6j73ERwSC5rXXZ/i1pmB/UMn6GsFEOpYSxEUST4T2CMn49
vEQ5myThtpY80OwedJA2XzLDGiJjrVCXYX+OBqBg9a9hFLRrSxEOt9/tKgq6daduZDlhQY5EWIUD
l2uWB8RRjMMEWhc6p1+XlA1HwOe2FJsVxuneVil9PP5sXC+TXbQT0evPar0S6Yn8PBtipdRAvLAS
8ZygQVJ5e4zcdSRybRC8jXkalSq2zT6YNl6zuplQYPDowkoeMa1ls6WBsqyAD/+/8XiivyQe85rk
w+QVpkT6/2uOMYMu89nzONXrTunaSJRIcXmdwB96u+t88ocuHLk89XTc8ybE4tIL7T6IcJUhur3j
wCtRiH8JYSNg52X8QgyNP4Bpjfj1IsZMoC10P1TJidB91qstCwfmxUR4oPUTb+lejV1FTyzMv9PX
X1ffrvl72NhqHUJm6Ub+Uqrp7gZIERjF6+UfUOsVgqupDr7X5vMbIdPUg/t7OV7WGGhmKqRUCInQ
iWzACMUMqmgrctgnXj55h7xGi1GZfovineYWCkAzfyGPZatTkWB1dxnlObxRMHfbKGQzvKJVIc3e
eo99qiwu8gK+avT9Th37S9prYDCE0jpzDQ3V8RnNJrWW/+i5cy2kv6NuRbLBGmZ6+5poq1RJpISa
JsdfSBRqaaResAIM4tDCtX3pHFz2tqzH+p0hWQgYtkjtWSyPO0EIFOUo41xRHHl2wNQ2fdwRqTjf
M4Tc/fxeWOFq875iBKctwHMMAvqN0dl5Fs6XzEKiUKjRirbMfDJfjmvfoPQYDz4CIgwv0EKZbjF8
bx022szLWnsj4ITZFmBP+6UVZ0UOq61CJbOOEiiL2TPuG+p7NdtRZ3S8xgZD5GrUr96oDsaw89J5
aFU3+CY2I3zg7uThjdxDXLgN70fAL1YKlTgS4m6enE17+OtEd3JxZpxzLst+BE1Cu907a97K+7T5
zhBDsrQXy4sRpfp0jUnLmA1x/1QhR8C8YXGnbOqZTzm6+94674AeBvVI+kksmt4Y8LlLyiMo56QW
hmFR7vBPx5LRipBE2jC/Iky7gPFmB6ovBo+/C8556ZfXN500hgWKbadhMl9AQGCnNbbsW5Zrs7Vb
aezJKEN45zX51Zt9USxt+PxqdXM7S5EnUtdTj2NCjleK1L9sZUY3KIeOAw4x7G7Hlqifrl9IjyN0
tpB7chg46/f+r8yD3lK8miQGC3p7etC3HRsmHFF/QWE7ijZ9dEVDJQfsFw+n51I9i9KQ9EjtjHDu
LQY1d0/q2HO9yhrEiOQYsJDJD3K8S6WsdYvBe3XV5SgrNWyfpzyitc2U7lbYKVGrpBGD0xfJHAkc
eyvoy8gnjlb0ci/GyUtaH7G8ZbYmJDqWfZ5vPEek6UaoOcvdp7F3/MpaTnTwvZOe4NqvPWi24HKq
iNjoXUWSNrP6+b9Z0JiguUPQdLd1nOp06vqJ89nAw+W0Fmu1BObHSslqxDZQyMdfavpnzasV8h5j
yP7NVhTiojod0fpB3E1vKu0uR3/tqbP981wSQX3PZV/Ph4FuO/xZQHgZ6NyC+lsZbOcT/RWrKjfc
R6jxQTF8f4wuujqgRRU1BTgTjoqkGyTSeVcN2G0vp4IQIdznRc4MKz//rXH4FDHT/M5t8Eja6VVm
sYkUvXnAIzFnmuwcM4vkejOuEJ2s/ChEJd8Zkltf6E/ELPllukeLmhztGGqxqEmJ1bzxM7awZkqU
o+/XzUqQz+Zgm0PvQeV+Z48eS5vNtdLXly2VlP0sHkFA9udyXfAJ8mtIXqS8f8716oFlR1ycq9Dy
fwYByM29zNE0kMGVmWKb7j3p5Y9OCSm3M8S0KFOpUhIR3GEA7dJzLk+55xciQJ97Jeqqanj9qh69
elsWl4WNARwbNlj7TsVgBeyoXftTHQmwanVIFcv3rxp8hbNRlfKFpkdwnknOPb8kBuSdOVdPewyU
MWXnBiVx7c/XtMtQdXImr0B2KEBiRReeKkzOt7/8ZHUi0kemxdZVHsg2jHjkt7qkx8K573qtcP8I
3K07JflrEeNL2BY9ZxIECmcN1g9R7PWF6zOQdR2PTmjgGw70zkcwvDQ1WYFNIUCbki9uHy9azAmC
EQuE1WSWEL3CwoKuS28Ibg+QO1eW/Q4ybDPdc8vmwrDlB6YTqW5YDCj4DuyWQ+RKRbhcuzKrOPsl
j6rE60z4MO06PZuK7PZlkyZUZHV0wHHFSorViMrzqmanXwaN7zMV4FOdt2+3E/AyIXlPyLrn9zwJ
DOS46gq3oJ7yvmRu+lOYgkrMd92Z8x+WIlWjoiPvWFmqVPtl3KZJiFRWN+/Ahb44pczWwYrFDGYF
9WMCjTK5hi9DWp0XUNHrGS3mCxpT3rqPf2T/VANaUYRmagY00Ig83TbhC/8ACGo+/Tw5OlNtgK6r
FWtvubMjM75Fw5ycGNEnQR9xsJCEC5xmJ8odl3ubrTdeP4jaxSH3sLcP42ya8wUBcW6QMpdhvFCr
9sMJ5enkxgBY6UdR61gwMc4mgjeKZwTm3joxccKk13nGDMZDfXXE1iZkOW9mocxSukzSwKj5a+VS
8U5jYo5OrHvb8jjdESsdCG+JXaT9wHxX7AfMJ4kabWxwa8n9Gu2cZa+bHt6z89C7V2GdqXEt8MGt
7NaPfWcbCTeiPMbzgp2l3OYTuGANuElKvCrUHVIRDPEFKB6780cCcF//qwav4Snajl4ewKu85JPb
XO8GQSwKuualhmIfMOKRqAJsaWVn3/xf5Rhn5SnWX6dpZGOAE5jlJ41ZsiQJiyo+qZOXXa7EjGdb
sx7oaf8ztxg1xzwmfS/3XjVVVbdXMSMNH75xH69B/hwXEL9GbGc1d1sB7OQPH4wOtalFcUXsm0ya
tYZCSEovP6eDBt+1BZi1qTY0v8+iJyxqRmKuOA7iEjiuPRZ5R/NDqHiBfRxLIHuZ/dQUZLTOCCcX
7BvUhbuvB0Nkx+jMA05fRTxTkeTQGN2Mo6Lm8cCp3M+z8g79qxP8di7DyYf0AEoZIQPgE/+icvs+
giiaSjEpBzrtZ/SmCU+TnFV/hvSFcIUBd3137CO6/y0sv070RFMuhMO+WxHl/ww9rhT0hcrw5SIS
7OY8SWInY0RJvd89SNTok4x1V/rWAEIio7DarqeASbN+ZKZw6GvCZSQDZkxrjoO7B8ji5Aq+K3e+
8zLS2Opd4TfQz8ba+EmRVG+gGMfounPncfPv9RLhDdAy6CsU4C7HJTFF+CTqp1Z51zRz3fPKkxBn
JkMXez3VS/weoBYKQ4vlSkyW0CmYPxOgEZQSARdLV16xb55qJETXSUqX3Ks4qhdSsJh2U1D5+z8j
QHrzY3dmyxRgZl2KMtDcYlbaogfmmn7w/DMMlrMYm8g1z28vDbVl/mobHZ2EhH0jaDf0ajGcaY7n
0nGNbfRNS8oMs6GgvwmRwPDWu3Va7m758Y3q8jBgurOQ27TOr7pOopYBxPEgJrEOlQm1yDMz0Pk8
fM16/K8fH3kI/It8WaO189g+0pkyFTe+iI56bDpfCoZnLMXVJ/5wXPjivJfzNW0wiO/DBHS6l2ZD
uOiW9I7GL3IydFWnFRfK8c7lzLLNDlAsghFXcY+y/VlTmDUBBisVnO6V5tcMblSeahgehjxRJNfX
42/RHSgASsUVu8VW8Ra5wcwTXcMH+zTDXPiuGzA2Mfo1re0K/H4z8KwwXglx0keGgkRCkLoM/bj+
yAtszhN41X4teQV61yRE2DpBA98+8QLNGmFa8Rh2gR86nGcyu+HSyx/eO7wTpx4SqTEcFgcSJtKe
43sO0po+xZUZFzCQPOebygl9feCifbBcm0AWnlkJj1Q5kYWIOAdzsp4XOMlSg7HEXLYH85h/tk45
X+HPBGOfOyEDwz3gAmdVDlZATCSQpHQO08Bd/HcIFJ9nt0zpjxJTamDfJ/rYIwkz+NJ4WO116XRx
psKZQ/78TVJIHBjuRSGcJzVXMBfUOkUpWC8AupNA+v644iQLUSGhhC7pXYDOnDSNmFrE6ghu0CWd
CL7pgp2W0Oa6A+9REHvpmRmsd/knhHDcuBQUdAyoC6M6zYw2DcB4cJywKXOKDy4K8gGPBVqUIutM
MPWbG9gQjhigz4odq0aZNpMSL3HqiOErg58eP4z09ggJeNuy7RGgyijngMJAzozbuoieP6ghT3NS
cGdspzkGCJslq7M366bwrfHGnUfrb4FxwFcSLYIaZTEHOUrveBT25ksHTY2vodHhwi8vReMRa98U
rDpMz81mhWBiq11LTrOrBaWvtHJvvrew8eRBxe8p0JODmfsZ5p//qskjvYB2/xE38nQpY4ikNx9b
8ELI+nGIAq0IPeEHn3jgA5etGmWCpPMlp3StiyvK6bUnobPWwgQrNDeGpdEQ4qiZ4tUBtHXzKm05
tGSvkMTB0XO8vr2cROAjooQR4HPeQr6gRU71hW56Eilgm2koEn96lFdt9YprUooNEJO8lNl0pdwK
UM/qWNE/omjPPpY9NDg6gSFwdinGuJHQD0ykAd7o7qiN5GypeOkoy3TuleMHUiIgvDW1IisKNGKS
MNU7FvAsTO0GzNsOaQSKL6GqYGqHs7diVl9hSHU/NcR73FVzAYUV9FgE97i3EPXDhgRaD+zcVPJ/
P3CN0Z/xXbxD3PNXSV5HdHzPOJamhp8pfHvf4WmNoudsTRdEcvYjxPGGM1E1fugGDunnsbIUzRFE
mFLQ87lOJYpONVZLa4v2b/xpKUi90meKWfBVYdm1AhqOdLCRr/vaosSdL1N4UR+AEvT2ymziuSKZ
/7ja4YbVTQQQUR7GB80Ha4TpZDvsgNol5BC63341HfoHx7K9PYrhbFvEGC06p77TxcTVqafv2mpb
aeA6/fyVLHWeRHNdbe559mCKO2mgR6pE44ns3aI7Oo3vEt2yA0Hbq3S8HuNZefj2gPS4DU6qDESw
CL+NpL+Cw/+WgYmR/YxhQfBSOX5aMduKU6MsB07G4Xd5uz1VEl2bR3m6vzIUcjkSAzKXC/VF59X9
vZjfOj5QyYGRwhtj7qbePK0HphzfNsQIWD8rOiaVwTAQPYvKS0F00vXOM2xPLD+XlvxmmMB32pEY
XuuoYcexw+u/oPByGYmeOmXzopxiobeyAuLXmuonQSnIoxiRl5aLnYXZNj/SP3FiSz++MRPHIoFe
CyFOw4ZT2rwbIp4BvLWqzELPVxSc9kodjvWASfKuniE8CtjU75p5RQ/J5Q02tB0DG58ctcrRrSEz
JDmN1DacdViFljNv4ycqnbh9B0KmKgDu8B5tVmztTQXVNo+eopswIaSXtn+SweF3ie1ij4CIaeA3
LT2XVo4gM0MgJIksMecR5nCIwv2IdO4r+Am3Ivsx+k5DXOI25FVpjomEdBL+Myqzb9AoDhhTturr
sNifVCzdqEIpTmcsn4Yd4LzNsuRoIYp/4w7TcY5oHDsZro/hiUa7gDuULKNf5HFdyA70MqiXgU5y
7BM/JWukHC0zugsR6UM9lWV74rVT3Mphlx4GHhfhS28wOiZhsXU96A3CQSsFYx34nxmZIAyDLQKb
Wb07zduMqf6vmxDTAnpg1cGS7u+ImtQgGImd5c5WgVK9rT+yGKrlWEYu8e6FTunnZ6tDxrSGj2EG
sGYtuMbJe/SdLgWOnhnK3MO2d4sFHbwdDaB1KiAI6f4xQRyTivk04/lNfFdwYCH8geLlXsT4lRxJ
RrzgP3aTFtRp8EbzULjH20YxoekUQZ//ykZGk7dimNrSURGGqmHZ2ITMhCSKZYh7RM71r4D0slq4
N8AC0FyTSj57OcrJ4v8i0lR2C+OtHewT6v8K9wSTevDSvRqB0AA/b2Dzx1CK5Z9ZRatxNPW0Ppxv
GQts6ZVDXcooWHjnOI8/cm7fuIfzDaqpYmknalNEPklUatnZqIf9qILIKw2I/WO1IuCuBPPYvLlW
4PR2Gz6ZWY2NUELDxP1C7Z8DNE4oRKyM29x86YdsoLQrzlYNxa/4cMBJDXuxlnCLrSpN2AjlY/WJ
wUiqkHdZ+tcF1uubMVE7UKyB6jzJGrPxTjGRKF13q/M4HEyjQp4HMckfDmf827v4lzjlNa5PtzTR
SO0TIqBE0FAeoR1wRkojhFlt2yNTEp77W/2MSRuQEV+RMxgSZfY3XwymDfNZDzjJEMqQRGtFtW1r
tckV8Q/UL6P63IELDr/6RUK3iqgeJbsK305EPArV3J2yJb3e17duFUzkyTYJ7XkAvdp4yzJl4M2s
3Iq13MAfPNi6ndrvm80vfmlchOW6xczF4kC/vkrA19v5DSWgQ6k+b3ZYgz4oKT6Aj4a9D0MwDqy/
pocSDIL0W5Vq+7mejFNBcVPY1mH1cmUtk3xU0GCd+EHQGOhdVvoYEXqyLW6xMMvsS/MCZy5ybAay
wu/pf4dWQxu1SaoTsTDW8gNlUMiNTSeomkM7Xlc6CUI052RayilN4AAJSWw9Zr1s4vmNlL+RD2IM
OjCoQJT0g82XZKDdQ7K+G+W7Tbz61jAqn5yda7hL8zUgFHxtcPvOPaapdTmW2PD9X2jDIUTxcWtq
ivEwipU3tg0reVhWdCtbvFLI5XMp3a44jvOgdJ15cSRJMRsbtVk21nDIuKk27cqsbJoOeMKgT8+N
c8FMg6oF91bC5T/6xFric8s+pwZ68y2HIt3aqTJnPAo8J/8rS/zEX6sxhBrjmMWYBHzvm6+9oIO3
dkNH+ykNpFeOFRUhgCh8Dh+GHCVDn2eWoaXBStD7TsSO3bB5xm9V9TErA77pPNIZ5m6BvCSaGYMK
m/F+dj4pQ6lVUKsGuT2wxxOIQz00wLZeF/1GYrcVKXQ+m7O3sAH0+ys+VDSZ/MzxGStX6M4Ro4/B
Jhj7s7Bl22QvZkqySll66GlNv3qHyBfBEAwKZbI8mapyzqaeoW27hm7bIMH9dM1pg8e2xumpEDDo
uztFE1MdloOGZQ/38juWW/bLZXHMjbhid5GFmGulK5tNrf8mgxaYKK5cUNpgGOOVtRzmgV60IMDj
EJQqQ/8J3vmplJlsmc5KmQCyJ3XB9a/Rba3ieSp8cvdHD3yMSvs45RrGUK5T2ZYKARD+ONEGBzle
UgaPW6o3bG5C+GFM9d+BWR8/+M4l8l4ULFy4Cx54pcxP8MpCoLQGKVzjQ5P69JDLgi0mT/8xfbTd
xNQDo6NKlBJ3NqNQhYun3AUUGjsnur255QAiZai6vqbgFiMs03RJkdKFRE+wNlcUlpWn6fB90ZVP
q7ZQdlpeQh8tg/RgQaZ3sGOhneirw5jV7jCa26csy0zX6YgXmYhz9ZgGucFEQenOmJs4wjLNkJCe
R0+fKNgk3icuE7cY0G8d9PKjTxegESxvQIYPrmoC/p9pywnrG9CX56Iy64YALtViQJWnsaVusfvw
0OGWz0dWh7Ap8L0yurimU1BOccTHL10Bja/D/wFaKF8hUwZLCQJ2s5JkRB5jqmw3QnmGIgDx4mPs
6Bb1bkjNSOp7WKiLedRFo8IT7xLCuqAClVPUMvxs2NLH2ehpj36NrAR4Hqw/LctobJZlmsj3YtKp
07rZLVLAj3GI6poUBQY83Smpx9Aw8UbXmrq629c1+8PvPZPVCx0VnQKUBE2xvT8SsJjNKqSXpfmQ
l6nyepk1UaPClG2SsDUzGb54usq/XQ78Rfb7PMXC8etrYIcjxJ68KSO9i4wWRnEipAR0KlP3naaT
AmMWQV0sT4oP8SqxQwr0OA55O646Oq/cAdsxBbqz2z587wgGO39IxyC72yBktgfV6zkVKANqaNMT
bnqjDT/SLQZqqEXeWiSZfbRPbB7i+9J3/0EA+UhCbgP1sxzmsJ1pBzxzzkIr2tpb5IegbSG7xqpi
amEWv95iD/r4U835kxnUK48su7i6pxHkfiRiAfA6HUFrtua6yUKi1eX/H9bWNCUvvtH4ge4kXHdb
07n3/msZk2P6uJnk2i5gVRCDNmiuHQD3ryybNWKYpBevOfLZhSfutCjKOlrUq7JRIN7PQzjj2O7t
9lxkg8vGohgPO8pFugE01LiBZGNx41DHPR3rE2ScOudGg7oXZNyqfdPI/hUh0VlFW0aC15OGpIYW
rbjciMp8mF/kzb+KUPbIWtyTznq/7quvlrOjrHTcJx6I6G8EDUPeWII2k8ptQj0mtmCQFyxSaar3
iWjeDGP0C+PUNui5c0sL1hH+nnuzSd9r8rRYDhmz1y8FUJVP4n79nXhlvVxbd8IJoX24KIyhdA5w
3hmvsq0vu0uh1hiDGpWZ+1bMoKmgDLp6CwBNpjqgIMjCMSG61tF0GjSCNy1KsFOMYiFAIrATqN71
9hg3zOxjIYZHU56MSUbTb4gzHn68BPkEF7Kmt2G/hBLjIC6rMAASdaAN7oO6i2RxBXiHUHS9Hcfe
2kqRCgAgk6sPuYNHz29L2Kxch753O4WtLoSD42BxEPh9BrrPLW2gtq2BfmN/MEE6byuZnpij+h6N
535g9U29H5xuFUIICT/f/IIXgyfFEnxJY8/GoUwNi6xYyk/Daa6ZlXh0p7FtryMnRUEFcOgk1OQ0
B/Izslm0f/IeBm6D5/fDv5cj1C3QKAwfhoG1KZ/O53EyfG2mJPmoHYieEx0xHZKNB78n7JKyIRuK
7z2LCgqZWFEWkilsKoKdyQpAP/YeQXzEwu8uHyDy5pgwTpQl9FJVCWzVjU7bpJY607gYy1q7HJzs
BgvNFtsWQ02/3wSsWAaNuRqTxzXWxMh7WziKtdRxHo8nwbUi4aghmKHdBb2pFJ1y1S6uzkJNc/W6
9IQtbO4QQH/Ov+xslrDXQvCxJpQs5f4r2c0XwSvF6bSFFnNR7qRwwP06sIilrnGpzUcjv+o/d8rv
b+S/GAuBQZGGCn5Nolk0CRTq108CP7VPLceIj56+Y/axi8egGxaBJJgw6UH/fBzvb/IGD5AJOErv
ITkyynioBnUc9Q62NFrMLaEvwjnr8oy/uKWRl0UWH63Z1BoOwcl3NM6C5E5vKIh4hlkhZNnMv0cW
spludahTiuui8FANMSoE2kxdVtkts8Xzaz6Tu9cAN9VMKGmpA9dEjOifOfMh/lMF7QDV/blnQAWT
AXZlw3AT/+acIzyyy4tJ3pdlzUadM2lG77Ghadlh/u0QukniasSBlXrT8x2OX2KzSnYwgzGDz6/x
qUW4MJ1x/aycBRHGLhngAKHIBXSO+qhGh8npbQehNU2+tUTojXcr2gGLF4PrLJkXOue3Cj27b9ax
QXJy/Pp3jidIGDlGcUHRcOH4QUvBbUAU0/YDM6hm8ffdb9DiaETpHj+neFy5y5n+gc8Iz12ZYKpe
If9UEhd4+t0AGQnNuYRim1IfHXCdgwTNC2nFtJ6ul5vxOHZ/eSspmzFIlaaVcOISNIUtqcd8YSfv
fN6s0udJHYw2BwueG92fjMPcpKpg+WgMXQMT9ors6aqiQBXvhU6XZZl40HLqPD/gGasYysjk6+UP
+Asr6xtaIhrO8Lvkqxs/zyoyyVNmHxNRegKTUmKg9GYHeIU6zPscM+68Vbkg2xATI5Mb/79Ux47p
JNc8nnl1UXpfI3tWx7y3kcwAJ/UxkG/TGBYSqyN0iBZbkLAqJHV/nLVjzkTWGR7p78vkiJgo/rnd
rDWBOAHnXeIkPZ7Bugx7xEMIgKsHBS0oOUUSqV4hIju7BXAE8J2MQUyklMVK/QQKgArVBd7XGaof
4FwVMBkUvh+YCO5kGSMQt3GA5xr+j8IThC3dS8N2348M7yG3KGjG+w9rIr/p96pyep1VZGNYz0pM
vqrEBhj2OQVO+/jaNgxJQ6BGCJffCR2Q46DJQ/PME/HX4tXgLh9IQuQ5l9/1TkpOE0E5ls4KFqaV
bwaZE12BI6ZUzwM+E6GkPlYOKlB2v/xVWxZwSNiOqB7+ZFcSzE+GHb2+Ovc62pxXV0dBCasxdJzu
+zQmL9cNuzXMzNCxkgIq/sR5BrYAHfGlFgXevDefGCJETqi24WWia2pMuLZyEUUtV+sMha22O38/
EPxfzTxLaI55Z3rbn5am2eNh9osarSxyaDhcGgTYBYY0FWaHdm1CvnNZrCjmmOIARjhJJ/L3qV0C
ijOrCTP1zQrYyNr22BiG5blz8fAWIb/zG2u8agLiLR6XriN5tdh2smYAULBf4VgaBMf3VKDPsFH7
kEHHK+tZEf1WNqPESaPyo7oumbMHBQfDwN4pF5c2y+p/ZCVYxLkwb6aAyrVXZ9M6rwFYGqMMzNVl
xs8VPAQSmsAx/yGYYqVXAGV03jMf62WOlguz19bT2w3aRBGsUHV4pzhrvlumNyY6vMZJ+m+2BSlH
AbcsEIK7sCDIoWpYyF5kCk/4Yg3f6UOYTPrvom4IiKITEnGGLYWCFCID4OYUDRLusvWNoWplSTM8
jl1qPpt6onD9WFAEdp8Hougqprzrcp5gqA3nc2L6m+XjlhFQ/BLVUTuDwohkaSt5TEK0yvN+2tJ6
bWAHPf2w2lM33WZtQCuY9JJ6+dpHaUWRQeu2OXT9dSy8e/Czwhvm5MPa0jx4VMIaTaO0c1rQP0Gl
BqWGrH/9qa9otLqXUd92VqZ/3jKt0V4QzedKzi5Mka5FhI2fik8qd2CBVmWLjlFr5XMOM1a+zqN8
6einPoZK5VCvqY5BUiiTR1+mOOl/tTzJlU9zFt2Roadv/t6GTBMaQYDOSIJPeB9j0Z6W8BQ3Ptc8
7mIgJVLIFENOF+LrC/aOilYZC77y/O9laQHPuzA8Wk3VQDyzZ5Teg3R6C2H+fQu2s89cMDvRrqGj
DDFSIkRe4/ACJmRc4FxKGB7k65nEocxrEJPr1FUXn4vrDQjXtycCwaLb4AdN671C17a6QtgOtLBT
/vq4WD17t12Av89MRPMz4SMq2/ZoQ2lBbgP2tvcR+/0JA13aV9YTlWk264bTcsypWD+O88fIfR3u
Tay2Df4UjKG8YiAuQLFKnW8c0ApH8lngiP82/2MVOXQ13TmpHxUvmQXM575VeYYGmbfCcnKIJjrr
gfk/auDhu6A4RMj4TrEAZJzG5+RWl6GPaMuyjT+4iR5GIGp5CT6wleR/7UDrDYtPKYaLxYynUrNQ
+KthevEofTwKU7HrtJQXXt5SnYBuk8h2PNAOVVCVpDT0fsOSaMzYjneNyA11jTxUzZSnk8YmUJg/
YLBywykj0ctkxcmasDugY1reRFQ98/Cjo2t87TnMyGbDiTczBuK8OF7mQGhoS2Vkv0v7z8cUzFAG
F4TApjJnpEk4GS0HWS9nLEnMjYUvHnnbt32A3VLXHr8posL7wFCy9tn4Kve46YMtz2L0MZOOF/GH
X35Mj5f/LCqvJdd5OVs80BcVCr2Tpc1XaSj98g8J0ja4UkJhjxXnY6p8cvswELi+FxVShggNDIyD
IXIggOyjmidJbr1hulwB/9ZQ0WlrFpY91unt/PXEhs4Ohwtz1U6VqV4pud+Pm1edsRDsqmzcrjcs
o/TVUdvQYpZOj5ZD2vg3NYHl3tmiDVsPP4GfqrsAgjd6ngfxgS4fWnvTDpB+IkVDflzbeR8lHht+
s1KDSz8qCK1+tsxit5XVUwDps1hrw/aiUGBSXuAGDwk1aeDHNalkAwDFbwfBH32uF+EQyILGF3Mq
ztZqNVQTjl3/2U8WxGhm03KJkTlkCpkSGhpiQ6f91IYoF4XK0SWC5w0nwsGRpAZR64FD5nvHF4Tc
y9/33SMGPg79OJ1LoIFLNn/G5E2seE7RtcPKEGB9IpoQk07H7gPfrWtCc+/CQvwvpn9D1YH5IP/d
BdVNkraJ3Ifoha8TI71ZSyR1QGW5n8ztKQOJyqUyUBK1qUojnpwtkpKfi16Bug3F+X1Ou1/FvyZI
Gm5nBIpiN4V+VJb+eMA/24HDP6701QhPeXMg/mbAvE1DNs7rArv49AIMTctNY7mReo1By9QUEfxO
WQ/kNIFQxVop7F/mTcftkx++nLzM4euz9KbAZ+SynJ9QZR1KlVhFbWnbrDKsZOfiQbrWWwxin9OB
CvKCjB1Na/AFy+BfKqCMsm312Wfk5LY7DHPdOZ6GbvZHUegtvfCzjXhkmCHSPOtokyBZYR484jUg
IUy84QeV6lLZU41IsOiTBoSLfT+dZn/G4oJv+Zq5ORwAsgpRoHEuOmVjK/HXq98oD88z6Zl6SBzt
uySDLkM4/e8Bgmw8SEWLLuSesVMeom869wnOTa9L85/GkLToEa0ideNSH7q1HiQYeaqWSvSw7vwL
YrcHdAC7nKA36Vs7bwOavHmVEy0NqQnI7soMTnNsqn7B6Og0Oqt62X2S6U2j7edr2qLezTlU5cKD
LMDZ/pnTtVviRr2Z4pFcwa5ntd+6hyvUKu0DGiU5FOhJbyKfF+6EG5+tXG+LsHGKuYDSsASe9WaM
N0zDqifq3VkYjSMm5Im6bsEAyQoqrOp2JjExzvt2LZLfgDh1tS00ZhA3u5VlR+JOH+ts9ADKfCwE
JqLoYDUmPmjbV9w/lRhnpoZx6TdokRDNvhCY4cNY7iznn4yLHroML5u+fpaH8p+rv0HjHZHsO3l+
aD0xmpa/ZCZThqSmFYGwVk8zJnjXFlZslyOebkoG6dtPCUpyzdO0JKQD9W4xZbzV086eVkJkEEP1
eQ9nzDqgIXMrJOP1eGH++LkwrwbQt4k72pjcjiw11PN7SvfYXkHs5gJl+g9cNBNIWtpL4PZb3rzm
RdforlPjsORlw6SXAOhb8pFFQ+GVkBEw4FzuRsizg7AJme9ini66YAoTDtUgicHeb1OTnh3ITFTz
HmOIJJR6NfSV8XW+S5ybgcElngp0YJzflgYYj6NcP6Y/q1I8F5VLUC/I/Avrs7SU9EI3OpqYK6wm
saV4ZraEY/39dONoHZd83mJDkE+RvnnF3Izd6ypDi+cD7rX+KTFyFLrrCC/p1wop/r82uznyTEc8
gXWFHpCg9o9t9a8Gl/KKB8v78YdClrKdMXAflZgkrXWCdKLBtjxebPuvnEGYI2n5yhcL2Z5FKVsU
j70Lr87MLiofGFkgUl4IyhDs6pQBqIkbH1fdUGEp2tfnruVNblYEYrJCCXrj5gjcpARnEY1n2+3T
iwM0bafUSqjr0WI2WWGPKWYMAMXw0r7dy2rlhNFJPev1DulAwbFQJUCgSwYW3l2EaJvHcAaj5py3
1h8G+DLO2S3LnAZD6zNWaoOa63Vqmc5cPUL6JtAV/SgKKt4L1rcZUzOBWbO0xZVvCtEr8vg1+HOm
Bt8K534mAkUDFQlD6rUM2p37X/P0P2lciHFbHOyu6ffUrOzygloVglQkLfZdyiSJqCMu9zr/6weV
X59VLUsODJHQYJXaR1Nhzbo6dQQCj7a/6FiO2OOHYG5ljs17qsshbfU/I7S6hNpCaph+qoWPXBVF
M411MU1PZmRykNO0plXhFtthBdrEgsuuFYuLW4y5Eb0XuFS22rK7JZVMEP/2xHdKZlvRqMRfRIt6
AcvbVzVR6fXH4QTHNPyim/4qLe4X9Xd7uCCEdKg/4HHlIe6OSbmYJefciWsdeJA4ZdXxsRSVlIdi
dZCq18Pkqxm8GFX6O610cMa8m9QXi0GIRjuAcIAVvB9llLflEJrm1S6U2MmXdp8kWphj3dfvaiH2
LoFuvL2endr9oEf/2m5QPjfANptsmKoj2Ydxf2gB96OwZVeYnsg9xrA7uYEeGpEUuF834+XEWNPJ
zcwmyLYGTh9sTf+LlBS/MHxL6wxTaZtqBK34jyTU1v/VunTj/5I+03kcw00ckLYtHprTgdTeVH3g
aBK5bRSMTWyYDoeYuYP06NrIUaAsqO5y7nO3yfQP5nQmuVigfngrmj204aXsw12jmRcA9Cr/p1gj
7aiIFfa5CxaTgK7SAx747fklmV5zvRiOZE34ip8TfqyciziyJwn6BQwCCry4fHx4oZrWMD9dt+/f
XHyz/sKybUlMpoJRAaplCDUUyKQtegXshcFnnrLohcvFjolMzEGQRTSAqWW/FOobS/rgFxB9Jxhr
hH1ojnBUzK82KmT+MlIUO9uZmpnvKYYuR9oBdZWC3FO8kDVX77JKHP16MuNWAHKJE4flOJZC6HLy
BCVZT2WuV1q+8tWiqeItkN1yEkKKEZz+apf/zCszvCYe857l2P/P95UdjynGUTU8BE1n/qaxM+q7
uC1EspHVqLm7fl2i9626kX5u1viUeU2/uDunXSEjDAMTzixQaXKtYFcEnTankTJr1N3zCqcVQrw2
JCT2lUXxVwTeswJZ1gjVkrh7A/1IqObZwjmH3Ekf45wYKwD9I1Urkyr1dNtSPCLzBoUrm3Ys8ifL
4yC2v40Q9nchPuX0XZDeI/157rQlpO0hMM/OmGYHeAmBvEtmHr2AQLh7mq4Zqe9SNVYYa665FIAA
fdZH5re3P7ft+nEWuGV5bj14052PbEb4iUiVevbel13ykpAGlBqrJ37LIa1N1hmZK0rxMoYai+b+
JMCTTXG4ialV+ThO3YfhRO+xmDOiUA+YiTDV7kBnku4rqO1k47CzUMexrKA2PDD25yvGUDbZs/yc
ZBUL8C7fnzvZNt7wsJ9w+Di8vxIPhzWVlXdS3C35MbYuv3HAOJPU6Q+/5Bh/unbiA/kc++yv1hEk
vTjUoVWpZAJbXDoNVpNplqUsLLZqJY8zAu8XXcSlSJCiygC6uoif2cvPOwB0gqxvJKAQiTPJe7qB
QtUspQKtYRboXlkHzPgAabNmRB5uUjsHo0VyipobbveijHOCexQQnmEapxNRw88LAeYUhmvh8BY2
BTdO8TzG3nPNNr2ATen6233cjFnuQ+mwNz9/Svaqu2z4/2/OOoV0lH1z7W1XJOZ8kEPzO+Zoelgq
H9iciGpFIU5rJDSSPx/gRxz7bX/8+b5rIpymyQKKkQMlhqf0ftVrDrEOa969sLBRJAyyuVVIQ9Oe
O3FtIz7iSRY8Yl+Y14M4gb+EFKO306AA+VSPaECCnaoaTH3lZf4aVD6Z+YeuRwB2PII3R/DeBn5z
tk/QorroP41qN2y9GMUqYg3HhsqL1U7dodKjoN+rOw3syiMAYm6gH2XtisDebxe9xKDeKxjfAau8
1TEL8HfP513Tt+pBvkBryHELtKOvHMk0Ft1rL3PNXvOKPs0fJxvSgvZmyp2OhSjaUVi2utHEjBjL
8exBoL3II1phHYE00rTNUFV0mjIp4Af7KG7MdcqfNG7lFgeVHkWFnxRjmkkMLfdxFqXk3jetTi4M
MEa9AiADQoZXwHfz+XPVZCyjIJClPUIukfMka2iD8pFbqVLW75EWYD5NyTh0J3/wwcP53AKID3Ll
lsFIXgpqL44ELG5MxeU9ILg7QKnRGQqFknkXEw7G/ko1oo4l/lKL1ysalysUj6FhZ3SBiGAEx2A6
egbQNbMOc9i9bL7GJm4F9GXx3nshUjFkJp01xI5N3fvUE638yw13tbNckQELFku8GMTC72HpQ0xs
gFVH5pEqdjEp/ACvDCP0qgMzYBbiOCeXkG74zfxrpIPYPHQ7WwWXC4edckaJln6mrgsx1zoXfhgw
sWbpzZrISiHw9ceugtzK0LldqEsOULNKV0tAsh9JAG6F1HDC1hNa738hU+6/oPQHHi2UWHX/At8c
x8eHNlQVm1ASYmge9Yrtsq/wzxNOmFzO67C6kimPMuGeeUKipy0g8AduOcCTUQfz9ZyB/c/D+ADe
BE1gdYJgklesucrHXUn8lPwl1KRZNoj1wAYAMubwMH2x8NEyimSPR3042MatQP4tcBiEd5Ebi5qj
XqqRiUysDkswBmKDd756l0DsxE14gnCWU+Rz8KX8Xqt3LpNEcEmg9J5UuR7asuHSS2oVMmfKR2T2
x1742edlXtMK79ZPmFGIIa8baLppg2Lj1ojGSVIHQ2Gn7k3qyALTgSNt+i1kXTHt1H8PYAFWwxgP
nDYpjFdSqRUg12YhtS7EMM2HBTsaUk7guPqxyX7K/JsO7H6QfR/zE497H+YQ/l9cK0YjFR4d/+ml
75NDJF6RXbZp/ZaLPILyDeNhYm+EEGsNVDbGFGaqa8fIjSBgBlKWvIR+R2+0r3QdD2lPmTXpGQma
qNHlLp4vwSM/yx1lqHVObsEKbxYYu8/wECaFtoQpJ+uKI+JQdQpx5hK3q6FKgYD9Svu5hs7g7xrs
fW7iQr5lEPECmIGn3aJqheEQoCiPWJ0HINQra+ogDBXbS9ZkSlmTYXq24G+rHOOqTYYCUFYEl8XZ
n/iyvzpbhIRugS7AurHnAxC1A9bFoL5VHocjtXXXle6WU6bTdHb4hb6qcQwicmet5PvjY9FDbo2z
qe9wj5FMQSdYeYoaYOmUtOVj2z4are4AtfguuLLECP/RBwWeTyI78gSjydAXTx/P8P+Z9DqqDQeM
ERkz0doy6cZq7sbpofNgWq0sQRMhhLm6asajOVYBm1V/nSzkrZVyRcd34bBy9DNv+CTfz3iIzKYd
N+a5k2DvRM+IE/SQbitFPZpZU5k/wFAmAhdmDQSuRBjTGsDCW9NuQDCN/q0+qO1bP0CSfEOvtv/1
uAnggmlhADgxDZT3V9KpCPmnbgLN8PoAXyJ2GoxN3U/fntAg6FeAFpmrkyKVu2wyqlOnKn557+0J
TolDauctuMGQCu8AtkbWETve56bW6DuCPcQ+upbywcftvQLTxvGFf1BmEjhgxD9T5D5CV1moxZGP
05LP+sAq+4iqBxyvG6TRemxktL8OeWC20IBTkaLtm4RDBuPoZsSXgFUqlH5q0eRk93+1rDkZVAUJ
9F9bsXWyy0CBeWSZcwsOhPAPWRI2STXDv2MOMRIjCkVYfKEKrrdt2Tf5VCBLxI4xKvp6iBWuZjv4
IHo+Vse2+IOZlj0RCGQrhzXR/s6Ur70adwyuIeT8fE9YYYCKGnkJq01Gj4t/swbWctY2MTqBfO7k
wqBLuyJdAwgkiuvolZnyXCSc0SeAWpWd7kLo0fXIN9z9HjCi73agT+2IBeJniCB6stbOJs7XIaaa
W231daSvnYTqmiAvj2IM+WQx/4uNc0j2fPZEBf3Nu7FpN7R7TdSQ6y2Py/Yu18pV0QKrjOlvnMsq
5bZAOaF7EoNgIcr8NL9C4gv/iC60ZORtZYsiUaRYKS9/m04Q/1o5SL2plk595Olm1d87h7LSWVUV
Q3xVo76G0cKgRhMzmORdrKNPHc2R55uYip4lZTQetEcyViFBzT4EwvEeAzAKgp/32wiFcRNqJRNm
yMQl3mgamCDjB2Yu29BOvKtACjVWdiCfCJ2guQ0/zw3QnXUhYPmOxmdwwsrgf8kmUm+SQcv36kBC
N7ym/WykFpy96odJNQqiFy3OaFTDGzZQZX2Savi4plI+MF1EMDEPFL/edAIn4ziUjDmiszXQOVN7
SFSMhD+MSVx/nuepeVJ/Ip2DzJs+wtneFLH3mpOAbaWo5qNiTj1zifXGQeA5ZhSxHrpe5ZDFwiFu
YatovnZ19/gbaXNCQ9HBeuwC689tXZWLhDQx790C+/x+ZhfgeVi2A0dBAejVRm481gi/3i28vkv8
hJsvtyOztvNn1IgbPVAnW9XX/PRejpRPIGnCYBx5+fQITEkIRjtKNMIjs96dAp7rEun6YJpHfLtt
TFQK1vHt0qfXlVM0Oo2/QhTQRzHKv4HIy1Ruise6WngD/hGWryyiI/kXLi4NTQAnlemQ8gxGUi98
MEwDcxxjBGyzAQLG92QZChC23Jj3jhQwngycFKTrBOIosAweAs9YFzkcQ76+txgx52Q5Az1srp25
312Is+EIFzGD0l5e5izwtPCtVtG4weLyIpmKVjskAyibwGuuZjrIhFfst4J0P0GcaNm9C/KiXkHn
KOurkS6xU5y7GZyMTpV7lm5cs+O1d0CmHZM3LLGRXChy/9JT1WlRld7otgbvk/xep4cugeL2W4hg
qh4VJuUXYcE9WJS6Eez8YxceU4uO8+5YE2QS5LM9ZlccxYXxmQRT5JzPKHg/WXLMLjIqVyV4mF9/
juMRFPLUAGl7NGpJJ/APxZOEMX8XxTPehIlL630lOckaj6ErV26/EX/HAUlDs+FatTEeTjGaJKMw
w9SNenh8uQEZR9AyJSLgh1I5SW5UdHGIxImTSwj3vPBPpPDCVkRa3Y0PpFIybVUv0bdBXsNvd8YV
IpPPoRmn1APWt9k0qEeEUuokeJLNYbQX9IN6cot6KmrO4H69/J5+XwZE6048gDLtiIBzXe5HaeDi
ok9P8UuAZT5IMfyXsyGoyhUTkxQLrB717JW52NHqkVhN7Celav5n/l2YSiRBtuFtWlqVzPvHO1bY
BmOT4is0I2SChuDQ6dt9wFL59JFsrnmGBBXCSDyWiKXtHJv0WN4clT+9gLf8tMuSq1aJEml/LYr6
RaQiAddE0EFHd9G2SMqOQ9knpxN2bvGlvkJr1BsUPCKkpexF8+Mqkawcdk5t/jnzKKyLAi9Y2d3J
1H8cOOkoLGkZKbIqiygBdi+tKrXCwrh0sDoyRdBWIZkxlSycGBZpvEdvfiJDpe7uSb/pAa4+Jo5Z
XVbDhR+ZElNEyOmak49ZJX7MtFJTOeeeGcITWoFbVs2t57FyH54oMds9L/PBm95VlA6VZhHKrjKo
zITpK9DLX1h9jsgCwu3dVMXTHuzEu5DP1bHEmnz7qxc2/jue92jZYURc6r6K8Lfz4BVO3gln1JhF
3uYJnEb2rUSLZ0Ye4ncesQO3RyHlO0kiw+yyGfiYacvSJDxEZTigi4Lx3yRD1fTllkzOgcaFg6XW
0ugz+jiyzIzRNj6OzMG9t15wSIpDAj/+XtJy5ZK8rBrEBbmoFmf/grAlkxY1hiTAdGu0EPDhDHya
HqVaZQBc8FKcfX3jbIj1rOBywdyTmjt5durvLcEkH0jiDibHdilgHyHErGsNjdTXvzzQu6Bb+PPc
skv2DHuTqLpi83zelIAWsKODAYYkhPeJXdsyn3d7iRu/kaF8K0URu+7gheO8gyZKmmSsfHQ654Zi
RY/DINCGQHoHlprVT0ODkNzgDKUqCLLz5qvz8cv8UDsJ+H5/2eyFXKOiWrs+qJ0umeDkf650UA8Q
E0RO6k1H1IhbEmlxUkaD/ORDraHq5tkzduwz+4PBpwXAP3FB7Amf3SxKbtBckKWNbRLjn4Y/NCJZ
8KwyR16aP2zV63tu6jK4HWVGAnkZ4c2Qh7/FVMA3QVLy9eYF6dozqlXEGipjNViyw4sN3HDaqC/p
MamideO4pk8cNdMyZWbTEq0hScFGQfswBQ6AucwPOJt27HrmPi9F/qp20jRM1BxpotqjYDTicaIU
lZIsPg78vPDGx69RX6svIum0yWul69ESl+t3RKH2FzW42gphnkry/ERn+EnTPbOsqnpts4AGrz3x
R7m3zO3vC35DGx9nGxb8uDAoZTl3jgK4tCQsL4kApBYJn3ewizz3F0Gl7u5EelwtTIU9Qqa0LCkD
a0kkfDNb3p2zNZZBG94R+y9ZNcYlF9lfCUnmLkOsSVU4bG4Z5Bi84derdwD6LzN5S6dEi/Q+IbDE
L3Mc4n1ZxRc+GWLVzVvY9pgHpu4ZFhAWRK3zA5GfIUd88pU0VjoNKVIbSH8KrweO5fJ+ccTtjSSZ
f3s/fVWww1DawN6Jbcd1HXtZ0OK2IbBQI+j9Q2J7GboEZlHuRiYia+zXl1R8kr6BgJTpJ1uWsPiS
Y3cjCe2eNiSZhB+CpAwETVLHEClTHQX4hgKWcaglCguBPfp5BxhVnNSquCJydKUWAQoxwFk55dFl
eioOIBRKpcLfuDi+SHWtsYUFPj+gpnTXEwSjtOI9Rg3IN8Qx5oSB1jdLx/S0mUF7aoyOMIZhxYhR
wxud4UZR6pU3Nyo+wpkL3vjEBSjCkeA9U+VQAO3/g0Uun+c+l4OjJfFr3kNvt9RpRTYqFTM5qOe8
wXrPUebJXKH6eiYLXEEd/hiY5yJ5mwYv4u/Qzf2H3ZTLipNhMaLevQBMKjDDXGxd6YrpwXbHscpC
kAnOWhgxh66V5JbiXkcp6MsSd3hV9Jd37TgcG988uT9sp6Wk35N9JMo+qPYh1BB09eqWmNERzbad
ZwdCzjyxVyK/5qZSvvqyg921ZzNTT3zS/UyGdU8tkhSO8YW/SZx3mkJof+HFUJTUU/9Nsn3Ap2LR
kE1Ec5BOxnlyiQUIAYDvb443a0u+EDiDVz0+GQHHsTII9QdiHOkH9NqSgUVVq6jsMS9tpDLct91F
2WnXO2xd4LoVxVcu37VM1vEm/dcMfuTdWJc/byhj1nEG3MOgyklfAg1cskE4D3ClqSU5LGojOTtu
evRZ3wy4wD2yC5YJ8dp2t3JmPHY7JOh4qO6ovlsnxaDYwOdvirWDBJQfLaHd6H1QkwCiTYLM0jQh
vsWrqigIyVQLv9f8ISTIz8PQ5XrFRE6zT8D+YlQAv+Pp+HUbsWnfx9cWuC2JRI/s/UDsNymdWTtP
RFy8xuZB4KqgiDIaUdNp74TKAO+pc/0YcWJloWy4yYWqNhrPm/1PLU5iooMaR46/O5yYgoCfjx4V
ds5+audQ+efn7VegbmNrwV7itahTY+25rj8vVSBVGQXL/YLnH+umwPA2kLhp0knlm/PRlCMnVcxb
7+p7DjZqdVAfU1CKjnffMSYzlWJh2Svb7ALQznBAUWaTbNmqlxnujZdKOxhL/UbuDjthysN29OXA
dTJLqBZq+HH76b/Mb+Uqsr23DlvGOxVTWhHtV8VzTjlDf6M1+N84AUHuAhX+tJkl1Du8M04T6VI8
dyVVC67OFgl0TLIsqS308bGqK+5Vs1xdRLXw+8idrK6R0q5OzizpQtG8bEbOKlSm9y2qB81Ck+yp
QUmNhTTMOEwDfS6U3cwXyYT3MBpIxQj/0LqfDF1bve2lsn2705wtMb39fVhuRbU8e3Ign5FWVtMW
c3SyNKRd7m5gUVzIxzItwSBYjTdPyjGt63LCn6DiPwEnG6ManZAdnjp6KHAA3BNa5x/dbXBQ+Qa4
9qXoMFq81+LzHHdvRmpvmBPhWxi2iZJdVEGUcYHHH6nrKqo+BBrk3FfH4ZjPON82QdL/Uzta5UqX
SW8gZV+xcf2SL9JHbE+dPga5AV6d1VZKnvzSIbAbE4iYoCPeW6u653labJGK8kMb/JyjlwPX1JzZ
uG0uAT7Pv97DN09Y5c+TLGisogebBI8WeK9IQ2efYu+XdTuvrKoYcxcb4Tl1HdzG+UPVJC7K/7un
zFQTyNEkZWbsNY35LqZ7+zg0nhpSkj0y6t23CZDfZCrmrUI3+sFm+qYKoSPz4bKnKLC9/V0+1UCj
Wl+TT/iUxV0uKrYNZI7FKqHCNBnnSiAHsbFbM3Pn4wSDLF3Aon7d5f/BqOs88JoQZedP+91L7BeD
LCtRTMgH7JuYFy8XygTxnlvu9cyJBhKWBhkhLsg88ui+NHrF2krFt7UO/ysk54DxEddCU7z4yPLY
9hMVj6ZMmM9pP8IG6yzcLAPiAet5+EEgXW7gFDnbN4SGlyBMMNGXmBuU8a7mtmNXzf83UIvbm7nO
+32UNp97Y7OiOHJCfTlonl6vH7Kk3RfRYDzx1yF3F6nSsqXumPP+TDejKSXDYUVHJvvKntRbP/E9
l8g8xGVPrg2OmtP2+T3pMVawwINwwtwBp9nt7XW0sCmUKWpyJZG/u6Jb5T6hnzqN/KYsYbdC7Fsx
0UrVPvAX5RNbfBsTn4dh1E/ZXaShlBCTpUesHDdHzbLna0V6OUslAW5BQyHn4bef8uFT72GWUOkV
VcC43bwm8Qptm7L2hZlYXwLRa+6FBXuQmJ89ASLhaEyZNEiNeQ3djAIf7wBOu9PjecnJ/CddGrhT
LRd3qft3yi9Z/1zGwGIybimR/oHfZGhDL6eStCSvxjXBfVGQE6Iw/AgEH9kBBT/iVGUrWHtVQF2S
FtuUobm6EsuhfD5eKVL5/xdY6tFn3FrsuBqbFuv8EgvKWUSd4POLFO89uCY6zQEgVVLpBsxlNpWV
KYb7KsEU+hr00OGZNcaiqFsBqbu7BwdlMP/CWy0pTaF9FiS8fTg+FaDW26Ek7RHriaD5xTUgTQB9
iGZlzX7guJA85vx6dNnFp1sWH1/vrmJE9JBNUk7GHj2K49gjLYHFO1reJHEPP7kM0T0SArMR1DZm
8yUSFrrgIq5xGou434nScerWPCxAQamG0Epdis9Agt8cABX82jtDHeFaCqPM02HvZwDDj35qEZ8j
Wsfgv6X/rvdl54PrIHtWUyrstHuHVmNdkow8owoLP+tcPKeiIfLkslPfbrqSVYTDMQGbBaegUSpT
tA6KZYiMwxzmtU3wRkl7iX71owhD8VUvrGRVlXEg7wLn/ka6Pc0TEW/lwTXKPDnyl5mVba3nA5qK
sR20mcuqe7Y1NRB7wCBkdZwL36mM9E8VjRBTb6HpURxje5kTBfF+GZDXOVYYPBdtTwJsA/jJn8rE
eKtupmiIR3MB+tsLgxDS6U55M0YvmG9OUrAIlewN4k+NIzKdG0jrw7ruMoOCe0OiWwklkr4Z99BR
UfM1yAxF9z/AgkT+pWJOwTd3SzgbYE6bMngeOOJLk3KhOXXngEFoLjWZbz8Mdqv383vaRikluojw
+j3e6M4WHdBWliMUS1HaHfoJWoEDljfD/LPEtQ7j8JFw1rSbdY4dEiIXPyQPslgIDqw8anFckied
+7GvG0asasc3HDjIcT3CUm7tBtk0AhPNUZH0GETdkliKGjYSChbkGMwR3m5e357OeraY9R55gHQC
SndS9qVvWsZLr0bupIBOMgRBwlSIS/ZPHP4ol785hFkGN52OS/F0KdF9O1I5FfZgQL79UkXCyo64
cbL/E22Yw7eZK9VGCvvUmvUd/pj/AoGN3nLFpEBkcERXYsnh7AXwZj+Sem++QLWP2tiZk4G4XK5w
RZusj0dOgNqISLawrMoLCVdxoExj/6ktGz2007+ZcJr61syvjDk4K3dxrO5W0LbT5L8Ng8r/QJ+V
/BSZ6jHVzjUOP6CFnCI3ObZn/jmKEnp1hCsjwv8fSdgZ0DOZMCLg0kJLE2z+l84o01/L/siz2fyI
O2PZXP+jpvRe5aApQOKX/ea3fP6YMsKrD8yHOXSKH4J2Umx1l1sS4l2K4oUnWKmEwGDbacAebNYi
weNKUhcxmadNqxFaf7LlNAEy8gEcCxlygakR8BQ03aRDkv7I2z+X+G5QaVdRwtV1kEiCECFMcPtp
bu2SXNI8iav+v+7eVHPNlg+7Rdq77ORJ44m0NfVqANypsn26OJoYt6+At0hk8gGE9jlw37tp/RJz
qV69Lormf7R23+I1E3K562ZL9LDPkzXR2xYhQW9DPnVSSTp1dmRsBmQumxQ7n5Pc+SJM2MZPl6Ag
308/USkf5aQ2rBf/t5GredBnYJPTLTlmY1u8r246bosBVmwCHK18EMdgrUXCL//pPio4ktqwz3/G
OiqtRZ+OoQvbThKwv2L10durkrCFhtySs+q3StowkmeAoWJ1xqZ4PFJh98nBYVf0L9tnGgwZW/Y3
0HvJ2xWxtpCARPK+1fdlqXp/Fk25poG7c0oDTHoMaf7t6Gy51LHn3Zq17IxAxORX67r+lpj8+gva
yT9/4FAzgPUPcbP46yhLs7wTWqTXPG4jTeKuhcA3BGB/7bEP0jPy1FXzxAs7iL/j/Xvuz4fuvCV8
CgnMP5dOC0Bn8SLXMjVfpAz+Rdu+qjD0wInhRIm/ZQ0SFBSOQovQBOxQmFtnFnU81ZoMkyd65Dtq
Z8stfFnOjgevOpIekJsBB1ZKjrRhS71DJxoGvIgsTwVeYPurQgZIrODvm4tqCG5A41yoqGXCzLY/
Hm2VmKUWTvLbJBlI6rEbE5kWVsHbynAHCmt1wfbjiFJQprF9aCOj816XtnLE2mqagUxMbGczeH6s
lIer0AIDoOWd/BqyUDh3DVkDLZUc5r5EEFOx0CsMsxwRKqCWxYDOvfMD1jRL+Ra+bFMEY/W+7L0x
kJPocHLHQziJRk27y+5CQohUvtclsoumIDXXHyo6nxzXWI64UA0/fWhNtvjurV4bAAATAIp7dMKj
wASCBQ8y7+IY4UeIqgg9IbY3dLZR55wkkcvAklHUYBY2s+xyQ49qJ7spGDuUFyQssOmnT+VxWkhd
auxWkXeXMx5ORPENhstMxmy9WIZbpEVd9die9msi5BRPMKTzezJLvcdQACNrIl6Ay2aR8qRnABwr
URjSD5DdOVEB35UVuar4CVs8RKWwEVaYdkv9MbpgZNX9e5omtGLq4dBwXpXZz9pJ4EweZ8q3++Ui
JRPXcgNGrnfqLZ4eD8h48gokvFzfpYaQIqfm3z6giplrdi0Nt/8hf0p8XkTLn6WYmHk8YUZmxowE
fr97h3vjCMJYFEWPoyOOnRke4yug9Txt3CVlN1KkgCnexT5DFwm6Srunx1tViJr+JqqixJ7m9I2k
7RZNmu6FkCSZmCLc2RkaAcS/hQgSEwn/OVm9+Hh9f6j0wyXH0T5yYdG7HuhA3HvMx7z2I5/FE0Lb
foj2vJpksjBLQ5iEIPBCXG+vDICHRFoTapKQmeY/ESdH1BzwbIN9IIM2LF114do0OQX2g+JLax47
cpmF5ef9nPjKGaWqyFotEBIXWd2csEQ619CoFc0DwITDyiCJjCIyeH9qU9VQFJjeoKmRZj5mqMs8
8FbKliQ8SxJFH3JhlWnEEfaVH+aNuqQDiVobMvmOdogr0adhT83oJDp45XHcsJsH3sQyM4G4alq8
sgmWJZp55aMn2T8kY5QXcSyRW2quZtcvaCfCbnbPa1DMKgHYmX9pd36ljtH4Wj5pgymh/AoHH0Jg
WkY1F8y4Ksn5kZ8YQ8NGEEPaGSRo0K/8rccc1xdF4T1FkgBSnQupYlLP6hHJmMCA7zhw5h80i35Z
alg4gqfb5+qD/LXPHSahv64ZxdnlRdr3uVz1NK0LuXkrgMOrHGvKR0uQLcP/vW+TFtX+w+iKgShV
CGqksUk/57edt66IrUmFHqLByAS0Ro4DOP4yhxW3whRaqxaCL5Y0gmJGNMMp1HkWJpbSvuiyAJTT
FX8wbB78O0G08rwCJbCiJFKMsQs3mTLfejNnSOSF/0I6P+qGmcpN18wyUIjXjs4xoEOIaJ/zoJ/U
j1KC8URawoIek0RvAUItlhklBUJ7wZAmyR0wKDVclLqHt5yLjBwAPiM02RSFrXZG2cpIuE4FJOB7
SqYgT5O/JXp6knr6uWKI5853CgL+4VVr2+qRFvsfg/5y2blbUmQxlXTzN2FjgtQWINrUlxVoSmcV
KkSd6QgQ5yFZctTqrnsrwJeyW6K01n5o/aSyW9QNlKY3ItHaGz0auWJtgpR18BCkMMbbd4Adzqge
RCzdQ9KTry9cQsLf28sMNS19C5HToZTGjh830PKCXeSp0RPTorzZBR4DZxmT5UHt38Dehv4mBqqD
0CNc7flBmEFAo66GvD0But67aC1C8+vhehiLfeTl3Rd3o7nV4iFvP0go8W/etF13/8FTnKVNlOGx
WHsxKaQLUTkXYXW6SB5X/Ou8wqiWtWlHc5lsdZaPnVE4O2MqMuTWPNkn2kNSJpdO6Xii9dPQKYqZ
17x2xX8aLKoLFWk3I0/WoWykb+aUCBHi1ENdgu2v0NTK1g+8mWrPbixv7oRumoPvQckRkE4wyMRJ
QuQlJaOaf7NGA0eHe9WFAzEVEkXz5PsGwKVIoKLhbW4NzcMTsYJ79ZWABBCzbsVJDNOVSlQNkmDA
PTqileNkHMxxaLweL6NitjM9/PP7eLMr9L3ws6fQrjDpiFKFBJuCvMp61EsolPPY/wjLGOAMCLOc
UHble0/81Rt9+EokEy4LfI8JgWl7IKzofgaoF9Tkf5UMqs7BdEt1Exz/FnP7x+DWwu4xgHbPmuLP
cb5MIzQu/yjXB9P9OaUbBKpOUBbFSbZ3Jrp/yFY4/T5ayTcK1acNDzbJ6VBp7vyrTZR1Ve4mxpEJ
gNJgW7UKVeXDaigE6ss89wK13zu+u2wRQnC2AirB11V3aeA0F6eufvLrwX9VGNuHDOp/5aR+sloY
zD9Tcm0FKBxWzJYW4i5IuCQWR5sakovfA0kCM7AVwpCULNkCPZYqXcv18Rv90f1Cjd9Ogz+pMSHb
Sc2o7GirmL9Cjrl95n6gx1kCpNnBKcAIlhCw1OXm6Z7pRTTLEWvPhz8vo3EdeMBOA8iparoisp9e
L8vcIbuDW5iR1Upnc4ixMLb2u0GTR6dmfmCYty32fGOaxEsvcorSDSxLSURTxzivqeRNQpShcRDN
SeHzGiWE2xnRyqzuoXdgiWyeZjExVRNgSsZBkYg8osQdWE9eDT29tl+p1HHJtoxKVHACtfNck9RA
eWeMBjw/qzXOXN0f+niDItzhnEHkEXMeE+gEDaOPF87hjhv0JTdDqsLDX2ki4dsSdQK2m7YrrgPU
OeRUDCrXKJvG6a8cFuJK6+rsft3uBE9sdhe1Jg50WnxOZ2cK3ygqM5XXr441s9+nepwcgYbYBAW4
ubTu5HiwEb0qYoxjQ+G3NxNzv2ksSD1M6oN/cnpoUf6cwbDECzZXViRn3FG0FHpDsQsIM5iiGjHk
X2ZjjY1QOJcYrIobdGPTNBZK1GVhkUIjLeRucd3dhwc7Iae0t20vbt8/ViXnShnHJ1fNdrGbJNV9
I9Y89iqD2A+3tDVO5cAeuCrKnNi8bvqa9xVgkoN3AI2gixChsbCfanIlJkDJlCWz1t+GmGMCHK1X
fHw5D0CqR2CByOYZ/xQnFwi7+DiMdcSar6x8jrqjCqV8S/n6M5PZJZ7+rFlnBpmOjb11oAJfG8ue
Q/leJK6XX7pcnNXyA+aHieMJq0KtrL/Id2pDBDs97ar4sEET5KlVRAtbvqiPgMl6Qmas2JpfkeIU
MDNAGZhv2BsWCHXWImPasXZrhVyStuGegEJVJbTRI5PkAedkbyIqAMcZ0lfuZ+VM+xOHEeGSisdV
7BqvgkCHUlMb6Kb7lG1tKbETlC/w17g4S9V1J1ju137Ss4Rkjr6a+toS1LbRPDhgWKC3ZVKJzBnh
rPXcTAdarGTRu+A5L+JX4wTbmfbm9j0E0blhSr5Z3kJNAep2zs7S49KFPrKwq/XOLbmF8F11+UJG
f9XAetDIDSEMDcX+DqZVHKFnfnW1H2+xF3qq3nc8aac+3zecjlP0oUAOW22qo48WDLVKYWDt4cPO
UL1xLzESYBTulc2wDZRQNcMaHrIFcBMno2HKoaZE26ATj+qUdy3iv7iYicwJuufSJ4d2dQbBdWnz
QMd/gONz08UMWnSrbISkPEX1mnIFRamnLM2sYqY3Tzj53bgDsOI05OM6s1jkXKpBG+xUb0vWES1W
iGUww7EgKRP+bPmYBtJSbMk/TdJxNBh9NOZtB0sI8oZkk/xAmQhObpJcMZuJCSXwvemeYMOowjGq
venNVw/18FgMggyXNgKZv462BIiuzXMvXm1ObI3N1JTVnbH31i7GYLAuDAGxGVJPCXqiehIpLTUO
R3VTMKnYEQ9ln7NRoNrLMQF4wz6PVt9oitqMRULMvYtteDMkq5MmdmS5DhuxKSwesWwS4dLtBpgQ
+3YKrW6Rq7I1eX3qEh7BXLTV14eEVOz1ceVjgFHRGDiIT4BXDy+oJDJ8T6k2jvkpjhoGuOSpX2RT
ZD1SwsIZK1fks2lEp9cGO5TNKRkcIac09wadOSFBJCwIe9zQlArSHfbyEvPN82eFW5WqswfaZEsU
ynV6gTNPy1yw6zEMiTh6Ljh9fAPm+aPLcNPq5ccVBImJxcBp2HL4eOdEbKaLovJgYW2o9Y4kskcx
D7N0EdyOlrX6dvEQGIfZDaQr2vZiTFjEksjINS7zeawTs4XgIfl2kUi8vi1FNLKh+yncZLmnVN79
bvT3G0DTIqLe9pHb3GhPCPccKpk0t1ILzZ4lMQfF7JVmOnnpDozRe8St+7YjMcMoz6ID+2AhcOwH
z7A27pv3kOWAlViMz0Z+cbVQ+T4WJGaR5fGFj9vx6Jr3qBRCM3J7K53axkSu5F0ZKsFYWPmwAo59
GH/1ILzsV5osMkUChcejcmeUv3O6qXZN9OtZr60XtojEX7iphIhIcvxpSAY1EfCUh9X191886rfH
hY5ngFlxpQeKMMz9HGdJOXGGZ2aGZ5kf9X67puuLhuYcNIy5S9iTJBbFeqHCu0fwE2FGpmcY0eLF
4jJ0QW6ilIcJNq8nvmDfgBR61Ipb399ULRTfbNnVcQ0cl8OGwmPx1x4irGXsj+0WvB6iZPJgJ3xe
TK0vr6bVKIJXKWESrIncHweKQ9xGddRvJsjo+F+EAf8UPtSdxihwamzZBKsMfcohVe+9jhDXnFpP
atYaeTl2PHWXzYzluPFSVSl8UYTHEdBKF2ALZDo5M4m+zf7eGHqv8Wbll2ZL1AZmOK4MlmtM0h5w
S8zkUMLNApArOPs+Wwo1sge6QS8y9g8fmhDLkFUb5dVd64vIb5TLWhFbwnoe8skVL6bDJ7lw+uVg
Tv5nxwNtoBIP5ZFizvtWpmtmN/GQ8M+H3+hVoNFJUm6aQfn4pgPZT46jbk/Ufl1s1T8m9GmSGBS0
c+77nQSYUPH7tQybuE/AcvISJld3svbXvBH75baMxADUWBXDz/CDQ6r8oJfpUJ9oHNTplp8sP/v4
JUZHvLa3e/PXINeopwAlpWtgsARCpHhEdnj5+QLk7rHYrzd04u5y7l+OXLV3Zc8JCbwO7rQ2yvvr
ZP2Tc+Y71BTS1u0ht5yv+msAodtC9aSFIVQXwxZuidznZ5udaGB2UqfqetFGRKjo75fzcD4M+RF4
PAeCNq6CSsYsyoYxsK/DGE4eKD3CUyURTZo4pVi83Q5SYWUi2ihi7VpEvEMoqTfT+vR+lCFuh4Y/
YP5VPyZYlc/oYQpZR8GtaxLyTYlDTlIsdp7RX/o8bB8UJk1Qxoxa+KpGsLJAoCeM1HGAX6ru6Hwh
J3BJa0O7X713mZ31GrMj7WWNsuvs4y7bT666Zzg3gwl06rjntvd7r/v4IL7UgRkr7p4kXG0Na4xv
iLCkRkOd7+Q0TR/gQUmFCKWfir7sJRGudBx6hcVAIj9PEjXD8Rox6BrS4hezxAqp1BApGkV/FCVf
fD/d90oxlrjhRM8A1zRHHyqPxoC2rLJaFwfbA4K/f2a9BxrSHp9pLoMA4fUtVsWMdRdqJ4Nnu7cJ
J/dbGdD9AT+dtx9adJzydMu6ZwB23v6WcMCJvu0w1k6nwBV5GxYY8Booh/Tv8zPFE4L5SkuCix0p
V+JxB+OEmKp3kClm5kQ8Pbg/fKF3wPY+595Bga1NHEt4EL1zc1lR4aIz8e4c+Jl0WTSzS0E/7bW4
tQJihdBcvo5APU2leZP7QI8mPekfw6qBL2wqZBRusXzbTTmrCdZS/N8cp6Q95fiQ5Kg9y79BV+wV
Pu7i/ohdlsiY7QDn+sJXDNTnjB4qAcLjDqeiU2HqBSVrKsVP/g943Iz7UsJ6BZMYkk6QbwVw8QGO
UZAUl+ljlT4F1uW5p5uiR+q5mXFq71KcbFFtxvU1xHYrtsaVh0nf7ogxs6mNpCYdML1CYP0XCwSt
flaqL0/uPASgq+WkNm03qcpxxmqHW5+tmW72JBw50UBS4YKO0hTbcv1R3WS6d5A0VU/mPsBd/j1x
ZgF4ZsSUDmevQpfJyjcSPAEKrb95OzyZfL1dyUiKcZGp+uUHMtj4QRtlDzbA/rgGPQmi5n3kax37
budU49T9LeV/dBVz7fIyV/yo1x+JL61gfTVNu8xu8krvkS2yy+UyaWcurfd5DEk7F5AnkP0d6pik
b5vv59iZJwVGviSISyxW2SauiEDZMizQKddyVjMNCt++I83lsGZWq++htIJ7YMMXTESijIX5207K
3pHBFp9I6yOr8fX3OuxXArrGQcYxUoObNDl51567iYyb7rpXrNWalnFMlYNZlXirN7101RHhO08y
XHldJTsiFgUSy+PNaboqYZflwFS+KlJ8C4NjBMuJvCYWNJTOeueK2aB1avmE1II3/rJZBYg+8QoA
5vKN0NXgsxt9J23VwBvjE0g+/djHdJqmoAsRTdNVojCppmHQtzqoegLISVtnAa+WeY1++T/k5eVr
/kzMF54XoP5ceFj3LD7EDFuE4L3vzCLAxIWbEKuDDlYotGxWZIU5MCRURK5SW0DMFbzAv9LGdTz6
rSHrrQIPeVJlmU6fQe/yIchNSkw1ALhh6c++O40BbskQoUdnELh5ryuv8TKsCFKaa6X16QP6pdWO
vx3lIUwGu6Hgy7vnH2Wlg7nDe2Lu8D07W3bWu7XXAxekNfBV1dT9hiIepF2CWltenN1lPA/NXxg1
fDUNwmS2nLtNyW1ocxqrJsbe272f8QlYiJ8XhSW2z9shauQLIpXUyHShoYB6qiBsvlhIdXRaqeq+
ZxULRi87dNpYSPyWo5bx7sOywHMbBU7nqjJSBI8u8hvleqtkXh1zSarGvrEBx1yDsrgGJdpZeX0v
mkC+JpounHmOkaZ1NWGj+oeXbICl22CHxYXo6JQ97NqqXIpNkfuomUCVr3oT+864uOBz3NNc84Hq
hoEBg6TffL5soz3hg/XH7oO9nF0KTbzGrZoazzmmB+530Ho/FN9SB/3FOvHlTaF2I4954qKdR5VH
6epNcmA8UeOo/EWz6jsfggOIOvRd94qBTgpufoyGg3xElbTLbZXHzleOrdj5kA5rQUZUDYj0EtH1
XX5WiqOrbBTtizTsxj87h05ZkQRWdZuZeQYSwDGxL2IItgwO4PA7j+JGDezIn9jfAe1s7Rtcvmlk
xHOvWl9P5Zi/SCOtfML207oSz/i7krr2+B+279wMN/pdf/A42jx/p98PfVvkgIe8yJp375WlmqWo
VbABnHbxgqG2uL0irm63nPT4+hl2mUW+slkHLjyJrygIFZmkRKIbywOh4qwYVO68QplxjygVE7lS
mwoXjW4qT+6VWfWmhFqWPy1AodlNAjzSM/tPS7vKbxRu0GQFT3bmA3EeO0MWJWYWd6qrOxOpU6Tl
Y0i8N7dxqB8ww4NZspeeltHfOBfVg3OPMd1yLDSi64GCysEjjP6erQyaf87RiCnXOeDPRr1u91Ot
D1d2Ll4Nv9+DKD3HR/AMGdIPZpu7zSwm6XPbzO3rGbL4rWW9atqVmkrtu9GgZUG6s+CpbBPv/lpE
C8d42Fu9hRi3p2v8DYCdc1OcOwJdrfvcnZH1v3VNzvrF372ZPKeFbZjd4gNQbJO1RLuRg2v4QvZc
GOb/wDKNt47oSxrVTtn3iwMTbvfuLQd30IitquaBvX2rR5b2fP0Kx8EcteSQMvaLhtcoQuK40kZA
Y4GG54Vr+mGdJAW9c9dN3mbEqhigX/92Qq35nbTeyAN5NsOlZWRMWhDcJzFYRYd/Aoth2Td1CXXE
D8gJjK36A+fu88z+Nud4X6Ipk7mOewguCazXwkknqjKVpt/on3P6InGpsMEO0IWbN8ehWlsdhfVN
XuEYXgQXUNiCupQ+Wo+NS9AFst3X0lJqdHmQc0IfzN1pqAI6YE38o4f0ix223i7Cds94zIBsut9s
eFPkIweaF0j8+bRd10Em/Yjy6RO5T440Bep8/Y1y17ye9s6rWsVQcZtLwXBBwtRKuETQBzs/Q7SB
UqUzX3R4l6bqrZtOAsBAfmacfxAhurF4e1s/YXe1RbpK5NkFARiaqxxqrPDMF5t9z/pvZZTP2MPK
ndGM45mr61zof3v3me2fIfHPFttiX+AvAdk4cLIY1KqfUKeB9SIbOsuWH+r0HUcOlcXFAF6Nmdoe
Og8o/EAnPTsEcL4a0E4WTh4fzX32xMW+TAmpbePQY9P7P3ddb4iQqFeyTh3B3kkL4x3jWRxvAeXD
g6Z1oFThFj4TgBbcf9gkvJQITZ0phLAjtTlYOuRMbEP8nGT1iiSFgHBoIkp6zmz4Tmx5OqQ8nH+R
YlNsVFCVhR9N8kCFJvKhWw/fShoQ7hH4wrtAUkBZv7NDIEkaq6br2J/6Rqm/Uv0zmQVByIyC69Oy
CnW52VNXP6JX8g//kOpjRS4xR0FnSFjGSnGyRbgTt6p9/QN5zHFYrbbPmflMPmvgbGuD0LQcF/uJ
TbpMGxZEE5PWUZBIWY1WKRpGq8+KS1UMhg1Ih9QZkqV5WwyECOGuU5P03/97K4eOT7SV8+AbZIq4
n4kr4iGHy8qAHYYtvpmcm+c3rnL6W7JqbRrm7UqB4hzICnTsvx8aaas6WFzl1XG6k1hfDIvdZJvd
lfC2brfvf1gPSIoNLI8M4PrM681TXNGUOaGSEB3A5vQhodluxODMU/D9+NU7DHA0HSrJmYF5EdSB
dP3ujufvVYQBAG4u6nx6S8aQRu1+sYtEWs81dOu/kxkDm11SVMiku5xWivn6/yWZHKgMk/8QtmM2
onJ+OaYv/OylXoScgHM3RMQ9MrWXCkmp2FRjNWquE1FS6jS8vkz6WHH+OAoUoiPK8qr57cBG4IoO
qRCfX9z67SlLwXv5M2Vcvlcr5UuCKuNbOqxOLezjYL6SjBGZimz3CG/BrYlkpGJiRryggT5dck+j
sXXU9eVTXJijMZt5w05V70MWcZgiECMORYiG1/BNL598Fu2KRL7EtTn2DcaKTH8dNTUFL2ULCiB3
M6hA190u+B0qS+inmyCmAYnkqI83fHMC0Fmm7ueov0PNiIsiDMwCqJWhXxnZt/Axmjc0PphsCBiU
0XMvN1lVgWTInxKTydTK8Yzm8Ob0y0eqxDen/9vdyeQ8mi2Rbi5zqybtInZiRBakWTHmnoRHL0Kc
VmLxgS63WCCrh4ZZJABOQrRKFf+f3ZL/Bt+OeJk++E2/zJt15YrkhhB5LOzti/vFrWsfTzSvYkF4
p4Dk4EBGBCa+N1/fTZYXSiiQfMQqFv2T6RVFyvQ3ZJVKD409y5+lG+FmqbRFrptSTxgytkeRYHGA
a2elNLyaFJ6I7pd6KuLHN5MJQMomD+W5WAbVgM0IPM/q+wa5CUNpXv+nATbYAd8UCKMClB4CiWT4
P/5zJj/4KzU7wU8eb7aDW8QggGHdPAIBP2jkOL7E/iNkZeNU8Lp6zM65ATAvhXgQXD4onxea+GcB
KZVwnGGlAEuUqEuABN8eVDTX9y7AqTyixVCaZDYsEzqHXietjDcVXEvOwCP3YtlS8zRz6yF/anTH
kPZyYPlsEkaD7NBH+ozM2+7rlu0mCFTkYAh71d0ivZLjWfmJncbBDj6vknC306rIqtNcn1apfu87
HgXUfcwQMpO9URPEKfhYP4AAsu9sMV+npMLGghlY17YFfA3mhvr1nZhFeHtJxiYj7Wots1yXdQ/u
KRCSg3uW1uykANfHJgu0ag/nfs0V1xl6LvIdreklWELBJW3v+jd1rjd6/eZ4wHfCNGSzwnAnmEW8
4/LFFtVSKo4GP18+xmjWXiRInDhY6ey4kvJ+Z1jTSzSBe1u6h/I9LBzLdgGqk9tFq0OdP1m3bBjB
X/3PdIq7IkyQ+3PGFS0ACrtuISu3lMnELz5Kk77LcUgE2lbx8rHlEd8qJE7cujVa7Nn6+jRcT002
Lz7rEcQ3YR0NqzvU0DOhVrxW83D6+NY1MX2IebWs/7Qs53dOvZodf+zootGc0QBQtAcJK0Ih8UtW
MhWW3u2Q+/QXWSv/EJ8hdiVe9fL+gUbVnQprHyM3z+IYEH77YW9DMRmp6WiJxbblQQzq1i87MMbt
vAfoNYAnewa35ARunA/0p5SHldYLmWvfRXnp2TqEASq49Ate/LpBGJWEXvy0LZM4RCYyDMyVHT9x
0AAtaLVbH0VkF53tDZh+K41kck98usA2DGAdd/ysvCc+QB6umvjp5HCCF8QJTkupjRhVBjMQ0l4S
6trYaOcRiG54b+WDoUJH7wqXgY3wQLayxEP7XXbsNmJ3Lj765PITtOYyNm70LEpJaMswSD2WYB/h
tdUAhLE3OzLLu9FmG5Cx8xiLLpoP/c4R2n3qMvBmVNZnbWOt7bwFxM+g5Fao5jMamcR3Vjmesrkp
ic2KHkgAYynEsDpkOE7/I0ZgyycL1Yvo+OEvHROPSqg9ima8KCTrk2IUwViRmk8SVbOENAlaSq8G
KGI/OK1lenYlZhnEX3GyJZAKe4Fu2WjhevUU8802dg8Lxb0tRG/e1xboKog5A+PCtaZFZGJN4NZf
vxhsEhcfkp+cuKu6GyqWoBtMjZ01GrRV7TNp1O9K4fv25L/6PA+XwME0bHkJiJKu9o97yXy/bgfa
8zdnwfWrEk7OKxg5Rp8upex5lvXGMMU8SxPFNKUGzsOMxWi6MOOdf7JX2z77Ip/OeQt3Afd3pUE8
uZtKOf/F5Z3UUaCNPDvntC4iG19LRx4XcL1krtexXm5yS/fkcWUFTZReyG8KnNn6ZfkroTWQLVXZ
IJnok7TRyVU8XovU1YaGir4pvxWZXKglBIdh/pR17/qL+vHf8lgMF0/t/EgwR2n1nD0JExNZlFhE
t4JG93r6Ru+REGV8easO7mcm0k7wD+w+N++JNh6P/ezaAfMWzDb8YM8AWfwmIuvAIc+Xy4vF8Ano
6N/DilIIDp/jPG0gTejFVVjd0nSvJZCfgG+tNk+MvW8nhMEr02mhyJIrfFUauMImigYlh5R15VZB
Uu0vM+Ob2R7IgmbDBMfhyQ+z4J399b2Rtv9iSJSOngaTNiaHgfsMdHgfQeIuspEliScN0448Q9zv
SIQK4A5J/QEDVSjMyyoQvC//gLthTysRdgCQGrVXljpbgMZPd0l801otdm/K2QWPslv0QBPWqgYv
dBXRMxmNxLoWhqlXn1uV3e6ba6Tm/jFk2cOzPls7i4qxfR7dtgn10VTygv3ysPdH2res+FQSPsXc
kZSOcp1BR5bKVOsOLBwCPpbPeiDE73M1hG2LFOXpllpEOqc5M06GJZeBHngMSrZQXWZZninkgll8
89NOGrqPpLWnBBavRuoDJ6EreiNSIbMaxk5NYBehE6TtpgEkxEF/I/8Bv8ErgbQUA0k6jL1+X1lY
2OcCsJ+n3pd5HLx67EnRFPO7S7BSBe74ACDPdhsAUkKe/qJM0am1dZaN7MqWnJI3ehPbBmORvi1/
9y/mKIPqYfTqLS+vi53HOAwp97vG8xwT/a6JUqXjpynLPv4BeizTffC+xPLCUjIM6+DNWNHAE+vz
Q+JmsRpcWz5ZGyzqYb1dKPmh6vslE2FSvFRZ0A8xNis6hgEyqP8p9tkMYrP+M/W43rrigdVa620V
iY6wiCcKp9wrKWKmv1Pr41CptScPcQX1wrE13Sw2GVqzlx2p7/Ya01W0D18f7P91EDdDrF4cpDZq
w000WroaQu6WjTIeW+XFvNt2oWx6GSGEaKebKWNiji2pIL12RPokVWZ2WIwbGVdSFcYWZEtA1DVe
EiEoDLNV0PSyOzCqrxcn54eZLQN+GDq35bxG0chSktwvTlxt3+uHrKMCijXW8NMRRraqEZqpfGIQ
9ngHntbjh3ZpderWbf1y8TRoeeCrM9oZ0IXCusKF5Ob+kXSg/dclwHL6q/DjAN7PormUTObo0rKg
BvWqWOa6x1n6pqRx4RojQOVk7DlnWspX7rxt8q21F1X8QTjH9MQpreEQ1+z969FO1ABbpGClkgmJ
1YYkEABgE9+tf8VIbAWPUZqkz4YGe+BTCMDwjRXNIOkj4ZdMCEhEFyxOaeTMt0fOQD3yyrKgNO2B
Qtaq42xVGBE6LhWeZQEkJOgNdMsXDLkw4HjjB3FYKnUzj0zwPRq2Xf4OCCyX/36/9dZtDj+n+N5a
FzYTnLYMNCtCsMyBSZTA5AGcjh5fzMUbOFttOVZbhOAVEpPSqKXpaFbD+dquEQaZ9nOV9gwxD3bS
fJwiaTWLk4Sxu41xipm4bvynHhVY+pTl9W1QeEUvg3/ZuyeZHqyuoySKDgNv/S/TIgLrrWL0LnPy
ZG/OEThS5ZfgZO2wuSotoG626BLM+36E3m9MEonguazCWcBfv7BLV1vOxUuQSe1LBfS2QP205Dlf
FfiFuUUaqNyXBF1S04Incj9XpvqMTUKVNg/xDT7jlDha/TfuaKvzMF84H+OkpeH1EQNy3uainzj8
cGk7e7gPwZ+vncQwUOb//e6vkWPAuamzpA91N9wVsUlRWqu09g3BUcYi1RXh1wo4SKVg1sc8Z9mO
K7Y1DFdguVZsBjkWiS/6AQ0ycBofOr44IVFAJ/LG+2CrJbOINPUo7yK82Oc12W7svLGZhbTiDq+9
JOw8xtGJXVL47BUvbmzkgDVaFbCBkUa+jxJqhYf1PONrFCUcZjdcJgU/+bnqAmnrV5E0DyoOOBnL
drjO5dM8DdlN7ER0vv+Ohlr9EGM7Evel9hzkqTQmsT23rfNlefB1FvSDMCf1ouDew/2z8tXrTgyG
zyW4SgVIyCoWwfRisDKlrTmY8FjSt9cPE0eacdlq7OISvH0aciQ3KKRxrrMDK+8+/kd36kESbuBV
SbkDx1BUghVdUF+HRak0A+bQ8TV/lDflREzQ90662inJ30ZIk+/R9xVmGSgkKXhPPhCv2fBSJzv7
Oi9SqCnTiEQvvmuEm7a9i/lTPUurd68G06holQJXilAdFxBRLnCgyHYHpSSYB5a4a12e9Q1TZWqz
88LDE8iVk94PkDj58a6Kt7Y6yo0krfCenf3c8kkEhjJcOcL8Yyq19Vioy+z0tGAgsLu72rDvz5Jl
6enuBU/6/nfNQRH9gf/aRMQIJfMHXgojT0UX1xjD9UBZ73WSISXJELJDOKuoGp32XI2ay3QVsL7A
r1tw/8q5SeQbIreVop5k3i3vtFuQgZiBU8V0FKqGqUs50tfllWRY7/YCFIat8OZa/w+/Z4dYRI1/
3Kuy4RYrrYk+w8hTYFWmwndjt1UHQfMqmlCwqI27rg65BDSoDMl06XF6Z4inJrStGFzBPkcB1cOG
E3PGYTxL5+iClWL0j1yQyyVZWFCJ818o1wvj8t+i0lCNwfyo1IAfg4pl8PRHDRm9SMh8xiOWdBf1
Nu0EJ9LqFzbfi/968SVqZ9T7Nd+gpU0m9BjJEpooAjNpuARP7re/Aa0Ci6cxcd9p9vVdKfsKfY0+
hjlmS7ZURljZyCF7ojZwbblCxqtrHxU5BEqRZqQY1VgY6aONuGdRnuEBjifwZXjVo86/w1uMpzoP
KOOB+H5J3N/fnhygHo9rCmjPIIb4DlEVn/UJJnUx+dxSJ7NYpeu1mAsXySYL2GjYzvqB4/TU/tqK
Q1j9EKGZ+nARy7SG/5BC/Jp4brU9vASX0akrkPzqbtiVweTgE7P+CWQIWLVtv+f63pqzshbBUzzt
0rgejBUgPu41PF2ydiDRdzwG5jK3lytt3Jb/jv9CCTtIq35n/tQ6OzCo3RasAPAiuUMrdBDhxARO
Vf6+Isl8edYB7WwdmajuMKxcpxw61Q6WhLim6yYBc+7zFFNEUPkImuSTip/GpSxFrTE02n+uFBgY
B1hiIp8wJrvKQnCZIsIpYFRNE5fv71RECEkUf0byQ4Ptkbg6n7Ya6UFaV/wXjA4nbmIAqpPUhwg9
wDjHwjcKLfyyBg56v2ddraSywYjrDf0IY2IYhU+KTVuC6zrn7eCNBfFIoilCZFdre9KTLyupfHfO
SdBNiTtTDx+DkDdNm5s//tNYypO/lThYAAQ8LtlNV2rkNk3GcAIHYDHFBgMETbEfMMcyGtI4oB2J
7cgkiJ768ZqsxY5Ta6LZQ6akSNzpdvPe3u3neYeO6/VTmWpHsxmD9MltK8+7YPiH9XVGZQh7v6rT
NqBNM6GtGNxit6VhFrOLLfKC3yi/6kyKt0j7LP74YuxwJhmkHXZ+lqZofOdJ0EhdfYBHaq1Q4Qrk
vNyKGOw5e9e9HHdvnBwffbQH9qRNa4Oh7pG4Em6wBSzpdSrF7bQnHM25NbDnzqGfBhyyVyJY7aNB
NDY1/Fk0aTQP1qboE4SiMpUVmdQ3sHjguTHaIj2eFHX/s7hG1FoY83aVLmOLyYzxukTzQy/7pUps
iNY+JCrX42nCXXWEHX1NIM065HfQ2j+/tzMsXq8stKGCNFDiaEDHZ5D4Y5TKRjgGHaSvppN3NZbX
rIWkwSBXi7ravTYfxueX2+bHkjKHM5PSRkqYcFDedSMRQWvGt0o2vCkgXihYaaaIHptLvB5UViIP
uhvRXA5KgN1lWfEwDKdbWH9YJ9ogAePZQTjqafI6j4eXyyDT0IiHYWuE7UlfKsHEsQBjCOV/LfRe
zbBnJ8f3TZirtorasVyETmc6H75O3jao/eTh677lP31tmFch3/BChCX06Rbw9klggjYUMS88LfWL
gLpRArlHOYK/oTzAdKXXj9Usw9DXgrxEUuWn5RegNuWumykIiKV3Eqq3QW+yAbSOTcjWlABM3sL5
zFbhzboa4dwnvT9Yp8q29vC/8Z5Qk257Cleg5VmAxwqDtDMyiDsRQUMQQKBmtWRDn+9kaij1Gpwq
9WwJGJijyqHQBOFKUwiMpbvrcOtvg0dqI1P2Dq/j2QNNQbGMKNEy+6SXHPGANI1kWfIBQcPsMXNq
/M/ksMmELHrVm9jdWXIm0kAWdlFWro0fLTNVBFDg+PpZIvbayeOurx+jFPHbG45itwflYSsDjj53
zMG9yWq1F8YtxxKvUxU2iuRLYWIo2257SuiL2wpHkJ4Vg6BMVUowNTdH6wmo/EOJTUNI+WxjYIKS
DfCM6bQG2wvuOt32t28IqRhg1xKJPQZWNYPP6UHfTBh4lT7j5vxo8kA/m3YK98aSwbl+p1gAu48m
MjJ49zpqDUos0ORxZZntD1JnKFubLbA4ECXeL7NiVOR26ye9+A/KB4y2QbYXqzs9hK4MaAeXyBbC
6y8f5S/5j7AvgtwLZcHrAYSUPI1wxYxUFicwttqiUbCOB6i5xTuc4Ssa9kOK4i5PBRMFubnFcTub
ly5ZV8X3juCHRNl4TnwPIajJ2ZTto5ZhTo2oVeiiNLGqNZ9d0whl//4BCA3y0FQ5jC6ghjoRcT/3
GoFnUmwVTpaQS4IBbaIZp5pdC7xWoUoop3RC9srdNyUBmuDKnwu+Pjkm87ZVzVLOufqKfp3XIAuq
O0S+jFnRLbecErsyCkSQwUBQDP6vbNrTEiNDiA9x62iOZKYq8zgrqJ/qRKIS6wu4lsbLCKFfFt+2
izAF40ld8LEiPmQHWVGhdq/RqNOp19jr1DFgdiW/JEbnlva2/E7XkC/eJKJWmwHYLBCs6rjwcbgo
q/6qMOSbwQf0F7iEp5ZoCrphTYys7et48sjzPoGAOA2EZ1IT4UgttoQELNIzrttAhpomSaTQakPo
8Oc7v8vGd861el3tGuJ4JaZ8hqBgJ5DcvrUdLamVW1uKToA6cqpeUV/UVp/5jy4yEvmA4jL2+bIn
4M+N+ScjZWw/HF4DxOE1aeyN/KYupPvM4Q0buetW2fIupOWum62a1gXqfTIGMzx2+50oWLd1YmXl
dDjczk9yMLzUXQWtfXaLpvdguQ5r8eXnhWCr9NlGarzBPATm/BuhNAROhoQAzwEw6oeMmK3ZqfWp
RKrmcpwZ7vWIHKjjeOR2FJEOswbRvqQkLH4P4MJeaSdbCrseATnDvsixOIC9qrgIK+hAKw+qehfd
EN3lsUDsD0biWASJdT1Ce4rOlpTRI4mZEmMuH43kbKpV61rwFRXuRi1KwvC/UJqrTCoLNk7xU8s8
YLR+OU9p9VEDi5eloTA3WDSkz0U+A5jqHgjkRA1Q2UYypkSqyOpswxiobJUC4nywsdbcgF7mqc9L
FG1lb1aN45JnhYkRnbtHfOqGvtyRA7VpGP6Dg/oci4fKg0zAc1SFxAIxT9KTAyzeXSqKQv7Il56B
xnyf/lTCGfvPYXe+g6dc/wh6ekE7NobdMB5My6ugAIivsz0PRwuiDjmPLNRWanGI7C904KSuEn23
P3dAsj+yLrFRCtwKOftxr/wU8AuV0ZgtCj7NZThkcEbhMP2lf1WJVLNvNzjIua9G06JhQ4tc8xLx
z0tgC6URxnODKjs5CCXfCbwQjEmy/6tWJBIpoaoMLtXJYGZozDjrJNVDWhfVWgWBhUM98Twb8VZi
PZMa/AD4dYf71vJ8DAyF/Svr1BAhB+RG0tNaia1y5p7Vng4L19t9B0CGeheFuhuxtmO/hdvdBsAt
AJoa7+3ClrWV+AbhwqNX5Rf9le9BSO83w8z534CgxpR1yFTkAP3NL4zwHS4cQeApbXBNnsBcqe9d
QdbTq67o6zRaS/VqIy3uXV2z2mpisWrhZ4tCyOIONqxN3F3CIVszdk6Xtai2LQx0gulLZj2PnugO
sfRh/OSq+Fp4c3jodaIChnIxfzmG2y3cbHIlV2mIWbfWgLaCOhWtsg+LrT5+2jlj9pgZXYWtGaBx
jlnEWVL72HH66dQDeMfU3we5rSF92wpU4mHBzljrV8z3Tx1G3bWBvaZwEZ0sPRaKxw4tzG4+fNkv
xwZvgntWNsM6z4Z2KiPVP2xuuw9DGFkCTavqCab2bsb7q4vzDxaCopixxLTwxrWE6qLfRaQ1evvK
636Pj1w51Gohjo5X4mvXbRNDcpU4il2mUbRAbdwX+UrXxyfcpqSzs34NjLasyTSnnPldTD1GtrpE
s1MKAk/CeMiO4MYtqdgj5V/L8TLy+PyszVE5zqgt+DRP/UmmFfO7UMA9BUpAcmhY4K5ECdYNLQIx
itQEpooEV/45anNBSw1f9fIA6ZbU4ZKlyD0ye/7CnmHRz3+IsJ2Sc85ACmaiBU0QhJh2qOkgmY4e
zL+6Bge7FSsY7txsrAvVPbLt2AXzjV+BfSLN8q1QS3tHk3g8OlxlTAi03TQOtX36k9m4purzTB5Y
u+Ud1OoulvvFioPsr9C+EWT0HKeXJOw9xFdrKw5JFvMkTO5x1R2xMcrXK4vGO1PGzbxjnQrlnbjQ
x3HNJJ1B2LbDh2Hrz6bV8WY0o8cSbr8i9aA1rA9F88grTyV1EsGsC7ntfmiHnDiVGr8W4DL+zg+O
ndiSc5iflVG1JvOMozcyGdpaNrphdJbgByVBRzegzEFGqGHAsAHB80n3K2zI9eHq3MK+fmKBAZjJ
J4Mw+uumEUqkhyQRb6YiqyYQrlrTrId+eL7Lg03GzPrMUMVO7kwKJeHIWIWcTW+3hTKFOQuwdjeH
AG1Gfx9ioGRNlDvUn2VJlz61SqghvBsl+47DJiJDP6ay9vrpprJmDrDr7T9pP5S764AnyCaf5esw
ZgTXqcDWhH36qTmJbjhKggMUaO1t+S3+wS8+Z0Y8wKPbcF+x3++6EkiLGjxfGwNWzlWDV86czKcY
5XNz+TGTlLxz36fylqbE4ptwsGRldpt/8EACRU62N/BeIWG+Dc9m2IdFH+/o8llVhJMx3qFD3zcz
OyPND5AS4PslMGTn7LQSXCnruVyS5IUVf/pPLvizLovvlyHp5Z4RUDmUWrypElOeqya0CFMVvrlH
M+ds209F6WjkdALOr2sOabpgjujRyPtM5GAEU1gz47oheyZB4rlapcrjAYrTtPK8pUxr60mLhpRM
ZVftng95dEEzyV/F+ixDqp8qL9fc8M4Z8h2hngt1ZWarRxkdx5iX6LYKboM4iKDBdbk6s46vGA7s
pPk/J7lxOonirVa1icjh7X8CzMQmWpV6LuMqWf3f/ZKuYS0jZhv1HnQX9PWvR002QeF/T6MrYzy+
akwzKLFxCBeYdXD5Snh7XaXPPFKuP1STJqwtUIseyDfZvAQ/RYlXpGsCE4x5L7iUgMLwKe67a1Nb
01veCN4WPEw6x0IM5qNdW7I5xs81Jt7utU8Q5C5qV4gLcEM5Pd5T/4z1m5R/7RUh7Q3+ydechTyE
ocsHy6SP5UoeXlx5/doNj7mN9sVxkWahRfSX1xlsb7LJVd4NLmAEgpqso68SNLPkz6KcRoSdDy4s
T7PQv69ZiZmxCEYk9bY/Ts3UjbpQzhpw/yyl7moL8PZdEvGQh2CWnJIEr4GxgAVWbJRzHGNcBvD4
h0WQe7WEDw/AnB7rWWFn771ZKl/cxC60mEiLGWu30w2SAX/K0djvMlQsZdmZY/StlV2FcD9rQAWX
Ba2pMCNy4/rom01bnqAPszHV3TA5OTlQhLn7wKujJoN9F/FPJDS2lGn901i/5+f82Yc3PY5CY1x8
qD95Os8GyUKD28P9+FWTiNESvCfSmSb6mki6HHrq8vmMyPAiLQcZnw0T/1EqW0MeNAXiegEy3SPk
JHVB7YCUU1xgb38+Jd1r09vB9x9HgxFM4IiJpiBkHYMCrfElLfC1i7ZA+l97b4/qs7rvDzcr21dU
WkESq8IBRhhylhojQJTmIhTLFlfvO8j2+e4HgkVJLphuFcRSjWC7tgT7SJq2dR4iE/66d4aMhSBm
by6ycThJx/jqefzqhxagGRVqClXaI8YkSv2cHG9+hgiOptAhNRv2W7doi7W2UR29J1SvCiDqA1sA
3wme73epxb2YXcrIXkS8oIVYNewXUAMl+tctSGnJtr+OTKpRI6gsVkdwf2Rvio3P6BUlm/7z6MZy
YBtlXqR+h9aklSx5U3u6pTNs11DgNuMg8+juR0lY5gdyOtJVDELA2AWRuh7PRSmLnlimnA+OXpnU
P7A3FOpUnGfTQ0zqzZO176ItiOCeKLjNhIV/xb7EGNCoDPGbmDRhiuPy3MkdN8UM4aWjce55gQuS
t3V3sh8HfaksavBcFfNG4F6/a4u2EAGnFzBb7MDyo0zhLsfvlPOnHuDPxCwWdeb9eRSvt3mvLusn
ZQUJopoyb7y5zyNc2tXdB8izXbBRtYcNshZmkJfFgcR5vA5yEZvr9cevrEYETjmj33srBroUb+D5
6hvq7I4y9lXX1pSzdM3pJUuorMNI6KWqaighUVEl5au5W1UQjWHYzO/+6E4AqVDWcpX7pWGUrNp8
2jDAgr9Fw/k/gFpWeTMvOsxTz5tLRyfPcGOBlR2x3aonsRcS/80Vb13FYRRMnGXusJ0jRyT+YMJq
aeUdmDMBzNs6znwEO/2u+hvW3jRTd136Ds02jxa7J/mvoaHmFE+yy6Aib6VYSuwRos4JrSEmd9X7
ZAi7IqDx1ibIhRFt9FqaD2p2PuwJgL7+tJji/lHUtXJKNIlYeh6IKdVcNN8HJ8f/j46ddiJY8grm
GUC/+BviYXFk+adAle/kt4Er77CUVnxQz0cujdCwqxS1NpmPNx89/IDjfxMPvmdO7zRfzzUW/H8C
AEErsZMmcpJ2HxKyfTMjQkJWEX4NBHzZRQ3zcc4GlnVTPHGkoDk6hiN5AJWcv17uK4yibvWQDFQZ
jZpq7JITrKkSv6oiWzc7+D4+6O2WJSRcJuMFNsAI4hKBNfntNbJb9OlFPLUHmH/CcU6pDHw01nsN
+BZYXyEpwT0qxL0MRA63CKYOpV25Y6ljU/dDLtU5niWXBbXFh6MMwc5UQo7+1EsAaGlsif5mGIf3
YRo66Lzll7ntE1YWCJdgO5F7yP77KJpEnEyjW3dzrN/LWys42nEE/64oPS9jJOmgedCkPWB6JTMK
LO1kb3peZeRKEHMBU/+7zRpGW/Xhb3LoWlHRK3/yKBk64bgYYFPOI811tQfwF94n1cD3AQ2c6BOU
IYMsfpFYS6PTVxZuQnyOrknEsQlPxv25JZTB2bw2nklAj3dlPhBbuBdgh5un7EZmwO1uYfzRi4Dr
TE9bQDbaA9l+HJDXzMDDA9s+5MauVsPRFPQ5IZo+O7IQ34x4fD7NvKYOKpt2qn5VWbwhe+ARB0c/
KyLB/EmSmUKKX10WWcvV5rlwC6WyuhwCoy0wN25zZIonds54Yl2xMV2pvT7970WOv7dSuZnx4kDF
YEnVCyJts90xT1zDSuyQb7E+Fme5lTUKZRZCRZOF67eJHSXc2DDXPLChNV1gdHapjxDB9uv5IejQ
wlM07tCoxT4fvA+/yhdGjaISlieD0CZL4++4NPPjk6nyXlr0MugvSXKfSFwDPrmCE06AqEzhYXd7
gyZ3DjuXw46EkV2cWVll4ePTzyGcYa0Kmq0kHe0T7ZHqtm3q2Es232FlBgGemnKV0oPYadKJnJJ+
9oepI7UvJoEVzqaAjeGiBukeAoY7Gdrpv4+Pvo+Onu+cp8WHREEbyAJvaxZz3fnhTkc819IY23/b
7/v8gcDKyKiIx68P4cF8JLydNLH+Rae4ZftLa8oppWgKiTyAXE9R9QtvYQ1g6r/HieAdpn4c763K
1x0wAmhacSj754FIho/DRYAcqk+kayySggZ92w3O07rOcdMOHCKUz6Not+oHRzoeObZwUhTukie/
b8cbMLtQJjsvS7LfCjOTMlNCa8bsTHmfr0zh2vkppXtsWP5hGRRbMp5isU3QpGDcXciWup8JAUWV
580enCFLckf+wjlhhG1BjF8FiBT92yhNfEvDVDIr5DrdBeFpG9DRnbfAtVHoZZ4f9MsDOiWpV9A3
veFoMSsIJjZgSj8LfXE+wszSBJj/tygU+drknVvmUzfHCogNd/43XvhuIDf9+a+hylbt5+XlKBYB
fpz1kR3IOwk3glBoFvOXtTYzBKBkm+YajTjCfzco3ruiGTCrgcjiQTUODdD9jW4b9Nr9iADg3jXc
lBnKU2WXERiAMNyg5ZsIMCzWGLsFWbtT18eZljU1JnS9NKO+Wq7nbpylK6MLMkZTBlqZFwqHuvKw
k/YzN13eFwKcTrwmEI3dZQAn2qU+3wOPxP5zGsK4dbbDFag7a/5zWBNwbvhFejm+xzayeb9UsffL
dXwcDkNChDFmkhZ6taaWa8vr+blwvchIobdHHJ2bjYMkb7x3RQMkKAH74Yc5wU867QwZt3DAP+Ip
nQyhs+t1WPvUg1cefGAJkCm3+d5YUUI7hRGRV/3RCwzWe2H+0E63n9CtnqrNMFUD/tarORRH3HDb
5+Ti1ONEspet1RCIFsXK7xD/GxGbq5Roh5yLCFQIQW1j1eQABz/VXx+SYe7u4hbNceV9wyZDx8/z
I7oYOHGgY6YAhh5Zcj9Mp+iiJbV3y+V52/i+MRMs9UBZMxWmIQRrIzlUY482fSeP1e1QFG7un4oh
0fgoUkBTyck+TnB8SYMYcri5BGxUK8QxWagdbDUVJYFs3dYZiDkhXpQW7LXlNrvesfkwRt/sXwoM
Rv6dufGKvTDe/8e9tPyY3wDYXCbUo256boLnMmgvt4PAPmadnrv8k2YnFiTOLTCjrzVr5p9fNuGD
TBEMQU9jlrjGb1udz1gFzdHQABKouujut8G6YNbRQ591Syv+aCQE9BlQEc5a/JPgROtsFUHAYbLG
sSXPO5EgI/29I38Q1lnT0cQROIB/XyYMjxEvbXAryXWDdBseZUh6FYqz0IeeG6cHKKm1V5u4tH/L
GvVZx+rg7OREhk9k/hOvOGhvtMxWBZK15mbdGXOQdEXyg3lX+wuBV3/fw4GLxTetcBmDjcefc7fE
yVHBkozghzvB/LIyDChMDk8N1aWnSpbawEKCybvARHpUIwOfB/pZ3HSMuxGWDiQ4uXUpSEqtCAQC
gYpfh0ZWFg6BgIVwKHjh3yXqu84iVOOX3eNH+1gSvWk9LBF1LQzlPQPakwzyrDdZhTXivZ73E5/k
WUITBeSiK2eZ0gSxFAqEMF5IU8Z5B+6rqVSFJvjx/rhXi0ciql4s77BMDm7YoIBw3moiQ/IHril1
qM4cKhLXJPQDqbkh2FREjgadfH23YdMScKPDgKypetTa1n66O2UqbquDDuRBuLseDeRxjuVSltMh
wDHcn3ty27yLtprKwzvvgK0fcr1pkPpAPRB1/y3uYnWbNXEbYyDmavxGl7e3RD9WIweZfPuBtWA/
FYRKIFTbwLESZw7BGTIk2UuZgMUuEGN+B+ojCLIc0dZmUmVm6y/B0nFY70QeZs0O2HXPakMVRS6g
xNxRQZ178YEZ/KA9Ndfjoh1UJNLZ2cmY22SAfSx2Oj+gf96D9/PmbYmC1mrIU2hAegyCT2+1ee2l
vAQpyMl9jukeBFGitI8n5wS/ElSBdOx1LY4I13SPeS5x3we7vBaium9NtIPxCKs7XanNyiLWYyPf
5GIJoNLORbvWVFUdnDTHCJVINIAC+lWAAgD+ic/vzD9QMt3yVRfuYGs8WlcfMeRuEVtboyUhm69M
ZlRS9Ry7m8h641TbvLe/n0mea/4HFQ+Y9fsOI8J/ORiIgQGrt1XusDesuc+djtxlH/YPerHLI3sA
kLRS6GIqghzq1v8o/sVhVUQ1TJPOv5RYC1l2ZUbsrp0GYWCZ7ebn3RjrMML06l039NxvtMjrK9pg
Bawrd7KqCKJuUTtsG+yWfR3Qi6u2YHcFiX2FpG9mmd1mCWvMBUoXYHj7+ucmTGpfSdFFYMiVgitM
WrbYBpC84XAxbnIdxXKKzIXjYnvwuPAWAS9uPckOsGYcfx6V+lmeOe5fqy0ctrxeDx8HtEKymSWF
/qgZssLGzp1U+UdSAiifVAynHnscCOqyzHYyDi/eAslMPq3coFQSQshdV32jV/0XISGW3lTM+PrL
Djgrj4hPPl34UpTAI58JW4LzfoIpzYBTs2JIocd+0U0rju6C5ZDJ2EllcjzITq3Ti6ogrsZvKIkL
gGQNKqfWKTxDCZaJnIDV1sivsNW+BfV+BGqtCXY8AbhLuhFcb0YY51d6KIvZKLHB8zs5yRCS8aEI
litOA9/FYNYh+tROSfmJfcI32AGCm22mlKXmVkgk7bkCmY1s6qiXAXGoHNeS9XOq/9GGRwf9z9TY
6i17cm2DpBmgSMKGTomiuQgZAtrZmvpb0NXs0oj/JHipV2GOBiuV5G/r0cMk2C0ELflDjNZHBtaQ
k63dRMgyPv0VrvTZ1uoFy/Kjs7Pf9S8GPQuTSL3PHNQvzeK8GRTOYO9mihrSw5dKwItB3jKm1OSY
9s9v8zovnfxpLOOI9fLsb19JqVUYfzNcl2HkJOkIhAxzmNp4IrHqr5sCHzMOoOYA8PzM+xEIVcml
+Uh2dOESLjY9IL3ppSaKO530NuoFLHan7bN9oKBBI8TTouuMJfELvY3TzXV5HJI0ehLyVuyroeBS
PVM+KLxUtslkXn32+mbzHUJfhluH/wCpuEM3AqLZOCHGoUwAEg2PWJY4kXqcdBjWEOI1x016tFs7
D7jeEe7PNHuxCxjMy4OCUkg1JS0gXmh0gj6Unxk2CfqvanvjvBQvGMvr5p1impnVFKcIlyrqP9hD
lPDqsDI9qE6EpbcK0/0n46SwcKMNjXeVSw8ZU04HiCLu6OSpnD2Ugyshc+IfCR8I207I/H1kvelT
yH4JX4MGogGowW++g2q93afqNNU7u3y4bVFNuI/hKgQep3U9yVz1p0T3d4tHJKkMD99OYuS8nO3U
73oD7rdYCQ058ixoXS1bfD0LJZsBbv5m0+i5SVDR7t3h08V6HdRQWlHqoUgGbNpbzZ1QCoBpoH+q
Ji1k1uqW1pAA7PvJUnmqHlC68nmazEqIo4ZhHTEu+kBtsjgc6pJwq5Chc0qwmFhGw9rANR/iB9Hx
y/7Ust2pv9vs3KUjSeMh5BUfFvSDnfp96eK92nm4kLFyAipWMs6AiRWkiMBVyCH7B9HHgzGSCTk4
KpiTLZdQRSPvtvRg74auV+5xcStaj9zwnnr/t5GFb112XigfBZtJC5ZCKkvd4tBIwCqz/8g5UBpp
cuEY41ztzfuul35kZnv7EtvaCmd0y28TF1xk8L6hpC37Fe4cIEk0ITS3GNmZpO89ztijMNlgjAw3
IowiuNDLEghlMcikuVn6Z9mve2/GHFN4Dbob+aRSDGS1mrllF5/4574T4BGLee0mBr8CGhcZC15M
IzTu3Yl0qfmFMcWGDHRCrLiYy5i3ckj+gQeqFx6mR/NKBxCmzHENndHAnFs49v2nwPUjWpctIIN0
QWrCDVVuEF6Jrej/Aua9eVf/YUacl+InUhZmU2EqbRJIvFREACrUU+zFSqc+pN7FUtu6iJn9GvfM
88U6jcPzcXyU1YXDE1LSOBbAzTbaVUrJ7T69uZQAHwH5Evd5NU5zm6HbNLFlUpPxn/ZeeNIygUgt
5TabYbaw8J8Ea94wazizbiGisgG6QoEx7Hw1lDcdk9P0+pzJ2vqq2X9IEd6eAK5YRz2Y7EtH9h/f
n221Xvd9mV3sn+xCI/6fu6qzgQIKlyZM0Qp4qe/yvnkBK6Hq1GDTQuhL+juIaTbgQd1KIxGJXTD2
5koVXgRDIHLfE9vtwyRZsCuxVlK0pHkuGzMiLOyV0y6krBOxoUnS7FOZKR+o+tccp6nzWg1vtS+T
sAA4SdgnaIiku5T9GjviTdnuKXZx8mlD6VuWQk3odsi6nHuyLRnWiHy82Pell8JScqtwm/7wmivJ
zic+5fIi6+yUa8YhFpDSe7QAPOcEML3pwayZtVzHNpUYXsUsSxC7mQRbhxTbGWHGGuhfqiwLcUrC
pLLntLAcSNYofR18FYww2wXOWHAh43Zq2ISYQmXiJiUCc0XRymbyCUqvX2HSpPlDij4s0FY79snU
sgMoG0VwTA6uiJ2BfKREaXOb5sG84XT4uwSbD+9pCKBh1vE6/Gb+HRvZBB7Atdp6IgZKym8U8/gt
9Mko6QvkvO6tkwJ8zT+gK6VUQwoPnSKivo+TdkMDpdIm+7u6JOi8mAQ1j4yP7Ff/JIAKaAtyP021
nnplQ7vGDNWZ8Hfb+LCu87zcwEq404CS3ep12szdpWJ43PPI8D+AtqVIt8J1Z5naUKjpoFiynsmn
2JFHTVTO4THjY2WFUsZtv34uBNv+yPWa4l8JU8JQqBt8wuTv7SsWhBCfGjWZtK02TGq1mLUUdzy6
RltS87kyhwBqcrau7Ksg0exb1O4u4cljHhHpTdFLhTdVqdGpxZkeXg2JuRjzvdYGJDANLC4/27ii
xTr678NbhdyZGt2lX+oau1LSNRC0zjbScobORHPbXMP6B5X0jHy2BPJxbChp3cwtZWwQjIU8q/XA
4BOApi4uaml0z7rONb64PyZqVWNgBYhNqwl4s9V+a9W2UUgtu0jHdaGqDKCMcJh9y2MrWwg/6oZM
hQKsmR7TYTAlGWXhZlSpwu0IOC26LNrD1jgdhNpXCEENKU7HxgofG6rBs4y/2R87zEUK92EmUrhj
o1bwKiCSaW7us6xZQkSqCxCuGPSJSYAnr2XHrZ35F1y0N8A+k5dQJBWWwDWw1bgfCqII056Bnxmf
KAjlI5AJVD4PY6pVKgJmkf7/yNBjjKz4UaafqIlv96daE5vD81DFXzMDDkiS8M8LafUrFONKhugx
x5NAuv1zOw7/rCCES6JUJ7fRpLX9/A2ffAzxcss/A4XyP67j0FEjTn3WD/33mP7WGWlXVk21JHE+
/b0nlSZ7J+PW44sdGdKCNcXRztTyF5eqnpVvii6KsNTHKpa/3f0PQIm2rOKggDGGMDUT9zvm4WFg
iS6e7NOndRwLHgZhNcdxLeXM1vlRJn9RAYWqy0H4H5HiWDFK0MWN/02iZUWdDbKcPkoclZxOfFgs
yPLhH8Vaq0QfJdrGcPKK3W7Fw13h+tzmYNQw0EjMbyww1QBsmC55Q1HrHU9QAcNKWBRkyoyqSYND
5Gahv+xSdB1vItrCg42qKNSfjFTm84LxPRqsN5ZHZ3AnMp4wDintA7+3byzDPB/GBFOvXeLbW1fC
pliRZBhKUsqwDnkrhDZ3v0sadMwj7IJZzAUC/NrCqNaw4j80Ab6KtLtkO5++i/CzS8G5IrD4Gtv5
VXb9+p9WJ4D3tduC3Bh8tpnT5eEubnSv5y36okhHY8WIsWFrTMkCUYjkb/d4730CBdAiSdHuWcmx
IsUZfaj/vl2BiCPeaHrcXLfiyRX9wFGNlZ2tDS7SdIAFvRh3fDXDBtcL0OTnVvM4u8Jy/ccHCRKN
7MmhiBiryymXq2v1tJe5rNRGhBOgazp/4bUzF9bGiOT+lh/ImK1KYkPJEYQbdlmJD6MevMkGZU/5
sSZ24BI8jrs3TT4L3uIElmGFKKumCpwOYXw659H0eaK3LUe82PPrtFcwXugoxwFJAxzhkJqkXx3o
wDluRxSp0e1cSaOB3tmdUPCWHbQIVan8xipsXGnrR8GH86CdBbeWWsK8a/PYswfMXchIGygxkxVg
K8GdhqBgjX8GoU6TwZ1CjnV0GyOoFaEFFeKrTt77CO4D0qnpEHCNFdcS7V/UPFR/zpYqa0yNbj09
8ukzZdwJxFMDwwqVju0YEJVYR33680PjOOYVl/+MOaEnGm3zfAwEDvrwKOknT9Gv0ap/MRaHsIMs
YNfaeoFmnRqNZp5CdixgWAKZ/j55qBswbLOpN4XrNfrL7OR/h6J5byDq3Io7ZHmJcxfUlsNZI2E3
ZZ7ARVduhACMfaLG8BY0iqvrn6qC0UyNS8RpAk9lkC92BPJIzAOlBVRjruUhZuy+OqZTXEu4lHnK
oNFDsmW/m3lo1X4pZunLjFU1dPMv7nllBD5Bnwe67wOYHLpvG64oizR+3qgBQQ8w+g0TFAOE6rFf
LC3S9phdVEGMfi/4seB3WwiaMMRjeEoSQqHqIudLkPKGQoI8ZkQUXm1Szs8ihKSEu6I5eFI2FlVE
9rFnKQGywYNdeURJPAoNe2OZYE8i8o8Vtp4CxBWfpT2EOsCeRroP7vUFYcOIgoY9PmQViE1NLzBh
RgmlU5Knf3lZGcIJWaeElP3HuJEfnEoPwAJT3JxTGXbI5gGX4jDBggDVA4S1bLKjra/e6PdnDm1U
KJHBpfI1OWOrswe9C3I0RF+BcH79wwS2zdwU3w43V5uvM1QyU2bFHBmNr13KpWbaZolUKS1Wyxaf
2A82jvPMfV4tTeTg8N9Gg7xvXDwtsi1PzDS7GuTurHGnn+2iahiU1+35y9okFRw2wRyUPhmfqKiE
xwqpao1ybOOl3UiexUonx5Eye9WGfHlgQneoXCvZI/eljWUs6DygdqxAvH9Aojk8fbmRgv7zQ2Cs
sbvGqwzhxwmfstCDzpFKmc9RRSjNp1BeONC0SnzFcoblKnI70qEUcWavmvmBgcwQSGG6cVZ/+un7
EZOUrPG4JK07SwdvtUZT9cbZcTjMa1aZP143SAMR4mTaNwFN4Ve6QlKcc092qMwhMCt5ZOgb3nbb
4KaFLMlKaT/C94Hvn6BmyTkjELq5PIOLNVC/dNvHCab5UUxEFMJEU1RuyjBU1oZkanyCg4tMl6x8
HLo50MfjWOYzeKzEbPxuTQ8gg5tsPNWl9lu/cX7LwodCJiwqCAKG5smL/Al+g/KUreYXLMcjLVvF
+kxPGwKiY5w63maJuM+fp44idr/rA1iFji/ze1FJBmtUYkjYcqF2Ul1Sw5GXeEmd+pYxOcUIOtVl
m3aIzuWbx4F/PmaXnpu8fETha9BOOYoWR+3kB1Tj789N8wrjv0GuQwYgWAK0+rsifk2l3DvRWidq
/44m3Sc1meMKSp6JBs2Fy3hF7kDp714s6jcWWwTkc5KmAAAj+Vj7hswZefwQa6Ns5qTMiK083aUC
RRt26c724dnR7VPf1IbNgL0Wo2H4/TVlJ9jdQD3js2gwATpOLJuRn0uA23fcDtzCyqc/FtvvfyqY
ZSMlo4B2QRu/n3dQLFhZfFUCLdWuKcby/NAjs7zcRJv08obrS8V39GJxk0UBOeKMvvtNPyBqFBYG
uFtjQROJENr7b6+I6zfXoM8AHhBmjqYAZzE798aX4pDEu5KGNYZoTACetKQYmlGus+r/mo4pRA1F
Yq8Fxfi7CSr5fTCwbGSJpH9+LQZXwiYLQXDfVqEd0DzYZDNjXzRn6U3tZEAM3LKrSy9av+7nEm76
0Cdetnd7EXiVFfo8uwU0070PdIAHM3jkBXVppYfvWtUMPDEDI6Q+srG3q/bPjk6gPgZ/uLdzm+jx
GcEEKatJzNGVd4oPuUpde0Tc1m4flcfTJkV/0TEqsHegXXtGGUHfZP2rmAk7OJOeBTZ5YFYjtAaQ
29b/Te9xKcv/SCCp7qaPau+36xeIzpwKIOmyORJggWAq2nRkUk5uO3MUkfanhnWW6iPa1a9BbSKi
YiVu0YR6l8RmXwXEO/NYbJFO8GLZJiksjvYm1s8kCcdc7it7C6Ptlf+rYiPVKMOf1yuedLTtnYrh
pDX9TBfsoywDhmch5ySe4fEqcOcemaSyORAnJYof5w6kqq8fOxQrAq0byQgtADiVMMLMldXE1h1e
oB2FVIR+441CzeVvwxsfyoWFuNR/tVRVkLTbciBnaP9q6wcII5pQsNyfWl1AIqD03oVgAJCZMk/q
NMWCsMIzS0SZon5iOSS9N16SjCRTIPvbzsrvGbrGh0/7UB5Ax0cJpaQn+6pupXwo+7NIUMFEMM6l
E+aPr1FP+f5VXs72FPxcMuvbWomJzYD9GlyurRStBne8St0NvXdkWwsxzrECeQkBL4hjwPs9eHeJ
6EPiubivZBTFVEVsbvF6vfbyAcBGUPAznemh2sz4vh8w5u1jGiMWnnsnIuvpCUfH2aoOpBftDafW
biJ9EMfqCcB8yxvdDbkq/DaloeIQrAOX6bqUgo4wCmTWBF6jh8AVpwno/PTA83sv3eRTQfKabU0l
o8s9amjqmmOxpfM9zOdTUhenZ1NvBJXPAk6DCs8+GD42GIRzY8zkzZYmgNU3p3LJ9yDw4MPEVII1
V1/zEhAXcDPiK0dbNLjThIUFz8xofjUowP7XI1kPon2Tu3BB/tebyq7bm8U82P+MDr+hnuM/ei9J
94IDb96z8NDLQpGbc8vR2teBe98BVohPz9anjWw/NNBaCml/hqqSR3UmASRq5FgXWMgdC4GtiVqQ
ewPPTabgpHyxlvYc2YB1b/o4QVQqGp8Bsf1pJXdkGt9fD84RFoNs1UYIrcqBTF+wFMQheekxcxui
1RoqPLfa20wb7JhmYpx1S/71MMQLWqzteERufJzPCOPFHO483C5e9P7zBigu8CG+9pEUiFzPxi8u
ZmdNPqT3MLdnMjRaEhCLu5ce/yRePjc6PGu/EAUU3S9Dl2ZqJmEhyI14lmgsC0KYY+9n6zWlJBum
yQDyZ7BRNcOj7i1k+3t7jYl3pcK97fzkRBZQ//mZyBT816Z5NQeqKuyPAN+R1RDptonZeQ3Z9ggF
OwTL4JLz2iUnTXGkDrsaCme/Mrf+HNzTl70hgs9i5Pz9DHQQ9NKSDt+HqMk87rRhUICNBU4Wf/2n
w20d30/vNXJuwPeGuupx00+E8YMoZPyRDcXg645pKX5x/loGBbQ7uFd+u+TVIzQAmQBD47h7FBdf
v8FO9uAEjSeCOJLAbFCingXFXKRiEdQpuLHhUgJZYpawAqWjMb8ey+J1dhyvrC0kMvGWVkLyUdGq
Ti0d6JSve9HJhvFDqgEvO9evZNGkRTH48545Z07c/jiNnlzPQA/1vAOgJuKOnhxONzENgO9RFh6D
+9bDZkaqRit8BU+qGwnnmGsgPVgvNHOALxGGq/kDpNe8BjOOJ9Mf9vpad/3m+MYCRQQvTNhZEh/r
WlPe3E15Fdc4zMSHK9O/lHTQu8L2x6vash6HxpfE5/nKo9jWROvRfRddMtirM/iqPitwtTpkrV9N
kdjGTszlltM+EHtmcsBkig422pVuLm+gWcZ0asMcxmqyoMEm6gToSJz92w3epEJZtDbkPc+D2sBS
P6/i4fFxvH9YZq+9kq6cZKdqpgr94bIfuEPTdFhALEnb32l5SdlUnZF9TweO8AKFXjzSoVMdJUu1
rrTsMNmIDML+VjEj+sgARR5xqDy8xiJYScm5MI6RaDT7u+hpCeITJoh/rh1qhihcUtEnVzOp4HnD
YPjj4IsOyyoTcYqy2YbVb/xxwPd8jl1fdgw4RRu6dBsCmmtDi7XKcml/uBFmlxd/OIBrHtal11v1
FWb+39kufgbyKJ9Glxig59SEYSUQpu3plWg0THJGdDc7mZ7CSgHMbim/0Dg0fJSGwd9LdvjiI9Z0
iBHImiXWUGC3vMpEHvrRJ3NHgsIMBaXhTWSmeJSzEkagFH+FEwx2HE1AYAP+812Lg3XZ/e6Nllz9
lsy4ewzhByV8l7ehp6JgACuZzAfCjBfwQT7IzaRYEO16KeH0sRf/cvvIQ4tnS7u1xvUmJplWqfGY
BaIkHwlNx2n6kj+ckSQ6vMHIngVJSla54hJhfcVusx9fOnq3BHHe2GvDlV/t2pqYXuD1MFubWLLh
Kw2ECI7oZEMvoJjtjXk+GWBmkv8aC26y0zo+Itwu6do9HyeJPcjokbpobn9w4fNS7LcYujyt/XP4
n4qzG8fFHU9xM2MiayrBTBPNEf9TWnucLIAHsPMJ3B6ooP36F3tYWp2kyaEoN2k0l2Bco9lNLcU3
X84i3fENWu9aV1+V8jXpR70yoYjXCPjLsQIWl0LJeMW0xWbPv7umwrpcisdByd/3dkuiEBReNJko
WYC0UN3hr22CFiIPuWnC3t9plKz57PSeGrzz1SS9UAluTx4I1J3+9VA1oPWKNb744JG/5zKZ6wGX
aI916Pb7vJEw+auwOKrxwFZkn7UfQ39nXaO8C/z6aU0R7RzhhZ5T6yORoMM4KmDaZqGkFIvDz8v5
lbgKMw6FtV7C4IXggKhYeCgTHbSoEzmPRnRk70UTRu0ZVv/YjPXsFutIYSV1bp6BXoR6veaJ65Ns
gmluclPPJVs0FuPsYhXidWnPdCr5c4PpX9+bi2kp6kfRcsgDb8Ttrue8LFED+Qv+Q0gumzdZFd4W
g0y5cpGQt59z7MLSgUFMCmYzSAqQBdm8iMkabmRgD67RUDi58ZriLYMrGRcu9nhW3ixaLGJQa6Bp
IJMQLX6eqngBwqzypz+fzG+R184LhLUhnk6L0ySZkMgGdMzVb0c/OR7vXgJWh0FIxDRUQH3D1AjO
sIvu8GtA5+jjEB1lZvJf4AxykN4kZZUID2okgDLYMWKzyR1cioFhJQXSVdeMCWl5/amfnMZpN37h
wj8dn/ag1WCmdD5FxTxc4SMCC28TTlysACmZ46OWhpJ5fyEQwE3FKuheKflqNrGeQdZfX2FyCCoj
aA706hXtUTm7dzMeQG2dzmBrabFVSyeU0FfNsUzid5NgvlMADwB+GOmlwT4Yc5HeK9v6ZMjfhnV7
BgMQSgOljsXpt+pf8wusdtsBMvxkfBZ2UiEDsfHXsHK+sH3EWEcTqzKccAw68MjUp0WxtRKnGXJJ
kXOxZLw7ULlxtjxYsP5To1ao4NdayIU5HRS1vP4FcOnvsbzYwEDoDs9o6ct7U31RORTq4xrwRmCI
G+Lkq46/2ET0YAbPd80dVG7gpPwwdw+OpD+3m9SngnxF4UH69j96j/NlOPqjpREEb2eZ1yCrP7/7
/ZEgxA2FoZ1ZZ6mYRXnAcT2n+OutCmKDAamF8p7GJZmOiBq9zkrrjl+yzDhGqLbp3m/sESEMZ8L1
exxyR0M1cbnmoaU3MaPZuacDAVMsOvomp5Va/8jTsJ6FyCt/hdIyKx0QutwylZZrWyLQKa3KPGTc
QZNGYGJEgyTSG5Jht+v4i90CkQg5j1+itQeuIIfQPlJe78yGeYgsvgnY3guylyBdAByO0mhPRq0d
NOp/IOj7oHCXz7Q3IHgqzeadb7T2EyiOb8gC2g4e08eFyUIEOsQbZdYXf1wbDIOKSjnfObae0qmD
PzE1+2VnVxP0+27JiYDGL1WO1BLCnagGbSLGk0LdRXt1Af2eRdIhvuBOEyuhI6wcDZjwz8TDhdcu
t4VqUomTKouhcUB0bxnAQ/ik4FCRGmo0D7+bUdU4D37ySqTJkZhzKU4LtiXam+xmT7nah9w9VAw8
RfpWkeH2pglYDwidhqYHbCO0goPM8Gz3gFrH0hUT5X3ovQcBsmxNqyr8ZV4ohjgqwDo3NdmYh4Ng
+8QKrYNDKOxZ/MLTqnJq8oDjSVp70oMgR2NyeeI9Dvme84WopSpp691xfXC18edUayPg2GJqKqGP
HZAV4U0Un6CaOaIKhqaYqKM7BIF9N5S6N76Suivr4J6eXYKB01clcMoNKNxna4Ais0RBrKEbQNAF
4RzMkTWw1H60Mw3lcSXGz2gTGUn3EVjF6s7RXrVtBoc5QZQTqRoJA/G4XjK9kX+qTALzrvoWGqpv
08fn+zz0YN39tNChYMdJOROwK0sn31ADwS7lC80BSLSiEFL84qI5qtiBDr1AFMqgMNjL9PYyMxdV
zagHODYaf+Beed7tO3pBdHMp+eG5cjJt8pqm9maA1XcwrpIOk/ZnWan7gCtbWP8DHx2rakiHlXHx
PBaPOulI2JR+53OJNZjnegEv+75PIb3ZzRpz3MrX8jlGvWm1yzTzzEwqmQ/yYp9TjivlN4a0RQov
noVozmXauiSEb7hYcoQsnFNxfv7jhccNUO4wbU6Pxka46UfCOUq8ghts7BdnaZzpqsbIBX3xp2KI
KfH6tAJfUlk+WaHWYUDu3GXvo103ZHk0QcX3m2Gu4+4Sq8V33SPq37vxaUed+o9IJR0MLikn1NZ6
7zPqq3CE7hU4XqJjDYGOJDU3QZ47IimhOsvhbT/UoyzezBm3UMP6AiLv2TD16+bl+2WUA6xasof0
YOIOnO5vY7W96FYfj2aSbNdil13+6MQZuNulUu27kBqBLlRhauYl8kvB6BevwSL3jtcF8sBslrBK
CN9of3tDVJz2znFdSl4i9Fydl86ftEBhflW81jJQ4Ph9kG4BjIhv50jXRSot4PoaWrCxczywfv8d
W2sBB9J8aq84xC4fvhEq/hhhePIW6D3p+E04Bd1fNJgvAKlRBwkALhr/satRermDKI2WOhmfGsPe
ybQxq1/VpPNkDvjBO97GYQ+wNDG5q4J5FgfMmS7iPxgshSC4VjI1w0nzCOMX2EWYft114STKOobO
uPyOUn9PNO32iUn5Yaxv9jRsB97bumyHO5H+kVB9JGTkgk6zYrBIOpR2LbVUmBLOOATo/25fDY0E
DE8+pYdVdYEf1imDP0pfqTAHxA17xYEZ+5W/iSeMA9BbNMx9aqOC75bbETr0z1fdUOkRSJw+o/Cm
DB6wKvFkStqbbfrQ+uxNlZ6f3fzvl9ReACleBPVT1z4kG/zF7FXo7/2fc4CxGMPjrknz2O2zb5Ur
06fNPbw61YG378mJg1OVwWLTaZHS/cUwFBndsh+rKWbSF2OzJMSdcgj4Q6rrQmw5L81KUTYJsU9b
4sk2k3UJSZONdX5+JdI2aMNfjFAzKApyQtXpBvklfFLOXdP8IL7JBEjGp5Bq9B59qGotMPpFEVwC
lpTUIMAUkaKzCac/uKmEtDtocWwyWK5VR3UItVTd4aabEWg6oYZA9AqvyCiVyIX7BNOuFHOP5w9a
qYxF55rkiOnC3hhdQhEENjdMBoQKPgwI4odQTBRQ3bn+sDVtL2e+mHvfIOSxTi2x7hrlZttkE1s1
+g3HGmtrVKfm8Jw3AmGK3S2nO/UPXypnNbVzkMstEVwtEeCIa9yQJSCfyd/nhGnRUf2+AZPi1zp9
HVlqYU8x+nWgajOMKZyDoK+8cgCIH7j+9dLRnvU2lNEsCBeljL8SbPlYS7MSAtXn36wYuJionYO7
fVSFhuuWKBK9axDeuUKsWAON6vahm5mV84zru7LX75WT2hGjU2SOiC/GwTu5mQtGZQojoWdbafDC
3JGrdVY/ghhV9w0+EmGXb+IqXrjbj5I4aBBrvRno7DK2PNdcLRN6B+1hlBd6bYVQlkyQOd1USKhL
mPBidbblD6cEv2oua5DQP9LegJ77xlOwCeUP/+0hhI0ztlKZdvj/ZvsXZBgbHiHi31xHk9QLGUu0
gyrfcR6olnaCdF5aovyJmgceZoNDHbK3IBqZMZ0M6u087Yn973Ux3lycZ/UOMNTE82LfJ2SAzz2Y
t4cEYpl/v9bUOtVyXUW17BIsxD1yIlqxwbEJfDIqJUcZBt7P2NWCHH/rAl00IP1tUtQ0po4WIvsa
b6c1XBi8EmAbyQRMUPvN0xKFTniPipoX3UE1YWjjP5bTdI2G0XA5f+BxXTqDnnRhkSkL6WG1ggiN
gjZNwFgoGvBFh/SSiFWmZMFYJmikq+hZl0crv1/kM7Du17pKArvKDXRvRvADhZ8JkI7E4k8go0+F
GTAg1FJ3iw7QrV/4x9PCAbLL4BL5pjJ37W4ZlyMdaBtftAqokQrQou/VC+6aZ68/OhQh9k/hygPp
EydDQLdEic23q7Auuhov00UQBKM7UvY2yTDTNGGz3vQMjiDoPl5FBh5uNviH61ENO4zVtef9IT/5
YZ4+1MLf7Am1GcthDiTfcRZJLWHntp1KiRb0QnXb/c85FAkNnTxIxycDFLqfsfCrAKLZETUB5dTn
4gvzYw4vVu501lgHF1ytD1wQ78GAm80CPAdgMMaxDZXzhKALc0nMbjwdaXwgDF07gPHDuhRnkSgD
fKRIpsATrJf1JTO+RxpXwdE2Gm3GS7KV8TeJ2lyoapulRftLr5FEfe2akutPgJ5X6sf2UkpdUImf
LRPq4OpeptcE5VzI5VK5Lgd02CmaLNBeVUBu34fmpXt4hm4JFxQLReJSEUtKsJeSClgVrKXMNwCG
w8W6DGkDvUbQ7fu7FLbl9RuYHDXixlj1kQAxln0aL8o45SNc9yzr/v9JuDZlo/cIMeSM7tgX/mxM
b89bs7GA2uDrryeus4ly1m78nSdnhE36hDzpW/LYdbcAvWNh9gQTauYzucHLoHMiiTRGXxBmalA3
ewaNB4ftbgMhAsnadTJpGKaSjSxgq047huKaP6MxmorFRQ1ZXtsrHnItW6bIFkWz/u4LUetECCmo
HrCQ+N4leurMamp3/bzIu6923LETUaikfiVw3LbtND9gW5l9W8RtMkCWl5bMbWzrStDCOV2tDlQH
82M0+Ccb2IPHdZDKVsBUEC43O98o7GSo9ce4oLDWE96qOBQApNWcTzgq/61p7dnC3F1Si8PPIfU9
epJuUBBFQEl5vzhIv+yzTBCBEJfV0lpKIbYfG+uvepslNQQSYCEvqTP/kZCidafjIfSbwn67hc+f
DJxFTR1nW5ge+5oMXwc+QvyXE0UL02SLN9dFvM95Hm/hY9eM5J3iviVgSoSRHbWV2FHjsK5zpJWM
IQvuYrPDNPqxY63VKDG/NEtddDSfWGYpcLTNsVpzLi1Uh0QlghRsochapr8jQciqIDrvUaluebRu
1EeMcvQxPd8vHGDrdH1z8dCEW5CGeIz9hYp9z6I+vvVuaD2LLo0vcJHbHW0mwKHclLySsfy93S6p
ghTqwNhYcss4fVGX9lN3Nr/dZ2q+N4pyfvOklQoMVWy7eMjbtLDMxHOIadLn6fiJQHufH8xPtzgA
nk7NJg19q2ACiyTBKFuUoErVG1FMyUxiUmDivUizhOnfL3XghG21A26Y22uBgKDyf3Wq3nJFTNoq
FJdKKtCiTnfRZWpGKzd5wTrzgSep+Uz3aHMdXnYKuD9daeby3itEc9TILdVk1Jg0HFjRcWl8lyhv
4FEjcz5JeIfpgdCzAQuQaeMs+BEtG4cdrTToiRZMypFZt9iPcypCDMNv/GLa+em1nmEhCY/L4BqF
qsqM2J70nRNwAJln7GstxmTRFD41lnb7dc/S5rPWautK3rMmID9A7qJ4PNDk5ibSK6eEvRJcPFWK
CI3/MUzJcEIgYVRKKDdguaMdHZsdtihoIbBGIikkGZvjQ+EdCMW4hpbuc7CYS6YEEkoeOccf8tjF
w3JV54HTsi6SvS9paiH2u8gIIgABdzwDcdZNsNnp4AS7SbwoVX1U3MFIMPo8IAE6aktwaB3ctFSg
E/31a6l6XuktrXqXzKeMmrAMOwcRkgA1MYwOMnPK49IYhPgsc+/6DsqaSJPgbsTMDm9TeHWm6DGI
Xd1kSPvybNN+4PZUm1b5ZleZjpC30uwZqoD24ZNbphX+tAD9c89CXnH3jpk8prRqupM8dowH1Qin
cbiQODjGlypY23Rhwkb1BJo6VAgisVq3Ouxx5pDf70Ft9fhDdBLVvXbkCWlfUG8NENfRSHi39fZm
AjPeDHNP9PtxWJLYmrBM0D+NlsEv/m91+NBbHVh5N0TmSsleGcolryYboaHueEbW/eIf/5Gc4jMA
O7hWjHmKYWs2/OyblM1n5u0P/xpI7w7cTL28mdG+c1OfG6+PmUfd5IYGnSlDm20U6VdDJrXPNOuj
69ejdh049wuItF7EXGIfbBAdd5fu6kAJywidr/WrUxCdDn+0P1D4eI2dPUWL6Ysf+G8D5ts73di1
IbEqqL+6h1DUTeWrMFBeBPTM57UVCXWQMCJYVDMz6gZPIT0ygnMPGQLyVGYgrNy+9T02o4R/wlJe
l8GQvQEcXwAoPHyUjZadSntCBTpjWTKwWhAGjqcR9qLCLDeGSI4f2ogx9lR7QCV/66FS19nzMmVs
SWgp9m7n+1i93xu1dvztGC5LD1pMbIrbrnJIsFfgg4Km49J7QJu/ZMEsIPfJvyehkLNwi5rGbMQI
dZaucQCn64vx4WKMdWkcQrXidhFJQ8lCH5a4IBUDcde5zMUCrW/KsApHykRn0XURtniy9nmgeGeD
vgYjBglF1GI/GY6C8+MJEXGpEtvpnWkImzj2GagYNoaeF8577Y3VqjaqZZh7pAddxkAbifhXsfuT
CHFi1p3lmGH8b60jbuzVH3WR2PElkOXxAZW2/AKfQ2GxsXlpCDVSxLa2w5eFuCqtPETKYA/j6RjJ
qQJjG1DqRWdHl0MaegoUtNp0P6+1HqqTlxpSNHNH6+97D7B1RrGkRzDehnzIOjv2VFATpecGdtS/
eavIyH8+st2/cURH+aEJhulkXsjGK+m6JuDV/9qPmYbaBE68MY5+dzfZizXQcfbAmQZN5U1JEShQ
BTp/a25azc9kTKIfzA6gFskykjZbZI0hlbm8QaACe0J9eO9BLABPIzbRXCvSzDAF77dt33oZ8ERn
+h8rxpKkAy1ybpWxpRt2EBt8xHAl4L667FliDV8Tr1gTiymSjvk6tyCGgHekWh1eA11uHAIIBKnd
qdEJLxyFEXbbdcpLLZc4o7ZyqiLR3CI073DQwTBV0zNRb4HhAeZ2Q9GbHj3aOOa0Tr5VkqbpxbzG
NaCTs331ufFtau8jF3KNX3Od/XBX+z52HBZh2IDjtekw1Sofkkkagc24kIBwtJXPuZWyFHtQX7nF
+aF9Q/k66w8ETDaG5N+q3qUGbE+z9s55766WLD++hBEgPWFgufniKN5A8LjghGF1mJxXKLQFjbqV
u8kwYxQdENmaqu5dUsyEF5JBerHKBf0X4XOsR1LAIhefKS0dIuDgHY8RYZ+Mg4qpPcF4nXlzNjc1
QZFI6ykDo6GW4ZpJN+dMU3BhC/gqo66j+dqla++g5677LFL2qRSQOLNEyTOcvRLIXNdk3JmkO3+h
c8P0sv5Dgc3kFAMOk0ZMRLTkkKaNAS8Cnth/CahQej/eWvr7kg1OfIPfMe6oi8jrgsiooaiKgFCD
KlvFiF09R/brpxQFo56AWXj3ZaJUdHVlk6eUk4kkGQlYWcZ1JcuuKR4TCt/Il4d7vRljkFDDziLQ
87LLMznAkmIYVllifRpIzILTLSDj/x2qiO0l215v3NwD2wHpAWA0DyPlPM6E/3VdyT0cCBM7Yh/2
am/xexQBP1XnD7HxsPr1limX0CVTzvPPeu1E9zpWEewUDLfC8GiAZf+fxM/2W2KPKmo6f2+3b72m
dZxL6CNxkzHoOWtuzjEm8l60IJ2rY5Ns0BQ25+W1zZmDaB4vqFAxC6YEaOfIOx+jqzMFw1RfW/Nm
K4Eq+qf2Sfz+XOPAr4rIGxCiALt8quKcGwTCb7lt0Pkts6BsZPUTNgUGpKahHBQM3iWrC+aYEgrY
KRVKFGSvI7Mzblyifqx3vyFLtCJEKyRTLFE+utWb9inDNbBmf1EIj/mIdVDnoB7aa0KD1hZ0aGKF
RdIL4Qstonu/rTu9Gk10khP5taF3GoR36lfyb3uNp2Skix+GkSyfIoYozOrbd9I/w6B46F/E/+z9
ukVzYpxocH8NRyADaCQqVUAwEtwC8HKJ9ipUFgSjRK7gbj+a9Q9uwNz3mfKS7KY2diQgcu4jBCjw
tnVT+U/kF44JjAOyzgT14mU68PNuQ/GFzqkcQR2nlTHbCRF5BkEOplXWb3pW6RmP79UCYgaXCMHM
P8EZVHYnlktpJ2BGSyP22iFb7Xz3NbO4qIt9EzbYJZ2+BpbDuYLXqrUvDGqOrxeA26n9df25M4rH
R8t6kqhcnOkIXXi8sNX1vprSs4z2r2Jq3WR7ZEE1DYQkjS44uXSSNb8IjoA6yJ7TRX32iBVpBis1
xV7xTn0flPBXFt2wJsf1S1d0ftFpIz4maGSrohOAQ8hQJqS2vBheulpBa7dHPYBbJu4IIQK9e6sI
aCyLqUAKZ1nxLTKVSs7eIruVZzRfsD9tC9rR+iBXn0bdvDDXQfUDwGiWDSFmFgijca0TsCicjog2
XNWiaQ/AX5q5TtzwlqY1gdZNqhn9g6W3OkUI7wTiYSTLnxpygUoXzkSC5FYyGkHbkl3Wr6hYSy8l
TBymX7kuxkBkzGvtLXXMpuDDdcSDFKoTHRWrYQzRSo11L1KfHacB7m9H0rujt7SIIqe4H1SZ/7xy
D5T4iGiIeeLZ/sHS2bLTueQ4YVUhcqvBsOx/3+52kbEE0agx3/heB7qc4EiVNG9dR31Xidsk/P2O
5hqWi5vhiSzNhODLbiHMND/afx5rFMPiuA6OOV/jPLYL8IwdA8pAdGtT+N3ef0PyufMoo+yVEN0r
8lv6RTZcu8t7Daa5XZ/INhj2lFSUxR18AsoOzVDqPCv8qgOznurjGj7XP+BFh2an9p8IBvsRwqaC
TXqv1yk7aQ+ec5UiTH+oKll7pdY83oDFfX0ePBkiye4qfiXA8f3eOo6Oi6R3020aIDG60gs7l+Lk
kpWYpwU8qjLu3/96zAmBwac9nk2mFd7maGmw/zt0yLQYqeU7Xb7NSioPE7hpkpZa9wsajs2uFYHD
61SfYfoHYH3e388Ky3MXB6oqahIhT4UOLExhD7H79O6OK7VaMbxXJXw/bwAyrxeW23ZKQLoodkAC
mUIIvKRGL43g7r6qM7dgVfMvc4pjVrr1hWsIE6jawbvrEzS8x0036vVDleUtARwxMa3TT14PnmfM
1vxi7Mbmqg3wvntspORCwqrdcz4TkjlZp/0ueFgahZDfnwzN1449SF0SR6wM9VcMpLSjzNzl6VCo
D8Atlj1MQFLsJ/SlzlZ2jm4jKt9/roOxDEoDzhXzOglJJlP27jrLsYDjPc3zH3POZhKY07Jj1Gcp
AVHYubxBLUF6AH1nJwtIJj5oeiC6/HOPXhQu9B/AcWSPqiVIfD/Rj3+yXhHzzX9iv1TfH9LqRM02
59e8LoDkXEIHh15+NVXt64J4NXv8mwrw8Y1aHmbpe4BNDyLkVC7nWjdCpvgclYD73jpnMNy35ukT
3XfLhVkpNFSBiIB7mauNCIzjTaFbZxrR5+PG6WJw2ruya5gH3dzryxuz8chy/PHosJDVlBgaGpGF
PL7E7sm7IZ/+t2PQK8WD2Ag2x7gV8oqVRXD/Bi0d2OmoN2RrcFMVEhDMLgXO5DkDw56ZlWJx2Ie7
Grv9fRmL68oP4Pnn0Y8Er5QiO3b1RLN+t6t09TUTeUZc8sri+2aLGzP8en5AFtDheM1EZSx2ioYY
DrQDdibGMaOPFiPQ2e0GMLVPeUbIsYtrhFXLd6KrOY5vejQWPpu//TWAHtz5eh0RAt7vpf2LoVfl
DBm/SW/i6kU0WHuwiaunwE4QfXeQ71I6g1eBnxPNDt94920kz+RX6SVhAgr61stXtFe2FgzyR7Sk
Q9eFKBdl1PjAXuLxwhNvN8tDD1Qihy9fv7DSXP6vKi5wAXgfkVRf+DgcR7PDUsUCB8RTYkWjPIkK
ZtXAj4cQmM22P1fiAlk2iFufHI9XOTHKDOg2AW1Eni4SzUq+mfcsRBVH9QlUf1XWOsb7h343UPTu
/SUtzi9dOX/g51Dg2FDtPbpUtQbH84x57V8PCyjD8/fDggThv0nt9G7bfJ/0GfYspCdDWE8lsu1y
zImPUJblQwNcRaBbV9VjQ4c3ctHwdRD4FSQnYyf2VDNsoMXgNhjHnsN308g9RS4W7Qi9DhqfNV4V
YQh2siVZzyak3oa4NPZFL1p0mFFuqaoBomho7SPX9ltaqGfcj7q+NO+t71PpyA5YRYI3d1WF94iR
WpRPDOruNqH6VeujE2d2Gk8mKBpWmVVPMjAN/Y5pbvHwOTF+YmcATAVp+hlA00hmpFG0G3jiuhpz
IOvzfE1IVhQhdVFJBibrJboC82w8onMdpKvyP/2y4U9xZV8STVzp+AQaZH+kEj7Lxxo04bma8Noj
r7dKPWzDeVywMpyfBB/n0QscjszTg7wlSawiGkMcD2McBnQdVhV4PIDPUeNg5ya98c8KIPsDmJPq
WzKJx0abYVt/zoUTMWNMRnt2+hoxkgrmE8CK6xhegeqr6D/pTPf7aKNVpgg8CXo4EaHXxJIX4gg3
4qJIKWpFgGmwpmF6SemlZUX+Fy2gnyiIUzQdCA/C1QYEGa4ltq9J4cM//Pa0bbO2rVXB/SkONB7G
RPVi2ozX0sZtypOO9hLJx3pc78MPOKKB5VYSlYiQ04VHxsDP+CcmY5LpWN7NiHXrbSxTt2AFxZfC
c+BroyCUXQVaWO4zrl2IZd/7x3yL0pr/V87Nkjf2MxbQ69/M/4F8IxJzD7LeSYtBJ87qnzaWPviU
9NpYpPhJ01Xw0M3xMaOFo1sGVi67kyvyMUlI8HY+YYOPBrV/viTqjV4JozCZNMyVdbq3oQkuck2D
Vgc9Ae2aHD8Fanm6T1RxfE9w7OC4sW74Zeok/tcvq9D0nouNDLYYeU2rdYdWFjq7XS9cPgtPtMkG
z0sjk6FCIWoWXKY4ZFRgxzztUC/ONpQVg0OSBYslLLqSFBEwU/Xl+x3hPYDiSMLGAPwM4avInQEx
PSgrMYQl1eXWt2iW2gi4G2UDTSSnKC+xzXQxchZowtJZziCQPBkhIYN4yKg2JEmRfibor+IXtckM
BsRmyxI9KFdUIg7gakjlEOdubRqZqUgxOpvn9+jxnZJg8T1tQceHJUpzezYwi5EnrjD3Xz1vdZbZ
I4NXduQMGGWYVD9HzMb4n5LPfs8TtUztXO14t65yuUgLHOZxVriowAdzH5B3/3ntW/0HaHGseDva
U16Rt9l9SeQO7dYSdQ7abDyklSiPLnIFJNwjydKB+gbMpega58Alwyiov/xsDxkFScSM7XfC85Xq
U8I9w7MX6Ca9843VvHpzFxoh5YMhEBDeZQYR/XSTsGjnfTvaDARbfaOeU5GaKpeFgAkaZDk/D1IO
JkBKMlQog7VNJPhr8pv1diPHP6YMF9t1BgfSnN4RX1suLPAZY2fnL0CbCqSdykPyhI1JdEJwvTO1
tZ8TmQqMtXle1k6WEEpIaLNpt89CkehmzrjXMSawn0RJtpDMCg4l2rK5l/St17cGer3JSqmiK0VG
+Wq/v4Epzlr9k2QyxX+b93aI3CaffjHIqmLFmi+Uz3vVSgo3FTjPquEXU0NLW49DHhqR7TeIC/Ss
gOIXxn0X4WpYEcYnzxa8bBvJK/aLv1NW5RfYrtXr7G8RnjfGwjJG8GPQUKblfW82kK+kE2InpWuk
rMaJOiUedWMFMR4VzLGVsIDIZ4qivmiXN6q3YBuHgJfQtllvQfaAOD/5kEa+56xjJk1d8shPxpAy
uR8uOQ/TYpsfMXYk4Z9Cran0h1qLLJ5kjNLUdymDv9K+r1eead2xugu3oYIPCk1uZv/FZaaYGwme
wCimE69SI17uFfxCIECzpcuENRuVb5Jake6HSHBUKG0DHoPs0Zybs91jyfGIOvNpWxyUdM0RQ1X0
N6HpJ/YM0dK5S54XAN8BoZ330Zh/y35RpaEzgF/MnSf9cJ6R2D+n2nqxnlz50I859z/9lqw9SCJ7
11cbpwpiloGwtzKJTgLH3040dQYKNFC1eL91fIzw7u1q2CDu66mckAZ+WdRyZ/MZmadx7HoYNbeZ
3Xuth8IMdrdbNvRM1/BDktmwDVbOnTAdbgIICwnnpDtS7uQGkIsqaarKoTORi0eeVHb4XsonSIqv
CGkdvrM1bLO3Z7Itk8nUXMnSzL7wazMh2JUXyMEf8M8YWvo8UyE7VwzBv4X5gdB7QGPLy1q7PQyd
llF1sBETf3vf1BFubFcrg3kaI+zLA5U8tWz2fOXvwE7LEEBcmcjC96r8dIK1ZAomAWfAO8y1CmDv
XL4aSafEQVGhTxXeDtPFOs8XdruX3Q58doEzM1ctN4yYfSLpIRmHg+e6/JldDHJatpzPBrNq73vO
1ux2ZgBDdbxVVUq4QHmmvZlJO1DDYmxQoUjR4Ck53PykXfUsnmtu3e0uF7rgEMBTY7ZPZ0V/J1Qo
hszg6Huyh94Qf5zWe/YCPEjHc3gyS+Pp6T0j5gAmcftzeo48h4RmWxmcEJTBgRGw0zlZbBg+N2lC
vWKhfeb7XujeKySxHsz8dsJRJH9q3WV1jWOJrdVwlMjj/mx5B2okeKki8U0JJvii29gh7XLWaugM
0df7wERrefm6JtWHFQEm7nA7m8VDyMJ8Cb15KSE1e/fCNQp8f5KXKBuHtGyY2fuexs5KEcCbIzPe
DX7/Lqwz2H1pTwmveYcJ434GhMCeuE1iKWOk3fo9quN7EnCr2V83uson8byI/JMl2Vk2+K6RA+LG
5qLWD8Oss9XdG8Qoc3PHIvVq24imUpmK/SBwYHnn5sZ/nFD/Z4zGOIP2IDFt+PyAg6gQDq1h0BfC
/WtSVItka0JK18p5UGn7de5XQeWrF0okkTaiwHOHlhjjS4Nd3ribqPEuRCkpaU0hfe5sX2yyHWEc
B4tJp2/v2YhE+z49C3PvSMz/IvtOBh/Z7kmbceJGl53h1p5Q7xxLAVDvQovbrEWZNGW80tesavcx
9J9pAwwf+/eI8t1Lv3c+FttDXhJRn3TlzXpsItmIiKN7U7HLqv+hxkGx/w3fyZfooQMjim5uhqhV
931opGWmhQ8Ol0rODp8kW2RruWJxAze2pI8hyrGKyABvdFi4ubv3wCs0xs2P1uiG937Egz94PJha
I6TnIFwicUMccprZrKdpTC+LavybndJdBeimQx9ogFw3KGWomU+ISxxLtDhKD0HFFOfdPMMqaTD4
FsGIdFmEeVRyqPZdV9d0hwOpSw8ohwN7bKmcsGmkT+90dZaBFgu7j0cOJ1Lauk7N62G/MdZnwAfk
RGbFu9o+aygJ2ZO8RlXAXBUu/lc5OZMWVyMilIi7Xm3fMWdFKBBehvP8X+ZaHm7d8JO+mhOZ4tan
Tcc/gMbLucxip2wf7V1TqWLF7xBQ9YuJpqDJ4rqDRYrTy6QtXW/VlfqBC+CgHcT7D15Naj1HIg62
PgaqY8Zs7Goielnpj5YKXl1ClwRp0ijwpCaQxnVtmjbZ0YsW/SmYQ1kM5yjkQkZY1+RQVqYzU3vx
BkBN7kTLEv14st3Q+yMX7QUf0rWKf/L1GMSGHPxi7UVJJyuDynr+3AGxHeZY/PdClCQY374em0f2
HqNDwA+06u/W+zg8QQaEEfew5HSJyPCak3xWZ5HetsQ4LOMeZ56dS4vLh9sz3o7jxBrWEqbMQfvd
aXUxbW9BSu65ojbwc9tUTeXaor+GvSJiCI6Gjk2H2Dl5mISHhVPsxsDnxkWb83CZWjNhH+8igds2
geZFtXMNk6WkGdfcpBxlyc5GJD7u8M5QsyXVNpAP8JE1hp+iFTiKOYDxAl1vqStNpXStTkSjyLWl
H8QH9gk2EbfiZRJgXH3oTWByQ2nl6V9L3EbEJE9kkmWCAIIWn347XQVcq/jzgva9GZsF95OzcFpa
hZOYUcKOqpKbUCGYKk2XKZBP+ZAiuWHe8/9YwI7xsG3csPrG8AhIaXgCfITTuT3eo7phosxr67Wj
rysRpGQX/kThqSaGMZDnjRC0aA9KjzPL/tp0Af1tDp4LpGDQEK3rnJV7FYIh6/K3UHkygT1ctq+E
7jFQR0QksO/AlFoYQ8275WkQJCde5YoEz0WAi9NVCna2KEc4luUI/CAWp43JiPA3pl7Er9BBp2ha
X7+lASmLTHkccqpwUrCsskfHuS0qZg90A9iJrR505gs0FwjGmdq6C5+nwqOKVT13bYozCQfvKE6V
/wLw9DyRnhmBYdv+flIKlR9QetIYjNkgOR8olYWILJSSOpA5ibVHeDCWGJiCaKd8i0OhsdBw8cik
a41UiixFT69P2lfsRw9S1Rhw2N2U5NQgnvDOlG75b+aqTsEJWdz+pTDEG6vn0H4Sveu+ZXzfemgH
pO2jdQqYUOwNdEZ10AZjr8HJ8vMSFrRXrBS7k2RpXtsx58/+lIftph418LmxtwcJCdi7s9Mej/Pm
MV+4285NI4sAJkU9Z6oIppEddBr1MuaAJey6WWPuBf/Xd+beinRPdq0qcDpEylDNTXCLRa4A6p82
7LKwR3JWpsb+4er8b/jyYhu9lR+XZbBFAlBCuykcK1ezHPLbIaHzVFM3tF++UJNjBwZ347aGT2mK
op78iFBRbEgs02U9NG8guYwZCzlK2Dd5Yo5nHshIZlcYOjNH3/+wABbsMgl130KiB3l3BjK+ni+B
FhspUs2GJXCRc1mbfpvb1TVCy95EhXvl72mfdXxaA0MdJiNwu9JvY5aF5x2ojmilNuGaHFP1eQGq
OuDckzloQYPwWUpOoCMw/c90l1kg+5F3EVcjb5mL96tv6SIBocIMzeItcOAtUNK9ldfuTIdYRB+C
kU2qCfz1f8Ipjb86RKIpAojfqAuQp6HV2AToAhXy6nilX2CC/qgwPRslE4qWES9VYzyuExgFIFpi
dY9r5oR32UBOHTwB+gdJ40tJxFQI+OE9Prdhe6jTdQCmutq6dj0sakBufHKhwufvOtPiQQzJfm/W
QP+c8b0ZmlK7CGyZ4s9+/ygpgNxbKZjxm4RUEfCC0jVULKSzohR/h8H+NsYnRh8SUZaqgRwlXZsJ
nmtuIw5Gzs1ZyUob/OGYPTPl4dfxrXFP3Dx5Dk41VRx98hdBNkPjubb49Tf9PKjd+gMOByVPuOEr
nRS8Hnck3lOmyY5buWDMIjUyU0FvpGEMx/5SkMMIqg0M5fUHaGwitFsTu5TA0oEM+tNZYS5TtMiF
WHy32PXoUDA4mMsu63NZygwKJJST9OD31rjp193UEpE6YQiOlf0MEqUW+QfAOjUsdn6jtKmOr0JN
d+5VAYyCv1I0KhW1pryTUHAZI8uFUgIqzCsV1VXR2M1HmEubGFbEpTodjhT2FOODn21e/XHHwjc4
ekbfSW0ABdfxVGSW4wU8/8pgCfuRZJNYYhunHg6M+8piQn4TSSSl0mL2ZCsG6xQswwFHf0j8pSKc
CVe8HlIVuTj9VZWgtCJKW19hU4Hgm4qo1p6wQ7BHkn38y0zcv+EpNhjKvR5BwDJCXN7qxMST5zoe
v6EucRXIWs/cx9QzHTX3EisEkL3OcnO6u/dTAH7mIUz3MF3/gK5nBsubYCmVl2fhcYBwP9UdWXqU
ctJeto7itPA5hWj5yJOcMOjg0eBXtyZMUutjDnmor90zSG7ryAPMnmyF3Aw54NxavcCWiVx5dQPf
98oyWWCrnmAoeAkjBjhPWWq9WQsKbhOhcge7NurXpKSGSYnaH0u5mNuYhK6EBGxz4CP9VBlt16PG
racDwtA5WVUxkkLwqfgjyb8LmxHUCB88rbjxfYhTotUSvCmWnW/QN6fcmIZQcaL1OPzxqTcr1tZv
QhWO1MDuVLWu5Dw4YZxPn6DreSNowCgvKyNdgd+8puxH4jv9r9gXa5zJMomHF9i+BSpsxsVhq1wc
x6bubkXzZX2Kvt4W2U3xFc/r21i2EJSxNV/+GSkK3QCbrGA85ecPBScR6GWOjkparyziht+1USuj
KO+Y8+B/kZ/zf0tb0Uhh57CV2+wgDs/YPapeEGuLHE8Z+Fk4s5lE5O04i3K1ptCEtLtyIb4JIi1Z
KYBvAGqcUAnO9cqwCTgMt91Df1DD/P8IvLrm6h6Oe5bAmHOHFXsv+dO+xsldXzERoFGel048Mbxf
fXWwLHAx3Xx/tp6k+VnEMtDgexyHYJv2aO01bxJBmlQtzYStTqOINlg1g/OYjwCRQ0AP+HGsPiFP
pKmacacOdA8vSDnSDv4fzd1oL9MVFLcEN0RuVJIUQb0dpvCygbJjR5kW2EhhifXOM09Sx7LOSEzt
B57Rto6uBS7KC3Vv9eCC6nVBKU+vefksm3cHqfK5HIjAhUVXYBto0Wj1/1oSUhaDUTp9OHsDcU1o
nb46N03oEI0NSsS/ct0uRuYHJLs7hGl/x9uthXpLa5hwsmmkRj3Q5hd/KvOa0hXQv+oD1g5s0AL9
JJ5Nn+Kwg3i7/1azasZnQ9IvqC+kodNZ8c5GhusJac009wRryHeKE4Ao/2Qiaef2NJTMJWeP64GR
Jc67i9tzJvEQqDV5Hhs3Av/EP0lh+eXXmHFH6OXarPwbp5uls4kezQNgRKOUrtVBjv81Gu53cm4m
bIIVI+kT1Kxc3DgWwChk3V3obXr9P9oIkBjUmOX8TayZM8YDijBjeY2mEBk1uJcmYtvf3RytSYmM
+/l8+Wa4ympOnkhuzMvXrOmYBU2zLCgPl1jjEqBHKaMU+MuKfpQbU+24AIG+HPm7XjW1kTcFjN7F
kJkqmHvpVIlNEhmMDI/N31I50Xbwt8Vn7299h9FKNhXiZspYAGRIMUav3dIWngranmo6xKgFTP9K
vLgX4G4L+6Fs4XemliMhpxEOExEnZE7TozBH87qA6xflC87vhAfNoLaYCj7AOIA2Sb3AlwN4iq5g
Hn5lYHE/2MSgq1xFEcfmQHB/oeIHglZ5R239UH5lC91NeE1hr76BX6HbOrD+Zm2RjXCJihOX9kNW
gMrWnaiTNIyo8TO9tD7odGqkm/5lEO+9ra6ncl9Je1lqcLBAvbeGkPUW0gLwrf9ELr9I466uUiA8
CpAWt+2Gqw9ly2yGwmI9GcTPzBEcqYU/6M/6VK3RZQ2WiTK25ZrINJ9dk8xpmlf7rB3nER6s1wyb
8jfL15Enc3zgKkxPHZ5zQ1KmdXcls53R4gY16D9YZs7wsHnlhP/atbYyi+z03t+Q65GNS9mMtsge
3Wg/p/6HG1+deKLEEep0IDjHm5dhUpPjOlrKCNDQDx9ooHLLqbgWrAJ93qX6IdQNQh7jdIkmhbHY
OFdpDh4ITAJ6Gdwsj5PT70ffR29SxN2ayaZppCOtu57JAk9MEXei2CroVdRbeTVOjYFLIVdTUyZk
Fm/S2J3id6vQMOffBgv2sQKUdw8z2p7PSrolmy8gVtABdDiRRlcyWCeCShDawmFBQflzoJ/z4t70
jmohDMdfcV3BGsGRH6upeCmXIkHTf9NifbgmyLlv1NwyTeBVzkjKTK97XiKI8ArnqCM60h+8FU95
V8z2HLDbvqkCTcZtgj+wbBZBo+8Q2QbKuXxkn2zKRFhAs2UdEhF+kV1Y11YfGOO5D+HAcZO3zoUV
27rFwFY95Rl+9gLcHky4ojrN/OtHt1lTY4BWMUxABZEEIlbdHREpR2QKd0O3qiVJ+O0KMtRzOhJ7
mva6UKxZwaKgmrnay5XnvYee5ojONLWy5X4NH4EB/9XmSOnRfSdjTnDmdOCY9Ovk3Htb5SeoMbK6
frGwNf9H7fmQKds1bbqGAs1AYqtdVw0BGyFuYow/AvYAyslPltAE6/w6NLAE5cg3EcD4mD9NWLFI
j4bmtM1hCsUJJRj3V8HvPhOsy9FsqQFClcjxOIabAoIl80Jrz6QcnLkry9vpCpX4SzN2WkD7q+nb
tV8z/oIqRJ/l/gTTDBL+3UKIG9bx2Tsvgcs8H3pmFtDtMtVFx5X2TuuJxcDkOmMFguixUow4Ucn3
mJExZ3Qs86EeOvWb2gFBQ80Vh/fmg0SFXintJvZfFnsL2pijlZjDCHVQLg+/Eb/SEHB5tq/4FJDn
kIO2XX1vjq8TAsAi8juvxeRjt9zQCFloUVYqt5hyvIa4qotVtEf6hw7qvIkls8m1j9yDfUkKnepJ
nK+lE+xUIUlnQz/t4ypnZYGOf6vh2WHyxaayEUyHKvISX/0ReoIx8GNL0fcSJUvYrFxFDhB8s2tB
5IAYAc72KVsXXlp3y58oiNdC474ohZI5EkwccpCiMGrEMeCwdUR20aU0nWIIEy9tTf1un35ROqE6
omwEVMDqPro2YhdO7s7KVzhl/NiAz0LI2kW/a8kAe2wCtMXMvTOiG8QoQqQ9H5+L7CcIScU3bSYG
/iRYinBdg34PPD5Uzgto3nSbKIW/ZmUN2GeB5s6w9v4sowfhSzygH78gbVeyffEWS+4z0E57EpD7
/z1yBhiaBJAnGiu0P8HfTNbFdPbuYA/jwuLvrnjqQeX/Mhv91eDdRJ6hdHYdfm47BftIeTS6RLBh
WwkA6NE3Q3Qe4Dm6FYpXO+afhU6NFU7XGSt90wCOgXdhvPzD5kEZnZQ2131a0lNLJhIC7FnVfwOY
p1f4i8T+QJxTWsLRghbdEPYWUaHFxjo8bqRj0Qx91RVNta+5pke8/cIDHYQb54LNELpVOgQ9zBen
RNiJZRxL4dvq+qZvxI5CAFQWmZQ/NB8xzB4tN8+ptI4mwSvCK/fod6ZJMzbDjntu9fTVrGL3k+Eq
+XFBu5t0BcIgl3UNIDfbSgEgO9MY73QK2EEL6UfeRfYGFnyjXRlO5NH+Wyt68CLeDDACZRO2vF3P
SbIBq0DMXUFUB+nJowarifyIigIk6lObvT2ywX6p8LY60015Tw7e2ZHZtq15E4SAI4raQGklePwd
P6kc43LGcnYI75m6MHTo5IKxBbuaeijrfoCgumfV/D/Ax+7lpfXOKzUFWICtahKvoyVoLtdkARXD
n0a5dJu2llGa8BE0N4STYzANShr2RQx4cKsTHy1xS0XN1xix8wR3VlTJsd1gzn02gjS4Ap6bwMXO
3+IDC7EpHRwUY512a7lrGB/rUyCvo2w9O3uoNcX7Tw92MgapF1LPYycoHO6w8UZdrlve4cFWnWDz
e9SvIWLvyMc2qxBddEhjTEVb4hyQwDz7WH0q5hCzNXNpEdtjYzTxxQi78C+3kj4bDlv/A6TBQsRT
bLh9x3gtg3HEbrBzNaF6Vy9haGrDCIxdpBxDMSmCVBUT7qOzJjm5T8tjmFTtlEOx+TtgtYWtv3aV
3mZC8Wc2txqBBxHVcpHkw3Y9/e3UhONMHcQvVrZBGkd9sICYCgOthp2zxIxnS8Fg3K80JeWosiCg
GAb8C66nPIfJegFWEfiRj2/uznizCyj24LFSyC1H4Cwkst+1FfpODo3KomLkcJxsvlyujzJoZPKV
VBoPVBE7Dtcoc+Y0E1U5405ys1cwz+LiRKudREBxQN9mvEqNosq9pI+wWOkRm4jT/yOvshnMrOy3
cvnVFQg+fumXnIVy8BGngxDaE7wh2LXBGI6h2t+0YaJ7peJibjBTeewng6PgmrvDSdWFupCH7jS7
vdxLzQPD8y5NiwzU6q3kKnGvIL7alKeDk3lKob4+Wxv99NbJftH+cjvqIX9YIIlmpN2HZxyrmg4M
5eXvBj9O9p5SxJdm+WxumYoZASBjXu6MP0Y5fd6Rhi9etpfm8j7KRTMQrT+dXl+q4xbhvJ0AU9+7
dIgl4FV8yAjPnsq2sqQQEZqkSTZuaTOVSrQYVeKZWNUvYiaAOmqnfOOUmr3IBtahU/fqj0ReU6TA
Q2FvycvtL1X4R++5LDntBT0P4EhpzNttgPqxwJYPI37QpIJ+6xckWq+Pn0P/6iGbJmICmr9KUDXZ
kFlL6LQhvw2e2clsoELdvF76oCyjeyuCxLQFs4HKnkpBSGEvxCDfGIJujcKxWGyWGTOHT3zNsjW6
n4av8TOgn1DCa+Z76lmmbupdankrgQiELUlkYm54FdrPByNHJFIjyuz1IiXM43gHRGk3gfwriRm1
W/ipXKxnjC31VT8O5KKlnm6w3epD7RoR119qSRfSBBs0d7e9FPPiJp7MAm0mJrED1ZqzUdxbm+gy
6evMopDY7IoxrCVooZVdx8X2UkYhdm/7wlHSsULCFsfOEiOBHaJcF6/9AB2SZem397G5ax4xb/e5
gzfiTBI8DTn7jaKqIaRi7xBfv2Ic/y92r8chimOpkmCWqr8keYDsb8nbjdyy3rXKUJqiAbzgQS/7
C7B0XBx1I1DDfJrMoMHB7bhFBb6ldqlweobH/C9YdqJdD8Tll1/tZOA6H3wSv+kz6FBNSEpVZO5Z
uYyM+T8Tz7U3ziqsnnjl5Zvr2qASJmLkvqPpjTEKwwOXFZIl9QInu9X4gmbDVpwAicJZLRYTaidL
C7PH/3OAYdRi25w335N3k0ehL2nh0JGyAlqS/0d73JUpz3/ByKZf+xqSiHByv61QHOX7ModMMz7d
8Llw8vimZG42s+ORQdzZeizSlFysjuPA4PXIHBeyvVHY90TLocWABXW776U+2ljjp3GNEW9cjthN
z/eSml4mv3UutoO7jj00NnsNJ0CS9lr7nCRMO1ZtElifavjxkix44AJXrkrDPuwEDQtUWZ6uSccZ
a1li0kyoV7Zfhi7uMOU7gl3RHmWjGsetgXHEmJcZolHMSHgEC76BB+Itt1h47u2QrVDiwWXvKC27
oydc0IQdJhs3QOPLCVURjv9rf9nsPfo61IOurU9idBppYiNpKEQxbV+FV9A4g8prnpZ+Ys9ay6DR
g9xbAwrW/vYdr56vufbdFxaa3b2LdVfv5WHR0dyTuamAWj/qutY/lDqluf9mMhzv9GsHGa9lIEyR
H26kcLGnMf/QbUmbdtDGcHDeHisvB6t0DUo6N3dk57IbFD3LrJ4EpxFoePDbkwe+5/o2cEhVeQVN
z1m4QbJLxWQEUVNTli+lc+xmpBewRLDVa1xqlt0UlTDOrgT0QhqnfjGiv6vve7QwuKpM1sdudrUe
az/b2e1276Why1BTQ2M9hOelgPe14BrWkN6TVgObX22IMHZBXSP+zopYoGhaVv/dI+Blf1nD90se
8Uxc6N+B1eNBL7pINzssUjVfsCV7eaYc7CJTT3vjZ6yy4Zyqz/ACeYw6WPs0uekO3/CGs7lhDoZs
pIp//lDsJdbqqu4rQH1HZnoOF2ZtBeerflT/wNpRgUxC2uvC7S4WB/j5lkhmPEEZrQcZA/EhfcdN
imZbuPSsYrePNmfnT0RziB5ZPF3qEG52EKjB26cAjqCWhoCBic5KWbnQZklak8aij44d2qb3ESwu
YPQEL8UoN2WKgrfcckZQ0Re0YGmHdJ47GuVcnn2AF0+Sgw+XPhhssaRhVxUIdxTebjhjRQ/m52oC
rz8njqG9CSK4T5OUYxtThpkBFzenXqLH4A4iWoy8baY4LLISXz9TKaRU3XhV8afY0ikzR9YGRcp4
Tryik+hXIPNC4HtcaWQnqXB6YGn4dR1YIGaaf8n/kWHCB6Oq1zNNQ2qA5uUKZTiFbL4O0vNsoqb5
nZ713uFhaLpMu5tEShEcxdUCyVHPukUSLaCFgSdK7eLDpX63u5Njdw5jCHzgRHZ6EiVS0vTHGUpq
HVnD7ZGyFA9xl/KBvUrjgbkF0NpHHN4kHWLRM0nzwzBQtByWXgYt4H9l9t/JhEX+cpY8XhdH+i8Q
mfV6Kj5JTGvnul3tGD3FPDvWAg711KovPO78WEd2Mp6FoNofwdpmjqZQvxH8qLFDMT7/vnNG9IOo
vmfOxIuT2xxC9WxTIm5MqYoPKDlS9mahjZ0QEa0wDUFgkMYK/yHIexeskEt6qnno9qxZZkG3IkRT
cWvNUMEfDLQp+Pkds5KNjvrLn3eyXhiUwpsRPyRV3z8e0WqAS79WfRK/1Y+eSU12Bx0qDIJXsFci
jDNIWqc0MUS9V5/r7j1GZ20vqxvrHUEX0pHWvI0HOwqVqewZTQgTRbf12mzD/riIKE1NaE3IIU/B
uiTlrFggpKy0PC4f8fwZ0S45QV03QYLAwG6vPnr3y/M6dcvBGfn7PwMOGI+IX/kes+YnUSpeDeeY
ml24L5rxUmerAd49FUpht8fOBvmb1ruoFghUu43+y5TfmwGFKYTfNJ+atcHZNEyD+RK79O9DW7g9
Vzk/pCAKXl7F46WIvcEdkegy+gyMu6uXYSHruA5RVIsoJiOggrOBqELy2huaC0T31Os9rwKTZa5v
8sQZ7iwng64bTtkwINtYzFtjkCA/v1JLNWW5nfjhs+u4ZZYEA5KPQ+Hnah51H1gWV9NYUqxSMZOK
ks7spAJbauVqPONPVAFoMoWcjAw1J7+l/wb6al3TXe1P5O4AzH03pvEn57gwF9mn7GdSxNoQRXXi
hLhXptLnJ2KO+AN2QgtKeB74+GnGorC/QaThNHCxrn2LjVRFRxkoK2wE7xMAJyiLUW0FeAZxT3JN
o4/7kXR4KcEnaZWbGAqOegoRacvTqt7NHGWEc0KkrFVhZRG8mtWM1/fS2ymMks6hn/fEuZqBCWWA
xtKiJEg+xoJcwcE71S5yhi842CluGlVVynXjHn6SZ0PNpp3+pJswR2ea+b5G2CH63u1noxszFWLN
AcSSBogtx0H0znQr6rCBPW+yKNOHU3wNdB5CDOVFXr1uxOHm08mo7p9Q6wmNMcEoNMHfV76kHA0N
HcZg1uPITyFhzmTnDqeoRDo3s54VARF/MbHy9TN4WfZW18wwF0PFzSN7UM7ycErC/eujD7MyJu8g
LD7GhjY69tYX7sD0oNeuJ44SVHLocU07TVJuhFuzU1fQzN3bOjtheOyYHcF1rYR34ZzU+NHxZCYb
PW6BMhZxTGXaCWDDWWkao2LJO+C+ZkGXW+Y/ojRsEUPLsnuCo6BrlR6VLEbJ/uc5NlbseErDNU+S
28GJEu+MX0U9VGjw/CwVLDLtQac0Ym7U0uHkIObdVjkq5M/ARt1lveBozRLr0XPwgyWnutLFhJoi
dp89vKHJ2qvhSLcmUUWrxUi+fAyiF+QFXmWSR9/RTDFJf/xj9/EkX7qkwA/I9h8xcvFBf90LKyMf
q5OkOE74Mj0Wu50rqeRdxgBHDmZO21UpyT16TTKgXok88guaL6tgOoJv6gC5wx2D1AcWSiz63Wzi
qj86gD+5Q/HtqwGyBMhwHyrmWLrRl4lJQMKVPJfJJj6O+MGROmKVXQYfzGXIEwqF6CcE7kBfCOmC
i/fNaOzLG9CjYVhfEDF6UYTErQh25P2CBIw48ikNWriE3DIRq+okKLbPPcpu9ffJ0Kt//qmE6776
mkpoG1DYYF6rXEEEGiI+dl/Ya5KYpQ25Wvgvpe5lGa9A2QWww0JQtN7cTPZqshwAtOMunC5HTIfi
nUJ4dlbY+sZ9GU6Uxp+dOuxMlRBrVXofmMuPoG71cfwSwPsKjkH1r76evRs64jQciaeomTHdgMl2
Uo27FxR/PNINE2M8GaldBoGmIrh58aVT4jQAc91m6Ctb5SZWxhF1Tc5JkWgSzFo5VEjdDI8Jf5Fc
FzV7DM1DPj2JkeK8vcMSf64KhuCHVRTPU4D9urshWMoTyDYIewNpJ/T6RCSzQJhVPTgdr402Ob9L
o6+ynOPD6Ti3V5rcouggoUbLFBIcjJHea57RuBP/iBq4+BeCADHaPtSa85+n8DTHFnlguVFRNNOG
ewWa4g5AAk+m7vp6iI2gtmWHR2weGutK39LopTYFcxpYpNx+POlVa2dAqv3x29Sfu7l1oCB+dVdg
7XsN4a8Ln9AVMOWhA2fzgxW1r4zybbSXgkB/waFFHKDpCYRhDGiHb0UC4xwtcbX4i9wzT0p/r/B0
bgT0LjFqRzWmxhjoDzPJyS7+VeIT5I7WeQIam7obYcMHF3mBlO8OJvR3t1jtMphIdMW3IkkpSNGG
NjKAPLMMN+DrPD9kxjtXx5gFzPkJqDzOdnGxE52/YwsOIY2RQbDFlJXNfq0OU8k6o/BWs7PDsFsG
ecxBW6zxQhPHpn7A/3IWnlgFadqYYdFcY+EyWS5ZKhcVfd/O1Aj5MeGhpdSPc++ef2XDhdRz4l30
s6NLHmFxHpJaCm2Q/z9ppm3ZD0T6dMQjoHK6mNTHRwraG+Ey6EDcgX9r3GgZyx13VSMetG4gdNp2
ta/6KrSaR/pPK2wikJRqTc8KJuWrVwTr6hIa+7/s5+aKomLplS0hAMu2WgR45UVGJmkN95/ZRbgM
vEDrtJ0U9AErmblRGPR2h4GQz2Xm6P1vsEfQlt38k2uKpWwM4FzStzV637cFKlyw72uHnC1Tqs7L
U+OZ2JcLULsCps+3MWKkhFlM23GMITWRMF+D2i3YUtnKWZBq42EnqSXv3V8b9h8FD+QNwxfWyndh
XJon8aKmuTRqmQO25NIFO2wElSWmE73dKzYLHB+0JT+7q8hLjHr31U4v/LD7+T7qS9Ib5FdrgYhB
2S/B4sN3ad5Mf9pVP1R4bZBWyT4LAWtYQdJedwMSZpE0TaTuxn3IUfgU06Chnthljc4nrqwNqCwx
yiVoF2kl7m2JvpTo/ms3ygQTDBhwnvrvvvSzHbaEqC/x2zlB9bFqJ7gDbPb5L8ba89tegi+rLC5V
biG0VvvCk7RXDp/geH/nOVjnFq4zzKKnDSLYxT8klwfCUgNORyY+z2ziTHNIUWO6yDr4N00E88NA
SIdMYZFYfuFCco414acJfzY5Z6veZEAUgRyNRF1hyHXigKkQWyE1cNvOOpNxvLjhfgHAX+cIkObb
kbQZQfAlxICghAtKxG7MfUgL52OSEvR4S7Gp/ldiiYYu/xQZvaRIr5Jq/thynNTQstGkc9YR19Cc
cej/VjlGV8p+idyLgB/KnHVQvN5qgwP7RjAaKFy1vkhSdF17TdyV8pq9SMkDkHbWniqicq14Vu18
wYuDmHbPIkSm9HQv+7GsLRhXNcsgifTo83gyif++s2DXIzZFer94HywnUs6moFRjdInfGO79de1g
glm+rT2FQHor2dezzMyd9ztn1U7ihJ0sb6FN2y+/ua0/9ZcKxsiJoVmgJMWmMsMIAiMZovhRMHm6
tPFEKUSewZnT/6qU9tX144tN9ZOaSp1ByD1PepnFrl0Kw2A6FqSqqEg5j0LZJEAXwHn4hlk+i7Vy
m2GAX9ecH99pY7GEhYfXK3YSAfEF9gMEPdfFp8+oIH+D9wiE2ohwMm0jVf5c57yMMR7e8DLtIlEn
8fKcFZB6fH/Ixmjivz+xnj36PFPm76qGhNvgBRNjRfj7OHPyEyt3+XHGWXKjKFYEBimiAaoa+ESj
6YbA+ZdqMnxmNs3gBc77PwZ/423IEAiEpk/LaW+r9O5XUHDx7Xv/c0Q3ApcJqpt9+yJDuHff9Lqg
1Yr1Eoot0WManlIgVF/MiRPRlrtOJDLE6P9De5vSOdCbS/w6uDCbq4q6ia6qjIiE48ijVMTRWxGA
ZcpvRIZlRgkFzBF7iDcTNUW+l9sBpnjZK2HLzGELLKI126RwQwhrIGOqsyJV8x/MxHR2QPjqcC7d
vB3LolEOdPrv+RSNGDkLsV/V/xqBnUxEX0S+Xx5NPIXNFpUvC76hxJ4DZXz5zb2SmWC9NO+9+QCR
8TrVFAgBNs0xXKQrUSVoT6z1vfck7MvEcZpWO9lafpQLRm2Wf4XAWQLP/2bkLUdDgXzUKdp4yUPl
Cs8N8sIOB/RY1uVvCu1RhuFt6Q2VXQeZ4Jd1QxszVEzwFMsYsSzxbfFAyCyMdGiHXDcdmzbGX2Cc
/YhX+/sOCrEvxdxRAnn1FGUR6nm9YmVHUSZoCyr3MOlmolQcxT9rqyduDhttLISw36s5chZ/eUid
z3cXyGFtaeSgDiIi4g0rlWmLfUVkpf2D3vk/CthXzVyZi7eTv62TF3DrbWgFhcXo6Ngke+jYrRe4
ZvkizaTLlIG+TpDPwBzpCUqf7XKyabt7SsUskwAiSpRbBNEwy6Ob6OUvWeYdA61PmwEIYdKKwTTl
VgBEocUvysQS3asbhWS/YxgwHwdknwuERi9GDZctMTnJWl6l9ucgPiDExkNDN5Uw1GEfliOO/TIq
9xXC34gIUNNciLe+ySC1NvJkaLBYyB01BY9ojl6ZvjGstyLhsIRaqNV+5EnJXUkwb59ottzHm0jD
IShu7q2vcbavhC7TreRBPY6cULSX04Zx/q7DTCD06e8cpd0/EgWbL/ZeDFkmosTxg/xawHK0w4/0
VdmYQJwAuCyze5RE4BaoqJ0kOcV3dPZkbFgSsVVYeE6uumDzNb+gpohvhhYgxB88R0KLsczp4mA7
6dtiznK9xH+YJxCHs2CdSRXFHfj20JNhG+UdFe2iCuF+piuCm1vnSj1jQEUJpq5aXzw9nEYpQusi
5CdfeIsPth7r0aNlxg74h42qVDWjTr3yHdpFoITgm8ckJkRhtch/UYAnTY43jqH3s66jnUkCq3JF
uQR5yeHB459RY/OLBde/REZgGRkLzRMnfK10socs+av7fUx70cwyomsgi9whTH9Lbi3pgJryfAUa
PkjwXAyPHz0FxBzN3Jf7EnmVHc5qwBv70E6izxkZ4YnfmQvaZkKH0PzsYgW4WwY4BvCEgUAatD42
mAEqEcvuakcmbUSeuByL/Jr3va2loq+DOV+RY8iPO40cmhivEclYIbceI0rAFy4OnJjQcEYZQG7q
ucB2FYMETCWWuU0hiebu6XC2EOZyX5n6tgZHW51xBLZhTU8dvtL9BxpMxM++TLV1cbK3HOhEYVnL
iUL2Tz/hFJBSvM5OmbTAwpqzIEUqLprVu91sC0Wjy+gfwcvcmdCgIwkE0giSIZxz/9qDVR9B4/1Z
dz9VgL98Sa9a4VqLP+zBrtfwoYC/Ue58UHPX9R1rbk+D7O571pvBlO7PLyuXMQkRJRaSVHw/7u2f
C5dY21do6RMyfmpksNdgEduYG5MEjqKSL5Sq3NksuppzKn3lVELGJaxlAUQR5SUI8eb4vKOUkMVu
KrE4vj4UAKQzE2hIAexu0qQnh/JIXJGnBbDHq3yu1LxlBdezjcdrR8usEsPwT0I7EkbyjTEA7Wsq
1cSFtX6MhwpeYa1m4vNFQl2Txlq+JF5F/G4A8TBvP/l7RQK9lHXGRQIZaMgbQI83Bn6m5MPiiDe2
UYQXTQyB79mou7hTDmYZgnnJwA9bEl3A8RYZ+7ZCqzLe7AS5VqhvdvDupQQYHwyhBg8WMT7ssdU1
wv513SUomC3KhhseqpRnp8Rk/NyQZJbATjp55Xe1htVETZadE7afBKPVfaGSUaR2u9ICTWYicE6i
PpC0y5+VPXnp0iii7GnO0IF3G4wjxAyeEk0dRCIaWmaE7QJ5yzSU5Uozi9Ml/E8/aOuwadXqYJlF
zZWf+zBpMZjeAlIHUBAT9qylteXCZe/q9hjwvYM9psr9gFYSO5Y8hGqXOFzyLDe7obKElVknuu5Q
Tej1g0riXQcGoq2iPVVJkmu4n2o9ISQZkmelFJaEI0ftrZD8mNAGnTvMM2705YITQvI9ZqcgIgoR
yaO548r1qEGu+As2C7Ck6xBybL3zvSZPPBc6rX0yZxtwYiZ8b2NzGO337zqfRRgeN85JXo1aOgSG
mF8WTsGdQbedm6VJTrEtdP6/2O+sOVjiDLfXuuEMN5g3c4Hb/iGDiJ8BRjiFAIz0JeIj+c21p9vb
4tb+gWNhK0URt2Ws/dILvDUALIt805+H9VaNrA3r+wWChC35SkQM3I0JuExiqAUY6t0q2TugAXc9
qLPz7Af0BWt4yCQTGrny9c18QyYemSbehZGNHPVV7WTKBkbGO1iPuqpXoqL9Kk4R2JQ25dGRnbbx
6N2tSRRoPnP8DnAojxMuDISOvxCCYeVnXNn5+rWCIMqJ+tJHN96CUVJsZ1IdXUVHN5w1ZgNHn/7D
lWh/OICOBfh972g7X0cLgTxNByFoW6MTfqYq5CrAS+LM4oFGUTTNo+sDe4FAttQGtEpcJLer4ymr
rTsBxuq1wcAcuzP0Bm5Vgst+jSvgB9jY1Wl2d4OdBRKDXB7n0pjclzpezc1CNH1285p8tfSxtOjb
KLXjenDdcAQWNWGupccZYc6VvWyRLZdyljoxEKCrWocxWrl3pseSoFP+RZHXFTq3LpGn0RM3LxUl
Zf2BRnnie05vFkHbQu5JsGhp1Owmd+7YUOUDVQuzTIjfs6fKEdHzXIlgQ+HgNXuwRpLjEw9gIPCE
ArkSJ52DmB8nUo6qhW2pplpaPlaLoMOXPHnmpxemGL5zBZCpxwJSPhSOrpc3c1lqn4FRKz0BQoLs
bG7c/g8MfVKGobcHIXFflV8th9L25sJM3u/GYzbtPbTiCVu5gjH5741kXHMOtpOUpq8ve7HP7tWD
WF4ul5riSN8KMBfYBNWq8QSBdzMHuHDtZOmThi0bEDDueuNwP/3xVzTMqRD/HeE84tA2b3V2u5Bg
aGO8uYWpi4qzkjSeee0l0oN1uglAEK2lVP0M+yP8VRkMiJYr/iMmM7ZGUZxcdfZMfu7KIKc9qzm5
+aUWzovw0txvJrcavGObNxgbB33rogRzGqfK4jeBLS1zgN+cunxE6WxwF23JkKiwrTWc+pcEf8AE
lcp2PtcCddi5vjU6uLbriTe4yfUyytUGVqhTajojeNNYrSWTo/GtSlsqqTIIAfQ4dvYpzUtZf4oG
H3+5Zw0rCgGgPj3K8MaKZ0La/Mdudurf25oD0oRtlbp+I6XBiRZ201RDSbsxyN5VU5ZQKRhzm+X2
Ypn/YDFBXI4ZUT3LvdBKujj2OkrGY6jVWhI+371v4YcqaRAk5iBM2LYXJxIQv6qtDt0VSle1qTzY
Lq6epvXkQSNrxBycTlQ8vb6rDZ5CyEJ+YrDGkshtRdIuOsydePZR052vVOu2R35P5kgog1nIhQ1E
Y9DiU7oWFLCMDScBiPJnvblyHl9hnICBnUShafGG1TQHt/NX4ggFGQ793vOI8i4N1QBogrOJujVS
H208g1CZERke5P2pY57uwwmF/fsgwbaAdg+cBQP8lzSD/Y4UaLowRHaN+AjPIY0IjIJeGgc90A83
Jt/JRgQR2EvP86wIOuYah2O1m2Cp7qZzUWuZg76WzL+/scXqnkbhAQQ1MUGV/A+HumF132d9i6dS
NMafFESePS1D5hSyCRAn2y5VAheAuSVz3y9eFYrVn1uw23KD17r5kx8QCj8Q7I76s849elVdWr1C
ixaqsG8iJ7ALQNkXJcnRFaA4zbuWmXG/te6INWgP4LMtX/h/Mca+LF0+Lcff35VmZQ7/HUOzWhRT
IBd7uwGBeUZT0USejcfo3jiFbikSFx9rmvb8uZxCz/RSj/0Wt/Y8gNXrU3TkY6ngBxTLnToqkc4P
Q6JcON0um2cblUBEZYKS81aO7IyGlId298Lq2qcAcxIAL1dr50me5MHCBP8Oa9SBuXa6ErEv4fob
wsgzMl1eXSPFnQnhPsdYg7GftSWpEE7HKRdGah4hv/E/3TbGnDpVbQpSE/vLnPUdo02RD6nN88tq
ODJ3A2iJWHetDpXKZo8cCUkW0cDFpRMCA+66YdS2/ce0EsxuOJqAEOCrQr7gSU25A2K3FfH4qeRk
BcZeaWrohjKVSYGDWXvgfKS77By7oArRGuLTtkt503SoKs1r2a1GfBq7mjNHdvaTcQHRQI0HPUUV
QRuzgjBrGSBkYNEMsChLCFdQvkpIiF07IIRmApy+V/lYZUNEGipDjmLXPFHEUFOU0WW49gI2sZGt
ZCoEj0JYCRVWK99fqrPrkMvQ7O9u61gpZKjLKutG0msX9BAQS74wo9tz4z77raKNWIy5KVkRHXkk
yrYQceop8CUBoG0u8MyWvwW4nLDMuvJjB40tgswzxE1mneVtP/1bBBcIhTyCYLKmtPB+ae0c6+7E
S899HrxsfTKJsKmtN2TjgISxjJnI6EBiPPxRDVBWKu8WIMvMUakvkscEJLOQFOp1BDsDYiLlzPad
J7qwNlKCOJ0qazuWocXUSUJV37kq6+1vwQLe3YFyNMhU0muBXpowrg5O4Zj0USDha71TzTOD9xm5
KLk7xoeQKih2Ki9RIeRF2XN0J69xjejclj3UQ8yGkUHBc45VV79EGGu/V1CSKJ2xGn6EQ/sHM3Ve
EVK80mIXhQ5HGX5HSGNxN95f4CYLrCymx3pMYpjeigVHzc7pXCuy3IRdq1jb45tmV2plD7s5RuMQ
S1PVkvXZwf8PSYwlpyET4BfF2838nzHU8/zq4gZTmjPQW4vL+JE7JRvLBrPpbYhse8d2LUuydZr6
p6Ji1Z3hdA19sGrhPhsUFXbctjpuvIJ+d93OB/OvwZXcbUSn+uMFKBgQpPJ3QIvuIUW8v6ihnJA8
xtkp8uBaosSLTqbnjUM99YmF3H7i7sVGjVEoDCoQTRBCYZJD2ZVEn1Cjnbcc0g8lmxCtbyGuNPKc
zBnDZpWXueRl7SggC2b3oqW2fFlpDtYtQKOU1JJnP4BirG/lKUPnyCT4PMrSSqiSVphr1anjHija
iK+CyOngzxL1ly/to5hB2xbd6ULI0BwYOMTp24NkCq7g1n+ti2u1rqGVOxoXzWkLt73PjXiKznlB
Cz/U8n+eQ8rMts/j/RxTUOiq/OM/MwcFITGYONVbfnuG2i/a2qqY/Bhgtc6yWMyRww+axVWMEU2B
+Wz27B0JoVrTjZU/xerS00oNU9FvBlreVzSCJK6j3puAOC/WJ/I8U/zduqDITBnUBRU/b0vSyM/V
Sm6j29tVXThmAPi83tHHEeQLBqSlMfd/BEGb6PnGxweBk23+gVxMgHY791SJrZ+OZ7lpPE4qc14R
NLsL1ySkw1JXyFg09TwDB53puHi/2ytRDU4E2sZc+292/9xaKaFXL777hQVO8UDxOnTDJr1Sgtd5
5cjTZoFNl1XmmCZWn1yZbrYlvOFMjAthIUZQTpDhNCsXTA7620cipCLewPHB7YBTpswRedxMWGFp
KzUD5fVPvZAaR+SIJKRNIsi9gbYNU+T/2hOIkmRWFiTRK3CQyev04xRcVDe1JtatQovYinr+v/0f
nhtY9tlN5Ijlz8F1CPMOLUAn56LlHy4CWqi4JczIpq2FHAI5YhqrL7E/DVmceRwwQmi7o/gdo4e8
yStUFdzBXGysDwtbU0gWj+FPCKOv3y/o7y6hgcytWsNF8trQ9iqRsqjnmAkuQ4QI9SFY1bURX31+
XDDmZGUSDM6FT/sV7wDfpPrKa1eAMosV0+6q7pWKo8ah5gNWbvuVx3qZitJpzxCEuFFxy6ewWAm6
1/aTiWM1TOswIfqQdhzQH2r7H1nP65n7ipELXoJh+VEJijneHNQ8O3Y6dbef4JpmJgZMllOThPxV
zgUBuhrYNi/yGQJehEk11jCvErj/N3zqdVXy6mDAaDnkXU04JiJzLmTECdeLI/HPZlQq7tY32Eek
D4Z2aLPbLbDQ452ytukPaTSojhW2rpNX2xC80UH0c3mQfMZynJHbRnvo2U3Au6cfulCIryRuLabn
ibWzAaWT+NLI43uS0KPYZPaoS5dP3CdQOQOVJdIfriYjUjXqC2vYFHijjtGYom3VlEztF+xdgygZ
G23KpQIBCil12Ik+q765VhWP6URkOe8PhpOjb8EBzhNgwKBGKzaIa0cbWcNJOVbj/AdVR9y0iEqw
ZGlF3eewjzd/GjCAqaqniV2Ittsj5efwNqHPzvrzen81K4UmVrZ9Ys5hHIjeZdljx2zQABvamfC7
Hq5zAkM0c0qZwnT6nWH82hkxKZIiTWvJvGsNX7U1pRpowjQAL50fyD7eBiX4Nx1sje3zoHPp32Ze
yW70Vgx4N/0kSpRfp1C5Qnu4/d0698uYmqPpg3i8isqHyMbf9Y3ba1KoRlH3kMMTbN9K1IEh+Af5
q4ZS9Kk4Y1xjkVz06OwA9jwDxjRBSZLUs8EbmJVcrKdV2LtyzN2vwky1bDo+PYgKjpCkKi/y6Ay+
nnqBctmvPGUxDZxBEhMZhjqTyJDszK7AbnYHJxLzBfrf4VYkaH+wYLp8G7oIZIaCiQ8xJy6iLyiK
YoiXySgZ7Yj1qPlTq7zi8/iTqLcmMHS06o6kixfc96dUEhfk7SoBHoRC2YpdLaA4lJuhB/8bDJuU
3mduIQSPrWdHjVfccSWb25tPEvUY1wGMCHoKYupFzQjVOEQlUBqaay242cOFX+TD/sHwYE1c4Nx4
bjY4X5V+GmNHv/ZONDOED/OOtlTaSNiUq1dldzMmu/g2vO5EtgEvcKOUgNat2r8TJN+KKmg8tQkj
RV/W1dALrZQe4wloyqmWmLATiVPPRlGQxuY17Dm6VvwfqeFrHBrvI61YQWDNVNdxwrcuwmZZ7rPM
WMuwTx1X2OJxDoQiC6ZbPOV9y2n0vZNg+yGnKe0FIgpQq7ZR8IyxQn8i+JCLRXhgkdm2irHb6hJ2
EEI3V66aHg43gdny9GeM6t1xJDFCA287vgE1sX6+eaEqq+WXreIYTXhJzEp6c6dNp9zdegSsJLTP
b5jezGXZpV8bxZzFPSXuq5MQx8GwvGMoG7YXUoq7JzhoGX1UBiCUGnZpXWzihQiK/Ot542B7SZ7e
jAyIg9ORM3am+MJrY3EnGBUebe/KT2dqqE0dbTEKw25c7UkffzW1gKV0WhHaezLIItUekyiptszz
ujQ+1wCOQWY70IVmbApBlGf/ifhsfA/CIYHPx2cDg9an8fcIIDIlRV3Jzhb1eQxM/JCN9DmlFwn4
FMDbVFaacHSSXGrXj196KWganvnexpkNzaUCxMG8Sj5qseFqwsEREodKbp2mT+RGd5uidnczYc26
sg7iVIIRLnA9oS52ROC68d6UAxQHDDqsGQT8nzV4PltsIX8AHBz7fjZYNe9cOJzMKg3O6MCGKbFL
sWnvdA5FEvHxbDsbSncKjb0Jz5zvx2IfQcrfCowQvpHBcVQRngFel9MSdB7I3m8lbBV0EzxGZOw3
bzRp1JwTpiySiEqeD5w8+xEEJ1WwJ9idrQetRxveN7q5eFJh7RXEw2yX5+IyZDODNpPegHJAN7/0
65XupwPhj7Wm7B74aEaLqlav4rT5T2yqHRH8ZjTpXZP417YspUUbFKzaiy7K5WcG0NmFXHMQ3c04
SdkL9K/7pCrSlAQQcSulIkCUOAUHJd8vw7/Qt2KMNhiqmXsLuQufoGdYKo9kKkbM249bhQMiByhx
6KqHGU5u7VQydxPE6MLzsQpFq1R4cfQrhYXBem6BCK3fMAjxEA9K8dluyDUUuj0wpwi3sOE5NE48
/W4c298ILk8pqbfwdDE/fe9hrXuyyWbq/JtIL0bBJXqHYthPypcUROYQy6Ahv/fuNWVSXsF/iWdz
a3lJp7ZpIdCgIQzML72y1ugxlDKZAbrgFyzwEombXEOy0NAXf3sz2qKIJzNgxRoBE01Un2vHRTrt
DU4Wb/n1Lj3oOndY5+OidLVFMxaC0S2sBxMnRzRQoQyq6hBu+3rICwlMI3ZZF6klB5d6GCb++q0J
r+VbKvVALrj56XOVshnTsi6p0gjGoYRRTFQEWlKS0qPPBReOwKxqyMVH6MC5DU01E+a6V+jnkVjB
pUjWfgr6KE3igniN/5Naf0/e3Lm+7wqbvcz5Lm6QOOQ7X/Fb5Sr6jKOCF+/fFEp/Fx+uqiF0NqA7
djsOtUptAsv5qCLxYboTAlwUJ/wuu1IRsqf/3xKYps/FPuceR499pXYeQrZ0Sm7+LxvinhOdYN/N
WnrhRCvvWbdEke6QBOZiQZ6Sjb9X8lSA0kwWgG4x62qm82UKL4GBPPGxY92jVOrt5NfahUdb+Cdg
tbwFyMoWUF7ozaIc6bPs54Yf6E5Pa11mVTtmPNZ+pgLE7WOV9vUeGS3R7rXGEYvUJEiMm9a/zep5
K5MIqs9LcD4hcLEY0yn5SQ2DLovj0AkuDeFOD8L5nlBBLxKOK9a0uTVZu0L1wmdxgyaXY/Ywwuw2
kxTXg9eWSEbpp7KNFwM9IF20zUnl6pMXJ8yxTDwnCIqwDyRSo527M6Knsnauz7091AnIEHPj0cjp
WnYDAIhTy8ydHjTMyLhGV/rk40bhLIb9EpjNR34V08wcVmCkL3fcVBHsuP+tmmK33IIzn2qTypdU
cwSko0R0ZOEkBIcSPxe4xdGg5CiAIi80x5vUfHy/1rDt0z4+8jPtMYl+JFGId93qJ+j1oqtRt3Ph
pDvXpiClsUexlddW+KeyZbkvAjvvb3N9ZgWCDHKDnutU5seBEGveTjKLO60aEvH40OAsYjdnJotN
z44xtHd3K66dzVJhSSlekWK59y0DQrpHU4+WZtQYViZVaEDSaieAwLImpEVUxjzK8LcLFL4+xMs0
kkX/bzN2da5jG5xJFM++9V6N2uMCyPaMMorvb6MXOOYRrPuNKFaa9WegM+rXTjYp3wFEIkKy9vLB
b+0T2IE4kwnR0r/BdNagRxCQZuXx4xC1N08c+9iE80ol+k71GmBu5LoWZz/5tV7iQavnbNIzl4Du
OOpcZ57fT934GdZRzLLDDwtpF6RrxyCAs2yiqRFjDnYr94zLF3Wnv4F4BORdqGiBZYXFmM6njpUX
ptnMD38S3zDQ+BRGrzKWcHnDnMma+pJCNenjHZNIMRv0jYu/e++dZmX5uTFE8jBFejPTJ+2BStUS
vQBXei0nmRJ81zS1jdQpzhZJWhp31TZ7rllX4eOo8vnQDW+kH/NbUeLZYriYgOGRoAl/pnHE5vNc
qexZPjFLz82n4wveL/qjRyfI6saGLzPa/5LyouRRWDwBfB1Z5rZJU2eU90Re9M2WNAtFK2qKZi1B
j4Uw/RMfGvGYcoqCfre3w73yKz/gjHjcK/rQt4kPFYx4ceuMFivG+2VfP0lfWz0kHnSu33bRhAmk
TW+0mrJ59Edgbc43SHJYaStKm9o33ttDQdnEn4Lq+o4diVZG3iDks7+b2rCi1KJaeArolC0O18vM
2Em/gNEHgpeLFFZfR66a0rC6RkkYW8HRmUnrbhvczc+26BYourAnlGDbhXJhjlhTz5I8+klVrrrr
z4+26995EmuCttWPo+CzQjTY+YFAZe+cRQP3yoIZAzqLqAzZMu5G4WXs/UcY41lSeignGByrYeOi
jzvFXxueY2cH6knDsz6FPsqJvm3uMQF1PRyaQbI6/gtaGCttWMWjHClxm9DRnmk/jym3hJSRhgUp
zALaTshs3vqUFbYud0cHFaK8Qb4yfYEpXAkwF+LpD0zOdz60+oFc5UmWqKuXWTOE5ceMj16KWaW2
we9Pd6gg6DMIVP7SWGSD4MkdOoLzxweItpNiHG53PzAvZZ5biBQsRuJYNFdrDcrdy9LF9W0zoX3l
+xCjJmwStaz28YLhKesAB1LWAfwzvq+7fKvtzMz0nfPMBgECLYalAoj/YBH9+vHUyMtKqZxbarDf
dgJOHzsHXOi/7lCb+lIDqRvbu8iEcCZRBCHDAC3bkG0FBnQhsr5eRmG1rAEllSSIxOt+KHZJKxhK
/CD9d/FT7Y1G1WT7JSTplGKP3ldhX42jpHnSPyb8/4SfJ+rf2o/EOSDKHBLtCkpFfTz5ZrY2ZIfi
9jqzqdhygGaz93w0wBHUXm1Eu+L3OHTbSYzu5Y7VLdDEsjP3I13FncyMlENP5jCiS/4TpoTfpFmJ
8aBP4YudyYhjccTfwIUfYHNvYdbCWflMbZJqov2PROy9Hjh2i0nMtdoienONzQaexbg3cv9NgMUh
IVWgjPTZbLewX0AjDUqmJ6bwUFksHHBBlak3yucgFcQLZKiBRQHPImtmmG2MXOgkOFgRSi8tVBvP
sMvJrmdw6nT8hFgkEJOmPnAgiEJIYj6bSIt5QB8O7YGHB7P00CIpSxwsEQz+hZEAaJHTx4aSbhFS
/vaz5mLgD7xKBsNMpVpgDgW7jgx233QwPE0KaDuEm47j82zGNoiNYJNEvjs/8kyo1azPzHFq5EnS
aUTu/KXK7wGlgZYgAbww8+ehGqAq7Lb8a79JtEXzemw9jRMdWfqVtKLt5BY82ZlpsFNwkWOA1aAQ
An2Kbh/WlEZO0DvyaX20oe4rVnvgQBSlzZCWD8MZay3OO030cyJv5BJ/Tgl9sBCsY3E4RMV+m4O8
86DS06z70FeIzNMuFzwewarnIklvlW/tQLMb2Y3ABLQ3jPUHpzq1xt0vdHDTwMXDl8FeX8iwhMXB
JPamOZV80idXfPErwIVIbDK5v7S5TPl1qWosImx12tdrn713pJswePfaC9ZLL/Q+CCag/n3Ig6Sg
6VSNMiLYdRGyTVlOk2ewdaPV7MevLEQYC4J47/Kn4yCLt3MkYskjeAIWc/MrI+7OnuA1Z8PNgydU
0NdRqioa4quUaq5GUxBDrwQJnTDwA/gYSUvIvM6sUu7GUyu8Hw4mInelgDZuL3OklED9muVQEcQD
s7yNm9HDwWSqqqehQkxnIdYK9/C0z/UsAr32SMm9qRo7rcCwURxNYa/IYr6xIkipu5m9hOFrTWAX
2hdbnrllbajCpQzIW4t/B8wP6QNyOF2lNfmCS3Idt8YqFhTWVE/dbU6oX5Nl72vHxGNE2jXA0ajG
G5RbW5SBxwrC3P07X7A6O9xccr1SUFFMloJRkrxo/zHrWd4tF78byVwmujMSDGobh8kUlcDT/dMl
UEQ3KY8V2AVVWLI8b3WwxMOer4BzGqZU8dU8snNr6jUr1qErkyr8ulTfePR743JGxf7aYDdyyaRb
9m2py0zSOa3kEOhnrDJ8HjuJV/bSMLDX6AI0vPDmYrafkg/jYMra7bTWMXZqTAeVIgJarCPrlrdo
HlTUkTvZDgzXb9P+9WNI2OGW7Tow2i+a5y7AztB73jD7k5CpIc7owUVW1rvV+3ip1h5w9w1bSgQ6
os03Iq1Stp6CQsJB+cjn5rwwRooUZSdXgvcLPGqZx8hZWHIioxucndVQAsPkQ9Jol0JwV01USOM7
U8q/vW39mnL0DDnvMxuSRrnRzcx1ALr3Bnq+lnskbhcpfVExgjztFDE4OuOgsBw/4n4SgqRMrlSl
WaBvNiq0jdDZ8W3muZYi4mmRjYdJmiG5LczQ1AM6jaWg6oig2iw7v8iKPEtnd4oS0bKPITl6zLv3
c7pkhoZV+dTqmiDcMxT4ptZSdzzet8F4mz1KSfBcEK99kzDRsyuwzXIdV1AiZax0Y/muWqukFIFG
9/8uq+PAa7mUP+h96PF/anLbC2xseyXEWq3k6OqPLYfaTgQcsEk7tMhy/YJaBEzOIZC5d8usTxV0
+eHQTRkZGVpnrLfAh+SLLss7juBsdXL6UoPn3hq9nqc7anXDAo/y4djw3a9jI+WTrmf8lfTAQFfi
49rbBFqS/Mk22ycpTw1BpO6VYOQoT3t04zZqOsFr8gPD0PhVM3dV/rm/51Ekw3kz17uIbxaPkzxg
p9k/cwRS2OC60lphgu6WdUEEQKNWYUFjBLCsULQtzs3R4cYQRf2Wlf5wjk2b8UNj5LI0WqXdpuWA
3pX4Ck2nAL3q12C01QDI56JvcCTOyaNf/YKCHZYJmpAEugR/Sprbqut/aHK4EdfwHRJHrfOapAgJ
i0qa5KB8ul1H3FLImx7NTn3ozKl7MTUzcgT759ykZHj2lvhQ2Vk0oY2L7IHR0GEDuI1gXm9rG775
t9NUovY8Jl4q9Hz68JL/wfv6sVnQs+07aDVzDF+C6nrTmjn/GGFqqhK1+sdyDHdsGWJ2LcmJYlmy
9+Or92Y7uaWoiAfYJYOePNKrr5kuVyuXTLm8ks4L8BMRXcHAOqAbAt+O6dkHjXA/p/yqbwG3IBnu
cIBnpEGZtbw+GXVDqMVA3UlsIqPbGCVEEyjm3iEf/bnC7/n+TOhwPHwlx85/Nlq4bqgIFZX7DgEG
7CXFXk/46WO5zYx7ZR8PPGgIEryenk0K1Ghn/QIZAe/RQuYxpPdH+QpFODbh4hRUPDDmJLyqD0Ll
WLsDtZmdVZ03tAIkSQ8DlZ1YZZrD2UkPrJ3V/OCS9JINOW3+wNfKbJ243Ogf5Qh4Ti1DbuLf3UqG
CRdg+hpDoVG1xS/8dZgbsj/w6fqknMyaJtHOgilkgjE2UNFfXrbd4LZTgwmekVmXnz66W/bFhvCq
nMSjXQz9afg4Skm+NyFTt81Q2OVyw/bgV8vsBuSgcOEQ4AzrsBDuyLfuu0KIE3ie71MgW8nrxQJu
n5L4xfPa+xMF2mVSRrJAnaVq+aaman5cfoWW1S3G3gFNRpSF1b9G9lv/Rp7Afa4YNmuveELJRtck
8mdmyxLkQVCUqivoiL4VTtng7kSIsOfyU18HhDkEiT+bEruILWhlOO9+dnIMiyWb5cPISLydqcJq
1H5SksgjgaCQ0Ejoa68jgMf2v4UXTuqQAskDx07pynYoJn3ofsiIhEku9yWrbQJVzKE7d+tzYm7x
+hCFjpnK0fgcmNbkpJf9y9QGTPwpbWtD5JcEl/hwY+27jq691ea2L4+uFlKQEPlPM4sulQPv8A2j
kAd0so2kR8Ql9SjWTBsKOJhK/O5h5EmwAdh+VMbztKS3vfM95+m3n7jjwzsKjAojuoasFRgqqvU4
UjlLMv6v8+zphBN2Mo1P6r3AsNrU6QLJIp5ZAYu8CZMfTEpJT7thLhaBHfpIXvPEOYyt6GU61fa1
kXAtFBYw4F+4uY362th8b6PNQgQ7Ev8kfXK7su+5qoe7/i8l3w+jqUZrh8HZuTGBOt26QeojWfuQ
Y3jP2ZI0kEX26ULPsGNUoKGvz/SvLRHfku3nExSwyKaOPljatWLLVVXjQbhsjodzKEthZuAYTHmg
jMvzWRZLlmlASjXW1VziylkPYFcBBF2+fVgQcAtZKcr1FBbo3u2ynVaLbSl0kFNM8ik9gHblzK0x
tp/cPJ4hhn16q0DUfMoN2vY5F/UarkfddIWFV36sqYhWNekZyJV429/vsT716O9607lsoLkKq0Cc
Avlyn+XNSW+Mn/8p9tgZjCRXpoRSsHTEX0x1oMFp9eoTit6ahOYUFJ7op7j835ui0uReaTgjZ3Rc
sa4xd1xLMwCxCj93EXwshU9QGup/O8gKC8nL1AmcqhL0VUY69gVjAs71ozEZFi7swASYlSDvrEhy
RMNdmuC0MszI2v4W2vg9uZW0/o+8TQwf53JMlwXQ0U1XUeIPCZsbrQ+xu8XURG8spir/ylkWYDf5
HXBjjWRW9YDpk4ReCj++c2KPbfb42uxvOt8bf2bCEGzuPThkzBfoGHct/8VX3IQO/CMNwKtyPJlP
PPl/8CzB8B2UyAzl3q9PhBOVAO2bVOwq2i1TzkQtSzMaYgO9KdEEvK+hDA7j3CbMQ9aTwnpSHORm
uJCarAzyZtRV8QV26E2VvUL3cVCFMX7FMmCkjynYBY18pQdLBdej+fFA9ND82907nFZ2ZLPI8KW4
neeOFYdf25KoNUvZfXJGBnqnofK/2BErVGFipKXNg3iff/ZyfoTbPqAU8y53E7Tp+aHdlpIjO4y3
bIuI2nC2g/tjP+saUh85GhZP6lTSr9shvxcWRVn/ArgiMxorHKljumaXTqNrZEJ1t3p9umwGd7Me
O+YCiCUZ3Taw6lDor00q8xmWSq8V50SdbquOM3bXmAXimjhdkQgNvW3PGSHfNHYtd1UO585CT4cl
C8OXjfRa1jwG+JAGwpD/bUATULozNTABC3Hags8yzSgnbjhS3Pq72aoW2I8GVRZGA323qvZF/Wql
LNh9ke0JZpoiu2RQlq6RL8pW0ugP1dd07yb5v1lP39gK00AI4jbrIENsm3WWQ/tDjj6/eBNjblst
5Imq2Law3slIyaWMeItcyBSO8tNppZPJhAS3VPYysFYZ1eFtDHJ2Jq3cELoNB5UijRa3zNiF4w5S
NGfE77vvCq1D+SEPV6wDUDi+/5OdjXiceiOiFvljFLvhbbwqm85aSb5wK3xzwXYEo2ez9vhV5nN1
w+dSiDkHRti0Wl1/J155gKTMu+pzUWcgq6z4OhFBJYOejLgcMwFEAvW+UqxNjR4bcFJ4WbIJLNte
VQjaFOjc8NFfVhEcjmbVn3P1X55YLeJmcpkIUaedNkJG3eg8d3Y3gzEZ3XPvqaCQ1duh8hQ17oy/
TC/WRqx4+Nos16/ADBzS1c0IuwnJuYhgW6wRqjh2W4BaKhenSMQhblIiooWwb959O4EDLTfc5kxT
OxyrxJSCEEzA5RkirlRaWb9rRCGi8pltGG/9qq6FZgwI4CMPpjBckdzVVAm1EKVOkW4rPOh93NS2
QToh0dWHmGVqpaJb2F+HD+Cb8DRUupz8mcf7kU5k+lL9/CacxYFiDLJ4O3HmsC0QLQe/e39NZiyj
VWURndQB8MTTeQp46Ntx6O3Vok78ozyjUpSBj9XlzhCXRcCcAsUZZXSGqdUBddUVwVyH70EtrhyM
e0OPVHf7l2o/kziPwtnEG++cY5YM5yrRC6Dv8JPvLyY7DIyz8JuYS3iI4JNVb4OozutgOHNcYTjO
8piDn1Ffc2Qcw4STV+psZqHQKJucnLqJ3arDp9ppV+qKxGHDlvVoynLQvx0Mf+64whIwYE4AMKBP
dvb7LGh2hv2++N8QJRiEqR4qTFuK7WNC1OKsyGGL7SiPwaA4GPUBcbl9AYkM3ECp1pVzOIPl6Tz+
8DEnu5Qwlk0pdDwiIG9+Zztk1wNbOo7ynO48ddJ01qoMj7NfHCQFo3yU/c4EHoXeqNo23QApkI4+
Z+s2G3mz2pnC2s2Gm8SRugw5E3fuT7c6XepMtw9u4yfwOILXOWhuiCKZAhQaPD6wPXJVNRqGg7AO
KVYKhEWGKChhXe91p1zqhpkPd/LOaKdSA74guSkabboZsz+SG34RjPOZfi5oo5CY6CfRu70sZhWH
CjAjHcd2Z4QoTmfoiY0F0/q9Bs7MNTEXAxZTqS27unBevkpGPrEpecKQsTohsiJcVq5xP1XSEeLx
9n687VMCC9eFizDOTQCyYA8XLDTWXnqctLy0ND8rhp/A1F0ZlqIRkrjItl4u701zfcwGtMoMX6eU
Gd1ly6Xd5Qhc0JMtoNb681DkJL7jYTeoY0pxuC7zoSeBN3MkbjD5sXUH38dAgtrn93aaX5xAcwGj
1ih0WG+6hAyyZ19IZsvxPQhssP3o3k5DTnZavmvX8+LqIXUScDeBHXJUVqj0ZZPC6Uzce0A1JCK9
ssW6QFgmDLKT7UY0a4hGhRSCBeDtNVo+6xQmSITxSoXxpy38f9K/m3WAcEdX0O6m2VCa638nXOTy
b6De0pPq3GxiII6Nd2EJXAaiTG0OJww5gAt+OwC6a4EhFGRsgzvpMa3698zBPCrHhy01jrvmVc4q
Ky2/UMKAzPbTKjjRBQgrjXZwBO9XdpY4j3NZoFj8k2o8j93s04/i8366YVXEjGS8nEcBC9bzGGMh
aBMmeu2w31LiY1cvMTff/h/lI7kul5WcSfUMKdiF16Q3faRX5O5vGicD82m32tIs+cTNtPMpp6G1
W8amdLOcE4jF6gRiTdKTpaD2rmbpM0FK+M6w5eJEgQhNNqzSK6tet2d6aQcepwa3O9xYoeYaNX8O
4kuSCNBZF72je0HDRlp9AQg2jMjIesmymfoWW/EN8OG7krhtgwrU+FL2o/ZVMRsjKvLdNDFNNdUo
QcV8hzXlMaV6Y+/XfjJa3raa90bE03NAp2XLz8pSeKHlLSZF/P2tXKX67egVOSoOf9/rDG8ddwlJ
3617kZk+EeQr7EFmmP62g64OqpuFOlerrtRRAHwu5bmVn/3bnjGykOjjsI3b/IWVrFv68zFf4Ffl
5lD6X973MaFoZQ1YlVmBBx2lORKbsBIshePwXYP9+sldAvTzHUXGGaBnhyTfQtVDcfvaSeFIYDoC
HyIWoIK+3nv67TpC+LD8eq3b1mSerITqlpvXMB0X2nC1XJtx3HO5WKclgKCezaErAzp0ovDlws3P
eVQDbnHnTyfbeyrxgBrDu08DRbBzw7L8o1hZeeJfbkwfTHunhkEN17BqRcvO99jPmOOGu+NL7gav
NXzIuo7kIGrljQSMUOHWquRGfqJcf39iikqbNpEkY4UQPcHHeasrS9Y1EZjuIlj7351zH2HGOgsP
f5VNf96tPhu6v8kj1Ej+d5LvFLbxkak1a+4aL5sLhOuVq1AEk64md9UTrsoEHq3Fcgl9G/DwyQcV
2Zwls0aHoFo1nnTc9/kLEYC4KOJ3yNy1IHYiSWxBHL1O+OLN8VRtuylgzFPnMhUSVpXHLcHBz2WG
nnxQsGPc3o1niFdhwvn1Cfg/DnUKmzXCEuIyeIAMTaF/F0WfSZ73XfxAB1waDL9mCA7e5njIi7MS
fZlJwNTBc++O8M7MHhPssiw4SpDOKiB4HcJSW1ANjnNu9eHuVQyy94u1FQ8oAf+qQSHGd+KIRrst
k2dDCqfMsr2V5xha6rYl60Po1FUQhc97QsdO4soMK4lu0XuptdSXDZjw4MRJ1v3m67Ct/Mxdbafe
lG/tihnUukEZTSN1aoo5iflFZo1bslwneD4tjVxF6SgX6pMhEAMbEOFoocaMBfTjbOZzlt+g3pkc
zpobyOvuIx2V21QJCdT3fiJD7ug8afWYp/XXCfvj+Z32ORhPWpN3zQ+sJZ0Ow+cXzd55U0YykQ6M
XkmIsRrwmjj0JD6IORF3jXGqLFXCwb6Bl7W70Mgk4j14zdb8SsHFzXtg874oGVvH6WD2LDGQEAd1
V3G4JyJR1uzXx418uQQVWyj/icHOJYU+NjsQArPcbNn3ZzAdscVsb01n629DgxVD8zFIly6R5xqS
dIb0sG9w+Gfb/dpTyqPsEgFT0pg5KmnfYpKjAYeFNEcurPd/ZIQryXlsDzhMdJV5T4zFXICpoRYd
VejaNyYW0dLWGEIfqJOGqFgcTV55l+DLGpmNBpDqnBscsclwqBVk3Rea5XOtgVuIBiIqbl5qUgAb
7slR7Xxzu6zFIkbynBSYRSbhcLIrVIBUmk+fu9BfjuOtMRkBI0bJlzuBuYr5pFjQlB+fCoy6u+Up
iSFALpQY+sERpCC3du+6dKpvJ8MCyZ4dgTkdTC8qdBlPJWH1Ni1CTS/j86kTEsR5YlylMe2TSEuD
I1B2qR1WogMv2nNp1itudgpy0/Vu2mdKWAey2uKPQxO0wJnbyVDGbY9v9APiprzpqnQl64rRlJhA
7VJw4DIjYExP7C6fb2ElLlmQlYnGGxB1da3PcVCEPtmWchvZFvLx7CgNIflBTD+VD4nUcvM6lycO
odp2BjXPDJKNaIu/Pwa3suFyqubD/2iyRcdnKhTCpD7z4kIzReDD97XEQldnPtN2eAqvslslIRcP
FF5oBPTcEGh99R5dkwb5oYOf+6aObkianOIq2odArCD4jeorx7gAYtzOnDeMrpcIX1z8ok+Lc/y0
3Q9hBy1692u6M8a4lDd3PIifyjMFQxSFv0Ps2PpAWSXqTafHO18Wf7d+i2MXziP5P4q1oYP1J2m2
sTUjj2Tf7Oe93dT4hdrgFvxZQs+/qAZ+fakUVFyVKN9XzuEAd1vpag9mCMiqlKxyxewBg5rrvXD4
9pByl5HucBxQ214vjAIXt4VSNL+iwGvigrvot62pyMyQ0Xd6vOs4Ry6cdxBIBdODwD+Zs7LBoXFp
sbhwIXgchq+kOWzPswclTuTSdp5ZmS91wgCoiBK/AQaxgGW8hIsYsw/BCsXuVEo3uRhcl2qDJei+
+73FpAdcQ9BHfjrWWaUtGfICkmnkIwoqSbpVJNlFt1VqtF8z0ihxEa+2/ieNIlIPEf0lomoo3laf
0sBgsa/2a0zrs4P/nF62Fnh6wBVKTpyXYy7OOcXeSq0ulu59B6CNu/fsNNMTe3yHP2WCzUOiZ30i
YyLGuwk68zZUVJkTFw9g2Akk5uwSfRvqSjWawBZBBTk2ryPhDrDF5h69bq8s767v1pxkSyb9Z9e7
jSbSEQ9fMA3ULI4b3xR5Rkbj5JgbcCbPKBqFXxwDOX4qw21CUGsGu0HJkB+6dxTdziBe5GJhSZoR
uORs5E2x7CI1q70BWkeShBNO+tUruEGlHBAOVNPTx64yUUjyNsaZhIWa4HKDrdbPRwTDEYtspqws
L4tX8K3ttRsSMnL3nTIn3D/fNk5RFeq62L3SjG8ZEpkVDujoRfSlQ6RDtQ4nhYXOag0Gxrv+Miq9
NTg5kghKm1iXbzam7V0TfAZREUfrwCPaPbFZhjW/gP3Th3z2wAol76WySHR1kS3MsSsiNHENH+2Z
4N4X6ce38F56O3GjhJVEAo5w548UTcs7EEIJVaOpDI7fiQeQCHtf3zn9UHcpGcgpqOLNbl9ERsAO
Bfp50NXnyHmCyzsD8fq4mz8unUKLGWiKCU/f+KiY6nY/nLzX8jLhArVqO/GE+7CA9uByKDJ2JAVC
kR8MRVl/TR69xBzETrJUu4i59BH/tK5z8gYnKxUmu6bSNJywCQfDEKRG04YD8SBz0M/mLZoxiygQ
mWSSHl83UcUiFajxFitP9FFZnEC5T6qU66PaqrvVAlC/CUpP4w5s3HnKFDGVZyA6pe+IhYUDneUV
pmgcwYV7HrRZieDwz3nTiiTqGzW/Tl4ay1WAvLleJGZNQ/PE/CK0ETbbbJNg2pAAgHhQJI4M2Zs6
KrLBuU9Ml2HUZx+9OnKdprMqgCMj6mC+Cw0Gh5LWvC9QB/5dlPuOOOeGx3Zix9kxZi5mzmAM3ZUE
MienYaSg2o6QSFlAIZaJa4UyEp8avPI73fT3MT0beO5kXz0DKbmQeOQNuOPlXDQQkwDM3Cezkpr1
C9Pd2hDS2fBAFayiP28nejhFct1Rim4rdswXsDd5qv5HIngsKGTG7d4DCty7dliU04UL1ls4R8CV
ro2wUZL4ztyFEZ/aq5QZIBk6xe5rA7uc1ESBF52dT2bUDJbtjXV44/0shXhB5X6bAgyFqBJGAOBo
hHjFOCPdlErFUzPV+klmt/VPN2X0BnBbzJ052r/l4le7ZrqZcQp7/c3KsnPTsOTeOV6aN+4cGMh0
NHmZIOVJ/FLDIfcbvBGd2QoJj4h+rtOM4AYUj6T2K1OMdTi3qQtUHLCYpDYUN2HCxAZddaE5A2WP
HCkuXDkzHyhjFe4CbZ9b2s2oANndj8KKBcp262De/ZF1icNrupdRd58hnli0SHp7ci7tjaoVZD4h
npZtem/UFakcNw00sDgGPSpRTCLZA15KkyY4qEEsz3VqY+z9uSRaEgxHFq3VAuMEhJQbQhUruKJp
PAGVauSYSmj4Rxm5mKyyrxuZ7nOi/EdODcAZT4bQinDpvBZDNa/urIwAhFF4/uTGDN/VXqnzX7h9
1bOkOmx8Dz0CuqHelTveo/Gq2e1PTiNKuw9BxNjgEXAKYG7J/+57yVmXC/rG8LUXfVand3XVizVN
UXrBXwlWyCXtSIR3qIUKJObv1WirRNqoq7D6ZO28RuQ1GsZpdu+WmmxJPYfwDAd3pGaou/DkyLvc
PlUGy7/UBvXyUjagIkzS/LuWp7aWApwlu6xF4kSfjEZyzf3KILLPZVLKGH0KCTHD4UAcMW3yFcsR
5d48XwTFcVOF/7qs57AJCh6z8PPGgLH1f+RCXJDk+bA7iAnYHsmkI3QaXasYs+aCCMOXDfgmTBKy
GwzcbEtlSNjFJDVxMavgz10i+mhr46OZJLiC2czTrmBiYiXACBtgbZWFGhes85w+Ou+c1fU4SlnA
a2SFm70rTxmXL/jGXdeNLsa6Yu0+iaSIgcLp0VXYRxe+HI66bwgmZhnjyI7k9ZIoLRPtDOpBv3/X
Pv91qa0mX9Bij7pnSJ+kia5rQXQGQlMfBMCy5YvBrkXQzQHUYZoPdKuQ19SF8ce96i3R8RvKjv1r
cMh/ALONhQTX+gpZCLppGzNWNFEG8TIulCeTs+SPs33jEejVi7U5yxZ4liWroCrf3X5FS2WPinb0
5Ykf0flJ1DhriSJ26IgFXLpYAW5b4GzgIeFYe5k4a8HIxxBD1FWtU51EjAterWQU4/rjELJcw+kz
pihdOt3iUy4rNt/3TsJFgK35TRfBLz/uXrcZaD0RsXcTL7hSkzVspoYsuRxMuno6QHGQWHswy2xK
phoLJJSRUt0qjM6gPbSrGHPOtJi4mnLvP+Rw7Yfu8fUYPnezbcUMEDq40l6MFm7G1xPwoChb5bH3
mSwvDEBzpOHNf/BxrJX52bSW8VMXJSEnIUFrUjx9rCfLTHJEKM1NOrOTwLoOvuZOHIrysrVc5s7K
/982PY2OW2+U47/is0voLbDrZ2RIrp3C37uCEnmNLYah0bbJqkSIdyey8zn0j1IZNihi3SzZf7Zl
9p3wo9BNjBr2IVGgEWHGK0XZ4KfIhQs3Pp7/cLvCEDXYxxVl6mIgiHZ7mfIpWXfXFiNjvOhEMrcY
wzgwqN8z1cIXrUAzTh/wWQvuMbril7o0EPdSr9z1ic2+Oqin4uxzXthQU14tl3LxZ3oF1Cak7/kg
xynGDCOXKq5lipcOcEnyvwsXZobQPrEDdBnnNBvxlgve4InUE/B1WokuKcuVhjbDcR7VRQquQFer
JRxTQ7QpwEsv4N0fFa9rfTrtWB73DSS1YjwwAEglhn1Dci5+dpymb6mYXc+nOS9IoH5Hq3VigunL
SqxjisvncBTglyIKwp8JK84yOqIjV2pP34dHaU0eGW3G6uUmW/g+ncVd5+szsc1tzgmU3tAXpmgW
dlLqOaL86p8leBpTwZLkDf+SCZwgvkFFFi03/7yWVcFGvAK6FYKPFBftMXGurM8phUzqVunDLFnT
E1Ep/KW3MiAXOeXp4v3nfsMNYFKdave7vzuesWM6hKVpQcc0PCVN9HMBu3gDuoVnEBGXzYpvPx4f
CDxlt5rMETS+iZVi4o3iKx4A/bJJVTPegnohYPJrg4+L6A7bPGtK5aW4Itx2tVjWAw9akHaiuNLc
/kEbHosVmJIA1Xo7h1hkK8y8g6Fx6uKLveo3bDpA0EqEwaUt9NSNNvwawY8MKG05sVYHc2gedtoh
A8rJXfXS8FeOh2P6aiOyiLUysjLGfQVHY4FN5/ivB+uiK+VZ4zPKLARxG5WNF3JEWEkhl4vOtrFh
hDMki+eAK/v6gQ1PTrX9njK4np07kXenUluSglGF3BSOUZjkzMUup39yAqPGMsfdS3luITnZby19
qmJrCqFdG8Kx1hSSV0PGaHdOF9SquKQ6Y3rdaZpE/wzgyjuwCgrxTU2EOwR33OCQHMtoj+1Ljzi/
e8b9/iU2jE9Yci1e2DIdnd6oNO8GcvPnq72lOqD2kpUqrSHTwDuuMdPDibC6XU1ufnRlHCIGj0gy
FHIHvt4G0qepUrfkjPsnEWBv53UaRH+lRmp1tefFWVK0xDIsE/XixgkitJlPnY4tcMjhcQDuLgWP
kWT4Ib2r7ZlTVa4Tbw+NSir10o8J0E1zO+4XsvKHX/ZgbjTpKiT5Ov6IpgFsoERmRegNOhFiqpyu
L76wcbBxvH2iLIZZ8qRBmcNlc/a1Cm0rIJS/7W1UKwc5Ht5K42iEh80/1i4WkhOM9sG5ur8zHY2Y
vTcr8kivT2XG8aRlgiugQBfPmq7h5YrTNg1HGzklT33TB+BX7LBkueT4ymwAUzx2sb5wHx8j31wm
TAIEPEsAL0Ii7vqVaQF1VfZM5xq1l2hnYZKHDOPvmLcl7AIJVgq5pY90InnUIRTIw418BZKPPPbX
VW7e+MI8fAAb9+U69zbM+GRDNHPlF8Uuq3ZtWVFY/4gP2puvt/BJ25x9WYkp+hSPmZpCMoZ2HC0y
zksl8fmq5kKmrt6eh2faHIbvPbpfBC2DWg+fEXAsoEh6DVgaIpvce6W/3b9tWeFOZmA4678lSZ7X
XSmVgRpqwlYWzIgYNPw5tWn3sT/DGl1IJF2nsUgDN68TZhba522iqiXicqcYSmErVBz1AchebHmz
ulPnAcxxTH0VMsnv/Vnaw4ZhMPk1Uv9XFYlP2zuJxvhJQg52gE8Qxl6QogxAMAPnPpVofw+OM1/w
N54mqn+QXQlZVeIVjNaPojeOPSG5fTz6i7tGSTkTB5wIaQeXS9h3MglCrbkPqqqjxYXMokhlkNsn
ziCUQ1M8LmyLIYTBOdzpocvNTVxg+HNM4s2WS/xZstyL/72VVm1Af2Z1jNB7Iqc6sx4HDv1jFnXz
bkjNH/ZCxaFYac037VgHb4Joioh8ZT+UHwSm3GNKlnqNujJO7VHrBl5NsErrWIGV/wp8sFxn83rN
RlmgZ7Va2sWSO55no3ldztS+A3kuQ7OhvycaK/eoFBdSDYvucqYhaW8uy5+9DnxT39hVu3yfZsHy
UUN8hHSv/CC9McppYipQBXUmlp6rFnK7asHvJYmVtFej+vXpbslj2Mt1UleCId6oLLemdBVnjTZ6
dqDC5dpgSap8OUx3TGvmGZHfAeTzXH6PxDQFmg2vRAURndp3nOAXp/2EpkNpLhwOFEoZDzaTwslY
aYqTu89nPQgJnM2l0RiAgZbzgrmTXfAtGbkQV+0FRW6bqMjmFrUK0H5hnNECzOcfUYmr+UZJDyr6
HYFQEnJO0GdbXY8IMq54q7s849lawIDAVAtFjpP7XlSSZPOCb5GawlSTNCf+s2th3wxU6xT9zrZr
Po6QE5xVXQF4fm0YwVQ4eojFCbQUJjdGUJtC/S8eRJYszIb5bIjx1522SWSIYMMrmWHnzmtq230l
w0xSwDw7+0TVIMfbiqA5FsphRhkEdF8qUiTPz99WTqVtZQtUdRRsQsz1dZNZZ6mqxp0opSXv1L/d
fWv3nxWZxmCNoG4MKu7tUW6KntRQ2/wSyFbHa72OfZGOipoAaZj89d6MdQ5LD2XxDLJfXebg+ahL
Kk4Myqt0ROLztFFnLMT3wvlccJeTMDCk7euUmpYXFQZxyruynSX+dZswCFYFKsdy72N+3RLRrMdZ
2mGj6JRI7tuvH8a1wTo+jG7WFBJBUKr3WdjdYitftNj45MKxd+anbYkwxggMpXvw6iNbwvxB46/v
nGDatkkqCp6oXatwSTVGk2seIFu5Z3x1zO5r1FYfz6hN3ubQvhiQiXf3JAeYx172RPVAytf1+SOd
H3AeQhqHBjL05IKTzpRfChzCtLy5pbgkJZ86+Jb5VF1n/2+3mvfwhGfHtRCkESq34t4OaPiexoon
07HXlIGz9K5MYiO9C1UwuoFsbxOTQUCZZLkBWkeaU9bGq9+jqPpt0edQOwyJGbONHKLFTSML18q/
gy//lp/uO/d/MoXkTfa1bXq0upIMOUq2pi/Kqe7H0B4ez2DiytIDTVu5Nb1H9jAIryjEAAvwvVJg
38pOsxjtKP9kBskAwHdHRLFVvSuqruJdHJTRRcLmXI4beQyugSNINPBe3SJ2A0i3bOvkynktCzeL
0otLn/rVQRO5iz9tVaq4Ns9UG6NgJxAH8hvAZVvt9szpAKgbjMZeDys8EwfMr/hUtqNHMNKbxYjP
ljUSu3Pl4Wgt876w8bTMtP8QmdjV7Gb8qCKU2h5xEMcem3xK3XawuS3PKZplJbs79jSD50nFKJ7D
FuosDHvmyWtTnzL7PPoaefSxg+zlh2snmfkFf0mzlRkoCS0USQVlz8Y1n3wQmSg5L1/JMN6EogN8
WAi0sLzSLlR8gQtNgGbViTr+mn61SMLu5ynlxgEOrsBg5/lbGxm5pZOki/p7a0YDMDFABw/0uWOC
oX6oRrPpLXK22rMgCB1pbXXzF2PomVsQ2XCqUYdyRfsA9HbrlQhJzGxCit9gwwoQlrmeGjymtoC1
JSTGVK9A0cfkCfaxXIaL/oVlHpTDbdQmFjwJRo0MZWEUHUk1K045d2i9qXLjyRDFgauqVu/CXf5C
nTCjuHYbDeMeU6nx996pm4y7Mh1KLzigEyo4/P1yecEvwsIwCEixXolIGXjUN9LBXf+WyuXi3kpl
yMmerzSZxwluOBnr2CM9QWegjLqq4Y7ItfBmaGZ9LQuoF7x1TSRhc5WpO2QaJBCUtMh0i/sVW8zB
LbUnOcmpG0no1gKRxmjwD9pDvO3JYGCCtqQq+VhG6VQ2p+rtqpWBBS/4Bm2zXKhntlXR0FUjluBW
YM5W8Mnu4BHK6fVbWA+mcQpas7rgNMszk38Qw9WQBp61BFLnWBcYhd3a0K8nnQJ+yAnr+E1j7NgN
kg+m418JaJ2pJSwqYIwQCvWGoysfH2oh4y1zbBUQNozqp1MfYFx/ckKLsCD2n0VB9TFwsXADx26t
lUafRvtocPz1qUcJQSVY8LcTFxqtq/R+NbRdMR1gK9m5K679PQXiuyKJwIllIBH89+gBb/7K2LkN
6Pxgje1xYyJo8bcQVdrajLYjFP/MnB1MAdE5UKaexonR23AkeHzSgRR2MRS4CSD2iOAcostbIT0P
znw0ei/szygmpSqlq2X/pJ+MjPc6rRZ6oPnmY32TjbJfrv1RFITNZgXRbaawMKyFfjiN+487yHxW
dML3ZYs/TWN+UcHCZDRD2IRE78QatfdwnBtw891z6C+idmTZyG73iJZzC9dkBSTUuz+A9imVm64l
XZf0Kf5O+cyLLswuwp6J7OKPuy8W+eWltrXWWi1aP7U29ezsBeidSof8xtqTIKWMa+R+lbesC4DK
u+Nsb6PFlvUsCTi9EXVJ8d7bfIZwnIroLrUm0P7KG+JWVH3PAH58C/G0OmH8qpteiNxIHISXbm5D
X4hoGxZaGivuKQQ4kysvYvAHp7iQYKdzGZ4kq069wHvJtqZ2zDoWLyvtXPdQ3aQXcE3Ul3cBPFS/
QhZSaPgfNM5h7jjmXSY8gZ9TVBD0YpHEhEClHcezQhNnz/keNbKM3Edf0vp4hAw7zMwRAWX2Lh4r
HKtJCbyC2bw1OEGvQ9dUi+A3yYevYMvBHcSKdQDNBIzKcE34n0SfJC4vXKO+UiN/+ISZFd0JWEpL
cEtd7653Kq97N25iHUlwg3H/OTjywdIXI0QEJblXDL4UH6EzNihzuXoSrEc74SAjD5PXjbdL8UNK
JmU+4zsojGP7ea8wqcGzlIHR9ml1vcNnu5Lbj0gXLCEpBBl+pZtvLr+FXKaBCYKpKM9p4iOzlCFX
s10D9mrSjUtvCTHfaLPcdg+1URoRxIWglySqA9h3h2hVd44nPlrHV/7IRbM/+Iqlb7PEm6NG6Opi
JYaiqX0KRQOC6+ek/B6HQO2vYu/dEFmbDJo/f4wdmnCp21ZMmO+Kwdhgbx7gVOX4MRcwWXIcbPIA
lubkIlWk8IInoGYHqwWNmwLc9h2khgr6oK3n4Ml/nTWR/lVobu2AmAdNo2OwWPCQ1fhFThDNT6HI
nLqf5H1C5NXoQPexPyzrSQ6skJx806vgNjAgRVT6jAduh2VPv6Gwl0Ww6NF4KKKOoFTMZ3oxdu6K
WHZAdRhTWEfAlqKOxe9yraNMiVrAD0YGTumMJVE8Z92aUmv+MvXUdGWDrQEHPP8+PcDPAZvIWP/J
u35SuAmhJSwamjWiEr3DSOFzzhM5zsGK3uZZDCNkfCHzISQEx9jb0KkUZrVrd5dXkspB05M4NAp5
EDKazjlyu4+ElVIE/OhKGDugj+EjJW76tny1u36PR4icmFor3sCiqgguM5ZjhSx6qiR2yZ8F3cAR
mClFClMtAU9QtPGn1zvLixJQyqdEoYqBfJh6Xf6N3UHtWV9tZJr8vnZKhbgVNguFjVI49rtiFqT1
6K+gR99UsOJiT3LrgCg5wEokbwEQnsAhqLIeFclnGmh6TFqeBPu84tf5oHiq6qGBs5Lxha+49r0f
xizdVPXwV7S8/N1n8IbZPPaCGQnuz2kvFaTZap4Bum0OvF3eCEvjmHeK3wdwwcOxT9dA/OetlFZ3
af3Wh7ZWYhIqcnZ8k0coWbgr6Uk8nzy2EBlizbmOSrsbbgxp8YZq2sBPifsSvgQipNqoKm7wUQ1Q
W1S1CSsb9WClpfY5mdmqveDlcWuqFjgR9MRsABp2hpoSXvWuqbC8u7meQ/YzFQc5Vaivv58pyXMS
YKqqF5UHNIQGcco604NGTn/HzGHnlyvYr0V31AD0UzAOcUsqxLD0RWmldsB7YqR9iSP6ly9/VdH4
5zfNcHNFr9lMGmt5wu4N3A5sCIECAcNFKaTQo8fgcAQtXvYdNGasy0VjoCxu8z3oHQ6A0hJ6l6jQ
hDpVDkIxCek6lFZlBsa3G2wpIVZCGvpiIS9uV0BLma03vbzxKOYHF7zdljaBXzBfvwCqxbB8Su+O
1D0xfUSJeYKXQBdqAmBwqIVXkub/A4slQo+EXd9nGkU3TOJz1Bg5tTjkvApl8/fSojqELZLOy0xE
zoXEJPOyGh/4ALIZrJvwUO8nyl30A9d3k+RvuQGUN/9oqWg0h+olKgZq3hSLVrbH/efkdLQLEiml
URAaD/tycHZ/+otjBzwSWfHj3qgyBNQcfPkkTrHAxadFvsfGX3r9QixiG/vsJ1t7pJc0NG8q8mtF
DExZ2zg4Dndps8yxtDF5gf9ALqn74dQMcuUDkBbPDWlFAWnjxZw1UgTWrXutBbV0QVMpMSAantao
ch6yB0Y4sXCMb54hnhJOC2O/6Yi2aFf48r0/18XxcxcVWN+sUsXorVx2M0Y9K7CkdcTB2ugvJDZk
ywvKIbxIfocwGL0skQxa0/V9gHDWtoDf3Ep8gPk+0I8kZGbdHBVaZxaedXkSm8Zcg25APA8MgaPc
Oit5oC/jGW3mO/aJx6lbagOecpDMHODZEo0ubLwgr6jGrY/imdFHpW6UOq6+tmyWZ/4OSzAdvo0n
GF7ba1wsonjt+XmdKHgFyiRIhypBFp01/PwBdVKxQqVPEha0Vm1udK2SRij5xstWboC9PEUqDBJ2
MnmCCUNKo5Lj02yN+dhkoUTKBynbZ1YJ3SDo+Q4ELvecEzt5sRjOfQw+cC8FrTSUnmDoc7MOWmsk
7KRp8WRpIQy1obAe+SC+vc+zE0Xuq+64gcPKiDQL6prMLu18uKsNaWkaTm0su8Mevbz2zTk3ApGO
Cer/OZaE8E31P/47SMaRU31fqpKyivLsSF7onk6BKc+ceyHeJacc0aEKs5uRZUun8KIoaK/EXiok
Q2cfNOTCFjMuJSkXNFdCdlDZ35cUPXkc8EPYfxvFJSK3hao1iGc7nhopVOee8WhBn7hDQdz3ircI
8yEt0DM8iaIh5InwUP7T6KPiFD5Or3Ckx3NLxx6KOo/CuUh37pamTy7wLUm1+sq29wpWWUnHfmAf
Y3y7cqfdABQddNxSfFRJI3i4kVb6wa2oOhEKroQ6Xx+aJauzwnmMYJAZj2Aje6imY3cj9HOgZMul
x9tuUaxQXf9Hv3DHOzQ0acaQdK04pKJtYxGsCEdUAEuAIcwCISajcx/B5rsff1esYAqNalnW3x59
SD5D1jFkdakKNoIQSq79+zTXFe1lUxTxoIaG5W7iL0Uv+ElVaIqiAC8eOvTFzND+9pl7sZ/OTyPQ
zRMCbBTkFhYRvPWWf1i6lixN29Xj30Ttd98SxpAx4iYD+aKt3BtRIwiZEQgpag2hxgxQQJFcdaQg
zXVM/dUW2WWf6jJ6FuAZNI2WCwdAdgGG7kQvWeejoCShsciTlGfPScUKjlDD0I28VsEIdkq2v0Sf
BZwqePWVrnPDFm8l4PPMN74cp8Oj1FNicgWxfbAGWdcmsxFuEXvENQZtR1UZtFshwcY9erxJF88o
Fg525oNXibM+pqlrJYPjG5K+aBU4tS0wtI5CAqTHnsvhkVTlKsDjhBlmzq7a3cXH3TIG16c7iuu/
vziMNwZF6WG2OtNf9ImS2yNI7v+l49t/y2UohBvCtK68eWZSYixS/ACFJ8M/NelUK9f8v9qft0U4
7paUWJyiws1pRVsP8B/UdxuA0+161fpFFl95363174qOf3jLdCxQgEs5VFK3ROGfzc70d8aLleqr
UxMqHv9q6N1t8HKseg7Pb4xln2IInNE0W/2kFozo4Gk9rr07bJV7pbrF7Pqi2yALWoa9czPzABG1
erdhj0PgQ+emWk1VQfGgt8m6JLyTbKGWsjYR14F198k5nTH6Y2Ll05zVdlFW/72GQNaOQtc1bgzV
diHlVJTZuIa6nYnNfyc1g1RXeE3bY9UwBymr2tF80G63N8kM8pK1dlH5GfNLEYh8lKGNb6G4FnFA
ZZrBecSkHz5+JJFexd/M8ZxNnqPchs7NVRzwPMsmrXxJIq2NNGvorrazvEUgF7Uu+FHRghp6Trcj
JVfPNxB8XX4mAgkuL0L7phTdNg276ftXgFCug6xnzLxNy91FiD4iVJIarcbuwDykufcRamzjoahr
d4HCBUj43kfUlY82c+YXN2VRyaj04m6QvMKgk1fQyug0gp36LlC+TZExBCCDzYw6fCKm2sjfVx1x
WPKcCgzP4tZECw28tbE1DG3rhc4o2ON4v5dN24Zyx0MbTkOGEsTLP/piCcLPKvP9Rf/N0ZHyUZLT
Df5BC24kTUCt2MohUPQl4GFVpMeTRZSH0mb+/clf2H5Z5+enKnp6XHl9jtf0zckej6FieLw8rDm3
2anjk39Zt9Q4MEZe7LlBDiny1896QsLy9KUQJfZmW61LfIXNKIuWYkrvg46J7y2UWexlyUs/Wpoo
LhiIpYpaZ9x8leTcwAJzK9z3bTbK0JcIg6V71pDT+ee2bLoTqFB+xVWE0dFsZwrTLvQ3lfsZX7p8
NRcTNHRKk2lNOL9hS+wtFU/nYL7QquSOu+iyYw7M22WUy2OP2x+BmhNZBLEwy1okyEcOFG1aD6D6
KlsY79zPWgWe/DRIIJ+PPbw/1YqEZbLgUe2fqAhvyXefVAVi4FceunWBHAfkIS/ATRE8HcgBE7rA
YBg8HBCZXyoOtBO2x1tT8fRKTZSjh1B5k3EfQBcijpeMGdPjbU8Fb4bRFHe4pwdD0UBvTLqJqisZ
gQeshXHRpt92ypRLLDL0oTS7DObrSYfVflaT9wrMT1shy0qP4UN8TMM3V/49GAI9z+pR+coV4Ds6
Nl09tiVD/6b1Q5lmQj0SXU5TrP90ote+pNo/ObH3ZHQu73ln9yCClRtDN/s3s5SeDsmoTi9TaWoR
7q8Q9NJMsCyYGO7RUa6QI3D2jlzOWRShhde3bfM3J+Sg4Hzo6nkFL9WCL0ixj/lKDOU/MQRjZGd/
F+4cSpnM726Uir7B40gjKtMY7RDI3HUsW4WIqPtX2+FoL3tTKzWywgAJ8ra/HtpEyAQUVmWsgcrS
KHzMM4eZzWgh2f/AVAsHzXDyYHYqvmhTa3rPivrB0aGD8iTtJhvK0OcDnh/2S99SIZBAgFOQN41g
m4iTNxmfOMc0jMR3yK7yWcb+my7CPCcQX8A520mONydxVYHmw1gqd55u7j+PMgYH2ov1SfM1EEVM
+y3FsnwSFNFlwLjtPAjJxz5/diQW5Pv1dDcP924cm/iUXbRYNUX6y73krbvMVu0aVFDXKYVjC54O
3MtJvsrvYmvkaKtgkuEl4/AE+v+HJ6+ww9BWxf1G7v1iYTLGwHiVG/Gp5UydAGo2itIn2FE7Uoet
kjXupG14bZ4RWNZ4WXJ59wJOH2FNUwlzKvHOI721pQwr/gCSg8mpfgGd4jxxHHvj8s3EEN7A46PO
qJKrzIx4o9nRT9cSAMa0QOaXFfcbB9Qls/sCKFWTECOZLwHm9uEj7wBn52nPDfTSpkNo9sQBkOmV
26tlBQliaIpVxXDApy1SuA3UHtiNxenahQD//LbmMj8dWM38YBSWEEuVHxMrKgaygLOjkq/yCK49
8SIyjxW4TmjdJm/06f0RnJGkvC/D7Jr71mNhNJZiR++RV18vtKt/d8MyVyBa3g+MMtZ/OGIBJ4WI
C/HCek3sP7QqVDfBRvt++WDE5Gy0ld8cFa3GS0t2rd5n6vsJx2puTAIJPfQe9HuMCh6vT8dzfp3C
K7qxmmSSV8bySjDlvV1FhuWgQ6xbGTssZj6Bw8a2xEC3jMeyldbh3sQL/tE1rNC8bsJukruoC87u
IXJ/WHEQC2iBAVUd9dK5yLJcbTcCv4gHOMBgPKcWtr37UqU4lm3NlYfAHLqpEUHxL69o0yc0VgCM
w8sybbtYPjIUEjYjbGQczcg51Xv7GO5u6g5/p8W+AW7/NEGbSq7KW/HQ6nhoUskqMDiCRsslaPlF
RyNv9W4UBGMpwB+IT0QNlJhKyJCjFo/7q3jKpQ7SbuDHSIgVLNDhcHvTgeovbcPv2dbZDEdkdLos
MPmaW47ICbMm5si5+r1NC2qEV2nKiXXblLw/is7PY7DjSU+lyVVO7EfZndSGPNPufS/K9aEuuw1N
tbLVfLRgsSHuM/Od1OZAX8TaIrAXaap0pXKwa0z/+w0DFnjKW05nkcx8gIpKnoHlm5sadSwylRkQ
/1rmwmkkwVFdnq5hgSvoFSs9Y8QCFBxHeEPauAVxY9h+93EmYHr4jlPnfAkSkkIAA03FlrjXb0Aa
CxpIW9dvFfpnFgy/JRVXn6qdaXk/B0gziJB0F4rJI43CYmLWEyLmmXCqy9RkBphEaOaebgYFZTBg
F8R27PXi4NWysgj94jz2GGCXvfKxMGaDykwC7E4QwnhuB1IiuAgh53z9/+zsEU9UL09qWF5BxZMD
RnVOfEUsgHVqXToeKbL+IjCtdUgOazGVU9nnkMu30pRoS6XkTH03KI3FKzzHweDw83oiXedDqxWy
sVlwndoYFVvPSeq0lwX7YF6z9It+rXEL6MIapxFuvgcZqmWP4Chww9FD9x48pJCTNrS2Ym8TkhNJ
Hk+YTS/o/4zSB/RA2t46WRSWDfQdIkidb1fb5FC2CVnGDh4d//oQ4OyvURS3y8Jkssj8cPRfIZUk
45TaP41JEVGupRNkc/u2cVB2b8KYy9Z0xCQKDOJZMee7MKbEh8DIuV4KkyeRDSTtcZxL70MlBkeF
761wayFmpLOfEWda80Fh1Ola6HEwOpvBYIzZEQh6NhxnXTpQq1+nrsCkpd6EhAEIXFnhLlPQ0YBW
d0wV3lwVu/vCYM75+Uw5ra7mfg9xnXGNS+kApjoSohmovaE73wmXOZy+4XKxSvXMYY5lfUUkRcj2
INHC5G55HitUW6DwMaYmeWbhnULsqg4QwsqoMgX2VsyTcVPmnGvMQrbzcf4Dt7eQUFLpRyp9mSCT
FLzpJTbFt2W//HQFohvnOjoPI7y7vKOEOvHMI2ejAK4Zs+6oYcFqRcS9ASJNXpgNF2PYLP0uuORw
s2VS6dGYiHc9zcdpXBG5TEGl0CZlmSVdvzSVT9VfOJ07aUFP2U0DB5h1g4M4eZexLvE9VwjQmCg0
+bQfRIizrqtnnlNkTHqVH2QGIw+i+GRMNBQlGQB66SIuFLES9mI+2pVcn2mMVHDEdGx2XYt66Y/A
wJDYPj9RIdd9e7eOIkgDLPkTlBQQU90lBuw2pPGliOErVmeJkTf2xBkY8OOKkWYy05eWjp//75t8
HfwAa0BSYOlJEn7o2Y0ODHuoVsXq1U1yf43gMOx0FingqyqDOwdZVGKaXqmFDsYkpAfBPwoDZXQQ
HKi/TR/cCnwA30zoo0P+d7jbMZcPoMHJD56soelQJUsy6UUSh3WCiiyRNwrlUJKbjKhGYDSEUwq9
Mjv/FBcMII6B+glAEHOZ8vi1QiV9XWRqyymbpKOkJlUPgado4Hem+f4mFwM29jkp931KRJ70i0GF
K8EXD0lPEC9OtYcWTB6u+7vEM4SG90oEk3aoj3q4z7PNOLTl9JzrMBX+ziqz704EeUV3bmqp6Q2h
3IJ5qH562cpTro76ar0FymO8CbQ8CJD+mdB2Qpum5c5/2Qh6t5hRyTYkofS6R9wUNlzIsLXMTc2h
UfsFoYlvNxL0+2qNmYShDP3VdYUtwEUeXFvLmkRuTSu8GLi7wo0KJZNiL3Nu8vmmsBGR7V3qNse9
KHQta6UMydgbSH0Mfwri5aBsNv/QFQvYR1AKOQSjYIAzOy5GLxTopoeQ0DBSLJK2uSXyFDSNS0xT
DbstyUNw3bsG9vcYWmO9KEYQbZDxhWhTkvwsiVra4TSd93nFw/9spj6WXhKBkFIQn4XZv825k7tz
ICmcge60xTNN9B+JGCFEq+WVKVnlw8/DdYmrsuLtdgkl5L2kSpc5GUMgCo1Uz1QHupyKHKrO4qzw
BDWOpZQhthM1jpXq1qtjXkTs7wUmYG+v9+KbdYZmTPtiOWR38vbUZt79lWJapPRVbbdzAauF95rd
bkDsr7ddh1Z9vVXx59X+6m/73wN0oicGpmX4uccWdY9CLYkWR+zh7QYIMTuMiAnTrbQadx/WKd6J
zK+97DZoLkdTySEvsa0CFmhgvCZq13mMQcHBDQ0xEYuKYn1L7qCLSutwquaLW1n79SX+yXD0GQgk
EFCPMbeQoMUy8JLQc6Oc30hRrYydix92yCzSSR2iXpQLu4D71FA2Xv4Rp1mMGNkp8YTsF38aI3dt
sSm3LR43kvoap1lU9Dbd9i1ehuz0+CIAskr7qUB/USMyixx2QC9xJyowWFlPmf2owXTRArtqfArv
gSko0RLzKAIovLNE24rjszFK3NRda7vS0ERIFXrTrVuHXCZXC2L15t4A2ckB4hV35X7/cmXf/Fbq
8U8No9+Jm05z2T+/6brz7NJB702XAz6X45zM3IcNkE4hxUdseE/cXHNrSgUcPcoyMSGj+wlE3e6v
MaucnAU8PpZ/6jSR/pZQThPkOOn6TT0Fyg79FMkuKtvhXFVl5Ph73uI7FIIq+uSf3kQxNBjZJbvJ
3WOXrFGCZ9jZy0dTRaKf0ESls8gN0DND8FkPcLn8IadDEIU/nw8Hlmr7ZH73nrRdop73MPs+daTG
MuzBmpS1GQy9kKGpF2hoockNgqUVklVKQ2vclIbSxBy3x4TU0ekjn7QM6XaAKS3BXnkBBgt0SvYc
LNrYRDCUk09bXYK3uWUtcuSR8l5SVDYFDkWMFffBhd0Jx/d7QlYftHJk+/OYtxJ9IWsXWRkgH5DT
5IDbKoPlfsy1mxP+AXxV2mxdIOq0ZJChot1ujXXRPhijI8kDn1a0y2IOUrsDV0M4VoNexpNSGmNn
XSqVqHpYPma/cC6OU55XJdH8vmpY2nHWtVjmLqFVu506ooX3DiQwYGFazhdFZSjP0Isqho3E3vU8
jYMOrMDCIKLeS/Xw6iFl9EoelYP73tL9KLIci/FU9IwzSDVnENSsLSmAj9n7fs/P3etLmk2EgE/c
9pEJP1aHIC9IjpiNc5JHXWkYiz6ZoXRO4n2x0effbyDmSpkr5tXjZVrTJfcFk5HBohKdwV7JLiUd
G+Eg1axXcOFBw6wJXEjauyejip4cG/RRKc7l9tBA18FzgrPQjR4dvqLkNU3gYCmp+3NHJhqJB3Sj
0SbV/DRhMfdkWlQYAxOJ62suXNzSUWXB8e2lCZk8VqkxOZY8cjZoLpx9FyVIIbb6lrES46fh6Cs0
Sbwmn+Rel7Xoqd2AAEc4jwkTFOQOSftu9sSNVBiUOPVGTJAHq0DtcW0Cdll9W0gGV2ysiy1c3J6v
9yG7l2HIjByESWBZqBQD4LLd87Tb4/hLBNJmziFIIvVhveFvcaBk6cpYnInOOJa1zTUIszV7eJOl
AatPTdp+PBMCILUMSibJED9Ppw1Pzm8kIiXaWaJXTvYxCHbRXYo4m7UejgBOZAaKXRNDEHETqJ04
UqquNVEutDljMQERyp+FUQWNFrRM+SZAoJpihfxMK5MVe9Mv48JnHDU2lgaqmmAzwyMMHYaxzz7j
kvUseYdpQffVdU1rd2m6OhkolKhws39lBoN/I9W01HTJuC6wzZbc7Wt7J9XN3tBg5rkP++zsAo06
BEIl4Eh1LlJM0H5dlYSFvW6ZxIhFyQTsto6+3kdkIH5cPH52q9p+eoRvWOXGUVhk5XfFFBWv5QT/
fVUo1cnmAzaqCHXlX4LbZKvp/wCFN+TmfhN/fandWCOjY2MzToKzJ6q/rCFCHqbLotaX7Xuyb2SL
BvrfRYcA7/ppEX8WsusQ7Tl3OGlFCKJrxzSPSdsHjYy8ZlatPPP8soH1YwmJlHngEsoLol9MTWwI
4OEdjXvVhhLiOJIq1+ssxtFwTw2QGwBQ5TnQUpIfTtzGmjYZJi2vYOXZsQr+1821uqK5V54B3HuG
XDvY/6zg9ukL73AJB27PxSlhDGRc4rUmB9VCn9+KZqky4Fb4XX0FcKciEvqWjqszP3XyUKhdo50a
3SotYOPwrXXAYrFwwMrtjC6UFzP9BksmQO8nSZ3/8IaL3GiZTIG+kZD3izcSG2T0keK4EEI2nLZP
Em99ZfmWE6/bspLeMHuEi9MREYCw29dwGdvwEytQ3iGJxv6kwovUzY0k0u81d0qxKyBWHXeda0x/
dA1EQEr/3x1E+Ag0oBbRn05Ko9t/2y47P/6ynZqiJVJxnLux4J2znbE+CMUX4Rp0pwVQY/GxtNlg
osUhpsEGFAGff+L0qZLHbjrzVwlAg6OGmVUkvDELtwhpFTtrhH9g6wtyaKTVb+jbgMNe4bOziLg2
9XlJfMisZdvp03z1196eYDDXKYSRTL4pKNGqU4SUN6Lmo4bd6ALCVYvlYNgh+z1wFdvXmp4FuyYI
uTrl6Z8+SiUEx9LGqownGvRSoIH2vFDmPDaoxsjFNOhp3Gug89rn1ZSSNbrOl/z0cH0r98eNMXk5
p5F6L2qOoNRsU5MmiLZTXRL2oA+P0gwQK4x5wzGlM5QCLDjbvJoT7q87O35brDYdhYNWlWMilfLE
5n8P8SEkWkLqBNY7z0SggmNv1TOzl1pUPQMX7OONXQ1BzsO2eplQ36dMOVQSjFzMUMYFY8cNiA4j
hlTYvLbD+79/UZ9e/LNpYMMYrcBqp3XN7vmwILQzraQgdbeBKOmpimBBFzjneZLhsxrAc84wTu/a
2BeMC9QGjOyJWvcDL7b4iJ9hCtJ5L/iV615DDJlNQMRA10BXeWN041jClDr0/8zkStBDzoJveUXV
h+09zySxdInArNQaIOUVWHgSgRHA59E1VU+rgvyMteLKKWs5vRHRbEWyoXqQ9WScztwTZCbm8h68
ijkzMwFuAg8vYsT08bZaxUPeL3mhKx7bSMsxghS2xaC9f3w51TT9Yl2BBAbu+/vdHBhupv0zKPNn
oRMPVGn5npzNfalT16vL24sDBLqb799lOxRMO3b+MmY72OocaZPuCF2JmiGmtxyD83rPIeiKteYD
SDbACIFw+I9RJ2wz9F5jb41uvzfGvuGcxpkfpkucRdUVSjBz7LsKFMihsuApoV7b+heiZzy6NLiT
2ehqUl02RFZJjS7w/2HJKsUilcls26EtAnYmUsih9/7zpDMlcX3NEDGAVj+9de3QVk65R+KJNbmh
fc8ywVRq2xNRzXLBddof5R4/71JgQk+0E+AmTq+LKph+MiahjO4jnRil+UHpiiwfQya8rsAAInqf
8RttLSb9verg+VzQF9c5nEf/98XaT6FSSOmg3W4wI8BuTbX7pwe3N7oaK/eUBXf/Gk+ndAumWcXF
PecVcdCZe7u8h+SVMAsOIgofkx7P8zgYFyOxbcc8yelPku+9tSs5ER9QX4CAKAi5yjMOuqmZbpfA
m40X29DY5zTrhQXooCNBASzoTSSzFR+Gq5FOUPJdMn1NW/Vm2+HHQ+n3GawcsE34uaf/rlFsyz3F
4DLy+U7akF7AQey2c47PukGklHnhduxS5rUY6i4D1uYHciMwnNGWRSg8dZgO0eltkTXY+ebZOyCL
KdQbtselNaMSmUSH7yvKKk3tjRZKttzTw6D/0cn6V9SaK9kHjmZ3oXx7uQRiIGxsPP43zV2GP0DS
3HOFH84B7xVWwitSR+1jkI96J8WE8mX20FmYIDF39EgYbUS9WivFfLdVwQCZdYRJen75L+pCH2cy
5apjQkIB9vKAl2z5QUlbOq3SEX12QRjWuO2JYAjSWPUe2hLaOuIPEJYkH+Vz9lYpsJF0Pt6Ct1Jg
MjOCu/mp7LKQg6+Mh4XA740wQpT56iQEyG5I0XEscsKVF3wKpvxYwlbcuyqFFCSJ5bg8jR/2Kek/
YKvuM6XV+cvTA7WCh3nqTfewIaneA5P3mcuZPDK219xyTGje3bAIlt4mt7BFakEyjtc8CqcEbfEq
ZVzRiqdCsnma2jS487ah8oRGgdTZusOeKyfXM5nXd4ROjmAvf4STO41mEs9ybf1ozryPd/R80WkP
R3ZnoEk8L+2i7spx1EkJ09YOJ/du1KSdhWFXBUg+YPhKr5MXirSeRhq/EWidoGW1N8FkGNarAiW7
Jt69HFh6cr06Dy7i2oJZc5/vm16GLkuKyOX/cUG/bSEcVMrftqkFs9bIxguOnp7dAJazjsKbr1fn
wz8YQs8mZFf3da4e98pZQA6JTtojcUuZlgcO+9c0G2WWBrQz/8bEWGPDT+I39iNsVA0f002NB77O
okCnFDwNxaFUUglhXy6uInT48AQ3H0bzAJU7fvB2jYqEzGW5YDnM/VPwzYYVeFgWQLLHxkWzqsRc
GUQgF+1PqUMscCA48Jytq6dxOxW++H7Olgs8IKFdaA7My6qDDKn1QLwY8INCTbv7HIpRNiO7qwjI
ClqQf9/ShNp8lPhqJDz1hk30Srm3u4Ler79M7IzT+IFEyBF4o7JDedXlK/LuDmXBf0+1el6OQv+P
tA4YcypHTnvRGENLvbP8apTrjLcI6BUgtbLr5/cGnZSy5rtxgzn20JG5Hx4EbjN0CdUWuotJz9HA
pGydI59rsn6p+5sYWWwn9F9+SpDdxdG+4dS1blRdjTa0p1SyBNK8E/x3GCWtXYmbOVYE7p0oKqHC
m31m4Lc6e1BYQ9phijgx4SRbCyOZ0YVL1zDmgXktFGHnT28Rj7XarMGeGcFhdi1yygz9zAm5r7uV
NnVHx2Mx4/0JZU7UrKOtFrVG1LlH14MVsDIZmxfIzDXtDaEfsa/SW9i7JuPYSMX4iUqYqriV3Gn9
0js7/i/M9am4KTzvwJX1WChbyW6p5Oz0Ra9bVixfTQ+WA/aoD2tCWxQAaJ2BKAJ+qmE5zm8EBC/T
rNtQccPaGQHjFt4clEK3+4F1wo/OGVVv7BTHqiVW9fiVbroFWHfsA6/lvbfCrAbGutOCd5tCW6rv
mQlr62sU/PyVYsQEq2gvCDHilQl2zeUEzAEv3uYki7hRj/firI12myP3PxzgPx6KnushgXhw3dbv
sZp4NmB3HiJPMYk7Kt1Wjz5/5TQYsjYA+TsrbMXe6D/Y2lxfDkiz9SEcpflSVdusEty9litD0QgQ
0uzzOs0nXs4Q2pBTPK1NMCGHerb1Gq4Yakg2OIEUOnK6JTJA2+JpkWmIZPTtvEtQBFA45RCtC6eS
q9+vtGouNJgf9co//9q1df/KLuszmkYc9guS57nf0UDeUPMpr98fjML6IrSyv22x44+AZxlPJSo8
UYnCsJIdUTzdeD+biH3QTmI14+DEHUibJaVn1yEaWjpOs0lYgipxxQkvLzx+ZELjY68t2RQ3g83a
bW+y4v08lAzaWgGev2m4E1DjBfic97ScKuQvLUaaE0T9r1sDFuYeATiyoFGJ09MrQ2OWLHK41cQD
i732rvxbi6MF5kcRb8LB2uTAxc/H9WQgR3d54zKmd1X+ecH9QgaGS44Vbdkjhp17GTAzqoTTv5N6
WTWLpZ007gFIFQAx6y/6F7LvGgf4TzY1zY+WuigdwRvmWHcA78DMGhk+3/Ow1M7F/wiefp7glJfy
OsYbp97eAaFWKchR7BaPPzIxXK+1RI7mP8eyengYE1eJiNu/V2pSNokrOHICK5AprA/8I1xoO76Y
8J+KcQkUKee8vNkoxCZFj80d2eZhT0aeTtHNFWFQNjI6VmEZaBH1xKleLXagzzVPIRfLRetyMHZT
xhJ95Kl5H/hGx51XmRL2s4ZyY9Bx8cA9nD6HKNvgcaCr4isI/IgJmuaFPoZFqqyHIWFHFCPeDlkk
kJ72vzIzBEDbDy7ONXnL7ouG9qZh5356Q1c2aGoMLt6cYmzGvyLS0xUzH14sSfe0trvRVAYBA1tz
i0h8C3QKGYbfVCOij7tLrLQQvb7v18Tukal4TFs3jYYQ0MkO/2+ttc3dg5skAzEVmlijfP15YGQf
DKN5g0BZbNwIzpIkgblSg9z7CjY6TG1RTpjM2oU1zv3z6kNLx16WEZ8FmXA8YoLs7kktpfXZmft1
EjOBAvhIE5KMR8xxMIUICikNKjKCysMWc9FP3MF1g0PQEtlxd7SBytxiC21xd3YUv7GCUT7u5Zf5
dy32h8usytdEXF06LCTp4LLlx4uewgFuWpEiVlMV+Kd3zbNe9wrwkB40X04Ob2Kam3nxbD7IIBWy
P09S3GBXYZXnbY4ysaRayD0d08dOyjJFMQAN9LnvvsUnGY6PSuPDhrddyC3ioHi8EAzawJI4V4B3
QUAabSGJ4i7nvSyr1hkDgw0TozhNKTem69lHTpzVnM1ChIIh64w/i0hnOd3u++KJTfMeo/REh2Ic
pyh97YRKmRLmoCbTKDo0bB3g/jsGnWnmjkVT3vw22Kp0rggXLDR2vyGsogHmrgfPj6o/MBkFjRzZ
zMO2m3BADMyKWNe4/vMsrwcfVBfX6uda0D9sS8Vdk8BmVAYihkV5wNLqS8+AwMhtB23GeunWv5Nt
/WVv9lkw02e/BusT8NlLpWF2JEqTwSM92O1X3JFZvdag1y0nzNAe3lCfwgzpMf9NK7/eqHD8Sz8s
XiSCKIs7pepz89IZk2UpvRMREB94xIlD9KrKVkOM+WJi8wb2M5m62/l8KbStIVLDp4TX6e0SclNq
82R3S6puwIOx5cXYu0uacKmebza4s0wpizOGRhQmJcfHRdiM+/kUsxEvaMEaYXn+OyfsX+xOuRn+
xV98WbQD4oohATGNXbMHI+43uhAL1XrcxyugLPqpIlRmh7JiUzEMqroX1u9tg7nBDTyhAgpm8VNP
LYbIwsVcxGEBNC91IpKFcSUbqXSru1Du/Evzx3GgDLhAa679S8axs6+/QnvQcYtzxxpFbtAZBL4z
jCD4c4My0XuT1oDzIIKjHChQAkkGsIvOzbKcWxzI9G6saScDcDcSFa8ZrcAutZyqwwTIEK+Dvub3
zUFK6dlqC2s4HUVe5WHLIUi/+iMsi99T9N9jSfCqTtcPH8cT/vfpyXAIVgfbIz0nwFf39ybOBNCo
Xote0OZUQpVbDCsirXlztk0Kf5mcZDPicIHdA124Q0MUa8PDxzFUySBJSkySj/5v7mx2Ktw9o4MI
lMOGBq58+rCMd4BaTQIgXcwB/O5R596ZdpJcvAARbVOpFuR8X2S9DmkdSxk6XA+0bSTQI9h10vmW
A2sUPMufxJdZGnj8znFjvW4H5SRKgi2AREnUgFvC0R+THRJeOJFhOAh+Ghxm5FHcLysETwObSWDx
jgWUve1zWBU1XC0e58v8gwYYH2xmiuTCCg9fpScw7knWayulugDIW9gNKgd2g3hnxdreWaHfPsmf
Jynyx8Kv6P4Jawqg9HMpKfWHYREDnLqF5GJGA/DAP7/OeXUEe9amTzqniLTlk/fakjCYgnaGjq95
XocR9NJCqh5dips5TzoJjzneXMYTwSCPPnUbjACiFGaKQiN911wG6yyjqMpYUJs12bXJ9EpmZXRT
8t4V/zC+0YrxnKSXeaurzvZ6sm4BN5j0Z7MLpQ+i77chjGDIB1MsO+tQfyJfAwv3BFQWFijqFfBF
Yh/ZFzJ64mda7cRYmV12zPKfvm1OK9G3MqJyjbIcUQweHaP/wn1aAZPkhNxM12NCe5ZeorZoRCBk
VIBu+A4gxOb/15mNC++Dbq8dGXD0pNdtdaWgB88FrtmlJHAk/eMAlFEe75aYG0PidwgkpJy9VUrC
LfhjTheR2AMR1GNe6rCj5awuYDhsVR0ewmnN6QSnLCuRgX1Xml5uNzBWXlIelcl9qpG0vq6D2k+m
i/wL69Qf9yPRHlygC/+yo/xbDiqJxknNXqAu1FohUk/nBzxMIC9SfEaO+91QCGQ+kJ7NzVzwqlFP
5orIfVawe9puJqQnl8QZ2JhjMBu8SvqDJ5sxcgVR35Gj3NW8+xyvZvGh0L4Vwbh9eBPlcMlLe0ji
px+Tq49CtHNpCon7TJh0HvKc04WhQ67WLphl0WtQDiP5NXUVPvQnzCLz640EhOJYYIRyAGBI5FMf
uPXtd9nfGENltFfC1UDByUD7DgVxZXloC5otAMKSlqGpQRG6lHbFTkxYh7f+uV25kVBfSnwaApUR
UHo75fXQPAPEhk9fq6cTOLU1fKzXRkoSM2uMBIqP3O91i4nJE6I645CCpyTHCP9yq9dnAnQt2KFS
8hZDj1fEEAvei6vWL7gN4AeeN3z8xcvb994mBE0P729YRKD9ahV1LYR+KiYrLeuJnKz+Kg0lw4G9
wx9N7eC+P7DlWJpPyZdiGNzy6RuOJxDJ0IidB3Xw9naiTJni93Esl/TKg3YyFrEg3H9V4pXaBk9d
QcdoFJBooo3lHovul4sZoXEvvMGR9tnoIpVp9RIT1loOu4lMSHzeM2C1RkGyjbhSjNlDoNw3KLi2
sTHHSb1KnObLORiBsfAIX1m+MM7AQo8b0o+0Ljx3vQW0lsh9f8fr4h1dBCPEpJV//MLw/230h6tL
xf06pmksJIy9sfIGk8HXekxGOS4PSIO96Gssk1oFNWNHR+aIXDiUm2ynffnN/IbBYKQ3w9u0z2x6
2CgIERUdeCJDodNypBWjqIgreSz5qtPYatrUyaG/r5D9arFaoNv9uueJYeM+4OwrDfJrsDeEyXR1
gVekMTJtiY9vJweDtrM5fOiJD7Yv2EmWfeVxlqspEqVw160+HdsswEVFDlbIT/oJllrsfvSUtAkT
tPMaOvBHEW8YKCC+/ujm8okoZYqhH2mMpabJp/a0p+eVyhoGWWJ9p11h2wngHjVS7bq6fw3iyUMU
/RR2a9vCGeIn2fgxWqlhgb3aEjbC29FaPqHLLph+2EZpVkjU3WCvFw5aD5JeJLzcLXz8Q16urVGq
fu9DD63mCxohG3QyLExRffVJZSWrv4KEcxHV8BqBk7b4p79EJnw0/dXCprL6aOY1CkyBFMoq0XbY
nA1FtlKI6G8jUmXpnx08jeHE6r6G8GmizATTuE9F29gsbSdSuODT4DZhIdwogUBUtcNTXLPGijEi
Z98UXLfCrFi38ut/kp5r9kCtS+RPIFJ0JeBtYDBjq5Z5bfphmuyOz6n+VsnnfjGxMhdcaaNoeVHr
rHta4pKOxQ4HAmRiS6gL/KzZ3ge0MqFwebGzwpOaxHzWjInIPD7ANJplmSsLWta5t7hYszOUCPWw
7FvocsKJ6shBWkrkf8HtYl4J2Hc5kqs4BbDhGBvM+qjcmQuT1lanp12F6kS4Q+G7+Ip+fUqDlTkr
4glwWW++5+9vDB+hdi7Orrxc53goZOlyCMlHUptzSsdbD7k/Znvl5RfLl20vwpLIBR777sBG7C9i
+V4YZSPOZpYJ2Jcreem6sBx50iQfNNwjZaqtRJg5HP4BD4319lOi0u1oKWoinnfhuxUvZBSnrcLi
8yGFXOYTz3xXexbjzcUYLt1qYdwQRVLHEzvlkF052SliDPZYP0w0R6eCOYeiJhUcLoCrUMi78GVK
sdK/ye6QKBLk5E+ci23brhd2sVsnNeVhF+KWxZ3RGgXU/EBE/URfTKjT+KfiPtDdtZA6wc+vkB7D
joQWJijpRQ9K/RzHXjLNxiyt4DsbmyQ4rSA0olTM+/hOl2HYkgaGr1EXdYPdoVA5XTYRhnNzVxW7
6OMtA3Gy/D+g8zLLbyTEouYypEve+6F/4JCWsKYXtfHb3fzc1Yu+QffN+qI1mONw/DScvHmbEnQ2
h3uLKMeVjLMUQjemgjwS55IfzFVPXRLMn0MYk250PzS2xHd9WW+dhP6Jfu3quN6vsMzdU2lf3pzW
RKPfizOCIt0SG+pzl9BGUcyZvd6CwyQx5Aj2ZaMoDvrrXftJNOPPLg4xQ5zE70EBsjpnhOdf0c9A
aGxggtfK+ehW+pgZFWSIjhaqebxFj0UkcWExJCkdkKEr9nAPiZO67MQWXuKW9wlq75G3yX1Y8KlJ
DWt/czdQSIqLCaI79emd+To6cOJOuhbZIYdddhCFGiQU2cyJoYMmegwvoIs45Bn/yiqMR122ziwk
QLinH6neganwYQ0StZug3XONRM6efJrP3x8TgDVAzqYYmcxDqHyhQ3kUpPSk1/eUuNZDU9x8UFcI
qOq8XQgPKsVvRvrlZf13ZWVMvoL/W1DOFUNdwOGP13txt7URxtyOlH2UhPboFvmHtbqSnCszxJy/
qiozdHJKmpe8LQa7zBt66kw4+UPneT+c/vNOg+QHYDOTBY7e6a7n3eDGR12ZStbCoiKme59nxtfD
mf2h8fZgJxfbT5ZZXPIstbPP8k36Ek4czwXWEmUPpG783NRY483qrUwAMpKlAqLP5xUrKXKnjkf7
VhABJPIiyU/RIuabOJFCka3awbI1Y505Kh24geiz16xRcD2OJz4UVCQsUK/qSnTyhsJ+BgN5ks+4
zuez6pCKJ/oxyPLUmRdZsuo1YgPHEsDN0Tg2sfIz9koT35F4cW8FwrwddDzDYljNK97HbVk6UKD7
Ju/+q7EHz69SN1Q/cUylkpKR4bHOZfW4vR7oimV9Aau82hRlQNY3eSw7n6u60RZlkxmn0p/P6/ut
4yN4Jl8c6hBswMzWw1qQU5acZVHUm8yyeWcFwwasFnWakLj0hpglYPuDmWCxX1RBHOZeHWDa+ETY
eUENIzfgAO9WzYfb8diLPX410bTYgiLxrnF6byWTWckUrGDYx5m8fdcEI1lJMawL4aRGOuMwgdX0
KiZ072Tqz/38XN/rpPF2D0uTJcHqw8XyeHhydW/B3TeNQ/XiK/qok2pu6BB98HVt1c5ocP3oEkmK
5PX9FwAA/7gzDvxtYt8h2y5O/nEC4nCukcXeGyncGOD9dwupCs3EekmQP4vRpwhv/ZwEg1kCem+t
GQhLKSZJ+koJbxUXblqKhSX0mq7orerh/Yeh6t+L3ewLCcKFT1U2t2O8f1NrLPan31kHBnh3+h83
7BOdA87BcDt2PK818v/5QJ3waQsWaP7AMYY/JNKOLeX8hEav77+EuNtM4/DMI8vjzKoDIUqYsgTm
RyCtZes2IqpzD/+mZGGkSE4lYnNfy29VX5zjdd8J7xGmjRXWP0qApmIUoum+GBGm9+bxoi5e8Osi
HcTwEH3FI/PxYBDfCxvwGECD4PTUUgog+u8rXpz34JqVWryvLSyG9lBHgXW6g3EOqmSsFqd+/fkI
EFqhOTtupyyWUz9bn4yMAgiSXE0vs1VkKMs/HVN1g988t9aPCxSF4TY5xzrygEAwBFbILJj5pdht
O+vmjoNArmdFsL+qpBruhTnFnK8WwitOgc/9zXUnqUUMXkfJM6EoJ5YrFwHHX7plrSkgyvxuOFWN
dgV8zXtIwnCy5AiNKPqoF08rXdlrrqTbQr9Ho6N8iEEiVxrcwRzbrhctcjoGIBTvRFG57WPiQffv
yurDF3PQTdzE9PV9cPpPi/zLmsKnAHIFhTUpH0aUSvCgdGD7F+Zd5gMR6MT6CZGPNvBStF0KFcgb
VsZ8HD+KC3cgKRsJnR0ebLKRYn0rdcb6cv91Qdm/qFyOVMXtVIXjwtQntqz4pRyqVDRwIvmt6x5M
rarkWIl3SRNZD7YgeLAO2pvmzjG5A5Wxz+oo3dsuaol3J6bEPo4uBzVB63+khoMcXARxnzeVajt/
3VrTuXQ2RU/i3MjWLqUyRRRY+06V+LTC4jkiDbLprUebKl0xNkXz2ndyJ0DY1J+q94m/eaBJ6HRD
JDDc+3qan+vKqMC46ooSPKtIv+LRCdamOPjdfpwjwli2vTBETLlUTjK93nb4puGN8OT9GHw0V++U
3vvEuyvrjbgcmqRkr9H0GWvVcGtT+Dh3Xc9JtW/wsNjl2358AS9Vc3C8RsjPdy+BfAdvBQV4L2nf
3Ho/xe+Jod6YywLewWZx0dX8Fff7Fpc91P/ruZBX23Jp4w1p0HdCrLkP4OrX2djliQmb99UkOvlk
wSftBFUHBdnpbAwQ+dr45gdIW6zmz23qjY9mQ3vh0VUnNJXntWNx2J1ZjE4a3d9OQfckqtnrX6xD
ZTiIbYuxyPL4Tcb1WDQnZFz3787t/2YIzQmWiaAs9wniRqhAErsbndlivoKU5Dx6Zs5X6o5P/46H
lm/1qLyv6rk/g+avwPHZVhSuY69+f/4nSYgg8BBTFX85RI5/UG8elL86FYOVAq8SPNrFSaXWh6/6
LewSdd6BNyJfsi9GHOjMMHXYc79vgfmLo19AYYMdG31OaoT8OH72tHFel4onPaWjhg1dYF0oqd/i
aRIx20knKP8EmXKdEVfCNnV9N4oq1FFs/sLZuOJ3ybwNRBde2TXqDbxBZiniUtKmeFwL26f+r7n5
ZFzJa7LWJhKP1Q2+xHDY+KRC1zQHoj1iC9Z7pPHJqecpKwSnThODHj7yrjlvmezVN+JZ5dVMKYJY
H8LF7fvREb1y1H1axrZDkGD/3GUTBW0nsA1wuHPfM9myn2zAlvax2jUHaVLMQMEHaJmcmoAyQYG6
LTRfWOJCBjQNwr2OJMsuALguyW5jz3oXS4OdPGn2RBaz2hYRp/PuLf/sNN75oXJqQeOwlEVS11t4
Pl8N3aqyq2c+lnMSl8rXZi+sFN4mjkC6FuApwJHiingQoVfGU8QW2YBLaAVzMIQyBWSV4EKNu9VQ
v9ckE3hHJL6aBtHk2F/pVUVqt8+aIo5i6p2N7bJXcun5LTqMS49m7KPWj0qa41q6YDZYvz1jwmpY
f5QdETarswThiwuCp7RbotDDjK6sXRfTaYT/m0PgkheZ2cmsNbi6G3dVjK2ve2pc6lyY0KIHgSX8
MtdW41TCrHjqyVdBMHjG2wtkVNyPupPI5B9FgvE9WAirezjsvSFnWsf7ViRKovi7J24ol540XxLv
Zx4Z4M3U8Qsfkc7KMk08ZH1rmScavruJtKjEInC0iYmylDTvcvqXz0SHdrmd5o15gZjkunj4esfO
WsC1Ip9Q+5ec/neN2e9cK2dcWKP/5hcdsMcQHyHwEfi4HrGK2LvOmuosYQFG6+lk5OFFqx3NiVok
4hB5CdF+gF9giVIWPM0KJ+6b+1SSk9nc4ca3NxXPMa2JwpdttNQkOFPg72CBVGf3lMSarTvTWXOw
J3sa57qAUGGOUjtupCdDmwZrZEXX0uaIRBPrjz/Z31KAlXJtWZY/D9PoELptqAcHqw8NEFTyuul4
5gBJWfm0/wBEzQwTBXR08PFBlmMmuuoRHgdiwj7/5vbcxLO8VI5OxIH/6jsXwszWZEqhanE3KaE0
Z3tb84xbD/eCfCz1qnydrgeYntCe5ItCmFvHFkl0tm5GeyPQFrhWKZey3LFHuJZ8OiPPdbuDdBZY
s/pDoiO5q+INoAnuvlOprVGpXvccSRu7YGcX9CCias5NESmgeUe6unnmyK2vK8FnR6fbNqumOg+v
hh50wLxItRxC2EJ77y5PbKzeNyKaaWy03m4I7GwA6WD2ASws+dZ+sKNwwsTmu6qdYRr8ekQkshFc
RcHExWZODjWpVYlblTST53zzbCpiHZCVKRCZRjccclFyp04xHwEu8c66TLLzNZrYbSBiEQ2NgKfp
B2oQCsKzBRXs2W58BLa0eyM80WIpl6vvqqGjzzLuAt1jPY95Rx7txwdpApelLSkRPfPfTVdzkzVI
CAHRVAC26AyDjxz3vf/IlmAJU4JwOBMczmnB9FlZysCsVB6gR06tRvxIOtqEQEvqR1HPWIUK6raC
jO4BAxgz9YRpr96UGtrzFcILcZhlcFGGjRhTRX2B+l+rZjVms0U0D1NNHb7ovvVMcrRezwHja/OM
yAS4mEz1ZDRZ4v1nnr9Hal8l73E6KOye/kx75D6qr/y09z15bzcKxBLIJhMq3XQVfU/wa0k35150
5sNNIMZld7Q63X9CGSmNWckZ3sI4KRsVds5UY3ykPdxi7XQzUyzezHvG6Kct4Zno+SQ8eapVE8fu
VMfRVmLkNma2Lx215JgE9BFSZmjBP0v7MQrOLg6ryAw2bzpTHHFi2eisYiKryImQDnozAXOUUwVl
K1n3hfv/fmbZRYHLHq0AAWTm8P/FnuTxaEY0l+UGIKIKvd4TQcQyJ5Pz03wxez8yyal7+h+rWega
6yHqFnIvh6IqoY5eXcA4eYORoBn2QBH+2cbvwtC87qlLA6RP4I+AYmFjPnJX8lT6heVM2GjKxP6e
sEZ9jPgRMD+0WuUi1xXhuV11nTxkboTr8H+Y1JzqYGJfAe29wGOOjgGEuXx3sQrq9RjAjI1tsysa
6M0/oJ55HnEwPdpbMIEBlGF74Y3BB/Qk+qBrcxLvmdTOh+ulsbzmnrcuXUguau38AVlT4Xv/tWZO
isyJKb3vJ9l6Ui+Sdt8Ka3ilsaDwB+uiN1YG8BxEzQRJBQQqkjUZqtudqPazGynfiqpo1RXHV3iv
NHxq/T6mVtutNj+BFDc/C2jh2pvS/LAGdEkZVGO3jM/XKR+cnPVE81ZCVortREo0grluSgP+48jV
ltnvLMYPQJnMZKE1u22t0Geq/RgJcjE51ScOCAkPLr7zaGRaQqZBAYVopiT2iFZE76ZNPTWLZ99A
TQbAt3vtddRyKn4XEa4jeA0mILIEU/cj5ZDD9EZlXyWKF+1C5nj9DKTcafyuoYPPArD3aV5b9rTp
PdT3AkNwU6fRbez27V/e3aGxtPMEllNBbZ6n+K3+JasrDBkIdYp6TRPKXYYOUcvRcWnu9azbB1zU
+xGEELJS3+KUWnhNsqXC2PSwDttEMGOWsZ/xcXLCBRdtzXNwdGSh64oxaxiXESET9IOdoqhZ7Dfg
G1MWqfpvlPuNqE3Avf3Jl3U35gKtGxIGdDMLTKv2MdZ6zQnaOZu3aF/bU+lSxMXUlmJiDXrlVYHG
C5To4/OgEsUSIbmDyA/PG1xI0Z5l808lOTSYRV7COwnAJZBp9tA46NETdJOeYlUD6Vis2KEgE4B/
QXpD1pj7hVpQjPfVGzfl5Bxzbu7vBS6cq330mt2szFeSPQj9K7lGbfhln1LV7OfL7ZqModiE0AfZ
+NIJUn/G6BkB3Zc/MUNsJpKq/4Cu9R7uBTT/Pgn6/j1N7FoQjZVDaqNXyAYM1v8FYQe4oaGib1j8
eO9/2b/A+UMhGFH+S+G/57ytNi9H1l70RKS3Tr6OZDf6gPyXyNe3pIWBHdiDpPuGQkG5B0XsFx8m
4eoDchi3MFQkfaofH9cEcQw14lOrL91/2Rpks4H5KK6F6tOT16VLPmTTgw2pOfGn0d1h7JmGecz4
tZYMQNpukXm8RTrRhE2NSIr2AkQ0qc3FiCFX42JpKTrhzDe8962HDxBHiPZjWSAzUW84WU4iYW3U
VVXH9/zO8NcWzxG0dLkkQWJ0EAdvExlOJLXa7XQav65nIWKb6Ux3bqn/UOJgrcksX3YoyDpt0B9n
340x2++iaC9YrXOyHF0yG8diPNFv56W4WUpNMUpA817OeaXzjpFlWNUnUdzUkCqjhlqtFRwXdp/o
8+AIRAwl1h1k51mE8AgVnOT7sQU1DyscCUfastNHEgClHDqTHvarEFHZG7Sc6AE6oSY3mkOJhCnu
YAlVf2JXRt2a8xesPcWUSe63DAq5VPigkF0OHQmlrXOmcPYGOyQ4j+AMo6kMvI0F0ItBsvlruTzH
Ejxk7M+Ufwhzpk4QAHF2YJNt3B79bxbVIswpnU8sTkL1jp01ZmuHaHNomU2Vb3G/lQjUVuZkYs8k
XpuofvSdqm95kiWeQmTJq5ATtFixm1NetAl/CQtk+rssDVJVF2taqADDOVMOygH9r0dKs6+XCWCH
PvaZ2NrNbz6FKuBfVhfJPgpekIZgrhqwB7p5YjbnyRgG7Gf/HLdPsUz9+qiApJAwF7wBq45hhWCM
1Nn9wXmxq15/f1LSEx9vS0gkeWHwcBYSbe42AdthvcuAOehTNs25Hv73kSkkcbH3G6DFHhIiy5Ec
UtRbRlFTIzgcCrPx53YaXA+My2JTwAsCRMVgj4IMdvvw0VR2e63pB2vKcdu0fmXTri5dnAeoDLEw
+ruJh5JuCngfxahoYXG+DWp0SuDn2atIdydsEsaZkLzrWFBw4gcqybv4J7/TkGmneYJEpeaTt9QO
XnprASzo0x5qRtdi/0R7lViLFfYE3N1MictI9YeWNCCFH1pl/HFktMTwZFdfn2JGCx7jpwoAHyDa
7k7j1pFMOJLmUbv/g0OGWz0c5k2DxuwGkHcMppzWAkIZ2TwOJb9GsC3c5TygtrCu2J28r/62HjLR
6x7OMzP98CbNCUInuvRHhgPZlQr+HJNc7eL/9y2W3gcpO11IVOkKG1RPGkgPWnQGctWyc+8/3dTj
PezBoPQql8L5tN3nq7+NzU+YuZ9PAcnP//B0t3sDkjbKz04LUnru2c3slA4aiwlVW4W7OBUrnmnR
jodlGHdmgzD+srW9pDMAJ5SXOSMwPjA0FaHXiWnAw/RJVh1t6wcC/RIocSQqazW/440BJyhXIqMN
eI8k2yHGL7eFvAQ0MGUZy9bqUjzU4DM5lf89b0jtDyiqyJN93bHmoqcZNwz+T40RbHtMJUrwEcDT
j3aO/kOfZgbYLdhL6xfH19o3TiYX2fZAFA/WyyKoiP4QC9dkbN22Pr3O9ugPk+nSJkRkZxX8u4I3
pMXccRD91d0ZSOPbG7ylFVj7slCineLkXrsMcZdvZ0xRMoCZqYfb2kO3HeJNJe7HjdxecAfNZJ6r
z6OUiUUy7qeQDCKYLcJYuA65ERVflTlhpg2sH1TddWth4u9gM3PhyBzMfk5J/OACsYiSwMBWkH+a
eVpoErXBs3kMPYRqu2Qs35wYay/SbGIaV6r7L1C+0Ysg/6P1KAs0Kiv05wVN+saxz0xh/hrMKI0i
Bj9vSdWbGxfWCKr+QkwgdlXX3LlFuAsbTxDIeTw74sftlz223/ASBpT09ykrRLpPZ3LLcKDL26w6
WQG2vZiBkOunYSC/aQ3z+DbyNqdzohcLhr5J+FLbqlWsqK5/Q97Is5aQ9xunXjUY89lHxRaSs0BK
dfZ81u0FtQWq+19Ay/ZGnyraaI+fZt/b6kn89QRszRVMTd4+fCOHiIVl0CB+FCZoClc/oEshfFzw
sym51m1p4KbevP2fRhIfk2b2bhtZggS20v/Y9atdAYkSKV3TsPmuuiBkNRvzJXtsTouKNYBa3H3c
mUMDTwRlNgC1DZlht7zfdXZnMGzMXiQpUhQzy+vXKnLMzXsxt4O7DNySmERi3nPlbBuhuDDPBd9J
+4pwg+HxJ+ofKz+hnYQM54pFSyb1CHBr2iA4Uw1pOvjcq6JVSZPyNwVsZrc6t0nJNM6bE0n7lrtf
0QdoQFxyBbG5UaQX2nZYCibDB7uHvYlFhybX8YOqd2nG+8emHdmndwHuw+sWVD4Rwk7SIxLgnZVG
uaExQSOEjrhULeGA69VcGWuuJq6mkICYEaHuSlOFilnoG9REpFVHxcrcGqybOYU6mNKDk7z1MMiv
+yQoHvKPG7gQQxIAFAF802411gglZlsLIqyAFRoelXpwxb3ipovI+H62uyPrUhqkpcLwaL/pw2iQ
0pkEqFkARhKjHuyVXbFoWtCmjz5TjLoL940+W3UyYVd8HdfW+odmFOei+WE3JAXiluqHpHsZihu5
KKYV1fAQpsd4DSFsVevF53blzR8xF/SadE3Zt6eB5XOJMg2e3c7t8qgVEKYZJOpId+/aKa/3HQ9f
pvT4pWCfCHEbuDQf9VfB4HpJooo9DusJQtm0LtHY5D4G06aMV/5hq0Klt9BvADMIKFU+xu4uB/4l
X6+7iYgzVWPQyKihaQ6lbmkPDMm81+CuZJ/l9M/bRdqQ5HG++XnqTHaMQAbMn/cN7HBCpfNUVhRi
WlE23edAQTyhrmZwbKhawKGrdrWIaSOzwv6bjzPQykOTiKqsUQjIxJ9MBsxwu/k2XjGDXOAH1TLr
VEfmBq2NhDn+1VR/I/nqUW0Lpud+hYP91W7erZEgpx7eFn0m0uTqGdtH73GmccVkosD/hmU3iDZ+
Wcg4lTNkNK9/QQD0MQLrkIL5BanT1ODKEEpxQdn7ciOUcNERsvwqkv3xxIr813EasEWwuSzaa6Zi
xXItiU78AMp8VdSZplV7WqCL0PLZ2cv3R3+ZxsUF7JaSLgza08AB7sKfCj1rcK42ENuYWfTQUEl+
yKgR4p1By84KVpqFUKcf9gz0BhC6JAz+JrZjG1Kg6+CWRBLwkbLRaBCh4yF8EektnRTNYe61hpOm
Mj120Q0IWFW30wu8zqYdPHZ4d/utLYq3GowkCJhTI9mGGqpW8Kt2p+0AWsy3LwjL88pkLnUpmK5o
Lv0XSiZPqKDi33dDWphwwUT7Kh+INsEyozSk/Zn06jc0gsQy2rbj1e1XVUj7f7ZYNMDQWV866qE9
OM3+uNcqXQoP63lhXVYV/S1Dg2Rub+cupf2EyeuthAIHcgZRk7D3cXUwCKa2ILFuWK/qbzBlP+sP
zZW+fATHCKHmX59Fl62GgwL2B0dbzEt1EBwCwXaiKAuDVlWjNGSrkv7eyJH3vnbyjw7/fQhY8tmf
VCPBLsV7BTGBn7bXvJfdI9OboAJmfHNJbylOdvrurlipPYCmoSVrgszBkVqwlC/ipF9dbYlfo260
gbz4R/69ZA2qYi0PQG4TfVHkbWVauaZIn/Jw+XWklW18MBSNWQSPnkMa+ki40N4VdXPc5hAoUjQI
JuYhgORJkwG4m8n61d2bss9HCqKk0HzF0jkoX8qSD+jB8dw6S8LxxuGOhDWIslMagqEPLi2vkInA
LUvEnBwbgwr8LcCqIYb4qDXjI0yy7HLziEu8/V9JrzEM3P3WNfYXZ+LOI5XX6qpSCsfH2ioxMB4X
6DXVGWJFM/ysYDtNfOVO+f99t5FKPlOAkRSo6qhovsMdjYhELtcR++agbKaDbnG8cMfYqKwEPaTk
qOG4NAAL174UmZj00jo/G40yTSMm5oo6kqhEr/l9Up4Inq/e+/YCcIE4ATkOPK2q+0NK6u1ia+Fn
EDV0eC+sNz0rF4zypl/YfKdSYP5UciM/Ucl48yySJFB+EZJr/2erNBCMp2yu8e7JJpCiQpRRJ6gM
mydRiJYlYhuZSqiVnHjAQJ6VKadXD0LupFnNOTlU56a7y7O7G7R1aqsMABBS4aFgkz9feBEzXjzp
bHmcuaAI4FAmGlw7M5E4NM5ks1S9g/dLjky3UfW4dKyi/f0hgQa/HIT2i7E8ew+Jx2gVyQE8r2tB
J/15JT8+4F+K7qX+x8DZPCk3V0P2E3W5PJf79f/AvwR0iKUPRyIEtt1qzuiB/Io6qBTcPrjyv8Ah
y/Z8z9PHVdCg7LGOOc0QT51uuznQ+Ctk0fyRHocsh5iP0nvp/BGp97DHya7InPbEx1kHvSUCQIXA
DvZ1gvLquzyW7UaZh5ECNxYLJ18VN/nDSdQLVRijTg9bNISP5VqgyE86dBN2fuTFfQuQU6TEv7z1
9baSvlO7UEK4reOjiG0kUJGb+s/GfZTwx86I4Ae5Pghal8fjB0mPCSaQnYiJpWOUvE+C9cZDnoMP
ymStuLMigY2QAlMQW0GAAwV8mIfwTpDmewQeHfnHpX4jFpANJE1vZKAbQDAKORMNe4sYjtmiMZyU
9unZEj5rMAIZGsRgA2zMjIFGn0NNZ8eE78MXupXw21id66+MXb0uEsfs0fieQq1H/v12dQkaAaNi
oBgc+91gNc/hVmE6FzwwhqvmTqlPDK0SndTVIVBKLQdJ1ao4wIC+LYb+XvHzMR+RzylsjFFQi5d8
70x4VAHE/sHcfKRdeJt7yaYRSm+DF4tSP9ipqH+pFvQfAFPubCQtjqFn/TnQvcWS8Eje3W+ne27w
Z3vJp5FnfkA1zJxpATc0HHsgekVKmW1CF8Aa0HGLlTLPlKfsoFWm2TkMhgfs2A1JbR8t5z58Di8D
iJPLGwhlPRfoGB8y0iC4oI3DlJaMc12tss+0RuDE6qrrQKfVJ0xsonBTdfCkVHn5aLxwt1MRwQk0
bpYHz5BemGo21emzgGxKz5ESxeFqxKrKhOBdYa48Mh9h9yNnOP/N+diNCKrExEV/LA2o6OnJTQtl
OeJc35Pbptsd3wqQpioXm40U5HaaG26grEaHQZccvg+ZJ+f/zUmB7rXsG0fvUMk5VwemPjeASRtb
GTisApm7wNvmtV0dtP5n00UqrkjIAq/zRVJriblTIwhTNyMVWegfhgEIfSbW41pTrHFY5yaBxrp9
G3a1Yr8Mf56w/NwfgoL2yM9twqVnkB49uBzzhCyuKeMwCJK17NBzz4+O99ukfu0wYOKIFsTu75EL
hg+ui852rxL673iaycpy0O3ueBu3HcqEVpIl0PcVwnnDnzNM90eqhFs7IXFLSDKXuASxwCa65Fti
LEiLgabDtUenWV0lS0Lnihh1So4gnsLJj8xpoXX55QZeU9lMr0ngGV24I7v34dqyp5BTnHqjrLq8
qW5Cq7uCrc5nO9/js/Wzb7yPOEjhnCpSu3bOhiKtf55yYmzJpslFjSwebJJgd7MI3fdGOfCBD0BB
+QftYq1mBOehqewZk/Ny0BdUvss//omNE6AYHLqNI41RwFVGQQZfFWJiU789C+iol2QsWV4ZDYcp
bJ+7k3/QzcdYSze2kAII6+6kZYONcYcZbtjRWWOe8CSvPPWJooe7ixBJhAZVtVwzT4+ZS9mHHTBt
dusUButhwqnTWPVftcwcJtWKVMPt3CVae6J1RhOQcnWQs+popLaGKfqwR84WcLRtzC/rNGusH1wz
McyK0F/SUCWEjo72TpDkHxcpXcnllm7RUJAYGh7pOmEnX/2KHamdzxDpTzeRObQ4udfkoS4Qet2w
lZN6XLAIaS8klu1RmRKdnPeMpGlO6T0u06y1N25zaSI60gO7VgcVYy8QtmnvKuRy+YZ1p2mS3Bux
zmb11AVcGb+boZ8BN0wM5pgve15fLxaT2x8U6p+WyhQajt/XSAJmmkE+yvwQjISlv7vigUTkxw0d
MfprVZBHMSNyEnYKvkcBn/mR4ZP+Ynk65gcY2rkn5Ypig6tzcFJdfKbwsiHhc5UMJajgCBYLMfY2
qvOoF/MJFWPMyd23AkLl0IyhDQvkkOhjA4FnKmuqnF4I5LuuN4MUVZLf1sdpIDRSaDgJEC+1/CiC
kVrFByyXzRAZX+yadg32Hr4OhSmVkHnDRDWtIN0kfV2sW6LfSF03h+2OG+aIuO4hb5QKm48mgLUl
0MgUHYWW9dNX71Mx1gDYtCLPZcy0YxYhcxKMV8LBuTJK5cCLtNj+RkDvFctw+C1GoCfAbyA1hl/9
Bvu7nIw7eK9T8Y4/03XjKDVkWYm26cKp/nPwZ27vrM1bxQ2bEGRrZTciT3ja41SJYsU5hxUFWWWE
lahoXnjpbIha+I+UpB3mqVMI7fL5T9FeNVRh3EdnFX+JtwjC3h3q5/ihtvW6rkcKpTD2xCCYe3Rx
K2kPLZBkHoa2OFyEn96szfg5Ib5SKF2C0Mum2niDgD5GJLDFOigr9H7OtvcIZPGTLFGD1s84xn7d
DMBCddlvXtrIfIChsprhRQy8OAnEWkf9BDbvshoAfkHBzXcAgq3LuWC4WkG8F/6233DkyvFOAeuQ
SyRI18Ha99rsWPv4mS4xTMBX0NGCjZSOQN4iro2zmjC1UG43rldp7c8KuQ50lv977h+3V7AUIaZ5
x4so6LgMLypk/ZgBEgfUOmaExvy14mtZxNrjJdU/zrCIGfHLz6yigt83OcTbGL1CmAhBTQjYELRF
NMbEztfpFuoyI7ZC+9/I232Jt0Y5/JfcRXGLnp7NElsmTzujPZx0AfEOVUhwFXhSHy3Vs26Fxxla
YY4+FSnfYMDGxP0dwAAOQNEPz5/H6IVMAo34NfkroAw3PtwWwNJ4AhE2izlseHhrtSQixcW598Y1
4I0VcDXgVJdtc6IWGe5ic9FGH0FQmK40gT4Nj5dT4vMn02paz/ud132NWez5PLVxkuoAIPiaI2sr
urIEfmbeQBffR/j0WZ8NuHhP7A3bF4KmzCkp4RE4ckqc23v6L4dBIFEDcCUty1qmBF/iNwNL6Rx8
Pk4DaHejBLPnlZRpCKjiXMOa5CGSWxmH2l0k7VivcCcZFhI7+HYQ4IgV5XGbFtPxpg9mbXpOO6w/
wp3Zw51LIgPVGDagOYpmjB0nf+aGUraTKNBe5uUonM/Cn+uoKgL8xTkoVxRIO6fALSS0WuY/G7B0
uJat3rJ3gV3Ques6UllcfLtlvgJKVGFl0zP/iTCNYXf3zPfEsY8smnX0Yfs8/hnR2Vx+s/YkpBbW
uymP8YQQPFwz2TLUBy8cVgXDQAEVRv+wn8uYZ9Zn+i82+Jobsq4Et4sRdw6+jzOxYNs7TxRP5IK+
X00bdCHv8NC1kNukPp/DRSiOQbgHtv4MA6uuBBSMS1m1rWASQZp6c3XDkY4M+HgpwdfViWIl2vSF
YCllIRyU9gI6CpFkIbNPTH3SWjeKSQVHqEqAjawyVa09cnWi0i/SvmbKUkHHtzpt3eAxd4K1xAPN
xgTvcj0ahIhHBaFEP5HVlsxe7K4x/+hktriTdLqmE09UXKq7XNu+DlvqCMhXDWIBULLffONC/ex6
UNfbDhIXoClezWykR18qje7i/SUjJEYDFITYJSlc1ZlEG7XEJoftF8ufTDGJWHjif8wMi0w4Zkbc
8KA6/hpEGkfJlZYIeimHzhqCAFYydGVs4pBTTfdsfC4vesUZ/XsXBAoYnA0yue8wjhUEn7NYnNdh
ahzvpYtH2JOplta+0XMBOIE7XxNlC5K9B2pvrj6UIDR1tizvi7mfgWFQzxuBXWDmI6sS485jDO28
b4dWsktHMycNZh5Iwe5uJqsIk+HrXJLZE/wV7/LwBghFgaNttlGY51WFtnsNzXQGKSmnOUHM4mrA
fMBHUCD3koiyd4i+Ak4PGJ5y0RT1jH8h0c6myOCQ76ptoTZUlSLRkfbXQFwo4zlFCCMG2XKlcy2L
AQO/Nw25UhYIpeRfZRZ1+YBOyJt12WmZLIXvHy6sZZxzOtbsX/nX6Otk1exv+G/0jd4FmUhfe6Bo
CCz+vIRGKOhe8qjfUNgyNahCgFt8CXw668biUiSPWBbwbEDFfYib4lMr9mkuVr0w5eXv+v3yArSG
xprECjNbE8lYq3mjWNBJQKeP1SZv3HnCK3UQIlgyU7zejqxKhMNEq+GNG8V5aLvx3yo6RIOFYdnP
cfK+4xWgj1r3B+1R7QtrAfOfbmfZmRZBwrSNe/H+6NHdCFcP8shxxBBzg01atImvFVn5GCjbpXYr
IwUlqXQ9qgtGghgDMkIaEefc7Tae7gb5yyVd1y72BunA/AhlhHs4xP4Gb62sOVAPoTCHZo3zRzpS
RoHc4fmq9nkUnYQL8w5jBsnI1mBM5Up5PNgbUkZdqbiIUHuNwEeR7B78GO/Ot0kfu9XO6XMCnka1
jJ934lByoProijhiSc5MG2pXTU68N9BHhVos67gxaRqq0ZeBApSkSnNozqCB6vGLZhCloxeRMjKO
99SJwHdlblb9lgzZxUU8PEQ4bb2vxHwZZ67rT7LzB8jwfhN4ZhSmcYhLwXVni0Tmy/gijFjU+mjf
F4FdL/eoy1dA7pApmupRD+HdZ8k7a8Cn+in7c/J8mXw4mdqicMbXR0of40+mP0fuLDEzb+xCorlC
Y3QVtmeuzVuZLcKpwWTZgVWPeQUZqY15qrSiykGLrqsAKxWQtW459Bh/VGRTK3EINyHarA7ZcL7c
114GHq79lEyvVNZU/D1gkA2dAVDQJt9rRwDLm7+HRgWRpel7fk2MzYCLETHeWtHEHmib31Yal0VH
rDp1zd0fDnp35xPg2WGktOnzJ6OuuEKQEIZgSsdsrFcpHT1k7ia8EhquhVRzeKV9No8Y0cuqZRF7
5TCi4vo8HWa5jRxpwV4wj471orgxMzC3jU6D3odfRrWp9JAKEl5Wsr0J/eFmUotqh9fMWuMJEX7K
eY+9M4azgluLZTc5uSEy4cnQ8ARARCZon48F9uOkVbXy4XHrhNy8aQwW5YCjE6dozvWL8vF0ovdT
aLw9m2ajBqg6XRvT8p8wGNQGC7mLqUfrPT0BuHt1iFtB66pNeCLhsjSxloLdryfhOPdY6l554FR1
Goaa7em7EKoCdDFpHHNRf7NmZ/POFNp4s3A8NPTGzkuFe1GwmSIg5yWnY+CSsbaDNh6lZf31XS8+
QJypO/rgitQSlsaprtlK0r6GkeW+BdfBHCnyxhyEzBBynzTpIWvin2epjiEaamh95AT/saLbxQ5G
f3TMOZuCtfGtYaSOnQZU7FQ5vtUbIJ85Jd3NW4QUw84QLFwE6YHXhoyQwTtp2ii7L35/KStmSadl
i1H1Kmbd+uULXg7QIxb/XX0gVMW5wdGMbevuDZje0yfZaWQDqMMjFGSL31l2UjgAz5kLSDSsOU6P
4lAe0AGtmO0mW5gjoGwT5l8RvwQ/4QvRUAh8FN3W74JUKWv3v5rfANr9lsuBq6V0xZT7A8QjWxQN
D5p7Ce5ETwbLwChUjgvOj3Uy3yC45bRWyTz0MubmegLPkafPZ+mgM91Dm4pGThp/2CRazlELsPuH
qXdzJ/54b5J7vI4DzvPoZYOJ6GbUjfXqWDN3ZlFSwAYypzvMzFQRL7aoKulKcyTGE45t8K5Cch3N
tiYQWWz64ZF0PGuXgRbw90MX8PvGxfJ3Fobp3oWI/YIQipapDoQdCTLFHQD4Zodhkepjq3PyyN17
HHuiQ0lrF8tAuoJ/yFY085tMXN4e8Wjwcw5XVPCBrF18yiudJaXoUsEc6JzuvdH+XD1CDFQW7FPl
5cFD7r0//vw8H4L44u5yoHfUcenNiOw8lWWgfdtXLiKgTBKR+WhJ2ePIMJuFB+xMGLGWAh6WhhA6
MPuPYr1l4F7e3D9OKbruQX5nd1rXXCka4D4p+TTFMe4yG7rZPAqarQomEsux+SHnPDmHHSkoJCAp
4Hi6ejh0MaFYlLAzyzNsteJTdaiMgf0O5cztsDlPiP46Ft4Wf4KYWeacMtrE3FoluoY61EFRcpyO
NAA3a8Q7VAPVPB+yg/ibhMcT77U392lVF+6/mHI4S9r6SEnTXWCE9CUz++ma2bpeiE2i+GKH0mP3
X2dZnX9ykP0HB9xP6zkNH2AeL3YZHCPHAGIDMDTVy1itaZ1Oko/jtkwQFW8I28+EF6iscCD7pW9x
ZdR1FmjOxFyPTJDwgAiTM4ZkvFy1V8qTx0vha6N1FxHZEKQGYBqYGaQqh+7b7TRIfBh3Q+aavhhH
u/rUc3lCuIXysAZH6cXYqtXgWTGvyFf6ShaWag1Sib81zFuCNVZxI5pGrzrFqhzOnSHbYa3l0h8x
hXw5CuQWy686hQUyPuNgL/Q1C5IqCpW1DgnGKnZN4UlxVQHFRP0vfyocm6OZmD43bRWQ+L6GTQEl
7Y+CfegO4KeFK1QB81H6jL/JR/0x6DwOPFvjmt/BJft4mHqOhnXi0ZapyKcLibAYfZ8QL3x2s3jH
3S8lL5TOsrW1P9eq5m0QoXxFGRgxXpEIaa4GPInTXoiKnUWawSGwRIlUkkr9DwlGWIuyPb3ihq+y
xwcnfC7HQBHxFT6yfrBHxlbDi5lVJjT3gl5HiJKogHfm+wKww2GOkwVBSBmWDEx0rvs3Ao/W+4Gd
6X0SzdYqF/tNJO+rM2w7Rd7fd1KkFTZ3WbnjaYV9uoMMPgzyanpAIOR+zFwX5YELZEkFzCU0ewfc
Xp7CxoG550dgMSnyJOLTzWckAcr3rcUiTU/biW9Y9G7TECCEQssuG7M0Rhw4a8RkpdvOe+QyWh/j
pKYvMQfoVnj4m7OfO/57tf/vGtNALGFRJGxXrr+hIQTpLHtZdUH8LI6PtkOeAUnKKFlAfQPY06Fn
1PsQw+x79p3bHhR2W9WljGWN2DesnJjfglTkETpcQ78N9Sr/vdSyfq5Td0BmGT5XGKH8G2nL3R9z
jwpYgG5w3jNblUwKTly4EJH2U6t7SMeuUsIycIkJlbXsbDG1cTKHdYBbA+N92Yj51RFkU9thizH0
P+5LEgLAa/K+G6VH514xnVcidnr51axTAh39U7VjeF6TRt9k7lb4sEII/a7zpcTGZIoeaU8IktET
AIrYqePA6DtAn57pLmduigmlHDASIVfZ+yymbzPFegEds2qCCUY3PRI9HUwHOuTkK6/w/XrUSR3o
BCQNsxyAo4R6kGcInCm6oPe2+ad85yWWzRFoeo39VEsdWkzDjsvE34mJkHrTG8JVa7NBvLF4OxG1
5ODBx6rQrgMYd1X+wAf4RDfiZaSxpG6tDFsjeEKRsqLiMBf8l/IockH03aXDms+zOdQ+mqjJsT28
EZ4SSyRiu1Dhk+nHxGKAo0TRIKUCP470Nh77UEGGJTYYYVvQl0A3Njck3bvYtlGWdZbcMxG9810G
d7FhjszN8WU8NrWdt+cBnQASn0wZsg0DtwnoLJ5F9740/0ij635I2KNTUXocQugkUdhne8yuTBcd
G/Mae/swQlavpqDTR2jLiCJ7mG1n2R0QD25Xp3ObGpgYWetkTml49nhi+kt7k9CBOerNofqUqjLb
wt6DnauxlQvR/1OXgSWHZD+dlth91g5c2QbHmXjMwJtbAL3nMl7TgzDCHFBfVxdfuTh5vBb794K7
GK3vavgy2As4oIRN2RHh5t5xew2aW3RdOShzGbK+MjJJBglZU3B2fMnUFZBOX0N7VMAb6MqkjGqK
GGq38oAf71K0u628h7U3nppePYa+ZTKwfifl1tkfgZQGZElhgaHGxfpd9imX5GmBwJSb32B0j0dm
p+ajR5iutGOyxtL1kMuTLYIqXsR76BlyYvLEp7814xA3hbAZEJGnYmRfOj0rVrgrpabV067cEt2b
f3PXsAWIfvMKKwr67J8rxsF5R2zQhVgLUV9eyXh0qtjx/+jKujP33tte03ijIEAWWwF2fbKWO7BB
iblxY6JNMg+BQuWXYTM8ow8HSQihgNT0N+VYWENDivKIOXlSZEnuQIFi8dxTx6l16xTwQXR0tknW
xmb8ypxjh5p3OofcV+uRGXhceKFua1Ara0MbC4sHFPWqZExFqT1Ld4n2aHNKyjN/6UqmlScj9aGD
2kSp/NlAxVXVefK79rj9u69QB4cgJlJNwai/bf5bZRay5LrvzCZsMNbuuJ2hoVbTEkTe8Zc8CF1p
FkNyyHbwqwr4ZOsUg50pjHYurLU7dx1t6bxetBeSvLk+SFTnO3E6+tpxtCBZn/FjWdao9RDkGXmv
FV2V9GbkZsIjO9IOoANP3GH0K5lQ7RgsGxrJxtf48NzUPUCZdiVO5dFynInuoorpu9ABw+EBHgky
TWdx72D4qHD46Gp+EAbAk7VVGRB1cAKUvwFOci1D/vh60N2h/0tPdxXSP1/zJBro1h5GK87+HyaF
1MvSAKG98fb4fZWdszT9TV1/++V888VshGiV1d9NLl9mJ1vQuwT8Ml6TMN7zIYPFyNmQqe998of6
WT2uYWBsD0Yt9lQ4IwUXP2KcxIIF3IGnq9KIl3PxQVqiJe5eCsA/Y7WuH9JN4W42NcokGo5xNBzI
KHf7BZ3xooafHlwNAvaFaXlLpvo4tyyrSj8x6QPQo5Ra9mywmXpiptWAndnlxxVkA/XpmigfLjeD
pI1u3g/Aw0ar1/GwwgWuVwIkuxvs1zuBbrZTb0E909Qe2w+JMPPFIYb5peQ24rMBZ2SGo77SDfUF
O2MU5VbbJ4EJSmMAoL7bMfG1zh26cqZ1mapncQfefT6v0eLKXkVUypwcBIsCGSboAkydDFajMwko
pv01qESJb2IUwdHnQ04uJy2P2TkIttmI8u6xlsleQqAGbhryXthx+Ra84OoPSMdi3NABksidOmsU
m0NuHheUkTzSySYxROks7VqM9BWguKq9ci+S20wm4N/zeq5NZiuUZ6HwNL6r5ObSw+NQzmmEJPg2
KrCaIekal2qMrf7KJkgRjJSkwFP56ABfwV9yBlh08EXiwJdVsBuX4ShTM/IMNvqB1Wadm+PmLOKp
JQaC/Uw5kI+F3JCgkJb1nbsJbLN7Vhk/SW7ROeGcEyS3iAtx6sTPKFMM7u3kW7BLLXPltgLEswOx
+wZhEGDUv5L7sdooqvdaOx+0wz4rvY7g5qUICPLkvMwZmPrBiITP/pq+Mxq96EeEJekdC/aHVoe5
fYl02Pdp5TpzWQTWEI6DJ7Z52J9DaavPdp42SyRLuxNzvGj0Ut3OSJn0F2/ctBlc74UFrXVSIt78
EZbvxrZUhQ1rx7wWlUi84HSxPbughe9Dd/Ax8FPF2AyrwRYmdfvev5XjDRY4Qxd84moBbAwA09Cm
pPQzVjWM9ffqwfs9iipCiN7QvFi0gFvN82Ak9DTrc5945Rc0gMlBUyp2USd6FbVTJxkkorgnJctg
3ADnw/jiFWiZqDch/gj5zFluOvuzVJFNDo37ZGVnKClToE7TvT4V1HbSLDksRiZddatISRS9rvOm
PJ267vUpKFfCUd487etZp0ByInOwzVhwPFFhr/XWXGilVVjFr/IeCf6eHJF7NwCI5wlubYeJDHh+
c/c86/OYaWmEvCtUxtZDl/AvlaEYRb+1iLdCui/f1Zs2XYOprKCeFd0zz+GY2l69Qg0SiI3cCmMH
eQ4LnXsNtg3kYxi+V3+QmeqEfVgls8SaOiVAxqkkepivOAhbLJhQL62les1lU1H6SCnZsWa4Dwz3
jd2g4oZcOaMYOUwMt9anY5WtLM3tlR6pU3BMpkb9SRsZ3tkRaXV4JskwF5rS3saSWf8IYokct0WJ
lCzQMJSo8om2Jl2dT5idnzDrdz5JPl3eR7nTGgJebAb9oNsbPeckyGZvXakjb6l7fRP5wzTgRVvp
rrVBoweR+YdgowuGZcZljuU/zchnjy+gSIABq9pGWUcT7GSVaKVm0SNB9IVqSnKUcOoDygmyItWg
kKGfDb6c1sPM0rLRFEwf9Zq+QFaYXUAnTRws/8K96iQtJNX+qDy/41zfoL4HWAAigsUg42rHopnt
R8T7BNciZjDwOlEG9gTQTj9Kut4hiKA/4TntZcSFmIqhbW5m0/zTpLoI2lpPE8fjbaYrFUlGPBfb
9SqLHXbSVTMdaTMzO2JWBE9/kt4PMvsideuLlqy/1Xsh9HYrNUVIzIKPXJSNEcLNwB5AVGIkI0i4
7de995QRVIFhCft7fpY/ICaVdQ8Lj2RKIbPROrU8LYcLQjUSBNPu+0y/REyde/1q0DUnIzPeCUL4
juUjaclr22ZJ/DoTx44VjEdUKTeh97H4a4EYRgDGfq7hHYk96nQ66Zg/yuEpVyVMAd0JzSawuVMd
0TC4Ud+BKBF0qcVk9d2PNbD9cJkst2Ex+SYNCJKS/wQIMi/YpHZUIsUdc0yyzBkuhLRiuF11pCw+
gUdhtzI3atSvyNGaBUMXZ8mMKpFnAxt1PGyqGtJiZJ1sQLGmYOBasIT/P3bBQs1MEMUpcFfk/Uh3
lk+a2mxi1ABwMkZAd+y3nESoHcl5ohG2cOf4UHq0ocwlUzxdhreNsiz/O42zBMA1BuuP/7PIYVgU
8VHKkHuF/CwiI9i+trEezNniAYnaGYuoqHPCyyFbtluas5U7hZ32iqbvkSqwDMSzlWkM36iqjYNh
JfWZGLC5OmC178pQqVIRoqOd2KKuICfd9dANWb8yHEyQH1YO2SrFVE4PUouf+XN0in04DyjKuU+A
SEqCjMi6gy70tYz3QmxvhwaJF91i/ytLE2CE43V9kdREfp4oSaDNiNHVArUta3H9pJIoVkEXDbOj
wYz36B+tW6WQBlYw4JVDqkZ/dcz9s3Q4SFIqTYfJ2Pd+1M+77H/9lpXABVpGwlSsig+FuMouaQtc
rNXhXQHJTJPZQDdnbeAIx+t8oCreb/E8/wbaMeEljIbDguwjRoJigBih7aCi8lZJO2nUhIHUoc03
1E0YGitEJ5OwBZLfhdgq3J20DIIljKGO5TOmQt9sDpBcTNZsWt/NOKfTgMo/M/6TwHyNXstrIL7L
wxndU5ha1G7GtX+7AEgCzIeiJmgViOq7EJMeRRj27flmiG7C3SN+iXFAiNMDAQgwmvRYaAVNhuUN
daGp1hbQezA4HGyQp8D1IkS35PCB1DU39bKYvrT+O/w49MbxlgyXTDJQ8eICAjps5Ysd3wA6T5AQ
gjCxu91dxGz3ObSu4TWP4TD5ETAw910bVrtyPsdQfMjeTlf1RDPQ3fsdiZfo/MK4+nXqioPUiX9T
N3Pi9qzDDX1pYnjKzaNp50UDa+MDrpHBigZHcj1A1GaWlsJryb9OlVFJMB+eP/nsOg6QKHbb5tIt
2apMp0fzFKZgVPm/TjsN3YBtd83LSRrpS8xC/ggFKIj+NDTdqtK7+b2V5IPb3d1ad3g0qc3FpRIX
QWJKodG/q2mcA/q2/F1GqavxLTeL43eXwBhm3umgoX2V8+z8+Dn8nde1RbbrEbHwv425YCEOhyRp
oklIg1SCrIF4ZQQejQS/Zay+/QBIJeizFBZoeLbAkRHrnPIcnxaWo0Itnm7r8Dj+cQ1zSCziRE4j
cg1hedzexxXVIC7a35YhoijMM6BHD+STP+9CKdWsy4LeqcbFOUFU3wqkHpmMM/vRrzzWvKvq7j4R
mqA5XQp0AQOM+40SncaLxRynYExumAKhCxRP3mxp0MJfuigBr+hu+4AiJjY0Syl+L50QtmfVC/Yt
vholnxMcikGVc+/TO0PaQUlAnebpeI4KT14pZiQkAUP0CBo+OBe00xiUCtpbXx7ARRuv25lfoKFO
kcBHP4wKf71KDUx9jSs9NfZYT4rFqsjWfH9zFJujA0u/RxOgeQe1jeeIbrIlYAYUjKy6NDfXVK0C
4GRhPaSs6+QGml+mQqS8Ietvrs0iDGofzAXCyuqzLNpGwmDHCbr1OAbko3SjoOpiUaYGLCGKgRfM
cQZXJmM41RnwB+MgDLqlFVTZHaLBC6SrJ8NbssXHWlr9VIi6KgTxh/rCGrMk7VntKFbT/cG/sbFJ
qfXhWmFC57MJ0GYw4jyTKYeMBjE54XD2G4+iuVFd46N0cKcnlldKvkGt/HIZ0x2jjw7bR19hlNRu
P3FaKv0+cCwDE2JRrGfHysaD9UTJUSq+uF/dT/fmCymCqKvic+i3o61xVzF0MegmSg/oGjBe3hU/
tVzGaR0z5aOCzmWlw+sZUh7qgtt6/i+ZxPhoFkPHFqk8JLPJdt0RcVeaOUxHiR23KwyEMDGmnCHU
rUwYSYNLbUbO75zjjrnzRxEByu9XIJTGIijStNh8Q06nhwzkTsTJgFP8rYzJ3wfdg8U3T+WCMMWF
0PKHrpJNDEKpd7mQ8LKryauSfZMVnDepmMCAQQAEpxneZ4rvybhRCUzapP10I+U3zNU9sigrNmHW
uI6usdPlhZFvh7jiXJDr3JX4Iqfxmm4kE6xrvp4skPfdhHbntcroyVA4ine/eMhPYe0Jg+0a19uD
OHzh/Ek5aMoMjHQmwCNvBwn+8A1+8jpPGdLRENEgwbTJfY6e5HzLdBAQVApDb6urYm9lh6S7KQET
FwNuBCxZRWxbj7xAciGBe1pFCfOS++ZUnCc4U1TF2pNtd6yOnqizk5QlFzg5SYv2L7fJi8QJ0N4Q
DmJ5KnzxEPu7OU4kCoKwssGr1YZgi+a5oaCEj/lXZqaY4EwBRr5kJ8Ws+NpPptjCNHiXMWJYkjEZ
e0NNykQRlC/TCs5CU+V7xg/sjGfCgNJSL4opYWb+Mk2owLWclUl960tpqbOGQqXg26ygTsq+fjf4
T2mYgwLeZTjb0p4FvKO9kn8Uj33M9tx5woFBHgi24YaYHWz3gKS0zR7vZk4Fj44WQbOIoAzmws8y
g3njQ1LzP1PQhD1Qm/MyWn++b3TV8KQ1yULKyNZ+c7ZYn2wVDLG0UcrrPJPpX6pvuEGTRm1mAYDi
qazneqg02wl8GrrF3iWV7OLyO2pfNNaYBnhS/svnrVuibsb5PVLt/31GPI+A3w+OJ3jPLlNcr85m
b8RQX2BAxRADaBsz60gN/XLPmGk1H6Htkx87QuG8JwlkUz235V00bjFWYImmuYtLAW8V8UTEWrL3
MczL7XD7rwo58GQkHOEJJ1YkYyOFaBu0ev0ezoMo6yw8YveOIQ5mWOxsoKAvYtWVKrDoCHnDjQsm
qkgMBM2Rq2WAJ8ulx0fIPYkily53rTZIjqLGHlo+KRgN3M8bGkjR6usLOcMOzU98KUc9npETHjIa
h2fsoyjt6Rvys4BBaJYPRGHTVYRljRfR5M9QdmhVujVOK4ai1gIx4UYwIlL7hto16LZZlAWzIxCZ
QFZmJurNaIuE6KuZNWebmAc1qYeJ3LgCRwAcEb5/FGTt6E0Yq8syWCQcbEYjUqm4sz/00O6OfCiR
Zc61XIndr02rPxQ7ZX8YlACgzWPXz5kHyTlUKOfPOoOrO4hXGqWk1L2mqHWiOC/JxCtyLXrrw9PR
ipUtjNDOtQN2pWsJUdvwc1EbKIx2i5eHq0DIMqdwRSIHKrF7m2eqJfg+qm9H34eHilYWWJdoyLNI
EvyaNyFC1QuDVjG7ninRk6CniFS4Y7ju/uMgm/u9dfYOzd3QKnU/LyUDrWaRKoUgfDetZ6w+6BI1
N87/BWjunIT/fHKkUqufZPx+ZCU/LU0p751XJ6walEbQHYyAUk9YSPIBx/UOi1cubGUXsaBcS6y0
4Tk9MOy9+z/urcTcn+OUJmNP9fB9LbTgIJHPJTObrl5QYt4/Lh28pooZlUl7hfa1c2R0eeNyC91o
m3/MEjmf1SjXVNudppaySKA9ots6ZLMoz6JHPutNTGjEasIVsbT6DHDdeUY/RCbwoGBmEDsaWHh4
gdu8196m3GEp92TZng66+19mTLgLhdp/nqD3cxkHWA7C9kBcsAFtRaxKmn2gvN1Bfj/jh1U++Jkt
+Z0O2PSXGz4mS8fTK1TTz+TJbyPbuPRK9YOasfvaren/1Qy30zcAdnRJqFXlzmjKMOyhf0DjseFr
JHTMFugbwISoaCcwtTrA60/lYiX9VxJ5GB+8pdtbIF61af4DpNDVG6q5x2uWG4NM379etKe7+c+Z
FOXeTqq1R3f68Tve11xcNAo+EeOv4kRRfS0WLRfGU9S3+Ovf7kX5ol0b+HxCuB3ZH1d/qdcmXxFe
rXScMJuiqby/Sy+3laVj3w5B4S1yeYO6lDK9YPOB6yeCml1PVr5GHn5ZuoqhrXUJXJgQQykPrE5q
EzWI8SgbsoBgEvsNzGtWdnQhKDEWM1Qnb9t9p6w1ocWH6UZkX+I5a5Bq4XZtmZ2U8PgEhZLiT2lp
3DQ+fZdRONgSG0kxC0UOukt8ezt8lGN7wGBFxmAZrlDTMDxr6WEIXMUyRWC9h4025VWJE9BzX+tQ
Fuk+0IhHxDrd1mLVyoDo/X+qU03+a3W3aVDKU/bCYdw8gBC8zHRM+E98qwFJCSZ8/pG0qkRVvC/k
YxE4QlgUJk+mz32OaCKpto34SF/f0xTu7HrpPn2NUCIwmRDz8PoyHZfYvQU+Zv01fqzJAfTpwfPZ
6PSG7hooFyrEZ4Bvh3og28NSuoVNj5b9+Sc79jR8ufjoWk/i8W27Z01a06UAB7WAiDmPe73QQguz
QmKub+aw450d0HFI9Y72HwDPjOEpv+w/p4z/m6tql4zXEkeHOtg1vGFc1D/4AGdNnuOVbZpOO1bH
jd7CDcillyUPIv33lzCR+OkelTGcJP1BtWMGfMt8PZv9TYhcZYlZhUzjA0FnTBrWp8Kav5EXVeCh
i/N0wOWb/gIWg3tVkmRuhWTYj+SVpWc7usIDJ5xUyg6WxNfRCFXcQCObCeMPV5YBqspW2xioNggy
wFyhcuEceaPFEjWMxN9pI91YzUXWnd7f5K5hzT+EKcNaCerAfBqYv9ftToi3wRGRPAVBbkAd2otx
omibkWwdcQYsqdAQHfw7NHXqWUN5UwklWHQ1akkHZJTWseMcZ3MGkKVDfxixbJF62wrI/GA1NUh4
YzByPfLATHCehYWpGET8ATuIM1VTfe2KaK9wuf+EVrDMQl1N3pamoDyipHwH1bYlyVxZ+cHv3phV
sZLl1IYHnjT97WrfDgOypnuuAfsx6c9qERaUueZ4hrbHtb0C3HkAkvHlxImzaqFXkRUjdFvqRyZ0
1pAcSsetxSAH+jkd7RLFjeHJ56NzqBEwmrPfXyD9rjFWxpQ8J+Sw3W8kY6kYe0CvIeiKs5tzoJTt
S1OXs1vZDZcx8QnThLa/O6FkWGnZyRPTLyzK2KBB4r0JZzCib4Kb0djO5edvyxiF9cEE9q7M+idx
x+TdWZVYQI2mDixp2vfprL6N6EzgCX0/9JNZ1+IMU+8ZNQ5J2RkhkB6t2BF8pszCd8Mc0u1y2jFv
TuMvo8Y9EeSo564ORn7vvmjc5UmsuzN5WRgtpaXnpvb9LXduEQXpChLpDQ5/2VOrXMQvzfqVDiUl
eZomjB+0QHLips5zf7e2b+OvqcKumM/tgOHExB6Yea3xGOifWNyJbgAtKVDfjt9K5xLqlh/kXt9q
QCU7DLGhxzjLJHAi20LNEUbyIW25VtyoN1xdHVvFrkxT3F2Gl+GtxQO6cTf5B5Ymwce38gZ2o6xc
a3n9a0K6aCTsAzFYbGAYo8Qp/KlC8UHsk4esTMeKGUnUlx5A36ceDKIiyDh2gKRNexnNEieto3ao
bpVW1o0o3ploeAwTMExPqF4f6MIFwVy8HAF0F39QFDq0Z2AkCSKfSviK+M5KzR6xtEl0Yj67c2c/
8C5tv+dx/+qDomjOXiA9HAhDUcOaaBEUoZQZkHacajgU9qNPFi2NIhCliu2TMPbJYR/3yooxC5O2
8Ww2hgse8YaXrrnvZzS9OMTGfsJIyg262dizeMfC8OYBrkTHSvXk0fg9MnBLC2GkNQmwRfaJEO7u
LYJJ9mAoqQe55G11WndtACTi2jPilelXruLtAXDEk3fk2QsBEKlFB9iNPi4WLoq3gGyUD9algKss
uiQlD0a+ej0AeswFifK02OcVZJ9FHi7NxpbcOgROo9TzR7ocQ6D3lAaxKXXlpqK0DTWrlBhy6aV1
9TqxZ2fOJEPtKO8Ewb1eapF1c6xJuU1CFwV/4ZiOo8usiU0xiesnmLXAqzr3IfI5bTY+2xs35yJG
y9sqmgrXi+e/FXmZleaDLTrLqE+LijgpwS81iQ9tIwRG5f8jL6FRjKeJTOHsJgGrhBBdBElF2QNL
rhshg1DH6m8dGBl53l6aprCrrLVjgQeqjzUtN70xmYuPwXggGdUmTXdPzjhSN3MH6auf485bhEzP
dPanCva9ebD9lxKcuANZVxD3rxEZdScFQ5Mxqd56HxQy2IUdia6b5JtcOCCCcPq71Xoe1mHDlmM4
4rnp7+rKvXOh9cWDLX74lCYsIosWMg1b/iW4WMwzuf8RhalEoiHqMAsFffHpayiCbtsxeNjrbUHG
ZziGjRT/VbBHoPWlu1qNoazAdwI3ASvTy3eZITQYvysq0lgb0aNa/yTkaMRjKuGDPzDBE8nHmyzr
PhC82sKYHnZEHMftXrW1X2Xbyvaca6115DFwLM58LGFlJIK38XBDTgfwoUh6eyBgz5cPRoQXU4BF
oR4vMu2R5iVbBx3M5b3/32Evvv0aIUa7ugt3IH9NgjRnR3DeXb/IMkNvmR4u4nqTBrWWmBV/DsB+
AbcOh9+Sv1msmWvt8c+woypxYty5SqozFfe45UYoz+uUAcRS/sRDtx26pKgKM3wLH1rnq/tV8iIn
gsdSbCS1kkSOO7oN757Tj0rq894q7iyicY3EbS82DtLHkwv42oJkAj9UaQ1j2Q2yWyYA2HslEbn1
ZSevFbyct9KZYzEBEFZTDT79f6lU1tBuh80BAqrVNGmKl1/XWWfDi+grJM5uS6e0+Di7tMFyJO6U
v/oJqTMedS9D062HD1G/2jofEsjZt+k0ZjyWfBpRu2prh50QVqDaM5FO78mW9rN9UnRDcFoiNnrd
sm/1KCOFGLKD8/Iu63fxwU+SYWT0jvlqSMGNVbYPan7Ehe6cdswl62eYOR+UR1IuF1e1gO2EMm4l
uPxlqJH5Sfn7PFzfYR7vEwQ6DH3W+xcJRrq6q3lMPovFY0Dk0cht6K8uzHjfRSSB99eWV++P82Ug
DBJ1jxvsGxAdhtlo5aJjrvOEfRJSkKxozgrG0yBf/2n0heW13RwCSjTnnZLLD9pj9D9GipqHAY9T
wewbw5ZQOqjQgLFb6r8wDmXSImjcGB9Msnl6bIFsHn+j2y3hFenfzihnzzfHoRcTD2/cGLkGnvDO
D8JTGZc0XmW6lc2xesR1XI3poacT4u8GREcb5ayLzWCIdUyYPc/kJSnSNxdi+J+YCaPo4nF1EE1s
XMwUgWHO6SxU2WquDAF0aPfI4XD7ykc7GgwFKClvrnnvbZR2RFxKaTd02eK81nONShRR5Er+JUEr
r1HAwoVZrpEZSs2XHJw9LArnMjC1Q1H+w+dbjtCf/WPr35Yj33YA+fJ2uEFSi8S9Y9JhwhTB2Pm3
k0CK8aTq1W+SGd6HHupCscKOYFbrw4Tye7vh1KtuW7dy6ImsXLyjS2fTXckL/nwDsO7wqxxXAURM
uJFvpvvkYAIOBtkdHPz5Fc3VLw9S2hw02AD4oQme9Uj7vXb+vy6+naMSGeZwiLkN4AJBuk9Z20kB
u66/f0YkwwSm2zV0CyLfy80Wn//bomSw2TgraFmwWBSUtdoy/pICANWovyh2tD2rYXzcUMDDJwKY
JpRypitmlME4cuR4Z+YTKW7+kQIqxTqaVtG+9y1/2xUppfFcpMtP9w0HGu3067Dg4/DFp7WOEUeK
OrKARy19v+vf0kp4QXrcfZyhNjUAlRwMB3wjvbYtLfvfLNlDn+vFvCsgCJRz6Yblc2rRxHV/0G15
hLY8mVvAhuCiOe1NuQlO7D7Fv30zkehdSivOQZM2SFUqmh1tOKP5pbcPKLxIZ35uwuBd0G77uBBo
J0ROo/dTXf8KG0mVZO5zhvHmIDpoppkWx8QLLmDret7IOYi/NVhDPEzx3wmtHdgSydAjYs6W7HEG
DUq+gZGk9ZDvgrAwpIe2o9PF0mHR/8z8pRzBp/AfNyjB38aVmXVgdJRVh7NqnmZ4Y26XEmC4X1D7
3pfhodPS/OT0QajK9nm+LzRN9L4gPsU94HmFdGLk9v6Elj4LCqyeXXxRDT5isNVq/sBpdBY8PGXL
kAbIwv2WTihB1KYNRlRQVruDwMpSobGgWLaQrNk3S0WP8Ai2i/zrxwdUUprtLSzQOuTone7E/tnB
P9wLRmQ3P9n6PNJ+pAqTVnZeokRItx+S3vrcSblCkVv+e333l0GBXPYFrtnVV3v3r00fKxyoV2so
/zj4fcTUSoSN8ZogHyZrn7+bFzoj0HLvctJOrh+WldMj1lECJb95A10gfzCkkEBSIWV3VqnINxfr
ZJuRn7xiHVkqjRMSvTaFaIsIWWizT1vDSSidJ67qtC1RRYclgUB6/DRJMLQBrncZflz+6swK5AMd
Qek3aQkk1Fpe3ZBmUppmikW+pSXZPQmqqfwnQBXssEa1zfIqQB9Nszj1mU0MYTjjA62fvpbJ2UTh
eqsELTpP9vWniOIN2XLmTPo8zVivTzAYFYhf7J1DDejVxJwyEyj81UUOBvjSTmISShqjUzUXhgKX
iDUGC4C23x/EoPZClk4+I9FkaBx6Fp+CxJUdMKJRtiz8JucWhAlF8cwtdwTRj1496TwlMHQxZv3I
fX5xlWYyAkwol8S8lKkmwuaoisric0GHLPh8jgVf1QqQd65OwVAORFasHk+PMi/4aE40tw+k+e6F
5Jkp+T+26IFcv80lxBv/w+DSimCUW0+PKoDuLUKZXfNfI5JxUHDQlFkdGnaDIOeXfBS6mvC+zuex
AOKoyZSjS3qb2FYDrsia5IITePnemYd6OUJpNKJm+1WdcKhgYBdgZLLW8bskdTJmFEnSQo0k3BY5
EfJFGXKhDSDumqasgjqtmV05S4JZEj8DKRMWBi+cST+M+S1X0ny34J1IxuxOK4Bia4P+yLbJCE6y
eOekkZZTK7+jSHx5otYN4B/LU5decjxtcD4mDq42NQ72caS/ND1d5ZNAeyei6JijD228FHGVrwo/
7wXvdzST9R/6LUvSB7iR1CEUZbqBdAw1WelaJSGNRzs9MXNlfwqslS/+Q8MHL1s/zOHA9ocekiza
H5JKSei/MdcjSAEo7N9aNU6nv/eHr9yEo04H6MTClRjiSmLN71YTE34RTCgZLd9UM+1keV7dg3b5
Txk2jYdkbQfcbh99Bh0MBP3jyDe0hWgva+LqyonXCgHwXQI6jaXqoQwMb24iNmZMqUS9CIXV7xro
W7YpBxdsjiTzoVNrTcc3Cykpzp1861KAMtWBG5CsCZP0G0TMeHOUgJFoX//RW/qNUFy6tbHEu7KG
GXIXW/vA3A3+Nej6UIwqSXVWh72eaP4Dk/EvwIBxddTdAsYi2wvQmQkBOTYebqXXlMI6QSq1qO7t
+ouTC3o2IcogtwwCa7rV5soD8wWmi/pJyT6PTFm91+jxnZrDbihh7fPtuVzXpFtlB+emejKOt9np
CJVxV8lpgFJsxWRyqq8jqvhaZDwjw7TF9cjpol+myKul2iYIcImf5FjHRIn7OF6rqBlml3eidt0c
E10ZeSqCRYUWD/XmIEP0K0KbpZb1JrOcCEgxw29+vM8SWIVVKzu29Q47f9Hz1BQT7ajdVco/dqCn
spm3qYrAnjq+0EoQvq/oojLQuvOSOWtFNzL8D2JEh9C4grYB0jBr5UgGxXZ/EX97XTveTtMsvCCj
pn37rOB2y2HgJJ+GFIT409sp4v7jYmY7VwD5vZC93YzNdfAlr6Sttxr1Ks0khQmvjkvgoDWf6gls
YR6bnwZ6U1gO+nKj6MKhZoNgkkYl8fVn6xPGlq5eK2M2e9EhEZdjHIpOZ/dtFQJ0E6hS4GylI7OO
PBVUAR2fqf6sjHc4LY6728qUIOWEwPzfI0UePhwWNhyVQfIkPaRGqLlmHfKey6j03os2jhQbeL99
4zpxwEPIbE2NIit9zDALzL+Jj8S+dTOpMYsy8epK9amyVquUtTUFsox/3DaKdAg3ZCq6QSenH0r5
anCRByNgYsYSUvbxAQuHMXj8ojicLQEJ7JNIBWFhdLnNuHHnFUG7K8E8RnmyktXZI4dZej2bbRO+
5A4vZ46UweSjXVlQaoa68TtVI6AKp67dQ/rnfu8iBTBgrcba26ltEXVvEP7R5tpU3ADLSPmr8KIH
0e3f0GLFn/AXGGet5e8juHbb1YhP+0LAW1HHAT/VQQFbFBgfRNo9sXpd2OAo1x7D0RsFALtJ7SSt
DRRAK7QMFjLrnEJIiwqtVviGx3UKVVgrOK0RH9tzX6DYq93n25NvTk4o5eBnK7sZGrCpIKDN9K4J
4/gjA+QbnGuQ5pqImvDWPBHmw6JBRcglLcS+jCQg4KusSRGae9e289tMfUuRwRUlqV5Ivw0RfNga
c9jr9L0Kp06qrjXeujT2TpmbwFEeEhMBKy9xT+j5y6qWegHsuYGNtLVzFJcqqavFvaEsFqO052Pq
Cxd3KWqfsTJz1DlpDikWVw0DI+qA0HWqvasjCLVIq4L0zCq9GNf4lJlaRMKotQo//l2qbcBSwWYl
Lvz5ZSmEpTzlcpbAdeJMlyyTAgv+6yitXkrnDXfO3Z7li244JuehLdoIWfSLi2qGAVkskOUBnqmK
3DkwltOy7FaWhh7AuHnoHPSuItrWHE2/b5HRkwcVkURfiPL+rwdTpJpPtz+3v+VKJuxfTdYnb5jO
DIyYI+n0PGODd/3KzKclAvpR5FwORiYcTxGUm1sPYR17/zW9hsmzc8aO8cmN0H3SL4pL2w1ehKsV
N9JKBvcoFkWf8QS53Gdl7AOHKXoYTnUB7Zy8YqFn31m5OAbDiiFbkeczrLnMvENxcMtGrFqqfmwD
e0Am/PC63se/fQxDuWTiSWhCpmpvc2XnwqaZQd3GCiNsXLyWCmKFnzUsBzMZXPl+Ld17fjy6Tbr6
RyE31l7VpG9oQeqwJMoyNoqanFrHRogmGyv++ninj4zExkuDIU0u1ENKqgkkI00H3CXo5sqjOGUW
2uHaiMR00IU2b3YD6Rs6kd1sL89apAFyPmUjesrn3rUS6JtUN5tQc2SgNcL5+ApWT5+oIj8y7al0
vDRZ3PGC/3HZYumZ4+CzKSFxwzQdgduYWpIIiRD4hCkoFAOAADybf+wJoUjULcEYi8SebW/N0rYV
sxWszZLM41Y1TVgZauOgDCzgROrbPcPIWRacuHOSQNWxQygHvdrJvUe/aQsKmLFhnkDBHuxxVoAc
6XrYsG5kMLwW2Xo0RIVwu1gQfdH8xkrQcaVoaYni/rTN1MH8uJuQxcoeE3nP5MQcpcSfJzwP9Ibq
AlZIH6UwpKH5IxojB7HfCJmJfJU/Z9Z67PrAbtKpmjcKcb4v0K2npcwlxKT4Nzrx48XNw4bI02DZ
SfdUX66KwrRHm++kaeygpOGjQX7WZYeWRIzon/ixMGdli5HarXwgdaikHkbwPAqDWfp8+QaKnrTf
Cb7sRIHsyucNfHL29lM71qxkta2VReOXjIhfq0mL2wBaWKUUKAEnc8H0vHf9uQTLv7nN+j4jA4XD
Ksv6UDITAk8nLknfFKYXeetZU3JubTEwuryDX5RAlTuAf2dfqRYb82jaRtX2MSy+GWxstjB7W/gx
EYcrKyyETN2la95AJwZJ7W5GC+v/8I7honE5wuEN95E+GBq1dMPYJ+aX0IF7gotK2wa2y792bB+J
G2L2Pw2PE/1CFZq6XGXVNi6u3DmZDVFmkg/bPm3dNP4Lcg4MywkOeezovRdpZtb0A7lPSlcKD6Mt
zkPt4dNCEHIT6+hQ3tgyMkjGIvHWjAo0GExd6LofzcSjeOhXGiiLtn7onY71nJ533Tdt+x9do897
6TVdpBwYOGuDpXeddjCw84YFpp69zLBgRJ5cqiexjKhFRlStOUPOQywn4+od3ZGyfJK7wOFYKttX
NUIp+SgomPlmdz4VxO9WgmskDA9q7DNYVkQZuXhbTV4g8lgGQIRNyzPoJM8u/0A8rtCsjxCfFeRu
goca4OyL4DrV2XFMmtxfOR1aZisEChCsSqw4dL1jNIWkqtJBx90BeMB+Ywrg6I0f+F4x1q+d9CJI
FiNqo3ye2lWe1M1QaGlUvNKTKJlp2xMHO27uZEY0s/0XwOKhvN+MhfsGVND67oG2xRp4MVrabpvz
dILIkCVdWIBFozDbAip8NN4HvizTzYf1pt51dz4DFFHHDSQFe8ON0pahjjuI7tL65Pf6Lbih/b/2
8MpIiK6Y986+ogbjupgXjPigA+0XJilburhIi0rOCx1hwkEUVyKvkuVegOd3ujCYtEjcrYFmenvb
LuganWuWmp355zW/CopsNaIgruyzNd62tuMOUDen1i0hv+n8XrCOfZ1zogGDz2V5oUlfS6sdnIsd
FxRWWKZ1e6Q4LDg9cbxM6SbE9IPEuNwBwRFzQsobuZwaGIHB4QySG0rUuLgO0slDNpZSg3ePKNa6
c4KzPXbDqR/44ZWr3ftyjFOGIILp0qbB6CodlexR+y8dwvbpY2pNxD0sPojQO/Twgx6kc+37jWW8
NgvMp+BUBY6hsD2lESIxCdsuvVVk5XfebwR2fWhnss7z5yJMR26TaCeUPW8ZcrVmb9q0koqRV6G8
m5NewwrgQvdby0E/PnlHvRC4dHOulYfJzp/OG5UdWpr/UQ6q2ylmeTIUjwdzUIE2haW14j8zp/HB
ai+oDkzGWpNxR1cAkZpKxDGUfWFsOwPvDM1hW0ZJU1wa613CCpBn2GP6VxLYvT3Ls134Ae4cnL9g
l3DA7YVv0kFQ1y0h39aWUDiYbHkO6bjMhPXKr/iYIFJgLAI9mKhm/rjAqPljtu8oZy33bfr0tYKt
mZSO42jiq1vOtELaQ8Yr+gs5DzkjYdgL6YVfN51SWujNUvAXbk2lsKza+buqxktH9CAitEtHehfM
I258qTCGycI9Og4lyQd0odCxlQc1WeuzFlUdMKj4RgZLs5gmadQLVYRz7ktZ8rJSKrF7rvq55nj4
DgkZvE/6JlEsLykeukwQQJgYhvx+tox0YyR3PHK9nsuu7zdmV5HygeSnDaVXDec1kPL040v7mxZJ
imw/l0wd2tuFY7EyOLWaLzrSXAOQpUq2Xp8QohgwqrIltxsXloVTRe6cxWtz3mfMutK+cabDvqLy
CzthGXcOA74EU06/T7n9PJe3GnQmq8tiEATnjBLYWuKfboJJQ7GzCZgxhkfrrBhebzvOfvDat1aP
1iT2O282E3KzlYhqJRmUaAI+IGkGgEAsTXMF1A5dNIVbyfp0n1dHZxzRlRcO7bMykksKQmrVNOnm
2R6nT2FD9mPWzXzIfpLJWgjCRMl6aQZo28lh3GB428+oGbTw2ssEWU2me1IYIaGGqyk+nfagslaO
pYdw0JZoeqTNHxDFwBq4EkU/2QlFrBPvTA+00v1LSBdxU8E323CjE6v8O0d508ltGvDGhlqFDOrd
SWnq+X61NFefySgUHaj7p/xx4I7deCKkjhdUPYe808NliqUYG+FnLqlMy51YySsQJ63CUJEAu2A1
FImhwoGvRVB9QbLwdS/zvlHmKbmCzQFprGDadBwAwnO2XTT3/kPfsxwaDqv4eVsbn6zUCvra6R7R
rlZMzzZR77jVOPZVwYUow/lgP8aP6J4rjKREk7vsOKk3GQx3EC6VCKVFax9CITmGnggQGuQofwnX
x1rWM7kS+VEp8az7hrSW3WVdR9Vli5IAxIx9M9zGlcg7Xb8LAbKMutF5pYjU+2nKaXrFExZ3tlJb
ru0B7/EpsNkJQCeHe6M7m6ACfmplNRAusQiiU6vpJPiHaQ9ZzLHelUeAoDb3Rig6ob0SJvZN+6Nh
BDktKpdLjP+FzUw5vUZiUKab9atuTH9VoWo769JLOXRqRXTXXnNoMJQENX+dEFq+Qgev5MHX6q2/
drBCltQETJJY0Ui70Eki224E8z6xFHFgCR+PUWTW+4Omg3yi4TMoH+sb+lX6lD8tNJiakbruwLyx
pVWszLNhLYBZ8ILmEh787husG5TXOLpkmFgwKIBKnEDdBFLUe/BBmPbVk0oQre0D1DvCeRVRJNtb
YgpvdDZkzIW8bX7JHiWwSxPjrY9QHYlouVLgMAYoOcNDuYpT2m0hB/wfQw24Gk1h9CaYRPdO7acH
ApcZQmm5pJLYzUMFCmI5sBFwoEMgnhlVmF/koBgoVy7e20Ch/sT9it7CQwJWxG2JYp+c0CJGQJK+
rV3W3jbnflTawwgcXS9QCW1pP25yd9oG5SuTMo/MLutGcY4vaKOXNg0B9LZoIwZ2ijHntBSdXMYp
DCpVfGTn+RBfH0srdAzgiM4m/l1W9DmLoAIF7sphZfCUrMtnkyP5Ggsqpq4WkJi5b807HmCVNw6W
hsSoADFYFYJy1dkJb4vejWClO2LrYFThm4inx4uzh4Odmesmt/vlIRGgn56wn+7rq4LYkaK4SJll
FjAfYxaqq5G7+AsIDwOHhi0uI+w2utXENI3jRkRvBgWDY7UWfJyNaugyh1VID5GFoA0vQa/tgXxa
36P+u5dkztILqbGoiZc51Tj3ACX3b8zidEmRmbZ6RDVoenvwt+cfi6yJ4wvC1RaYPs9hk62SNVdu
DzU/MhuPcWJKsK6pmgqfeQATYbqX64e3X/HtEWAOGdmKXfthnK6EmMbGDT+7LjgE6ye9IO0Xhwui
9eT0uoMLDEIZ//Z+EWne8gACjatEUG75iM7HIjgcRBMdrXBmS1FyReQAK17U8cNAy0anqXBBsK0O
rY1Ci9KrZqZUyQjCDBQMP6310PPFDBC31UbUhtRLyOruAoQEpxyRDU8wEQETCySsLdWr7ictP3DX
U4+bqFUBjU2U03v1Lvii5WZxfNsLshpq1qCC7bOQyma6o60sVvkZuLjbUBrLdbDWSGO90S71RLXL
0Tp8eP5PkYK2L30LYXuMRk2QBv3EUPU78ZJ7VA4hvJfPq1OEckdmIhxPI2yw1WUfUTxH8rdWfWyM
ZnNqameMOBwAOXhjHQjfXIW/pPrB8Myffw1D6M/mta74zkvB2vmLAPaKkh4W4ZG9mTsY84s4SdAs
M9uzBF+i6pu9Nj+TXmWuIoGWrADzbAlzwYYbqe1zRgjuxqtI6kLJzNdWP/1U0FVFG2dWclNNMgYI
ko/Ywd6VVt5PKAGzvvoGHjgV1tyrXDsUYTsmNMqqleLtopwIB+I8kNzj/R9JtZoxcHX9/1lzzpt3
hMnWEO4zWYoo3Yt/zgRc2QzTOrb1ji+K5/7y0RTRQOpjOdLntqAafIAg6CS5UrkUo/b7W7+2Tlvg
kFPU+P3h7Drah+DzSOHp6Ep01zZ9nUwNPR2BZCHeqVhCGvhvXb2BuHRzL7xcn/gIz0H4Nj52Hjxf
qmJ6AYdEI3rBqZ8fK82IOLM1xpGxLOT4oBvY+/WvCgDSczKfg1K3BFwpQbfqex9YpDhKkhOVPZFw
+GRsooHOqNs0Oe/cHu+/9YWm8deyt5wdoEfAWi3GB29CXt8yUnaX6B03ygET9645FiUxtQJ88dbI
e8FzQF6+B7S6Nj/E5Tv0Apr3/uR6mBDDg/GYWmc11ejrpT9P8Vf2szESEKgr4pE+j5fluoCEYYV/
DKva7Iv5Mmuo4Wh5Ppl8mDCHn7n8436stZfEDAVUkIkYr79+pw25pKaqf+C/6GxQqnOcY9XcsvK9
P8cEeiRYCILW6z4yTb7k421h4M8ZTHY/BBegGBoDGSvEQc21pSXpRqV+rSwaC/GVsDaF68nWYDdh
t29Oe7qf8NoTFO5mKupQ1Ccc2e1OK/VKcXm2Vf7Z267kdYyFr44BZWVCqimOswtDTs5nGc/G0Zcb
Obyv+CWdluHaDzl+t2ETRqqgpkrfJvkNlZcm5RUXT4NDue8ffbEzqzzIKXYev7NnN0I871BDXOLs
1IPCzqySoYYhN+t9M5Yr4uAY210DMJjSC11Gh5H2s9zz2NY1WMFbnZMfISaRctcMyBXUplqSOiiW
kHIsXHN04+t7405mEweE38WX7vPcXeGd3ThnTwidahQfTYuhEEPQFohzk6qT4JnWDs3CBphdGaZT
97JFrUp1zWNi3E8dr8zy6Q3XUQmlp3A58O2QO4u6IpX/zFmIYa1j1S0XdowaOZlQoxiQ152nHVtJ
FrONOqSGNt8AMAkp7t+CdX/QV7kevWjkgCZWYl/tRc406fAGOG48L/mcLCVwbYidUx+NwKU7sx0g
nhhK1LKlsyOMgfiFyN9ME6sNUROT3gJLHZc5+rgdUdgaFB6o/YiEqKB+n8ajsemZkhl8jJ3MA69c
nkbbZdtbISoJTVlbLUumcUo+GO6oS9FFhYqri6bqJOOWy5gisPnCtr1y5OelC37yERm32QeRY4cH
ECPfupXThq6NlS1A5vJG35I+Svl1cZeK0uMozTjgWRzL+Qf/NFLHNKtdIpcR2qzH7kYOAwVmsKFY
mHkA6J71De3I+26wGFCLx5kpwXv7B0Vl5CRezqr/d16c9agQazLNodM6b01uhHE1xh2kO5yyFcnl
mK+Fv+oilYYyMF8UxB8DzcozhwETxyFsF0fNDpxk3Bi+fQF3eAOaiPgR4G6Rh6sXEhu5pARwfh/C
ld0rjY7nwoytVhLypo/wT8zczuyJJcutBs+K/wOf1L5oQSSR8o1ByjmB+FQE3e0T64V0htHSPl7c
bNkiXmAowm8WGu135iQJgsQuqQb1f6thwMZMRBtijIVwLM0AXDBIN/tRSTrPJWKGXAl1wc5r4KdC
bNiHYpR2gT9lPqUsKoIMuRRosP54Ocys1FRWC81YUm24dK7YnHB5KLhAXP3cKj8VMY9KcXAgISjY
9pfqe2Q//lsJLL+o5n02zrKPFrZV4ApmQsvh05C03emrM/peqQ4oq/JMZUFo/u1SX5IREYD2iP90
n64/VU40DD+l8Wm8+tw705h3qNPEjW6gcJmaFF7L0+7WLrUf8gEydCeAWIzh6r34r+atEVGNQtHK
SycOKpdS6z8XhDiEH9ZnaGDv2vDYfQbnXIQdHvqxlbzGL2wCNJ4MwCSnCYTsFUF6uBFphrgm7G+u
BRnt4smf4CLSjVEV8B/sLyHo7gOziQ16A4iv/IWqfqCAHbXa47LhV9Tql9FbZG6QJZ6THMRaO2rh
kkvgRBcD/8bXrun7dmZYLJBDDrOqbhp/xf57EMZcLIuGqkL9qVGL8CSlAA+n/msUJ3JWsuzn5SSY
uinW02a9Tpgcklw4MXdkeJqRRb+qKmX/oHUqbLxDWx/ta5F8wKjxqADmSqBMWzAjGzE2EoxlVt41
0zYwQ/RJrWiZ8uSNOS1J8bdP7wzlgT0ckSBglL9pP7d/a+8fBlV2ix06+fNEys9m5GhcHYNlIScE
my84+ohh5ufxoAmE9EyzynzAOemWqaHZ6PvvIVm2LQQbcpzgBdy52rJM8bP4gnrTSJX+PyY7oJ1E
dDMJh4pyDEswk9mOz24m6fFuzrAbIIvJMjN6sAbTdDZlvvUf68s0uamoL49vcKUtaDihJ88vTJY+
USujx8KEPOntQv3oDO/CJESegi+p2mF9YjAsd4cKnBaLqZSXgIqLGLbwRlU6TZ/4DJvkAS9Kgvcf
7pZh5u9estznBWi94mVZp0Udly08tt3GluRcizPro99nh5CAhfA3VEeNA/P0Gk6zILz30U2mnkLb
op1tvZyBs0JbbI5gvCzQW3iGCg0DLNIHUM9Sp9mbB3UTZk5mnfwcdNPdQhWSI+FfOA8h3l3Y1fal
eifyHD1XEHb5dQjxxzFOhxXRfcD5/WZZ9VGOy79rx8OBYjrAnZXE8WCmW0q9GsAp3YuxHe27Cv41
K3InsqdqFMzp0xYfb2r155sd6Fc4bix4zXRsS29oF1iKZYu0Lqdum/neGOyuUAuBErkDIRrRjMg0
mrT4bQ9jAwa0xZzz+DPkGwhkdaW2kF5UfPqaxUp6ZBwAoUmassDEZU9gGGvLiJWYCq/zIuIZ/S3E
TYCOV16ENB5C3tYOJMRONoNwys6jd5Mxon0kIp+RbACAwryEKFO/URJGQguNQzxu/BcJw4+TFUJl
sorgYTPgFangS2KIugiTGvj1awo45quIHqPoUK4xGwHNg9/j5tI2pmve4ZgWHRYpqnOEfsYAbFqk
wUII7sIQ9YclSAqmafPjCVCnxwysGw2LZpyKGQaWd7UwrbfiA6+Qf1vU+MbNbiGfO27qrhKQ58ze
l+h6yOdK0fVeFM3mzMsld1hKmsDLVzQKe4zTM6YwhI/uiZuaDn9xiQVQSeHXsPTS6LF+PIlguYXY
7cq/Wnoepv88jvc76PKCnzebfRs7P2VmIxfEYQFyOLZ5wnS1K8Dht/8a6RAELXJFPOdGJOfO+xhK
b+o+DazglzRzrJ3KoCDVvuUFrfGfY5xnwjJP8y2t0mb5E77jyfUD6L5WMHa+nH+3DobowTvfHlpR
QpXsvNSk1NOe4DMy/2/70DwOGYhkgbK+vIwAGe3TZ0QVevexLTuCFnBIgycOSeI4gNLw0nGRY10w
nBbayDC2+cDmo5KCmtmLl6FEroNO1Ip7sPK5Vhbn+C7Igf/6pRqWRdq0OhjbFnXqVdVUIt6DJ5Tr
1BPzlZalRoIE1gfJqMYmIewvhoSVtA0UjFwUbnpJ9fRJQKQs6Qb/SGmuONHjt/4/H9C3QPB0D6Gz
nwZZorKJkolkJDlvlCLsgWYaM20E66K9U4wJC/VnczommHqXwOHhVskX2CyETFoUbtKVyjQWstHA
9dSAdhR2EEEDHqa5K/EBUEtZeH46NtchyIZEZ0+Gv93WR+HwLkiuwD0Ee4ivs13Dvmgth7MKaKsv
lWMB+Zkx8Od9BXY9dUkVE2XzRSPUHN6bma3sgzXKpovQoEGByE1Fuoz3UIHU1eZOUPVEAHKpva2R
h87yHwzdQlzaRS/5mGekUkLkDRXaiJlrQJGp3J8D4anGTYA9KSVNynxtip/tSKEG3w66D0OFs5/R
U4fTTsE/23Xn7A3v1SBLJgtaqJHvVYPtiskZUC+9EOtPqopN3kuH+uc8p4k8lry36r4BZyzcUagL
Q5LnQmTp8lJJZwStUQpSbnjtmf65GJMotw5Rr6XhhEw0mtnKsMqP8cZwnypVo3tIDB5j98ICNAzB
cuvxzEiDNtg9GlfhRFyX0/Q7QAcsKBKj5921GO4l/eSBNijb8fUFPG4EB9f8itadnPAdBz+zPw6T
q78+4a78gFNGSAejitl+LhZQkOoZkVdMAYJsWT8f6+Zr/ZO/9luiL3Qcb6SzNIYX2cDRyBccYe6h
ccm00ZJx3Vl/sEcCOypO57Sx8AMjLu9oqyfo5EhgMXsN6mj56S6cgGI3apFmksfRcBKWddbByTNC
o0aYYIwGZ4VCGvPRnbn1RNFQYyr29+pwOlcyyCKusy8hDONzb5bCqgi6eV2I+Mmxy5OC+DL0iRCI
foE4B1SP/crdK3Co1bElJGOvm8NK7gC+iBfvxxxAza2dQR3TDS7OXvtyULHRLKvCJltWVqEHOkK9
1FrZ9/rc/4vC1LCb2CVUqIV+HMSujd1F8XH8D2uD+4T9q2L9t69YU/lhZv2Bmag4v6/iEPJDhDe0
Myw9WiIUzr+dkTeHvcEoEyGrQYMcYtMY5aA3++3svKS1lvIeVb/66d0pjeulfJaYe4z0GXVXn+kT
IsBA1RTt6SZD7lescx2pTcOQ7R7F1oGcW55OdOOZT7Ld8txtfLM3fSnJfgyQjusv4IC5oPRc8q3Y
CGxjT2uL7BG7P5SLmzRq9iKbndARWLMSun2BN0SllQXddQpwaW2i4zdhWndfeib8JvGSPhs/Xl6q
NVg35n9EzGNlMgrnhRen3izVxMPS9pcUlDRKvmupnRd0fD+YazogIyM78x1CaiTrbYo3uJ+m8QQ3
4/USvGsM3hiNLyfmvxrMJ8kmPeIdKA5TfrSahNNmbSQ2nFpTIdAatlIflvSdXkoGGgFsYg90WXCT
qsGEUDky8/APaSeNXYzic8IIiahPWFomTSsBZd248nxQg2w078Z+lnksOB+WzrvVSg3EMSKyfqX0
NhnzryvF+PoXzTbZ6N11PlJ0GaN2sUNFqyupdlIg353e9uQLW3hyMW+gH2AHSDj1yVYfL7jvmKlB
0bM0x/5kD7T3SvQvK43S5lvTJt1bt9mfx3GUmMV0it0hL23Ag+AKLvivXfNf5vuoUc6gG0cZDUBY
OSRjkBXyoMQ4pz/XuWuIz9ir7WtK8ykVS6BUb0ar1MUdL+8bvBji3BK6nic8F64IdsWQkdokojbJ
aSpN6jmn4rsZ1iqACfhHP6DQs6tdjqxlkIcl8bXARxQ4+WSKMU4IBz2qnHnUKUtman0Mum+sh2fS
3A4XFCuBuskyKbdyjYwNvkY9o4vdtj7c9ufcZDwbYcw+StykmN2Wqv3ex3QGeU7TGwFQ4abWuqNx
FPtveIZL1EKJZbwINdDb3b/vt75+K5Fk/kK4CazeHmihyABH3ynf+VdqPajLhDZebUUsZeYKYiof
ESPsKOO1nWclLdjv5m6gyBXy0v9cIoEVC0RaBXXMBDO7mitkOJ44DBVONK0aO9BXAgmDMRiEcCQT
UzDZlmOf3Jzy42BTWScWAQJRrWXiZPBhoHiV6DsaK6dLNgfA1V00zKNPSkc7C92b7DSO2qFpBv0d
N9Xq2xt1FFmsrrtmvgIAMCYYAULH+V5pzCBCkqX8SjHuDKN2sdUDGrZGs7gjom15OOEE3O8IpJVf
9hEOZ0VmdmzESswq+f5CKe1Up+V41Av3sLuLTTdTN9+HuB+h+fSlnZFQGtrVvqU0I5t1WyuFXS2+
PYT/za1TBvEdmZsqfG2JZABq1ELKh9tHk4KU9yCJNhDDiejB1pkViIji+Ae6G11xHv8uMKbPaFkg
8fMqJSnMhx0rrLXBeKCVB/bWQ4AyUULHfP8f8OdpdvzymTswVFjLqv4wyHaSfEoxYbmJvTHhWIph
OsqqgVeDUL3glva77vWpBQwDfPzv4f9hafGBf8LxB4/Dw519xgg7UYjZ9LODGCpoZIuEDiNIQQ5W
zNB1/+SYlx+jCwez9+7353mC9F/ZjDpEw8XTJbFyKs0x21ivKNWBwT1kfXgo4+mPwQX6nmVqVOmz
ff7C9c0Yc96Z3zirmjjBfX48Twyz+Sbh8xvPVuk8UPYsI6saV4X50sIJMrhBVS13RdwmtMtgzuMJ
1vmBoe2inrq2iDpN+UBzigPbk5i7QpPIgzwBUWdBSNBzbIfrCd241wCSZm2mCYAju6FFwDDFqiPA
X6tzKSdwMP4oIQLBaze1ShZv0h15CCGwYlogb2apAcCuLXo9tRAe5BEQaLN4DBnOfD+aWRWh/++S
TBKx1sRygBWNDf7bhls3CCvaOi2avX2mnfphmvlDchsqcF5FWF/ViCLNPlwMDicbZVhd1QWGZySr
NudDJD23z+sOVuyM1ybgG7t1I0sf6z0xditJHDnorX0T2p+hekit5p+oDIVKTGohvTmnOhS72Qu3
1sF9UVoHmdjKPPgf7d3qWnaqWQkdAbS6sOao4N1i8acYhvoCV4G88JPJjOwufhPd5z067+zCRYGN
uSqWAN1aa4RjjgW3YDYic+QlD0r6/1v7go0CCAJnVqsk1w9Y7bwpTfq9s+8efeOTmRX+9rA3Oxfm
vp8upC5PekAXvVU8xetHS3aLBlwSpgT8mRxFCJpiiv5H/0l1LX0Ud/IzvdJJmtA2ostGW1QH7Qi4
a/U4MKmmcV1ofHSi4hgtySIXmjgWUfbPQR5w5ABDYjuRp6WuQ9k4hmBqPv4o/KK+WPFFuiQ3VRn8
56yf/CqNn2eN1MhIZWMj/cXtrdimsG5KjU8C3rbkBi8ub8l/r/33eR98KtQ5NwyAJPHKtMIjBAVm
SBIUJ9EwZnWcuIfQ3rRREkyeK5U9t0mT6Z9x9h7U6FLxGzh9PfO6U+xeQ8wxqiT7gs5clfsXC1p9
RrSst78Tk9k1q7nvP64r2MfW6Vcv6uJkHws7AT5ENLIpawQP/Mjj11Mwkj8yS+hpYYjFJz7554Gj
+/Hii7UEA25YvA5MXpqThQd6JsSpeL5gNOnWg+B1QGrpJVwhBWuK+nieaAI/HdcJYlgv6xoVR0Xe
5Ef2xe7mGilXsRVguHUO5S4Dk7+hIzlOBR2iHLl2TJAHCC1lAz/FnFlI4pjw7OaAgp/aELH9PXTx
Sfn4gHONrXFNaI8oF50umjAYi5wiXgFWsZs7FrQ/uQ5sLbLx+cgGavU30FleXedZuKrwWLNHZ7vA
qS8ZI1bvIUi2hIEC44T3mzKlWnx1AWBN7rySUxK9892CNn5XHBCfOJek2YsVQ/4wtingvmi1OE2s
oEUCDLukwIlb5GynnKyniTs3uHcRVgP9M751GCn0xwTFTTVcdSuQfonIG+Y01cDYz17ppck0dgWN
bL4+2dkiSNE76ZZFal6ifYZdxV8pmyO0XVLhXRuJHUsFqoMuyEgmUJ+xaxKHYu68/G4gc0gCnOUM
BbVWGG0g2JTAIhZQxCG36hNA2lj2xXf2Z/lCoiw9Yyw1/E3UB3u1R9eUydWNM+XXhoOUBRxe52fw
keSpi9keIJjlX9NEG6GwBg/b2dAXMK7LiRVvDyra5xjtfqGRPMONGyNuz+DaaeM4h1uw4/yFyRTf
zu+VYYaTT4GbAdBDxB4FKLCugmvnOsEsq4mBsH35RFaauv4ICYqFtUOnPCF0oqDVHCoBF3/vWWmy
DETFZvrFH9EbbZbiuhsEsTyNFO/4T9mhZkZxWLBNSLnt0RzRgOaDaR66OILk7HxOF0QVTGby54c2
G2bN2k/t2n+7QHKr3BJLFo9TsNXRHXuC90AmR4k+B5ExKzUZPyv51HJ2I0nMWKg7jN3NLb2jYCpS
sceONs7FG30TNCmqO+wuKQwMC2dM4w41sn6+XrKjoobvlRvsDvyB9V140HZx+wQ8W9JHef8pOzhe
HExAPc4uSxmLECeAw4UJyD7L1F1+tIHTa0YuJkiHioA5afhWMXLD5pLBJ7xxwwDm1cYKe1tz/+hf
Xgzq+dK1MBqfD62lA3pbPqDcRA72OtxaWZ3sYkk5IWndr4CTz6ANkLs08LA5Ie+BqD6wWQmgwPYw
6HWkoJ0CyQOdfhGO3HCq2CSStkHfcDVmkWDY0Ght7FZNSjwiHfTLpZRluWQEk7F8med3ykLdupVX
h4NkLk6z75AVdZATfAUoGF+xCgpLGRsTMkb/6M6945V4/G1xkniPOHzmVaYxCx1rHDQoL12fOTop
R5sfY5B2VJheX9XaW7bcOYSff6bqkX38bCAAtWM6YPItz28fXoGncVIovqR2xbPtjdpPnFLem104
LSriTrX0/UdJNQDD/tJv0g6fKLNZGkNC7HlXIpfJeUXniNtcPEo1WxTYfoRN/Z0LFqqaTpqRs1dH
nOViC8l7T+L6cZRhyLSjLUW3V9iOe7+QiBnJj3Ux1PreUnqxXdQl0hkc2yi8YXgG3f6B2CTaKkJT
dBVaayM/lVCme/Aw6h2RXZiPGiYWweyYd65wB5PPbGtHU0PcisdQuh/mguueg8p6dtaPWrs7fSAR
gWI2TYAbRyRwmRi0+4d5gMROuuCiCfB+ZocI5DQuYLsalmiLQ+D1PjZzY2hPSRAruU5nXcKXLyWc
udXEm6hGGB1aCEeLrffXWAdgaHj26EyibMYAQJMlOi9BR9pwtaon6cBdYssfPgV0IpTSHKXwiMrP
GI20+cHCfMXqUE2cI+2L+cnFM8nQJ7yqmYlSDLblhSpwQebFVsW2PhI09T7SKluA0wkz9/zQTDbl
tJpmc7YJPto1VM8Q7h0BMpQv+wo9z+p0rLnv7j3hOVIe2ZHRDTTpwuSWvkSeNeDeXMVyMKXnvkH+
zzldJYfzoqirPwFrdjfoNc6pQCNd8pPWAKdJ8d/wWdU/uGzGgIVgdjeVcRbjr84+CZCTXsd6lYNi
jo90bxJtrJBrP0Mbxmad7dz+BHoLapi/Zv52Tl3IcyHa5wS9b9K7wtzeagNT3CPJlRFc3GUTsvYA
ZElK8TA9s6ORV6XPsYqqbz2ERlq/7h3Lm/c4aw00bbgp8NvQp3aNnqINyMOkvy4BCmhkSJFOFW0X
Y/xVlnW13qC2lC7HintLsSCHQaW04zioCO3bwuETuGqaSNgtfpTLG5txY91kxalA9VqHMDHRCT+J
JHGujFUlNBLyVT8lA7kHN40U4FQvQF2mZL5SQ3cMcajfCJKoo3k7zE4lOpwSt2a2hxOiMy/Z6yHn
Vrt6CzjGunmBr03b4dPzItVPBjHzSarWHHZMoZpTNC/kLJyGVFT/eVtF9Gd3Yye/JL39nnqY0cF2
3IIJIsfwHGNJf5Zt393G9CNMIiKZaLoUabLQxUvpEUlIzZXw9BUbR2rA3aXlG7LjML4o0M72Pnn8
kGpWvcxQOY05wDtIh1PaZmDpiQJBjJAWelNl1fV0m+X8hSTLwSF0NvpGezJRhCpqJ7EhcLPaBqwc
RDJnfrVW428JLSu8BJ5zQ8gLt+2b0zIuyPjoSh6A7JcmcBU17IRKNdnNEItEycpF2ZSSceFxXK1D
jFAXfBeD36IzP/OwTq5Q6AanN7R9g6WyElSH9xEDTU/GflOwpyg87maDE5Kv6leX/8mCBpatdkVE
OzGfS/CzRVBrueuAUNNDetXL+oP07IQ8E4KmrTjM0DnjIHg783tViFYRDOCxNG59+GpojEyMNTzU
SA/9LBq3hobHLGl3gfwQBMUXsejV47EEEcus1dkjxO/BOsDt26YrOMdbCMgsapLhceOnGJqog+m/
TxU+fYnF7G8vyz2nVZxYjROPZm13V+cVgY50jRgIGbuEaw37ong90RB3UoBNqMpOg0b5UoaSFD0F
Poeen3LXjG25iXxDBL1eqtRRsB6VhOwVOz1YY7jIv/ekz1a1dGc/lsVeIGWnWAcaEFsOhwmTiZ78
7cIN1Q/x5BhcFXpCKl06c65GYjqPJ1M59YPYergmg/oOWwMPDu2TqDh7I8SVGuERmuG8Bz45p0pT
d26K1blqTbin7i+atyNknTvGBtCgnLg7F1563raPluSMTsjMDSsSziMbja42nJw7FM0HP0NqrRHH
xZ3ALk1UiUE72HGBs7AU3hMEjCxshsIsULUBXVmXFkEshfcFf6Yyne3ZBYS76YuOqlVsHuJ+7+f8
Os/rtF6ypKlenowYRQJBsJnFz5L3MKoGfWF9t/WsPJhNdplSonMXFuhS4YXRKfLoNiAKRHultvq9
XBdJOJYygUuykyPEiXY6kYRYkmaEgGVk2UOnQLzoJTN2FF2KLwwocZ4/3LpmfTqiyHiYMEgSvuq/
jupHADsscKi5bM6mSLZC/As1OgwB735N2hd3cawsAd9yb8rFB16OqK7ei+a5ktpSXEe8ouwf9Ins
WZxvIxadQpTIa91ElWvBIJd3XROQGvdoeYhF8XnJybt3Z1tmPlMsgXSqKWBSWdtUIXgQL4IcVxkK
r0oRnNoFg2PsxEqq6+AfeiW36pRChOTBuHd9duGpSxYDpoBWNYBSP01kFisgEPOmEy1uAT62ybY4
eCM8bz95WFjYxVJ0dysBgxnAwzhMNlUeox9VHj0JwM14fo4F6GjrxOxGhUFcHAc/9xcGo9IUiQ3i
NT9s8Yd30mr11QfGCUxsu3+8Z4G3MgN1GXo2lS58jsdUtXg3aQmDk9pho4gb1kHZC83DY4Eq0sEi
DOx3tELQreelJ+77ceLOWsP+STuAGUMYE1SjkKq6wpeayDMWrgs3Ir4og1aVIEl60i0NamepjfVq
9bjziLjFxYZTGtZfIYkXah1/ikIvp1KuuAJ7rKFWrirUBwJxZDNRYhG0diKY9cuIVWakmCbR5a5a
OV5HEpZgsR4gDde32wi8caD0c2eBsVqYVe6xc5kFYY1mS8a3Eh9JNxRsoZ9sxyTCGLGevIhd/z4W
Mu00crywfkh0hRELpksWz9FiAlr+1nhzMuCS+esRIsu1jrCsYbjqCk+O3fmn6rPkIfZzusQ1CYrA
BSj1QQBxE5TpvvYrXS0knZmyWfSUobuj2ZnDI5NCIlUx03vd6NsLPwpqyQZcc8O3rr34Mp96N6gs
Pdj6pTPLGYGcGdREaTO3P8DchwvBkePeRBDeTci8tw1r930FOoFQJBxI+tjChXFl0A/UiV5mnI83
FEUVLIQZ9eb2rYKNgkEV648dZhjafwywJuWLr2WH7QcWNE1S/r/QF8XoG2ZUj0mnmfy8VYLsUp6A
jJzgGqfIILU+fIH2lPKjuFF+S5B5ox2FwVNzqs3iWBZtmAFyZ+cOJVv0BmW38o9JqB9yia6qn9ii
2Gxw0ptQd4Aye28FdanVHyK4Qzds4eL5LH+3WWUbzT3frh8i2oEpIX8A+Oxpp9b4w/PARwEGiDHX
xCAr/tSvZUWhIOdHKHrAXm7jhNFbK9b38JOEk9Gy9B3JxvRNllsC2qajQlfqw6z5fiUWpiRMtAjH
DigLPIG3mQtxtmK43YRcnHlwWf1uY5lQa4rcrsR3pfpta0rGiDrD/hANCpFMc+lBziIqUe3HAazx
nEe0pAZ8/C8LvvRdt4+mghVl+cPaGAi0NOoPOoDb7hZNWrPPM2CbKyop5xOm+kjhonvm5/hMzI0R
Z6mNSXgLdWNHWmWG2EYaJ3hgdR3NKGgmvQskiqpbQdH6KGqdztXUDp96BbBHNmwPJ5ir1OJadN9p
7OlV6n7A1X9FARf6R+roDAO+cnsmakldwkQ3OXJRKCKZwmTGOsqxmyx5GvlZoOmUcWVWUCqaO+xv
FGAVbezwEVzdQDRSf57Ehmblbx9uCQvoW8d2Hyuj0L46MaXQVRGnuzUQcfrus2QIIz3FGXT8QuPm
9LVRr+RKO5rSpIVxgRlH+qEZN7Ryq1AB0AzHLy5XRvrfIAVu4/zSlAfWh8SY0XUD5T4Q667CIUiq
2PdhercNM8EzuauYX5OFonN1JdhBMiT3cos6Tmw+QMjCY0nxkSaYHkx2pE8sfF+DsFXZVtumbQqx
I68hd1LMU06JeES9n2yyaB4P8xnMVP4mtch2qSqYdTd0libXU9ECeu1/YUirw1Cb3ph2b55BTxXQ
rBYkMJUQ8NnSDGoqOo/QrBvEhEuMsfNzEtq998G+NIeBHE2LKvnU7EBy949tS1cFZBQePQBzdDf0
T6Wwk7EKoA9CtI1CmbBe81SACgz4ihXNPxHIWdwHPICcjQ1J7X9fBz+YAcmOgqARMHwMPRw+ickh
s6Xhf/0QFhJ2Ny38Gnbn9WNClr5UidJihnKFozCgU6q3omN/9H9XF5guyw39zAbg/n3YUAv5XSrP
7uKc9fKomqKZIWknYSh1n/MAn09Otr4VGnhOg+cPMQdG4IaRQc2/CY0uFFDTL5NtWIcbh13a7MTT
Y99boEoZ7WtIWp738vRdLOoVlBIEtXx9DEIYZ/HRf59gWNJdUIH8lRyeW+He+tGLPGLDyHqm1v0t
N/2CRapwSW9IUIQ27yewuDIOwk86G1OTmSDnfaJitqalvghsy0V5ahNdo4+aRrFML9C8C5Wxm97S
LK+6VdLcfrU7etb59JL55Q++ENs5RJiiMnhCeFp5wia24t6EDDjr9dBcnSySGtOI4N88qtjbIEwv
a2dtLvVne+ca0lzzqeDGS/9jgEj37G0keZJP5lZxlSrGLYM00/TdPH5MvoMMz/46cLKGcHsmLvnk
uAk5DDR/tcmiihfA1Z0lkNadxWMi33Nv4MHIja71qwYnNdROmAW1IY0L8ggioID50cD6KMF75NR+
rR2rX350A7rpFELLy581CzfNO2SkDfUNZhzvox7fyOwBem9ckUDhNieXW1aJi9ldAaY/tvwUl33g
mstzo41nSaV9wlFbub76TX+SWyyE3cDpkKtX3QQlWGUVUNRecekLZq5cIxCjpTBqNewdLJpg5tmx
HC7xcl3kgCiss2AtjOAJkccIEzCpZejailgZXxuy0gtjAj/aUEqy0gY3yAp9a7fUdt939fsHgafg
ZlE0JBHxqJOaS6V4tZxbxJwygAFqPnZjpyfTtEvqWVBcLDv7ijJNjBJ3eV1JRntvE0rX9dIc4bH+
8/976JyMTrxvDRdDKv4iis2A/hTIXZBEhL0Z9g2AC2gkNSU2zxzoMWXqusESEU4OU9XDzKXVEO4/
Sj6oyrYKQVhYwXhFCbavVRpLypTN6JoS5wP4wAZPgtOof8iqABxUFH376JtAwytX6PHU5HGF6UmK
7ScXNtvn3wjrPzW5awGquDL6zAEwsprjDpy5mKHsknkgvkIi2n62I82mog3AwIseekr6TecSIzVW
BMdivctkxG4DS2v7b+8eohmoxPrDZX9p0tr2NAGVBmMNouYtqBuT8rOa5Qw4c58VKb4H3tSYQBWL
vK3PMKYVgJvzyjmRaxw6kSXJIha4sa1Q8cR/bG8yp8nOiN74cFJn+UCVi8edvb9BxBRQNMWizwJe
RUlJyHGQjvdE5wykGZmPR+MH2pIJCCc7qDx2TzganWn53QW5rQ2y+5OeKIhsC3d0bgVkaMuaT5Hm
zBybs/NRvXAsfqaEVgEcX0Ff612fU2iaw1uAaEZoYwoU31/f2ZCoI8TRiETw135WFF5eV+x4gdLl
cwaJnjbaagiNXhLoB5qNlaVWuNhggnVXezAh70GErPlVwNCmWe+8swq9aQgN6vqWVfXfhG9kUgIL
vCYcH5mlLNpzrxYZTImV/zrvUWjM+otQGJOZDDVFj5NvUnnyC2f1JizBFpHAOgDlNnkNTAeOPWlF
kmiQJXJnatfhtjSij8Pd6EOifIAN0T2xreouPNN4miycbCqZ9jF8bA+FZBvcvHbDHP5u6ZK9LeJ8
sZtC4vu5dNpB5bCXaG3skFNF9axRniH1efW0dKu42lV7Evj05r1ydXKV5cZlgAkNJTuNrhGv/VYr
t+rWsxz+cc7hl/ZSgHJqDCL0VyqeAD3ShItG2B5IQkVdMF7ZwZI9nX765Lu0mRJWxs6Dm1CvjDcR
eFWvn20O9TnOabLkAi3S2BF1XToGwZ/i3oBJ7toXQQ4W6PmfoLXYx8YSQU+R0COUGH+WJmkkXd9j
XJPVqxkv0kmh9RPTptjs8F+A08Wr13hxazbFMlWOn44/q5eYb2fxbAJJrogrRTsaF1ht+iGH0e9o
CmoZVBtcTtnW7ZwX3oASlz12vJIJVFYMbzFBLF61po2mt8DGwwPhQnwlCElElOFfgDG1q4QDVhvi
30BqVMlODC16rFy+8NRopJCpCqrWXSy95h9DykBgjSdGejhFgEEr7yUGBljBTaWo25FPlhNM9+b9
tI/p4hWQ93kIwDDc2tDl8uEgnoLNjNDahCVwwmWa/P7GgvHSQI8XBCOPE7bkIpzg3jZTN4DLqbat
ayODAIUUsgv3KfMOOjLGBExXUyd0wCtzp7ZuyuvhBb5jf037CCDPBnSrUCFSkiV5zEvkfXyu0cSm
9DuPB61dRj75SR60OQYQ1IOfTaVkQmht9pxqyax/jD0BfuulzgT3rQHegCBu2eALP98Nkka8lEuO
dshxjZ5mDlJel1Q+Cu5j0k+/XYOXpaTiCu9DKyuJwyQxxqJlK+mUyoWRqcT07g8iX6ob56mhtn2Y
dFx9wvq+iEOhWsl8wsn+PSagWWr4c34touytCSuuO57RoeBgxolS8U5iN8zJfoGaVbgwjBd2ZWXK
ao0sPuA9egRKxCoOxba1KEIcJakSseBOzYlXcdJXCFkXLb+1p/u46dX4xi1S2d3+HK3grtbm6nTE
/bCvVlbPGWiEfRxpzWxXFq7Vf409JDOHQZKJMzEhSk3UyGm7afUuIdHMCW3jNSTCrMj8zNPoFHto
iMC+8omUKEFLD+ldHmzKo9zH2hgJvfVePi4Gcq5VwEJYKfgTjaMT0wv8hJOFvBGtYVR2K9uru7Ev
7F6golo5WW/enGJRuytREN98VBq3Kz5UQmXmYGZwONEscRSTH3XC3dyRjzD7TfS/VhH5WcmC8qLw
zYaYK8XkoofRVj2wFM8JE32ptB6EUY8Pq33jYdzOM/iuSfo0kSr8EoIBihQhCk5bNI8MSDQDrPA4
XjemLBJGasY8KwdiBPwwY9kPlACvIJZHMLfPDZxjnU/jsR9ivm70HwThCycIDyqAvu3bzsfIKoOo
O+i58KeEQVIFpe/oL99oi1n/+r+iSEFU6uKxTpUNfn/rB+KzDOgC/gvFoWHlONyjW0SchPqgnApL
EbTjQ+4d5r+9yr0VQaJQRnPpgOeJSz8ZTHg5kWeKt0LoKZxDoJ5ksyMfHbQCf49bQZiPrtRiyfx9
Dl0pX46Q8/7pQgTes5GLzYanVQAu3SVfSfBOtT2DfMN8+rYHeGa3MhDFu5nJiaXzaGQ9als+MVhm
00lzxTQOZrcxWGpsV0MLVarAiSmU3MbrvOI9kGIHfPoJseV6nhwlxvoUaUDuvZLLx0Oxmvt1qiRe
Y/9mc4/hbHUsS173SHKZSAp6qc+x9WJ86X+jfZ9XgTtyXRrfxOQ+CkUs+KI/RdBT8qKTd86fjttb
LbvdfCh9Iu/Q/otT2FPDo+akeyrEvXMFI0UvC98GiYTrcIJ26ttXH5ydplDp+UMwyeXv7Pv6fV5n
Nci7fHIV673xcY9AArrknQDh6VgtCCisbC+Hf740aYYdD7I289pwNtedr5622S7uLjr6+UDeobP7
udjwICj5jAfAgxMxBNXvwG4zPUGEakGHI3L15AMvlO4yOL1L7Na+oGea6sItxLKMafI0U2qm9JHl
tmA2uCa+C/g98aezWQ/0RSsSOONG1WaHF6D2IpEFT3YsuiXH0qwvEX6yTwWxJDanRuoGu/GbaMA8
ddiLiWSI+HEfkgAGspAM3SyyJ8Z5hXCy9S8g151GbLlsQtdMW8VgFHvI/rbP1J/dgvUJhhmRcHrf
tvncsctG2WhyEIbavCJ1VnYOb93VETqgv9+1BnSjb+DxscIG+wXolOegxj/XKg3R1AjFfRRroU+k
bpxquPKmdP73YhcZneMin1B7xNi5Ztpmi7bDNBa/KBZaPq96WylYDVq9TlsXuJJxUPum7rWqBVQF
BWBYR0nuShMJRp9zvSZWG3Vgif2I2E8ss9Di6SpSzHmvXlv0jXhGaintpXKdtxBaigYalx03M92A
nUEwwwKjbNAhjKdJOUh+54Sj8R6eKuLp+XcMpzr0Omnd6iaGUtWnU9TzwXItvxk3mg9s/PNzzV6d
b1m7Urcfw7HDv/0DSb46iCXY/DXxk6q8T0QkS9Nbg05F7/sweyhNi2HoblxYHOtfAF3rxoT6LCMA
ArNxZq2jRcp7vLAykPnb+XccVQtvgAAfprCl/x4pz11bH5WTJMlqSpH1pRb9jd6wTSgb7ueyo8dm
jpajg+bBw53Qoc7kDUCxhhloySJsxOsLxBlpOfC+QobWorVWNthzCsx1xGajVVj8OwYJvkckFgid
g3NMXm6X+3mPvSiyQ0EXtuKOGz6pnmW4EqnEmJVLUQgIDrpPcx8ZeQOBRlJsucV4wz2jRuZn01aK
lsVQquPAyiJTIeoaV9H1kkoapAyKO8fXOsAMchdRo+aLO0QSVjmlO8crIAW14V8aHy5ONwsAFsdq
Cl6+ETimD7vdbDJz3EIaVm0jb/G2bqdREMMtlhfaOlXLBhbOmi/2eb1uJWX8qpqosO76cgkTUlqT
XjGmg6W2JEqXMsq5BONnsKZapsJ9q0edsRyT4++q1fnu8lTrd52VyPUqHQSH+YP8tbspHJsvgOlc
celXNM7gZU59s6ckT2Z3NlhlT3zfCLk2TLJz7jHbxHQDPgWRK3fqzTFB3rsoUv9HG+WfRFXuH3+U
DR5VMONQfamrcaxBmfyWUBoLGXFsS7IBjUi7D5UPnqQjtMGnofrum8x1vzlLMehUs53WGP1n/vCm
nLSMb1s2aS1gcrKx6+D8+kt9UFK6sRe2z8BxK2Lr9I4pyDUOv66viWGNllNsQdlbTgjkSlL3M7m9
3czYnffZ7Jq/ETPwi9dU/erxJAJsd7JzSC9Y5meNlUnsclQyrAtbkfAFogr4pqlTp8WNAhiLHG5t
6vr7pLpIfRyvFP4lfY18cPQgEdIqsNrN8NBBpUmoxtBpgUNxA84paE0L2v39+d6MNO67iNu81Urm
VS2d69WVGW3D5DtInlixFc2KvjQyvG0u26Sc3PvvCV1deM84UXjXUfXmk6JLyR6L3Kg/VHd6rlrm
T1v0z02yvKOSPE4T1JWQLcclSsZjx2+f2uj+qAzklPzqBHvDK3SHYufWufy+C3lG+SCSsoMxc7Yr
hVlTjII3z7cw1cGkUL2G2ZjbIvaFq4ixiDLmHMYzQ90UJV/F/mxjPBI+NqFdUW21p30iRHJz2xvv
DjfcU5dKjcOQn7aF03HgqFcU+B894t/zytUc+IYfIX09CnL5QQOTPUKsJNLDrOuVV885Uh4R3gpS
8Hh5DjlLYDTNR/NvThSBIuGTeWpcczy+2tEyhD7D92YWLK7SRlEx8b5OzKXuHyIZeE/kL5xLy7i2
9MekMGITdxEkHT6lZdbk6+BfuiHqBQvkcdJVUFNfKWjI7dHiSopa+rmOyTxbIkqpRIEc7etEfovN
Jgo7/akduJI9fXEYPAjblPGYkQQromHP9OqqEQbMF7x6JXgj3izfv3WvQ9ekrEazSeBXTdxOY/LZ
bVEekvQUQhZo4ITR0+eWyZIG5RNaphrfuK4UnTMz+xb70qfjQtOw18qS6mX9CJQnmbxfelH0YBVz
llxzks9qRQgrTYdMEQ0ZKH4ZnNKurYTErLc2tsrWCACVYJ+WXFGn/lGAMk5LzCQ7qiILZuahs/nj
Bo3EKIf5nZ9bADTWneuYcoyKRScoOarfLL7NIxz282qct2v82dy7Ioi/15pPbqSYt6quFET3+lGo
KYOyPfMaEsEmyLae/CoHjdkBa+EX7ENbC/dce9PfwspxNAMOfW3EY5GRE/YBSQjh7bQRSyywcMh9
Dyas/qvv3lJbVu+Xf1Ejt4PWoHWpCCR9KJ6DboObpuoawEpSE7Hpog3TeSam+9xMXBV4fr/SU+GM
V7WJRx48XmLpBXMxlezSOxeQUpUsH5cBn3/eOiwT+TES8JUhDLS5BijfayzU0A2h5K+TJBbh2pBG
C5tfn9S+kMC47qwaSA+D/yKW1KYDf+8XhGS/qDODHbb7nSxUL8Az5Sj3f0u2E1BnOumdS5s8fuAB
j3HyT4Z01EedSFZQaVUccFJfQiReNkuJZmkhquW1Zea9jjsiZclJYPC7PpZVWXSorURWibl2ynGZ
Pf7Axz7coz97QOyJ8/3N7Sz6Maka6iD1xUsWN3crjxvW6RjOJXod+f0cBJRtYP4+8CAjt6xKCU/T
Sql5BOVBfoXuTGuePDQcau8NbyB/iM759gnmtNOqtOytW88b07g92mPbfnMeFBJ4PVKgjp6T/sWm
Rp81MFxwkqCYZcM89K+ToFYJqFCoHPScqoX3Ef4cagbD2mKlNdkfbi8zguhPxmV1nUVPCBuRStiZ
BC1Uy+4sMZ2rfxSrWCgrAslaDQqxJCb+6eeVMQDGHnCAaP9GsmYxnjJCV+1JayW8KvNAtrazwufy
Jhd+Ot3IKl0KHOZnUQrwuLWlImxA45vCdZOZ39qV4iVtI4zMRqeFqDeNdeTVlydhycahMiIlRGXm
rHGUG5WewGppHlGlwQh3DsyI4uFEUIAs1XUqde/NZQSG5E0/GIVsOQhLOK2cyDbGLXGv8prOe9QN
Mn39u4e/oSRw00jOcU3ZGbZJqC1FwlY6Dwup+hYQ6U/JrTnQPOstuqD0KcLZip5bKqZLa1n+/7jX
lBlnYR1XkiUuyPUPIzzz+g0R3heEt7ClWdptBnuQ3L6cXN8NRpO3Aji3cIK/De5E1SF3qpXVZlpS
6fORPdCWGLztL+4QJD1gzt26uKxW5ur0I9eU0YxgymXZwPBSjwfsm7jBbFMpUxPefQSJ/oEeD6aY
S4DFOLroX2u0PwvuAFwhbWkdBzWXGKvakVN0KqN1TgTQNUGnFTbaI1eBHp1O/wN7geUZhzviHp1j
JiqU0XLN0xngruhjKL1zEVG8X7xHtQZryu/FZAKvNYjtPI692hu6CC4/eLArY2dGegMoYVGJHiCw
GXyDSEZB4MdTengFzVAfzI6yiPn3sBzJP77g3rowEGOvQ1SdutHpaDu6mAdwx5DJcMi7bcytgy7I
Ai/qrPRdUISIA5My/NGJw8qU9kEyOrT3aZfjHBVY4TJpmgl85wFuqcofIkmJQI5P160CQl72lpI5
xYb7IM6Cu+j52Lvj4lx5qwH60pY0Ij15pueXuE91GmTsibknaGu03eGnCD7WW9Odbawg5Y7Do0tN
wKZ088zTXoDUF+7qv/gAsPgVWg7MtmU2OO08V8ORh5rFb8F/Mcdxgq7BQxaKByxYvHROjEGWxk7r
uDlYu2sLs8BN19vuCxgqmbqW9QNiqzhEn6pWwg1FZIHQE5pa/8sOpjeler14NGY8EgT7nL7qtnC+
FUSuBGSi1fopTmpPtJEvFbUMm2WyStzS9aAH2MxbAz1FPOYplviNgZnU0XWcQ7E3aeTc0nxRLP5t
iFAyINawUU5wSCblopMU2IEY1v2qrMy4mR9Wv0m/9aKnu0lQkvJooRjg5y5WMmFfAa8JBrNIsQ8U
ISSdneVV54iWXpqlIynwRx+qdx9PloXPOCVDHp8yC1+GLn7TRhUqujsi+irkQX3LwS4SiA5OuIJW
g9rIJC2p/5ZxyE6R7jeMEtNNWf1iUeLxM3wt3gphQqi/KWET+b1lvM3pjKD9TbF0LH+Uml89jOAc
JkeWNZ14p+SwfBd7S/hPTL5mVq16xLaZGtX7FzoFKxFKmJQMhC7tnRioyCTUz1qr66D1kEF1GLX/
r1A6SvV3rdNPEQjamQmEaiJMBzhXgWcMzSwd59/DIvyOkxgnsHZfJWmvB/O+k3DfEHhRCua23SZv
2eSI1re0o+NE+ImylfQqfVxzHW7jXZGLhkM1tU4I8PUcWgghpviwCTR2UkxxTcfuG54zDMX4tMca
iPLSoqTWF+7O707u9wXA/ZkzY9VY9JQpkjv9oQx56/dLTgin/q7S5x0qHCgwTPfAGjyS+mJ7cj2d
emWfl8W1sLFFy0beJ4jQPn0esdf8j5nI+6hUlymgGExikJ5MhxnaXF7TG6VSetuRmyoTY/UPDoMY
Y9fG+KxkHeAK7TmQ/myb5QMvMYAsa+aKaUTFRiQikVwGQB2Eb/SiR9DNUGLULqZ5wmu12rmdBxRI
8Ro2sQWl3z/Apb44KliKyfep0rkULalSND3nsYXB1+EFLDddJBwXVWYafePSt7aAJiE5e5tTf91P
ChnCS+5Q17aURLl87NBchyE5MdNQ9mXug7iE5yC6K/S+kV6S9nvm1uGovV2FKPufIQ2/iFGzmhZo
tw/CUc7XNJLUHT87Y+FMG4OzUAZgagWBer0IP6tdBvHEjFwHomM0AFHS7LQJADRxGVzI1yyuuFFV
PR6zQ7CVNBbnPAYzMMNMYxY5ync/ke1D+y1PoQoN5oro7IliEcrbWGC7akJcQMYYWhidPvlAv3wj
Sa72QCjN5UuljIzjNKRXqJM7qCtGIlymTyhIQ6H1av3WvY3kBYLwjHTlV356kOL2JhMKKKHftP36
8CTax6Df1OuIu0Gyn95JjiLf+J2c0Bi4i/ANOddXe8PMRNhFFC0zLa3c+XAM9Su5LzBjv37u6BeL
pU9uZujrVFVP2p8EqDFfVD7IiGPm8zabegjZb71CQ3UC+v2mFX7tBhplZcB0+SS1svsx3Kz9gIiO
RDSI+A3xhm9kDZAZT+grPI8LCKE4bHrtkWA1btzei6W63k81Jq2XcBHmnmtwYRBUMEb6O6oGvY5x
INvgaR1srLA33t16OzbZtMpiN3FtkDgLl7JdYeA45qvejLTCm+UwBUb60JyknqpdYdFaP5bNThrl
oXhRufq2xJ0GB0xgj8xxpWAwYyVNcbTpQ3kEKAYELXcGghDD64jS8bzvfTuSa7N7qFH7xiR3BZRg
6urTsCgi9HUbhz8Vf0cAYdlqOqhHsiNfgRL6Jnw2gWVjgG6rxCKYXDacaLYqL1YfaUWQkGmo5nSF
u+v6FaGHdfT95CjgJAJp8k/RFhWMVF+WKQeuzzvGPAquhLHtoSAJqy5FuxZqbWSwT60cs0f30YtC
L0r3hycsX/ZOD51v4hsfcY9DQ9vxtBzRW2yHG2kgmcXx/uB1HgXCATr7RgNdF4DsItVJcoKs6FSN
wWeV8/eSxNSa8t9C4sNu8nJcC82GhF7lKh1rXBQeq/tDJ/4vJjlM9HSuI0h7e4+sHtVJ1goF1jZH
ZOby1MY5sXW+HMZcJSHVUZgx26piS5STBWXyd52k1m6e2MR2Pg+F3wu1m7ZE7ybSn8IWs/T/fSL4
D3snO9h6b2+Yka2cq/2//uH8HdMXOqSHYI7YGzhkmDeqJwN035SWOvcTHlyiB/8HaxqYHhD8qa4w
A5C1+y1bhkLJ9q8s5lph+qad+XRUslgYXbSvOFDDNFjYwps1avGE74HUP/qRMiTESz9o94gHCUI1
41+uFW4exuhaQ6u6ib77+kl4wBApAhvVD++FRXnL30LnrlYhbIj5b3ppBYksEJSQxBxi0G1R4VmH
/KwXhJcYJlV6PbHHXvW7QYiAge1HvcxqG70lnfSS02A8WsQ/z/MYkgy+E4ZNHfF/vuPHJ7vXjgRC
Q2esPXSfTy24Uc5DnyDd3OukaKZ48ZA8THg7aUjQkgeO9e421iHfS51OL72cyHWxO/dzvIfMN5RU
6XKS6o/2httsQVY0OM1yRyGPJSVZlv2v7bvrFa2mmgXb3rmbZGNsiDP4BguYFka734josrqFcxf/
5oh5GF0qhpRTkrqWPBnyBpuRFn7U0XIGWPCidHnwC32Jo2Dqs9LYUAkj4RxPVnw4YtxD/lLbakWo
ejEUbbFwlaYxXsHCJlB1d2Dsg/EO1kDWG8meKJz2JPkd0FnMz4hNoXb+KisFp3riKdweJZHIPg7s
2HbFeii5irOQ5zAY6v70DH+v+s+NQnUkwnrWG/4+A//6r7sYb9P6Own9kTKMj/nVGQ4XEe+A1o8N
qvFmHsSs1IEfI611cYyxp7BHSsf5xQUrYlK0GKAEFbWneRCwzXBlI8Slp/BAXW/jd9fN1zOGNC6b
TX8a0xwcKDFoFXeeOBZzAsG6MgxV5Hpu1iGi8nK/A87QK2oLoACqkPHPAzulEf+xOFsNkjnvJcKm
B29yizZouYl83YUIWD4qusZUSjs3CLb1zq9aAu8fXcqeohtkfLokjC0hgBAtkyJjcHsWS0sY6c2J
dHXXYFDB9KJwwM1bjqxbmlAH55CajarR5WvuF69SWOsYsPRaZ6Bw+/DZwibQpMse8WIRPsPIuqiL
XxWSXBu++3OmK7Ucjy5U/NX22H45s7KBJJJ0o1CIlK/krLvKzePzUAy00bw+nN+2w4lKD5ocgSEd
RQuS/FIeUebBFmMFysQsh5ja/xTJlznX0ZfjbV/QRH5mxpbutBmfef90y3H6YZZSE2NUxbHVfP2y
//J5zmRID1ikOLUpB+yHVcaizEFoAOzJ5muXIg+TYIti6f9IiqRI2yFs1+3HaY6rhOsrtWGtxcwB
/uP9GHzqVMd4UYWhHgbmaft8rp1kQI1jezbT+1fiO2J9gWM8Zt69UbgP9Xj7UzoSfjyNGSSHaWtv
G4otm0GjhhuE1hUxRb2tW0ODKWzQLkDGsfMxQ/ewq8K3O3o1oAr1thQ5nUjM0pedvC8qFX2U+Xh+
FREQ+JBrhGv7FXyXdnW7pJKZDJ8FQHR5qo2Jm5zQK4r9NjjlvXhHUqidq4wA+6m8W+4Lkj7+toTK
8ILbNUl7nB3NgcBkjsu53VlOG2jMnsTk4Ap5oz1KFJF4RXZDQL2BQSH3UyZ1SxynrP64VdpM0GPM
BO355Wj6GHteAiYiEAnj9unOYZ5cb29DniZ3W+itCRzmSkTWgyNaOiWo32/+b0QeUE6zTOUIFPLi
iRpDXVJxzD0A5ceydmc+ibJJO5zYKNWqS3IbA/f21MoNSPPSJezD0v+0du7mPp5kCimdsdg8E8AQ
4SjXtkblGCWvydb7Ku+QwlS4nWHU5ijCTwTKF0cv01ALf1lowUC0JuRZdbyTgjtLWN/uXBoGIWp9
FE0oQvly5UawVsIQO1gZ5BvQWoWirGvgMzgK1ZrJRN6CZZOl77MXTadxh/vjQZ6YUwKHXjyFcWbT
Ih0qKf58SPTIreqAm4ipu0+RN0ShITMSpgB9dlA88cHmnzSFA72W49QknR7xbDwo+zdnFtG/8H/4
rw1OXs+KtwRKfGgqBoAFh6/r03QQ472MlcL2Ozt/dOUp+TNIEqex7kCzjjOKanSIM4y94UqnUbzc
BDlDCDUjjOASR/WLd9l1Kcv2yTvAH0kWgMEgIMgnm3GHVKYyf5IKiYt92T5ERx8ucadiPdhT+dvy
FV1J/TTRwBX5DfwzvW0oVxFviN6ARlYMUeK3qU8Z33WslZkk2xe32s57mDiwMTHLK6OfZa6pj2+p
sdAEwlHo0A+LdsAVXB5ABddcOT/OpFCVsZWTvXRbVQ4DvymAyNylrBrKQAgIxzgjyKMDNt+Rs4uA
ImLwGKcIAVYXoSolzbpOOE1oIBw4ORAvHWjXPXJxi7BmbDob+VvFXlUirVa17qLSbog9KKg2A8XD
5B3z2ViMMs4tsoLHs3W/t6so2nQeoTHT/n0S2KNw6Jh+lxncuszbw0GddMYUOEmgR9lL0b7wNWN3
egX33frpSjBrqNqexCZ2VyTvae4rKhOJd+FqzU8kdiU8doW4R4vz5e+yiEWl7XY9czOc72CBhU3i
c9ZSPTrGqziC/W2zJEEwqDo9LJujJEn0vt0hwBcyOwFK+mEmrmJb2d9IwTAcXAvOJ9aQ9hY6Lsnd
RHBLy1woOWx1bkI2p8AmPNi42CdwBc6dK+LeTlN+jMQsbZbAn6oL8n3Nus3KEYE0XwPSR4yk7Jz4
T1nfFv4YIvSui3t4DDOZoSRxGm62oH6YAy/tXlEPRZcsIG49BLO/Ref2HTvKyQACf7pDLJhdyGTw
qbmZDOfWrKGC6Kyie0qTWK/dIvJmRU31gI1WaxPCIgvdmuQhjiIwIGTuJEdxARyNvOLzQZo6Jbcw
hMCiwYh9JvcBRwJcFe8z7jHK7WJ+ItWHcKMRKgokdMDrwTgJtbSmpAToNIlK9riGBIkRHKYiRe3f
a9ZjpmwtGlFEzaDOsGVLggnGKS+/BetCW90GbcD0MB12bGMQtKexzfQB6pZv757LrcZmkHXzrb7j
RURvzxLF3Q7DdUwnNTJdOtVS86bYKR96x/zKHlGUmCM2dTu3iNAwYZl2LS7n1vUNm11q35bCBkdk
mAg1t0GcNIpX4EjGCl1qMcaITgO2MbYXEoIUbLYb6EekcNg/Hz/n7yaChDdTeSHignN5YsKicFMd
zpTpwJBxvvjZyI38sK2az2+n6AtADxP+zqn8odL2BkKU3HtOFNz/txlmw8HPdvEWB2Q0LeeWbNRy
Ci1gBrvXNgLdpVinOheS5pbr7+0JD6nHQ5q8w8u1XFWbl/V9H/0jTgav3sb4oxpAVkG9a1COVmxg
PXHHs/RHjDTAs/9hss73oH0T5le0/IFWBRXrN/PcxCp7WtYdLsuMTLVhytf0qDRVpCGwDh4s13sX
zQjVuIBuh9oI9DLOv4rjTjFswMmBlq5EJe7yHvL60Oo5wUwe7fZPuepFHipohQuFEYGjhNwBZTMh
Drz+A7B1DgXN1KXMMfylbkP2BWcP7liaaSOiSS7vTeGSb9JUR41KLZwPzayTwGvhnNC5w7phLtnX
HUDLcjorykGvkY4ddcjG4IPFnG2wH7cmSSXbwHsObovj811wROQvlw5r1BRQ5+0ONszSNfROTJB0
eQSrkDH7BIL0QNLUGVsUengyg+BhqwpBVIfCi0Y4PGHoaYWi6d0hOHfxWg3Gfsod7PvP4n+HskmP
G/6moPuMx4HNm2lLydmQiwQ1PxMdwS6Niaffl1Z+39qeoxLKb7QFBX9gwyo1fSM+lT9UT2LBezwJ
SMtpcMCWqlGq4zgv8Xz1jxWT6KRWSRaI7kmDEO9ovlY8DZU3/Zo1kChWGfLxC+NDeWxr7t6rA3MB
Am6Bq4UP4XYHN7g4juHA+0+sS32zKPcQdDweFrCOVUjjiYx5d+qbis+JgrsaXETVOHzgs87ccCG7
MyozVhfmw07LN9fKBFu/Z3/0El213s4L3U4t81usWsPVg5k75kuFv5NIKKtukhqBuHzot7BDMJkp
htRPsM1GfzjvhH1yiZvoSCpHShHVOZ8HvL+P/Rgcd7dsOuYTHZdBqCKcH4MIcijKzISkSPxmiOsd
FwNYFQF+RHgaMo4yD0YB1eZ+1GrVV8kkf5WSk7ssFA2V7liCPL31w1qC6odPa0/lUbLHwrSIbZDn
6/EZcO0lRgVX7NxKNMgZCmVvF02y36D1ElYc8d8gGQJQd/Sk5rXX+5f/xuyO4AdcffUYi7uGtyUF
QgHlCIT2x+ZOqBEZGCACrGPtFe02H7XDQAOc52LJEZKZxsw1GVxcM+lidI9ILrDNik2izLwx5Il7
FxJwpywPXogwKVFwn1tBoi9hSDPs+5F41Ux5OXnbbpkv95kcnrLxdx2YPTwlGwNgokI4BquesVuN
nV6UoCO7FMp9CEMxL2xwHdFbpG16fzQPn4wzM22m4aG+mWn/ELzgpCBIj9kSR3UgKWzWDkn5v7VB
vNPi8iOeeClCjCVObK5zyTIK5I3XTeCGZ55pnU2zG/Hd6Gd82a8offSYPbfpjQwKZRoVOv7CII27
ZipDAwLndxKeNkoEG/e9BxT6jLEYGmUrYS+B61xTy+NnLzDGTLPjnxCoyUFD7a+2uhQ46wuUO1wJ
JE2rsvDZaJrZ5BfznJOORzUj08s06D9Y5516s3tORXkkpJySic6/2Ijmhq23lk7tFNoJnMTzi6x0
kBGqnVdC/G++YhvgywP4ckAm8ynUFc/tcR1HZq2ztj1RAa1NkIgsrVh1NjYltOv8bMy07CIzqNvv
ME6PVkNGUQObubkORRagzEHVx67gsbdpIf+ifvFCSsoVu7g038iWbnXPZ+FqPrF4tAf/+Xl3Vm/F
nXUOiz2Mxg5yYAC7KTo69h/gi+Nd2SUlhHtpJdq7ZdXA4xu2UHbc/M+xCLVHvAEsgcGlKTHI1ZFa
Agm2iuTjAfkPGPgvd98Q075CoW5G5lJRyq/nCvy9VXAhtSr/NYokUYh+gwMW8xDhKoefMfLQ7+WI
v4anipRmanILkQreOt3IPDA+XcHbOloGLo88UqumXs4n8mYWVI/98gXV6knOwJRc8WpmQktsEWxG
IUkgE4HyBRouX3wCXkU1eMz4EwkY6Oson7Sp95A9MM0vTpjGv4FE1bUx9pKcL0GlAFTA7f7FNTIj
wj21UHBpvg1HlaJ6IGdcIRNP5ToiJyiILzzSrCL/5tvh5yu/aEldXvQt7JmyxrP5A5EhCKuw/MYs
wI8+/DplH4wNcFNKHlJsMHuGkjX9S/bBGOBRWKgtb2bUllF7Epva0Z0A3otqfWgh7lgfPP8YLFRz
0TfPRGruY+En0RBCMaQxDwhY6PiGk4GwNxypalnF9MrjqtT2BwfXyaX4xpIiwVVDd/qt9rpjX+oI
5NzkGvN1MZT3eYuO6Mepf1jE2FaVNfDta9ED/uiH9UEARSybnbgFiM6uhGBte/1hG4euwCTlTJQl
oQZB2+EF+Y/Tv0GEe4mkelAXD8TTsVU7RBykGP5xCd5AzMehkjZvEryCcSUFJH19wq1mMydSzVvM
ZVP7zVmIBgInzTjKeXGCPxEb4NaPCmiKnhavv0IrDX4Xbz0r1pXlMEOpP8TLa9geWlUUPREsm4iD
K5GjW24dN1X2pl8cl7DSNKBJA1P/42Z9nAimdD2O1ybR8CEuJccKfb2+yp1KiCmRHBXVPrKVIZVg
0pT4Hj2B7agxAH382ONEY9Veh6b2g6JOf98IZdnvojcAW6pQKbuZEmHaS+dQj8k2ImJ70EyGnrIV
et5IEQBJ4WJsGaYHo+GzEkx+lpYsE9gQoQVfY7OmSfYxlHtSu6Y1RoD+PubYpw0qNiLrVXWid2t8
O6u+EAHvOt1qVNaqXj69Tt0VHbIHumlePU9iAwCPWCSl9iU5odzHOjQ946gHdxSuTEH6eYSDotJn
kkqSrgtmW36l1NJzBlRMLzdLngZ/bcMbaaZlKjYVS2JuyHzbGXSUCYoRjX585BJk5y+ljXytS/vg
lsRZwN+Wzou2S75FQ1NMvfjyGOu8WmT5ZBVC3+ZDilLPoTpWMavqCrcgQBCNV78bWvzw4Txj8wBG
tfs88JrHHeZ5OFtR4q/mtFQbFmbcsKy5XrZJBMI2paz3rASgOLUN6S6DpqV6St9gBmOj6VmjD7NU
Bs75tH2P0v/3d3iH5UBftZfY5q3JH5nOCdnXAke/W59KAjL1i5c5VqA87PE6U5Pr8EpcEQwUHU/q
zAt3OSdXTK9G0i5Ahu4fZOdGO6Tttllzk6SbB1SvXnmeSi2bUACOm2ShWDJi1E4xTNBc1jsmN+4x
dR4xo736ymShyfqSpgGQKppxFmgD1Wc9u38aFzm95G6Qa3IM283IeJMGUH7rEeVczJnWsWkNTzgV
fsAOgjuekXCVugQ1/W9y+Nt6Nym1cwmP5hZdKMJvgGBQUiqjc6How5g6zc+7BUbnyjrY68s9PzOi
AW1rnoKTLY6w8UvCFrsgidDnStpV8yEDPtI65EFwYLcJDiwq8+5xouJadTRjACzkpAlILSL+3psh
GNvZC9RNfO6B9DqbFUy6viXX/96IM35jFTTiaT2dXPpChxndi319qvcBEflFjxZgUXzb5SDqO+AA
TrJkZLWmRHupw44YcxB9/gPbaHO4FcSH7r4fZSvgLUe8CHooGgVCGM/TvGyEL9nXcq3Xn3xtfNBp
t7flp0gHy6F/ay3nE380YPgv08z0WiCgf+QOuW1yXnduZFOuYs99S0sd2Xtokb56kvpe2QB467DG
M+vNsh06jVOhYWxfaMZdPA/Qyu7CqhaQTkQ6OCrcKftpHo7sPku9czNLkY1AHnRD+ZtNDv8eivCr
FqiYRSIRe0bQc7AypNxYiH0wuVcnWHpnwm/bfeYNcwtw/NAHFWEr0CRuc8+ugyVyi78XURGEQnFr
x/LGYBBBmxVo8ncFbUsqoh7/FQoLps0Kfu8uuF+l34NvXlw6PBdrW66MCZUGoE2JXJ/V9wq5HqTh
y3drsdIFwIhLekJPx2FbpS/ZsvYnBQXEtIBcG1hi8mP9AQd38S+fRiVgBArq1JgEuz3T7ONtdAKV
QloEL1S/CwZpcVm3T2L6bxyYdgztJ1C2fuXQukuXiN+kmEkPn+H7rwvNTnkq6I8N6tzpqd8OyNWS
7aSulGWp2XDzpWJbdhkmqDlQSM8mOKI++AdNT3RjvHod3XOfS60yR/zxwU4ONMKVoSHGauyAbofq
OzGrGFimhkpsDNzvaTyf3qvUa7oOyAlXilVAJSBF2D3yB/IHWDWJPXm3EKygqysQQk1omDdQg40I
vy/Hg0lB+uYR+oP6n4Qxr33STAnOMcsEDnbYQ8KE1o66W9a5axfhYc1qcinnQ8kHtvHc0APPat5o
ms3HwZl1AeL1zeVgANTk6DBxVMdU65ctnGXey59+YfkCFpYZZxVkv1pTyE3hRXnP8H2CvV2Ww55U
F3EtI41WhxN4pZ6894p6ZNsYi5StYXcItQIqy7QxpgHMX6fMyphU/VMHKAaJ3CKpY39oCYyQhKGn
wZIQ+lhGXnpY5KnUCQovqAoNs66oWpQDYJ0auyAIJOT0Rq+Vv9VVMsgJghPmRgdg8nqKUl6X/6VF
p+F1Avj1TOWzle78x3FxvSzkt0Bk2Rukek/PG4CZ7u7a1sLyHEaDKv0NqvebaFxbgvay5V6lU4vz
afZ4NhiahhcdPLwQrlPhNxsH3LlLDLJyd7637D+b4sOo6jAws4VfjO0gLDZiE9PQ4nRUWs2WuwqA
K9+4kvuGfYPCVD7nzv2xdFXT36t6PUM9pSStWVHok/YpbbVAWnGJdiNeDnfKajvQaL4wb+k6uxhd
GtkCCGqDw/KvolsMZ69g9aQgnu/EJ7ngzEtVByn/q40EJUB/Nm6e2CTQFNfg0sBUMUkqX4WvBDZk
49RBZMJgAgoMWOzn0/ec32qqUXPzbguMZDB6FOruhrDq9Rvu+cUFeQYuc7Jon1wqYcT6RcgmofEB
utF79Wg0Xn0WJ1L1URo3f0+PsIW09ZPz658yT4KpEGjFOLo15UTx2cmivPKE+OoscnaJQMeCbY3d
gItvN0xQO1gMQTZ/uNMHCoz+hOOSR4OZpjppz5yl45+Bj+BjVAjhKnt3utP4qts0SsCi0aoMtzVw
XcBvUH5XAE5bZNokWlqty6r1bkHDDspSLfuhZUyPsPIw8ybF9Tu5YA94UQUnYJTsQcKGRsO6si+U
AFo0cxEW8twLeuHPnBzC4s70y3mcVfZ/AudlFrYdhSiNJ8F5HkUJZKrsJ846xTbe+0pzmxFLCxGN
h7YDgmRH1EK2xtPHmRjpsWB5w6g+F2D/gYOkVnPYNB18F1TLmmHNQTogO/3d95tRXad3T+Q4TYfd
u7/54jo3kUnjj7VxGqlaxrgKU5T6kPUIsyUkY6yTFmv5iDB40s7McsulwBwLIXVujMje/I+0CkTs
6vQHdjdnahATwBpeDH6KC021BcKL30ka4D+1CI7zyk2xgyOZCohUBjl5np9hJX7+kHe29w1Phlkb
y5k3cRxuxyORiX9h3z1HSQHRYnygqwIwEQGWE6w8npv64ZEEGsZIS1yFD1vcbwo99nab4oLQ5cVR
UVoZbPImEkAaCaxm5ANEcbrresMVLiAMRhD01ikwdf6J2xuy4QBxUn3zMOV0yNDqmjum8n+0NMwR
RlToGNrVj9NKY9dj8+ht4VC+JNreL4JYh+nd/FgZ/8Kch0dSG7FCdqQgxMUv705WfbwVBF3dTTkZ
1qst8QDBDJu6A4kkcqe2Jg6OONbSN8HkY434ELpYcaWX7d/GG1I7CaQb+Q2/eI/CuxkhIuECMAXu
axBO8MMCcj4k7cbMkGjNuI5Cf9uF/AIdHmF68TpjmdsdMlBIiuLxWQsgs8rPZNbWWPL+T1VEktC9
Y7GTtg/R+WA8viFQawt5poDLsdvi3JCXGMMNlsGkOq//DcK3GFA+a4QH3vlBHEQNbkpKF9ThlAdo
u+QLcEulP/AjFSa+5M5jmeaFYppT+fkZhkFVjXEN7L0xPUFBATvDqHtCepHThIc77cnfrglJBVHM
cY0vPTMltSMNh/5bux8iATLzNceCf95ICMLtHoPndE+Ca5kxkghJwY07ndDaQldH5YPt1RD+Z/Eh
7tUV6wBM7ydrbr4FshtNXaqR5q1hU7/acRLiXyhrbwV9g5todcJEmyBbnzRBnzb7a8oRZOuQKf/j
28KgfAHvp7RIYidi1+bAn31YpUBrAA36puZksGcGVcpRuH5xoXChLyOBySbl4gcyGEhzaY1B1LRj
kkmG7lCkXHxYr9MbbAc+rsd40SW/PTfQRkwj+Y9Ko8Lkop4AynIL2m1PUp71ZiguNVhNmtd+NEcA
nR/2f8Ng0BsdMDG4ySlynrjATYYU72xR8qZV3OliXV1mAKf7Jw5lCPACigDv55EgSizP4BGtvZc1
alVAwZYVxck+Z7JAUdsdtC001e7scEYznmdapqrDxjrikQBoX8a4bzHCCt5ifs/RfpX0sq/gvgz8
kYB9UFxhhKFRrndOX/9Nf6QRFkijKn4KSV7x+RC9mvIUTwSpicS8Og4SDPO2y/n7DDznQFDZLlHt
/pF7XP2tjAs4JWm1qC+fKpd5AO2OQ6RvW2aL/lqhUbFhZSJ7FRB+TFFZ0HWWq/ovMlxq6JGntMUy
VCE3crA80EMI6b3oX92rzPhHKAkpN3vzWIswcI989HTQqBIZh+0lvNAge7Kp+5LzYurue5HLZLlP
n9l80t9i8JOphJUTwsGNc1WoSlLXiy1AvHPoFBxP4oMQxIk6mYxhWCaO09aYXLtGO5vOTzGTR5wX
+BKs/zBVZv/CRP+7qUHT1upBGMrfatW89CE8fxxIxHVrfrjkxD9TqebnOOYjUEEvVWHiujgy3tZN
z6hINANHJ2hPNTpEfQo/tApRTVl/knYyL9Mfsca0N72WvgwoCBrztF+qQirVm8w0AYFGAmVwaBd+
XE1HogoVHl+f+YjWL12dmwpz0ABlrI0f9a6LKE8dioxce3aq6BRrgzD3a0DASjAWh6mhrLeB9BLz
yvSrGhiEC2wqAUATRsHA14pb7HcrNEtE7waPBpIirVwFUFsvm9jAThk4TmCRSEgIyNOrSLHytlJA
uSkcryuMN5mHLuwKEs8CEF57uCcBdxgiIc+HrhuYVydt4ZmWmcACXgHvVmpJ9YUHf5nDIWJLmu6y
/dkCawfjPEx+eZw7VK+Os/+r382OI9aG2rWaRl4cfA1KsPq3FC5RjQNYGJeDLBd6diOcID2kC0Cb
FNy8k4qU5pnbfJjOV/4R1aQ6KGGDr7y8BFtu10f/DtYnLjDN2zmgw5TLXFxyprzwh9hvshiah4vz
Blv0eerLYa+8JjWegIGHNkF7iHC4V+rZyKkMnFEzNoO1XxukiuHzN6JlF9RqaaZFyXGWVxx/rIKK
Z7Tz7H74pjSgE8Zor9VKqfDziIV9jFj2Ab42agAbcCZYF4/lc+BtEeej+v+QFY8KTTGq+o+uKau/
6qOfKfEH1YbddExWzrBTMALq+fTX8tMEJ2pKfLtHXytRMiu+tgElnQnHoiZFDpFYrDBSo/HCH2C6
esmc0zhF9/vqVulC8YzD+TgmrHmDkiu5XaRkvwrwYK3AeQCmBZqlqFvHWAwTJ/9Qnf7Sxdix4ekR
ak5DkiFXK2CHN+++bVrllLbR5nFW8OOuppgT5OO+BZJYRnJVIOxNXxcULtyqfONSi2DCavN4TOAj
Cu5jxbAILMXF6/A3p2Fs2piCsLx0xCcUDrbBgAh1o4BkePgoH7pclfZ8/M20tiUooZvv10W7GqpO
SWjLKjjZEcSYOIiIwZif52whiFl5a3g0YG4ULakOScRFFQNAWSRZUZDZdpbxaWtkeHV3Ffx5GRwz
OmPY8dRnFpJq6vzI/a9zyjen+SqyQ0DJcljOMox7aB3w3o2pGbm1lhwBl7QSxRW/x9sJS9DoIRxO
zy7zAr2ZxZU/kKYycMEYFDM1YQ12oFlPqeSahQiPcAc3DVIhiiCA2ETviK2iOyAK/UznWMbz8+zT
7teAP4rl2uAtt3NzQO0d/Bw+iOr49xwz8Oj4LbSF9jY0vjKWWXPyQSsylCgbfgxFp6iUf3J6bUwM
X9/BvUNztVoA/0DzXilnw8dXvv1Nkfsx5IDVy59MxVfAOAwXy6aG0xwV7cAHqu0vN1wgnP8tovNr
G+vlEvPIHHFYz7gTuQfsejk3mB0UosDdiGuyV727W3yq3T+FMNGhnsHniNuPidyvxliE7QH3sQRl
nID1QkPT65hk/NnaRQE0ghJZuj4d/LwOlnJmIFYB1PaEkrjeM0eiTiO1X+JcrkBZX4w2uIMhodYC
yKETFNmq1gDiznHVe0tmLn/ndyUymBo5Ft6tNm4pIoqV8Pd/hLMEDoeb+R/evVix/xlrxGOdCxo+
GeyzqivwlpFr7Li+00J6tXkIg1jY8ZqhJHXXgCRsv+3NnhUTXWYAIAl8MRRsgZdqh50yEj1TyS1W
JyUZJf6fpu1etKIZn1Xjd1BdWDpwooQG12lrSzCJ32Soprp0/DjyVDw7VxpStYIAVpF0gcMcDv3Z
/terl9XGJuRXHjNic9a2Cpw8pHjIl/DIJXkdKXj4+xF+NlSNZw9I6o4YvI+4kQSbgyn2gqQEEYPa
oJrOnoNS2QjBtWCorkEv4zJENgDQclm5koS5SecywnP9tDKtO3a9OhMzjP3DI4wFM2BIejKEUbAd
OCBiIqzAN8P2VhstLKoM7DpgUYWArkINlww/tXXwWS520uoWLzni8q5hEF6JI+TKvM3D0pgUM01u
s3Urjm52xbG04Wq71Z9cSR0v4/4Gv+wIGr9M5Y2EHwnRVVkI1ElflQm0a1xBo75t/HaHF9ZzwcCA
t1hi4y91EwBfUAWjFQqoLiJNQE8fNAHuxkZecH3j7QWftUVBEpg7cKl9IhvaE0UTI151ASOgeW7z
/53b9Xdw4chaGOLElpZf6hq6684zbKhQhnB+x2dSV4YS6w+JSgv0GIfglwo168K+9C4iIQxJi2ZR
T7Nu9fm6BGJTCn51X0baLhlQLC0/4xSgCx7EAZAZaJ9mJNbKN3kCWNKBk+D2dM3y/cWoonQbfpUg
INGvPQQb5k7FohjQj3KenS/HELTiTKuu/LqgO1ckHlbpKzBLu4z9OpfkorSplOSFsMpL4ypSpE5z
uyAhB663dGFymEhjuioNE3AddFqLOatNW2RhLpb2+TN0n4kZsIlE0pHPghIr+kNS4fSRM4Eb+lE4
v+DO87GSbALHQpg9a7iLOvcR7bFz6WT/isrq0P6r45t4+kYoCjuYQP3rolYLzl2J6t7h5j4uxJsV
zn4eE35L0UXwznbJpXqGDToKD8CjBFf0M84b6ltczLt9ltFaRM+UR275PAGVztPzndIz5pRkaw+l
ealJyOxsbGRJUDgebbbBiT0cPT+fjQz0Okl3gMoheWg8kh6TXubkOduJ2Lg0Meq4zbbYzcyPudIM
cHCC/Rcfm4v8P211UJtD5jnyqchxhr5lCbmoU9HgCrN0pXdSZhv5uikKL6Yp7GGS2KJGp6zFY9Z4
jXMysqDq2oBYmubJgFfHGA8ktjaqghDrhdwahmMGTI9St4W+q/X3ebPiag+SweThek4mKH/4Ulcp
U0GCBzrA1WQThidPVhQxVdgPYnzjKjbDKijn6Zxa7SovnaTN3rgDLLjk2OKZ1VEd137c9RSUofhe
JZiEFtYg9kaXXHm+wIbTsZlc4/PymdlD93dETthWkoCMy+QS2GsUJRG9cIjatBJFKbXgeFV1rsDh
92826cfCKRCz7JWC5Kk2slDADWdyTLmxeU7DVvEfWT3+NsylTTC1qe0l832GUOtpjalZjFwCzXGf
rwZIj4VdF6R6JSY+fH8E203snhEGIOXmZWnBkYJdf7p/1HLje0bsu8tre1Rf0yw/WsAeRdfVL4eZ
mpDVD/oIbI7vAh1IcPba5Bs660xFuf3hOdGsKwdyW6BW6latbyjKSQDYUYG0HpaUbr8VG4qJM0v4
FdRi3ZzQpBI39KZ1nxl4annUnYkcEiMyrebI60dgPNnflh/PNeGbLGGu7IDjVzXmLqgxFM8tpRVC
xJz1FIX1CNURHF4NJa9NDCn8MjiHjLpjrdn6EfjbStqip7ayyBRplHwTnpkxovPhwjdSN4jxZiAS
byv/IRDh8YAdlDbDCB5GeSgrMxnr2jNB15ByzGcDsfHzC0azUfO2gDoigx2BBu/cOzCFTypvyXTr
mLJlZCuqdvc16VITX8lF3aU1dHY7pa1p5DV36Edg7ZTeRDE4iV5P+gMxgeRtJNBJIv0/xI0Jb07P
6LQhLA/004uiQEGcLt629Up9l94OfEiTA8yk9I8pukygkHyAkqNmxmttGSXYiyJXWu+5VPMPruVg
17JXGkgfdr28okPhCMVAV6Nzsrs8hb2Isj5e/ehadjxzCmcjosJJfOukk80FT5OItXSxtVXBm134
Elgffmk+jyCD3jhq3aDWP6r+1NJLqRP93aWMzAf1VMF8fizh4E4fxjdQQcNXCGzIBA5oxdgXJwit
vdaIm+mmiJe/7FRpwtpDgk220VW/isk7DtGdTUhVnyXC4FHjL9cIbf0ct+x8DH9VUambPvC3yZjQ
SXYinPJbiN4+W6XioFaVz4ys6/WZ/US6z4XbeqdC5+jU/rwcSLkYwq3zN9zceDpcQcfaZzptfOo9
kau7phCs1a9McGWnj6d93Hi7U32dwxNbDKWAnNnHuArRcYaKi+hQgp8NgRG2p5PniVP3TBnL0HPl
Y4wbrwsH4+z101BAIaZqzZtpe9dXvOX43UnCpAp2fmiDtIlPpNUAkbHgXkjGV/qD9PWjtOWQfivF
mmjEYMgimRCzo9TzYxaQKKqwmsyWUrTFf0QHggY39HeVk6E+RbPgkOb+L2mdEh/hob7bPqFo4TZO
7ZoIXd28e61rn4Tl5UQVzZ9S3iraeYGYOCQ4UomVRxYMCU/OisGKzJkZPmo1yMPMiJAgDKSwSgWT
jh9PUnLo4eOdgcBVpI8wpHrwJP+zmM9DAwvS9Q/RHyfNsTaTPCvwFPG9RYwJ4SWSo98hH+LQO5Hc
9Kb4iZxQbdit4tWOqWUDeqnM45XMGGRWwZJHZFboLJnO8qI74o4qYUKE0eJgslTF8bxKMrS7LOgM
WScenh/G8kRnPoTgZwpAW6fin53nNMfmI3Xo0NJsWgGv2odQMG43qqi7I1n/xLCCrP0ckAUjg2Fc
QUsM3bUmWtQfn4u9/G/bfErZUFamvuDU7QzUopF8ORo/QBDKc0zrS63jLtMyEjXtWM6g9pMlLuxb
sRz/Ex7VjAysIT7azgU19xIwFfuieeSGyUSWhK6/bO2pWZVTAM6xXsNEb0RdE/Vu6TV1AdIuTjm/
hDfLLn2r0LnnFOTcMbE6iih13yYG0Y8ccjqwexvwIyGXNuD9TtlK/oNY9EmQ6le3XnVEX1OEVTA8
xCppt8Be3kvK/LXNGpd40gS0CMsI+3tBDnNCWS9IGj+lPv+L582KB7HuU+2aPjYQheXPUoZ9VWci
1v/cnnr354yAhD36qlFG9blypksYhok5UR7Ae+QaFbOxZxPbQAxjxbSorMSCaMLywjHLCxGFVKwT
vs4TlcaLDflbnAPEsX1zu5kVNRJA0OTCmikAtaMYNLHtjZxMR2fvEMJfk5i0RJzMW3YYbmhiB3kB
MFYgZsc48QPXrG5jF8BU84kT9Up/ajjelKarNW830vAGSg5m6ywLKGOUBJ2+AXwz657tg96D/GWm
XSLfdSHIYPp63T1qCzP88JujqV6gHaxVK6WHMrWS4ocp5VFJXD3jORy6o/PeGuA4nE3mEAA+etWo
8ZnOuCWocEP9nXN/YvoAau8jal/7wQb7oekwSCcBjMLB2Zk7nYgGia0vcBQsIcnjcYCjT/ahtKuq
3eEfS1Jy9FYmngl9Ps3jxAjf+JzZ0Q21SIGKzZP5R8gNogPKdWupeSGBllK3+v0/VpMZFbFoX3js
V0HTbjDdFrL7Xa5kAdE9Rh5TNYQ+kjT2f+rOV2FcDmsmfXGJgw08c7Qcd0RA+cGV8XaKV/j+dm2c
AFp/hRYwekoBWOzEl17AcMz6nfnyUJZRhRPerY69UgWSjvGOLGiyZGxYvDBuzesVYEAvUnPnE+NK
w7esdms2r3B3wVzMWUHLpnJeCePijrQFVvdPwzknlSEsVCRich5UztLBZwRZDgBN1NmBp2bdIoK+
mxztjEuNgJsRutS81K+aHJcNZY2ACjF+bYc5IhoCekRwdCY4SQXLgI0ogNdn+IYJ75aC3UK/yTQA
MyRC0GyBjLzGn5i5RBzHqp2MWQ1KQY64tm4GUIXmEMoTH6WTodNwAmOFaMjiHreLyoGbau2nb1xA
baLUwOOu5eLzXV7tCycke8eVG6RFJlyt3YBxbdh3cJsZG7EZzdpjRJbj9C+F02UKk15Bq7rxKB9j
L3doYZZZ/2VEFk4PnFlV86l7ndFXBKQ8g3a47tDqNCygrHHBA2suTAC6T26Yow5ItKgdtyPNz954
uHwd3c5WrWD8tv2/3SnWl1RJAU9NVmcAVdVUSmNC/wC/uL6K16fCbZ/OUFrdpHvEnPMhLfT4c9Sx
wviuPg8HeRIMXJLupUWQBTXA99xWaYjDXwmg6LZlL4Eqo/7EZRLsj8wBqS2iaNCiAjH4sNUzP1Ex
0UfkQSHve7xZy7MT4P69kE8SUL3ydFumx94tF7gOwFDavqhp/5VJbothGAEbtdJAMZACMB/ZxAPg
xvCkYye8f8/zJ8rC57XiXOmyY8Ru1fWwwjbAciNxK8xyNc1NT6CL1z6rCT/OvvQG31s87xWRJqRC
4ib/7sxXOYmiPxtFKa+UUMUp/hyfD7VWdZK+OK2dRmiSjiSeYc2N7qLzW8bKB96qhiPFeaJQdK/c
5OVB2vq4wbyUZKppTRg9gq19tIb1gf+FD8axkUwt1K5N98o+1cDxAQTiihZ16cHoDvYif5ApY3vk
W3Tv0tpWm4PbgSSUT4MxEBFKfd5LSKP56CKY2Z8wmNi6IhEWtf+yIH4eaGKIvuHFGs4TjbiNklEA
RWAlIAcdoTahPG7bQJkkf8YUOeorAZdL3WhaFwOtgAvfP9RDhF3MOkJ3J1UuiBBvz3AqA7xva9jm
kZf2Y0ksltv8UGGWat9vU24MdF7A3lPMky1KGq1Hd4/oYkJtAtvKNojT4qKNKfDvrflzFpGqn7Ip
3UCjoLtXJdMQ3Svr8ucSpA3zTPEOl6s3K7BS62d8Z9WfrAWqhrknYvCViLCyzbaeDaFHqAD2dAQP
dcVe3/fndvz1DW5Rch7/vo56ntP1nQrDO4vlwKim8NhnZA5SEXQTbKNK7BGGkZ75fiOJLHciK276
G2pDCxVU+YhQftqCct0RDCBnbKzCz260sXVrqAFxczCg8tkbw58CgdT75jlEsrI3BsbuE9Ke5Cuc
G0DmRWji9qhrE7BicEuLBq149rXg53LYfC5Hz5Fd+M9Xv066xTrqXsSudlCQgB7EuMjybYlYO7uA
hwVqT8ztBj0AdAPYxRw6IrtLpkYrG8p2DWY6CVdfrky+Ibz8TqvPhAR3Zt+VPrkYx9vD6OAglB6a
KpeznE1XQg1w4e9bYRXorjdWhP/QoFFFAxazCNm0PoX+CbRrlKvOomdcebXXdOyulHp4FWdz8s0r
IU3G7w5nceFb1ANlwcrWqpq9jMWhrpYA+KKf6QwcVzPhptqJ1k0cQv8twh2B5JiqXO4kVZHdo0BI
MU9LJ1aABoLtYStWlE8PwyDrNszhrk4A2eArhIxSXq4Yb8PaWa3uHBiWHImhNyKRJNzJ8RLP6uN5
J6S4uNBpj4aMplm7M7CeD87hYcwNQwYDWDC2RVuKPGxhRzwGe5KrzjIuVfH4o8FdA9OxamFhEmT5
Nh45ojpQQAtaIxacxKfFkl5xVxOgs8vKQhSFGhVOsatc9AUFF/3Dgklc9gaWs/LOt/a+WfJL7wm+
OqhXCXhc51tHkdocxhesCdCZqkaan7rJIK1wtwUGjJKHzBi/M145Dj3vexb7+mdB8awVq/C0MvVV
yxt2OJCP3+NMFmrwGz/E8EQHK9i3zDZ5rBQdPrWt1JqUkq0GD5oPKjpVHlTJtzssHHPgrEXF3VQ8
aTraEL5PXgZ1+flCWlJtO+9TIlzAdQpZWLEIBMIUE26Rkzr+/FtQWkY/H6sE7J29VxuPNynFKR3x
Rzggsh0uK5rBHv6f0nMoKY6GYkBJ00iW5IPUEo+sUJPXgCOgUzgrUOBPCnAXIDGsL7/q1Oi0ckgy
js7MA13pOwg0y8TFynyz9HRRiFhToPWhGTSiY71sfWcWTMIOSVIjDuU7l8c7PxH+rLSd/bT3uGz4
KEAJgw5FzIv+IxEDepKzMAz08pPSjPUEO2xQ3uYfF68qUZj3dbRSkCuU1JU0IBp+fdDCkEk/ocik
BG6s2piRmaPavL9G+Xe1tcoHw1cwKxX6VcTfXvQ9XbvQRjYXuqZAGRLd2PyRbf9SulM926AguNuq
/rwRueOrK2GIMZ4ZpTrxNytCL806AOLi5ozKcXAhhyXHKiU0pOTsFxZbTcFeHlnkgerpTW6lxFPn
RYGlOVb/rMVFH6AZ2W+X5DBewlS4krt57mm0pq4R476bsgJ3P8gTFGaLj+kmabjsQ26Gmq+cDR7J
qjCbQQE6muh5UJdy1iKSFxWHCY5kRZNCjvpW6Amo5rM9mc8DFU1mjWUcgmk0ySUUfBipElrbOJvV
plyUiXYuKoeSZcOLVGdrasfOfgARP7w8D4PwjOsAIl3GK/HYLRMF+2qh2cmUS30ePkva6uiQ6pXc
C6HiAugOMLez7iL0aHyKXOv8rsXqB6VOmrvPp9aGBOAtbkVAt6RuAUh8LDRzweIQMiNfOuVckAga
IbhXzRidsyiQRs0wuFUH+3kfku6z0D6RVS9SYbo7elrHWS8jPx4Eg8fOB3khItk9JKz1accZnYzi
8KBWYEVshU6EIUvhep2d4O19Tuir7zvN3QmWnRJQuKN3MznQtjKxTj/TE7fsshg05VsrljBtxyrh
u3oe7RomQm39XM5cdQ2p3LMKtKsdwK78Ds4BBioikrXEfEmHaTV1+szjr0H5rR5TfN9RQ1dZEuyM
4D5l/hFVVUrEUaXccPZ/l8itiEUOQWWRsvug1XK7E0hePGVj2B74kIUq0+8W/fYxpIKqVDlbnFDA
cBLAEynCFDa12/BMQkLrYFcwYml9M2Z/YuJwGONxr7tZOOGDXKD6UJWMoaROoxbEzFVGXJ9qP9QE
ZSKSnu3R3mzomNk1RPijjZD/u2t2opf7PFN0S+7Xg6U7MtG8UHDp/DnQInHMVB0AJICpMUvsjEde
DgPf3/V+tZiliY6uH2ROxdiazK+BjM+PK0gWaP05fs609NBJwYy4FaCnTIXbQaY/fqOjVOkKkj8P
ZucMS2bKa+coNuG3kpvbjodcnVpmoetG2mzZmfRpJ4r85kn/tkAUfYIbawsGRs0iu1weB7vrR2Sm
Dg2h1twIHdfpG9eRIO5KYtdqay+W/stlqMGeFgtyhSJ5K6vy+8rX+JjhWxSdr0NnBJHIlyui5a+L
xjys2xVPZS6Rp12mh/Y9myt1SjkJdAAyERFCl944XC/H6aA6oI8EuKU3rzn2W0zkLOJPPiYAws+X
5+Y7/0GwzgJ1SQ/InUDUFzGH3ywiKo3f2w4pjBzFGPqp6IL6VvfSP6cdY4bzRTPzaACqqxsjYRIQ
znSCtTn1sD6rRgjc0008bjBM+k1FMa1QofpyD4wZCagxQP0O6DHgwFfEoc4nKNslqmyyUcNZNKQv
FT8N+1d6BiiD4dQt2eG0txaV3ii2Vw5GwtMSjSUtP93PmmnCdIGHoaUv/a6sJG+2DuChua600+bK
VgYkFdLLau6NRL7ApYtD7tZkFncf8Oc4y5b+KDlCtn9w4wnEb3+CZBBDssQKXtqbjvFGUZTgwRGK
+gJTlQKnfEbcq/sTkOXSa0qsjxKgWJpgI/oIEF0HI9WT7Ed1i0EKHc3ogL3bxWt93y6CTuzQwwqG
b6WlRNz0tOUCjiwPI/pMuNk+hfioXxE6eNlI6GevfGq16UZOASmz30afEl506hmHI4qW5NPECPRO
2GglBzoHLErP3VmJpczECPYyCenPq9NbrzYciLhZp8TLWqS4pGj3zvqRAD9H09DTYaENXBwn4rCj
IoDhAQdgX18Tcoz0yL87UgHgrcPNiuJAs3m3W7WXM8tryLWNAMas22a9yvI6W3UTbKoUxx1hbARi
dByzF60pdwRimh8iO7FRutFD/BO5xo/+z9Ui57Y52jKgO91dkYhNHPrajq1py924OLyvOrKuo10N
IMj9J/lQdf4xXAwMRxYGzNeMliv29VduMQRWrB8dK/XLyrfxynkXITkJOKdwvO5aQLAaK+gFlfaq
qAkRgNGeVs8qAHdEhTIsKhgmSUgDNp9XCrNPOpImovSnAkt7oEUlSHGBmhMEDs9PVZMY9LHigmm6
qQC8PSH2ivMqGOapv9zBxHtcr7pFi+2hm9z4UwI8R97PNvhti4FYbzR+ZCL8lqX17kxr5clQYTMc
BJtPZ8BAw5e1XRYiYyj9yHEeXmCzT1jcst5oyultHKtjNlGVN0zgDOqWl9KYfCh4JltFvvznH1sL
94290QD6zsiBN3Pn+OfbF9eHCSWkgn30ZD3SGfIuhq1agRYBOt54gY+e+wRyW2/0NN8KOCxOIiJY
d2Enzlibqpn3SzeGAj2ge9Db6wK1kVcsazk3tF3jl2RIlY85C8KywotaGOu1JHWAtALfhN0CCdkO
BQYXaYTAem+p3RaQBp5u/bnCtZvq44OMpuHgfqggNivFX5Bs4my3UxYArHRe8hZdDdJI7wUYUEQN
YeeGhQm+s8LauUsGrlgLem/xoz8GKXuTXs84y4Xc7TxfmOCkDDyEf8qN8QcNNyoxCwpFWSZRemDw
/tqBK8zjNHrmoomAIsM0329ZCsNRz/03bKgSTgbHlecJtKPbrMp1OTbEyvEJU/1Dm3S/DNBNSkmU
GTXacaHTySd8p5UoM4eoMZyL8bV28owtzGydd6GGpRNoUy2yd9lYlT/XWKr8L5z9rCfP0OQlmF0M
8k9h+kwp2Led/lyk71mV7HFwF4udjlriaQpZHIHJkoetckFtHBPgOY1ZQWjwWY4j8xPKX1bqzrkc
sUOG1Rds4CDKkqd1Krp19EypP3E4hPGpaC2d/SGcqgHsi0UhykLeBl9mEcByVxFFfhEYMpKEwPAc
fD6o/oUgpUNNW5JgZu88Y4Q6w7dHcJTeDVpGHRYMrtGruqOdWha7Lu1zoJFxrdv9BddtV1dqTS25
jsFwWAgZMBbPUW56AhHukaTqDMNEJidRPvf7dPAEumqR2rmyOxH27TAys+uis1b6HS69dsWvJjkN
LqxSmIaVvn0zrjD3mVsG94UtizSHVDCbdsXTlhXelioOkTbE90q/mtWiQ/5Ea+KAE8F+OJx1G1OV
yoO/8VhKshuVY8XrbsInfS0QMZE8RwFJp8YKCHpH+YgQovz82aMw1qrp08U5MSPwBFaWVK64pD+0
WWc42NmBp7yJ50rEFHhSeT9K2EvDo2+I2iEi5YMdm9+1fUHfXmxZYrUZmTx0aJiRda2H8IPPjeNO
RcfdPuZPogghNl7HrpTOELo7vS4bm5H9It1pqumDD3IeyIIvFi8xv/u16qHAISHIlL3xZL7pZ9b5
+ubD7TEt1691LEiqznR8Vl0OlcexDVPp5b7zWBmn89j8DOqPOsf0fqrQ3fEXLOrE+2bIXO3NhgAN
sIbkbLeE3dCzILV0yB3+NF3DAkIaxLubFK6h9tbQQKC/0N3bAfdtH9ToLHFAshAeuWnBDPgFH0rD
DidyM83lfYuBs4IvUUwrcyEVJazsqb3wnTFRV94Q3yyQ6VdFWmvd3Wx+pLY2pd9RRWjhFD18mtZP
ZmJGVO95SI8TJZMmQDnmDBDeUpfqyMha8cJNXjraO6J10loIxc7mqslXdET5WAXCQ0WO/Q9/APk8
Oay8ik6BC/n/nkgMw7rmtWI5UBVr5QD8PAyYwSPpbBWMKs/jNLXXl88kg6gsP4KpcBdcOIRMljkE
b+7272HJ4ZbacM45ZgOcg8S7gqX5zEKxesorzuceJyDR1f4aZ5HFDf3hUGf2sYdw+dMDsLz0eSOv
4VKzV+6lSlGgplKh3AM6QIfwpjEejPzaiTnXLHOwcXo5RrQ/CSYFXLYGTz48BTddubTugXlmuZDg
CuHTtkKYilNiTBOYu678n099WS6Zi3m+pkcQhO0W3n/Duu/3fejr31p0+pcVIGOSto68cdmAwofJ
dYhCWwcwMzz802TJSnRV+UKPp7TGJ7fG/T9BGiSnYUovu7x+jyRD29WeDFrGT0BOthzKkBCe5GgR
oawW1EACuZL+KTIC8SDJ6F04XfHgoxPArz1yOI5NMcSB/NluWAd8137l5pSzuGUD4kwYhPPDgSrj
z79ox6M1n6AxUQPxUZVedl4GGVxNg5cobS4753SewNtp121gfgcSRUvBxyL2Opv5n23QjsUHhv03
B1A1uVBqkbZsTsrcTaKE7a4QCB4YiMzYf/ZjE/d9F5aGwPZKbNa4gp71O4WX04kF50mrD0G/xYGP
ZTIvCjFmJHnPvVKhxXdsU89NOnZ6tg8wQsaUN8FQloaCNtGp835MPpxwApt8mXcP1So86FaEDMkf
NFQ6YtWeTsAFsjq5cycKRZ9zHFUSB2SwRWNNpbj95n8ceZCk49q9mJTcQLYzU7b9SNNSFLYGLvJh
/OgD8IuWvCEmPPj/dbtWBEwloUOeFExd0LjDcZww9EJqtIMfTjCe++goy0kscKz9eGIVCJG49CZO
gcnHugqi2B9mcBLYOKVuv4tEwjYYmMrwOaAwfHRXJUugeKGgfPehxjA6urvksud8qqQbR+YLIr3+
z2vGPONL9b5RXWKInF8LQzxy5ZPBUl74BcmUi5Ia3SO7TjSFUxsUacr9wzuip4DYvk5LvuKT0jiM
8qG4x0Nj6S1wjzj7Ya2YFaYXmW+DfZoNDs56ZxHO4LTTdeOjS6XqTVDqHd0nFvEAmc49JSOMsyS5
kbBK5ETFkMG80TrnNcIbAHliVWtU3ZgLPwXVDbduW5OwnbgM+vK0J/hFssKvP4KtZw+KxoZMTKy6
3YoGOASCpEj4nhnW9g7kXw6Z+UqMhbgI0nvOKkf3YCEGVeAe5nFXGh2NoQ99+az+RMgQo2zg3x1D
Uw3D5f97ydNuT53R2zl8ChTPT7sba1H2NO9+JKMv0DoZ7hN0spypVMRzv9k2NSUA1RVxbAPmUR3U
UaJHxpUW41ZbkISk7GJaudsSCpIQhmHojqFoInlYEHFQjqKFTe0hHJvZXJpP0pk26fk6hu/B//2L
acqhlvxgRjSwnwc8lRkXnlta4CFmgZiZbo+Ss3JzHm5YYdfpCHdpL7EzZzKeou9+ro+ab0imEUXo
EGWrF1oN/+nH/GQWyOowaxLhuGCF+tuVoDt8nooWIf5QcJhfqnQz0GEGkjdscUt5+2U1NDy8/mzW
0uQuqUqd2KtiZdXySFRunmlwZVULuP8qLV4AiwNmpb4/Jq5oeF5zSsziVH6+MucHRfoUclzNI0jk
XsFBNuJ6t+YkNb4yJIyp390aP6Of61gr+lOZh9W8Mi+Ghp/LfaxTMLLYeQdbS3FV+JjP3UZkG93y
2oPHaAW4eMAEZtp7TSknVgGkOXnouCRcYPVQ3b+88EyEyC0sPE6A9amYt6YhI+2nD/lsLNn8kBUL
d5GOe0ocfMM3Bd50XMUTh3LT1dfb2d4ZnJVKO4w2xY2At3g5Wix9pUCzNKkvmzL2sCZw+1VC8NcJ
2G/ZzfkU6oyo3+RbkzNa2EfxPzlPquH8FpyNcIxC+j65qLIL/16oWv5M7zOQOP9CM1zg7aGLrTk8
3Htesw2HPsynNkkraOhBcJB+iNZXEPi9dpf0m8V6NiApc80swWgXw0p1gQKd784iNsfcu9ttUN5w
L9xsKvExoRaYSudalPyA95CFhDR96GpnJiGSt3YlK5C7d4hTDQE/+BGvrefV2O3CsVxYCz3X4WIF
9u69ieAz/Z9IccsBvgQYsJErEZLcEoI+2uuluwsXQ96y/5QnCeSnZ8ARe4Oca8OrZP7zWazPbysL
AP78sAXcGRiWWCKv0CvW6+0S4vcQoDG3OjzavSHhx/9Ux9PDbVFidW1MzyrDkrEYxPx3Zx+E0L47
6QVvsGYDtqcdboPaa9H0syEiyQxyhVy+hNqOsLxC+8XNZ4uMke86zhgSpf6yWYlhCTIc0xfbh3Wn
2L7cPGG4ZPXzYKcGV4kI1qYYlJuLkLYhwuxmytIClRXaNa8D1llaJPTqfl1zJIY28VL581mlG9ag
Y6ArF5QEYsfnQEvEEPf3YddeG8DFX1UABnky0o8v/IPv+sJKfW4ua6csC6UR3x8+3qbISkTa30eZ
NGEZjDZBH+P4kwugwyGK66h2mjDC/vS9YJIv14lBZvvhkmHAhoIWg6rlKCW3jp+X6RBJ0FvkdVTv
rYcKcGNnfO09OWGPtfrTJH0a263elmGZKnEVJRPdzOwjcV/er+mZpPeYRJrIXo1CTfl1HGaq1u4g
ZxhnnRvu9mm3gbraOX01KVPX5/pZP/tg4cl6zWO0BqSlrHlmbMNrwOnzzgvGQjSSdI1JJg+iSrv0
tIoP1wI8yWQxT4f4DjkgjTxadi1mDFK5PydiZRwhP0W0C8FhuwzV04sBaQzWm5txCZJ8RAc6krsk
oq6WAZ4givBC2TRssRpb6XBCdcRg2MaO0Onr01Hz3YN3D2Z2n6fVqBiwfrlJoT4qHjLVgg76Srnk
CKyMW7l08nnVsih3mvHQbBNcBx1+VeECxQPhOmaJohkWIy2oNNMCzOEi+nQsZRwpJlI/5tT2yE4S
5f+lil1A0i1lk31kM0OXV85un3GUkdpO637D/NB6AnKo4PwfbkmLn8CAP0iDD16fCFi/RWYX8kMC
fi1cTna80n1Df4MZ1Aq0VTIXGE3pkLv1dT1DIg8VnRHOHcSTvAlOAWMhJ0/aGYFn0FBrBXv8aWoc
aL/6vi2wF176z2ojbh8bFUNMj20i0IJJtukaS5SQzhDwr/3LcVB1MRYTxHilI0OmVnBBtuCyGHQH
3yAPpJ+t0/CcapluaKt/cgM7GjKfKLtZP/OR9mUbQh7bIVatvofhI4io0KhwAbBIfhYN438uRo7D
mIn7Gg1lDdbrpVEbRBif81ceXuby/z4DGdrCYyEUp3+Z+Htjb8DWsc3TMoLbJorYfpzqT0N8SKtI
6+HRmbGlyut9FMjQ/YZ33nuuNkuoCrD/h8ThSWEJadS6XxHwrfgwow1L0h4S7yhhztqdgkjCWp4V
nEXxh6DL1Tocp+W5YLsWC5ijkpBsAlesbDDz7qBnJtM6zSSqDRUVTfKXJrzXvp5pafyCScYJL05m
hdsWkhcdRqcJeGCoL4NwcPvTEOEkAUQxosEKFr/QWkcUol56Hrll+MLGb3xr8kE6urtkMPqB/br7
HjxA+DXsMSZNfMMxbMG0KMg5hp/APAvc/DLV1tMjS6l1LV3+6VMk56zuTwZO5yCzpQASvxRqdM0c
IMfbvkY4MF2AjffxfXT48LvBFmQcPSjpIrMrWBPXVwDaq1zzeL1XOy6O4caHCCSHPh0wB584/gwp
7cr9wZjl2Vt3GcVMqerarpPF6IcPF1+vqq17ZhNI04KQI92iE7dTuRvFVdoXGaEzNZ+pW286DpaY
YR0MURMNLLfSsvaSE/ctrDKwwlUcev329IUI5l5q+CdL3P+qKxyZtZ1ziOzae6zFlcFuCSJsJrIL
UkyiB2A8gBnn2s6fCZBBFbO6IJEiNIS1WEtGxk6FFc+AvOIjs36YNQMNAdWHNbsWNcAItYnsqedI
bE4AFmRin0zuocW3D/EDnPeJ4s2z/vObgL1IxNmdFXNh/jtcEbl2JH/pQQg0uIAzNtRBNVXyCcqr
FmbVr65x+sv7uQsIkmmv8wqjvJYif5aD6k4DSC1vfy/2BtDTLtWFLe5adzwDg4hESb51uQIpAxre
8IfkWYSLR1n3WcBtep23XP/qvDc38rm3LYYuvv5AK6ArXfIXj6bNBgbYhC/4BOXVuP89qLJ6EP/B
/H83Gltjys/RIQ0qK6mnOTQlg1xygCWL7F64sZFPcKsAlf6w27EPNChqLk3WeRe+aqTE7AFndOrZ
q78cUFa2yvORdj2Z3sXTH9Jxra+E9na0scHQez9rLE2sq+rf2+YoSUjMwXQRt8TOzc36XNHqR0Bw
AI1YqLQ+Ucy4rj5a8bU2oQMW9V/HsHqVQofxElB1odmG4sSDNs+uZx8/xzkTV8lNxRlhTB54Jf/U
mVKVO6farx1RcLphjor73NFpE2Tcnnsn9xXd6SxGl9QVJKhrx42l24QQ7XafHEG+sRNSUnK3x0H/
K69y9q/tK3Gb+m4lVYfe9vHQtUfAQaggNFSfnptr1VkT2sZK/iaRKK2PpkOzxfoIxSRLCKYZBTaI
uRtrIUSovF5KJLI7UVsQaOpY4KloHyGQmmOxxHiNPd3W/U8b2BpvGP8I7EdUnEeaetEkYzAdoMze
mKT1dcUlwMuukO2KSlRI9CrzItmaZMvx0d+LvNQZId0yV/iROmbDrsJCom2N9jUlZYEO13Ae2AR8
/M961JrUDHkq7TIkb+qmq/ejlcMaLFPUUns76Vsjqh4Od8PZuIhx3EFTX9myw8yFH+Xea5UIvoyP
snhC88CHHNdPP6TP24EXR7pX3oxlfudUH8C29SsTZ+dDOv3UAhFw9EP9ynjtlaeKzf45tIUU0V7u
F0YdEAC67dd9R5QQ3QK8AfnPRhFBxHB5fKSAFpktkOqsBmmuJ7St+6AIeRd4igshjAUNstM+ojQ8
ogwlBPdGBztHheo9nw7U8uN/GSfn9zZtHwmfliNcLJkwYDhUep3+E5Zxi34h+iZmh8ZlkHLjumKe
QH4bqMZAJdEQP2xngIkjKXoguifY6BtJZh7jUxzsZIIN07Sy67szjS2rZZiE/GacYg8xMBqT0d9z
HzkInYOF5Y9Hy1NGh4ylbv5AFBLYyXmWlwkA6P5S00ncqYoMm4Ow393DOuOKthgOACbNs9hO7+21
Ves/XKLMZS2dgJqW18tzov7/ogfHeISHUrfwE/xn2eNGprpNMb4HSmCwzRPFvygN0HBMGXTW7+xo
e7J9qU2OZaboFIYSuzvFs7vOg1p4N3kP020TcYD63p2QpqYUBRi4nztLX9jwBQj09oZVSS13UKob
znvTgv7MxQJ5J2Iow/GLvokGrXwU2IUSOydf2JiZgvjDcxp69JrX7PhkZV7QrK+zfhBGJhxaNZC+
tQewcXpEs5EdFsC8KiGoP6CLXGWi91kBo4QnJwineJYlEHQJciUV/ACoCsJefFrxTed0vfN0mJ4A
sgwqlDb72yUWkL9rrleLgcuBwZxSEwiuQTYVAbp3V+kOKMhGCdibOTEO7ydWeaciXDVWveqGwcmM
UNj87HF0idypFVTsIGFSq1ik4T2XM5oNQkW3zufQHrvf4QtLfvCK9zvsICU6V5A1I+AWgaIom7+i
Jf5rNUHCwP0iH6bdSN3xdme4syq2WVFglZqIbhVTAhV4VEHEjfGMabCDUPtsfPOR02MpHksXalp7
trvSVXPgQDhQt9yBY9mXkwn+wo91hDTvTxYyobLePQ1eLBfg/CzWa6XFOjVsoQpUikpw+3EBXe3h
tQPWa3HPbk4i+awArikOmpRX9Q6T2ebq6LeUysGBF7MB3mM8kSySoURIcs1tAPSN/4D/Nt9o9oED
ZAwUGaFmu301LP8yvrCXekW0xBydJuziVT5ML4dbCFH9jXv3s/lVtA6gbgNT6K/Javqjoce94rYh
WlG+AHlzyk2TcqRf6K3L4VeSSaiYY+pbL3D4N8SPBMHYH1CPt7RN1GGjqWIOGLdhfwmTRoj+Cgvd
gWSorY1Ke/zva+yJrU2+xqEW/BRAGaQXwIwmKrtpVRPe97AUhnmwmYyOLiocgE6S9fsHNnFUE0Fs
0cdO0+6wl3yBB3iG2kWzEQrCKSiaGokoQ8Q+0nozEFwH7sijqvxodvi+MW8PTYAuifpA9k8lN82k
WV6vW2I0aOQMhOZOg3gp3m6GZma3mg9rzmvwICtZUomvhdbq3jfPan6lOC+uX4g0zECqCgFSH1lA
0h55sUtBG3L7ZapgM1Ol6/nhPW4mL62dl9Ecmh3YHc+tHK19XhTB03bTwNoxDSBMcKSVTuLoIwVq
vd4i60LMVEEx3byNcXSZoS9UA8stnrV5oy51L3EoSaERBENcCPaMp5uVehsVuQ2gPZ/s7wBSwEIo
amSQMXHsWNo0z2ECpWb9DrJja4wnizWTLgJ4WIr521i5xAur2fzHn2TvSuWLu/9TR0ohn1YdvOLt
RZW/x9K9mlgUX95MkLgsUyqbr74ysc/W91vpmkFPnbFfWqXWDz3JYXNP/36QfwwTTpj49bRqhw+g
05e6tJboEEgW2bZ6Nl4kyePFAj825TWHDdvbCLXvE0A2KAik9s/YISe41cjAf2T003VvBuobttbA
3Dd5POowj5jtgxBYKeudwDNiaGSMCcf07dzgYoPiYKW1cKByzia/746JDMEc4ynAETWhZLvmuJ96
JiKzK7LEGVd2I7K5FC35A4t3k5/ik0EeGHJxnnMVS/fSz1DI5QPxT9YXePAvp6p7Jg6Rf9Tu8i05
I2gvCUd3x6KDMWKNY8f6PWdXU4cjt5ogn6SyoD+VWTZgsFeS3rFYCa1WtMVRnr1SmGq/SEkXWSbo
J49Cv4GiD3OAUYMo8pb2eUv5wpwK71D/8fluV3FFYbQtUKXg34cOPNzL2/qmdgCB1nZGkAF74n9q
XeclK4H71NpNZRnZrNKjUUz3kVGI3bLiJQdu0X+flSvLSEQQlmdvy+pRkLWIUkwOGeC5ScZXSZ/5
FxcdDtIywVrnNNx7ssz5wtCvzN+SgpY+gPm+x+fxBgjjZCnK9yFKuNQpNbqQrErwTRDnkcYrTL2z
vlLwU7KjgfAQqJ/O5kK/B68oqWE1GcoNIncCT1K0JOCBNcALQKSFe2vZ+v8FRoKYZHPDiOBv3QYf
VXsRe76JNGI+lcz5I6X1h/cI+ipAvRMg1Jledda1gCkTS60ke0XTAkL4aXyAcddh26Yvvl3G4gcG
jRv9+SUWk91JOMVb23Xs29cRThsN50/5OHn3vWdEQoQe2kHMVz/OYUEl0oGWuWEWwwKwelJAxnMc
Z7SuJQziaZx3fQCCVs7m7B0acRrJGZ2P62bP/6vEWYkQXeOn/aA0RAyuokqz8weSI9Clt4Hkwbvm
4LkPM1rVJuxTHdJ9QkDiF9Jj+7bmyx5QPjf/I4EgEyONFBStixGMYrGf5yO1Cwp4gFicmaliMc4p
cOdieEaBoYu/ipToon7TQXfxTayjpD/2hcPyS9anjTbaAI1gEL4ck8exW36kMvaMKRVG9xvOV0cr
XjZiawVFt/8vliKTaEdKJtbXXdGfl+4xRxbaccqXejo6iOOWbK42s7e9u5e1kvZj9yfcvCwdY9dd
MYYtQwFHC88U8zb0Fo+JQSbEuS9eKdDdMuMY23O44vdP8tlBcAwe7yuosfQotIM5bRNjgrX/jgkA
BBqm2SPibPjctKQiPeU6St9LuTEn7u3dZy9+Zc8B0AgrznVWqA1SHR9RMSqqQiKfM6rgVCR+79EL
HPMkSRd/RRMGPCf6PIFEXTJGLdwMC/3jHT3RJjvVZeV9d30fAMU39YGeZ4mtVG0dYZLIeCGif4Zt
H8SVbGwLV4Mv8bhUPKhGjl4CqIxC8BMFD4yMsvqB3GAPlKEG8VtZo+i9UjdbwR+MQpGEjmQjd0qI
Ll8C9QIOqUNfMdFtKijlYDefMayovEBwrb4JrBXmQFVbi/PTgnyqPY2ylROa8Jw0gyalSgjUOsAf
6HQ2wGA2+GflA+4TgovN/Fvm0HFkL8KbJ1wy3V0JJsBL3NhtEPg9eKLUQnPO6ICv+8WPFU52L5y1
wPlJklWvmBbah+65vBkPKjcIEP6cngotfwap2RrTGXGBEP1whTb3JrGEvmSukp2tpjOdbaZxSNjI
qJw8DEaq0NZkg/8pgxCutP7RJe/g3PeVjWJUHYhQ9WXhAVAYJ02EC6/9FVHkn7QrbyZlX1GATiF3
cmp8qq6PPNw/JqmEvRhLJpNIqnMpweuIeC+QZ5n2Z4yQ+AUk6QXjYWBOfYkPH2QRR4Bl8h1Qq7iN
EumOv6ypxR6RGEe7aYjKm0QT0Qgw2Dq5IpP0o12HRFxVxnBkbI5ATPJh31/lo5RsihnZB7/uAdWT
vYNn3iFXdrYhYN3ne5JL/AlDa8MoJxGwX06STI2I7v4s5xZzBDPr0RyYpjtKtMZ6mWR3REbN5mk4
BKyMYTeq5FTBgrcm+fSnHNDTmunYLd8LhEzC33qidWYFmFjuwNwkN019p8wIkS1eQgK7vb/U+b9D
LgSVQ5kYCCcnphmzEzYwjbpMJOZoqJX7bSIIJsOB1B5IK95Q7KXOHkutC1OpcsQ97vwhs04eauo3
9zF95don/5vwM2Gudvh+U/XEC9yRvBUAFlmimQAHLHssGNT6fOvfbcS5edbARxXhof1pUFYeN/Wl
J17KalNKigGWJnBKLTTyOSuQ6O27MjBzpPUwaE9puWLazjXwW4EhAvmZOFaxVbkkmfOhQePfkukK
r1F7uY43GQPd47c4MT2ep14EssqXo35Acca72M/ukT4FUDCWZKiQ51N4dzSdxErtHuvcMe28tDUA
aGOGAbHuS9awT/MQjCsUeRInQjkHXzL1VQHlCNYNwIlWqIzqlNwDaOBvpHa5Ys06UNXUTSOuAQcp
vTtVGCQ90gp19+u0Rznc2t/RKnItnJsPWL+9EiazEp0OUUn3/vFiStGEaB5iT7wC7e2PbBFrL2VU
1tY2TWsMtIBF7rnB90FyOHxgAJQRHeODYixYjrQAJKFDXqzpFn/jhW6vWFd+GtS0+UAA0TYzHgeQ
PUOzXvaSYqWisk97ujPPyAJbNfsQdafnR4QOMYOWUYsN6uvSPBY/q+oYeLfk+OGoTVkQBiOYjbXY
t4St0ychJeSmikTtE8EUquu//5GC3AT6GNKddrKGRA3K2UPVuWeqaDL3cGxyXwQZAR4tj4EaBHuU
o8hvNGqcpUwCZKkbI9qz1Im0JhpkZemqm9NKVlBeU/7YTFeqXML6Xu36TpktbPyU4Cr3w1waf+jY
W6UdClTl7+IE6UyTjrE5LwDOQJVsrnAPQqMkxdaEOBQnxd0a7l6rKrgr/LHTPfBOlwy+OspUtxzC
0y4VG1+piE6STH6zzohiUWMDSbaLdHeLY7g+wuUW723b1UPuyOHZYUvlJIRkN5fVSKcIMNtLC9cd
upR3ayTU6AxIml+fpmrqns44RAXVv8/7rADdpHMKRcR4eh8ywXX/bxNKolopF3GEPMIudQ3+6tHp
xZ2klML+K+iNNtyswwNBfp9qrTlB0RqdjHdefbF9RUXHYGWuj4oPsrVKBo0Q7JKdB1GNY6tUS9Dq
uJOGP4uuxAEcy6G8ukYzKBJsXl6OLlsUtKSok/L7oT+sQl4jBn2lTh6DXSbD8Kc+3vtvm6yI+gg1
6C0ZmQTl6vxhaQwdwpRnC5EVI71wh0h3EQcxDHAFsyFSfJO03LMCVbuzwnEj281mGOTUkYAz1S1L
4+z1qicoNtVZlSIu+V+Ht/cZ6iXnKHToGmKh4vhOuODdvBLZi/lCCTcv8sx/yxBv9NKzMqO65qcm
wNIljJA3b+rWhlo6EvkE61d5j1OY2NIJIS5NVvZtnFHMz6scAZbRukErnS23rZJ9VNSuMb1ArwAM
Kmgn9Ho7RXboaxb6gcghbQNcY5egeMOXBHGiEsyUXTBYv5rGr7MiXt0408YwZlHU62O/IJV+7CI9
GuQiv+Ptbe+niRquZNauaZVZjZ3qpmIsJp249II1XaVE971GGPXAICMGAzT1BERp+SI5yIpEFHTG
y5Q5XBln3QjriORvWzAf0VPx3O0kevz2JlOr9J/SZ2rN1TWu0A8LBz3gDhIhryGR+h2JD/gWcU/l
hGpRbGLqGaZ1WEbxRDmO8IUh7Mi8+uSeVuRKhQsKghSXBZ5UkvLERrnDk0BhF9CFoseYej/sISlY
mvkL38jJuwYX7tCfm0fi26RxyEGg/xTUiPwLDgwDAqF7bYtw2zeR3wgYMPBEi/7LXeBrpeBAcAdX
ljrakbHzrrPit0ylCCziOyPEmzw7TdyX8MrKU5cVZaHVjCzOjdz8tuY54EHfSHocGnjmJ2gkiKRx
RgmJB5gut/79qvkCJ5rUVSkIIDIi4UnJxBLSqLn+WsJvRCNLvw7NmLDdAgme0HYVaeGYdKrtWONH
AMx5gxYv9LRNgCPITDOax2vytLEdxjPon+nI8d85mhPD07nZSRltN3Ri8RD58vJuDej9mGOudjIG
JdWRB59M4qwKmyCa5KYZGPWQORBanS7ce3G6WLl1ungSLqhqwN4RJfnOTDJggZHddGYtaRkA36Dv
1xyZhdVPtGrF5gjtMPOvnqlnjVdNbYdLelCW6Mt+Ww7x66UzkD2ETJfGl8g5nSYufe+aVjnqaPzC
IJ2cz4ym0GWjYxaMJYfOYQ0JtcfId67hu5hG92D8cStG8vvl6eCLUfQKDuxBWK6es45tUEmOcrkH
/2eENp1mk9hjGWXnDPw8cf2XxVyRlKqJq/L/64vdQmLKuhquJINhgQ+wFlZBVHVNJBCMBx2YqjP1
YItE7rETlfNnJ4h6lohBBQyRdFrSNH41TQ1gYklAvsIfAJjydFYufp7/pkW6DJTXMyeJlKRGuYgt
TEwtQa19Vj4bi2K1sjvsn2HwCMmdl7Qumr3om48oG0Eb9Wu4s/TbhE3uezTg5WYLaf7ytBOUJljU
um+4vZZyIJyOxeI3lV6amFvJbAeNWFOnIeNe9Ad/2JVEs0g/tzhsJQpqlV6FJPeyw7n+d8LhDpLq
V0mPr47I1/g3mO4mEuVIxy5HWoSU7RmZ4jR1bX6cQ4gt/VZ9QUwkKYXoiBynKsIlwoyj2x5JUz0l
+tILHD5NZPgiyTWFJddMKv8OKBkPGlWxZv0oCD4U6+7OLSme1fWHfcU0I0J6Ny49UFgMgb/Eb44s
4Yy9UXs0vX25mKjp7gsOYXNT78ivct70c2IrBi93eJ0r7iwUgcqoYcUnA9c+LxY4AM8+HdZnfmtO
rAWcY4KExZpVIsk2w6Ycgj0rUJHjpY49otCBS43FP88qgKesRuPE1Xf6Ru7jC9FTscePbPT4/GmO
t+4vHZ0BSZzkeDnN9WBd91CQvxQ7GGbyp/d51BZzl0QEfDK8ind1PcHE4tATS0ld591j8Bt75kwB
W2XS4cRqUyWwhLNjVKVqKIoLVbmksJwwIVveo0awNqKaDZINL+SClqYwHoxzLeEAdbkItBbn4lOB
+DnnNabM/tJTCkQ7PNEaO0kQBgqiwOJVTBY+IwwySiJi/UxysQJ76piMYLH6HCZOyyY32TzEbmkP
xOQinwn7tgIO4kTlA7yhH2QV1sLPgDzXFvrlcIff4GIWCjfDFqxgX0L16FIwjX+WA2vhKCl3ZcPJ
PZL8nLPwERS2zT0WiJaT0YHRlddyo82cCTnavJxgSt34z5BIbK2Byo62u+bd84htCDLaMSjdd6V/
E/OPp3q+TcBazTyURUO7SA9KHKM816ga4mbR4G1UCM8yjlo3dzRbw3adbMNbRpaTRTCGyfVhIEqG
RtLQxQeHLL4EG7PFy7qwXBGxXrpnnOg5S7IgjQyr5XE0RIo6HfxADQX3nEemTzI9Q5mXHfM4fWw6
j/G4UQlDe/jRoF3eUeMn2FK1jpgfsIqm45n4PmD1wD6Or71BAo+4NkObCUS6lEPcaD4ogjgvbFmf
h/Wr4Jhx9z9EKxplyubY+d5q2p2d6jfq547u7h2CbJKCUAnF/y6O/L4XhQSTOQSsMuLm5PESY3dL
qC7Hs09Krrhs+LH2H+IdBJRX2GuStmShOVw4/o4265Gh29nFJo2G7EZ4Ovnmm2Weg1mJp+v83rIK
/5LCt6ejetHW6sLzlfgadtPcP9NWdAr/B1efUvvwS/deYdTjkyWpbkdMRNyAfZaAXMvxqdozoL9q
k1Z3SJ86nq6yL0sSgEzs8yMFtd+pH5ugBmGBTeE2Fz+yNRp4hvsTPuPQ0735x9UlKvUBiptmB1M7
SpYglKxN6TndL8kmvpODj+Z7NMgYVXUXtxblLp7D6cckKs8Xy9HWefX9/g4lCjeSVp1mQl8UBJsE
6wZA4FBxqwakamUbvXC3fv1LjWSQGOjNt7L3QKkII6gbs7Aie2IkVEF/hOXiqpcAE1GjiDMN2sqJ
fypUtfZNNHRkxDXisd3AIToYUvMO/G2lzmV/btonX3a/pvC3gBsctyG2WC/+8GSVObcQzUCgAH7k
rb0GdQueA6WV2l3n/q0iQK8IBidraEgj/YZVV1iSBZXTSReCxKOGnnVUP8CHf/eEqp6AC22F42p4
y61dstII2QNJKxL3QBFNDdxtbfVh/0MIvUye34hSdTeeR+KRHxPEWYB9djonzvPPOfgLYaAtPmbX
ASDSKB6TJMOovVqOgwFP7nrME4uJH6nuMoWQDYuGFf3WZKUkFy+0e/5ikHKV3b67KSIVIGADEilw
TtqDoYoHD9KKz9ObQDEHbgdMPHM7507AEBwwYhZ65CeUG4vqlTEHyxvurCZmMC3WUCudPniOMLUh
s9Yaa9DN/tQp6zy3/3pg8s3CBPJDbrcBmnVb3k5LbkYkCm/SlUDC9MqR4w+3p4QbuQKi+dnxwykO
igo7Tp5PJ+rVg6QTG9ErZdn1dkMA/ww7xFG2rbDoqEOyf7Iznr85QxHT70PseZM1FoQUVazbwF4J
YaXZCKuTnKpUREbAoXp+z/t9pUSfmlMv9oH29HSIf2u5qFHMWT3YrBiQii2jS4e8AJ3wUzsjUIYe
WN3C892xKl/CdX7Iyh7UcUNzZbxInMKhkIV+zKGEn3Z5BU8P5uL1o5v++7OpWoKRWdyKsofYcaj3
jDEhzCZR3Z4H4UKa7UMB7T2o8MhsVTPuRgYF5LrntMibRguF8IJ2IboacitDtS5C7mDXdBZ6Jfav
tqtcC35ZJuZZroHRbl6koq/RT4hpKepTyW3tp7ObrSU9/wTaRrY6mWij9ijdtLTBU9JYirXcGIgi
IbHI4jHzycMrKbFvLs9bPPTRh6WAcO+HzBzRm7yAwwgJdf2LW2P/CBJMysJgE635k7FzWzbIrz0t
EdpabU5CoCoqoz4JbVNcjVm7Yr5mrCFYEAf+t2c7kmcJPcR1ZWhW1yoNNwanyQMu1fqVd0T0h8Jw
aJDZFg5CksiYZ++z9hYnSyR1lV80fzLd+rJRBwWSyPvUg4rR1C0tK4dhXGbQ3UaPhpj3A+2rQeRt
VQWE6H/gvKdaKksCddaicG4lSMc2GfBp9ca3tsT0AN5+IooyKiLPDhMgcYmkAiPkuMs++dVKbCBI
g2K0qG9HoRxat27hTUqzGYoQPl50y7QucRfYpqET4nQbHLxKl2JCxH0yM3Zgd2UqyGBNaK8jUA/A
/bMzzBz07RUDEAVyhM1QTSr4uVU2c78HzLHxPdlksK1r9GIYJP/7R9VE/ZsN4mEkbcy0iaHsrCiQ
kg/pIEiaxRt69R0udqrccwZJMhJzxR/1HHRHqtHVGk96B1gNKmveaH9AKvw6ZHw20sEZA6OwtcRM
unx9phtlrCKCUbTYdp8xSNnhNt1WCm5i5+cddetqyipAhl//b8EZwrqPAIepqhwNYDHuA+5Hyo4k
PI5X+DFkupkhN/CBX/XIdaGR/72G7V8fbXdohcaGwDF+W5iyGmNynopKxgcQ6WleQJOFJtMC0z4M
2DG2+SRm7A2XCzwl8ykgxD0CGVkzu7/nUIrgzcm/fmA6HeprjSbH3KJsZw77SEl8mMM9XRApIUfI
j8sknSiMS4lOVAbdhlz7kLYeCXSIjhVzNzExoSMWn+uWr9jHtrWMeqVoee2GXLFIX3vjrdwCDbf5
VX06nxBYVwzA6wuMrJ/2Pk9qU4PWAddFMs+4gCuazDrpANh29PkYo/nrsrPVs3zKjo3uWMu9/hzm
SPSnLpGFH9uaDXAKCBO7Fzdm7cS4z3a5jURIMGbjuXVsQSyB1AAeluJhafTCRYYorQxOkaQXGSeb
zvoR4sJV4+3REi8j8pNnCkvoNIkImpU8eLcpXMMvTSgmmsFgexlD1iweKGKFdOomuN8BRTJsWcVv
TbiigpQZmGoxh3hjvng5FqVhpny5xm8iCFRjMvvMBA52CK2eeDz48XvpO7VXcsPux1kX5bQCwGY9
Bq/lKxFFv/BVEqJWfRd6X9VxNqWVvCWDZKfOakYWg6+vXBj24fCloP5YMaxSd4QM2t779Fd9aXOL
c6Cdl268xhuSpoP/6s3NDodHJyPORhy2LOrsQB7i6BKRd8DbKjjLYrbGzjn274Opgwyva7gs7h/f
1uhkQG2M940PLbB9amPQ5lJLIfki2EKRF6FfaF7Rlap1PmdWFHQ+lTGl+AfI2foMZIlpkR9ZRifY
CRgG7n9Rkd1nrj79lvCONZlxM1k2HjZldbJjT4jkWB95SNo6Hz+4nwfjgYVfdo0qo5AiVVHf4wf7
TRgAtZuY4IFCKDs9gjXhW2ghfZhguaPwoi4qo4CPipK4UKEUWHJQvROsjJQ+iavNn4zy/eCFaHqL
1Wmv93MaFnO2l/YrROMI+0SaTtZETSxxq+T377Ok9vTig2pOd7vUp2fTUm7JKsKN672p0TzcMaIA
LOiiy3t9QkDPq0gQXaorm06PDO6Ua/trEzFTEab6rcGJGKVhlCLxPmZPpKZ4O8ZzPgSOFJzZThXP
ZwVds33OKjch9oFQSeE2YfMvlllJnPqxCDNN5kIZgvXfwlL9uU97nIa227FJCbqv7gf4szxCqZZg
5EWVSVJWnGASo/UjpJl8D3YxVEKGfCFOTeNl3Go5kwi69mEYnWlcwJ3cNsyeSCMcWuuiv07tKDzU
4XFXaRc6fFslw1QFrdHxcZFEKtX5DKKpWoUfTcvkw7jl5LQwvd2ogpmHuc2GCLhdForBZRE2t69m
oWpQpgeFIQx/VKQo7h9ZqMEMF2q4r56ABJW8dBkoFVo+cSM6zZkfv1RsfqZ+iJvGWgZaMwooD55Y
kPsXL3S7/QdnTfM9YGtHR5hVR7DjbM8xk+9KnIIsdELPBoZ2Tp7yFF46E3dNzbNuUhVcVPfH3hHI
eFvlqrncrMKlvVH2L5WIqAeP5JG9tg4h7673eplf8rRVVNxdWPVom4sRA2g+PlFgn7HtE8Kp8Ooj
MDK9lCjDcDX4WU//pK93aqsRZptwkRUJfC4wFrfpSjdddpPFeaYYuhG1z1HHJmMnvgc7hzbu+gQU
bBhwfgHYOFYqrOMuf0SIfOqxC9auP75GR/Dc1l5fJ2pN2tl/2aME+8SEd7MyKNV+2uhhThCzIZHg
TjfXvMGzkF4gQTNeNcBQmvqgL2t1SVVSyqa6yAD7lqTJi/XyvWY6K8PkrkQ6W9Lfkos3Qj6rVr5N
XB3N7vgnAEdOjpc+Xpw8xC+yvVAeSFfuM9RTfRvfl9kwcB7sNAWuTWYw3+Fa3F1AedP7w5sFotat
xa0bEiYag23XgBENEL+bddWuQvbT8TgxOmogGImofi4FgQejD27YqWX8T7VcT0QoAoMQa0WVRZ8X
VxQliLTcOHeg72bkQXNaniMKK/bWfu81kvFEH6pP8oCxWQJz7SAkxR/7lwmujdDYekrkr49sqaWd
9VzJLe5Mroc/VcW/V0QmbQMIyRieWQINpg1Tahcb2Lcq66MuVAXBfLBoZceLbNK1A7pggTDh7WX3
CYGk1T9XWetXwRXvtqJl7heyTJvxsPPBpR74liDzyxkmAPtRsFiC3kgOPK0h9JLUENniVthMPka2
RyMyDi6vgRv5bBu6BZ4/TB54PqOTR4N1X9YvQFbWlwAj4GTXBfRzDgHe2Tfq0+NFhX3EjH9Gzz59
PKeVUyfL7AXCDT3/SPmRGxBNuSAj9Vg1btfylPaZUNrtnr0F20WPNvTZdwAoxLt/GsPtZkIRTqW4
t8M4eR2A65b79DZCTY1oSFGIIeze/ynWb65SrjBpmVpLGYG+SyJYircJRb49Q5YMbpZP4TwIruAc
ASGQBA3Ki4Kx5aBp2fcNjqIaaaNjkwlwJKS7ORVUCDDaHv6CxppJtWvh70/0xZnWJs6KPI1w15Bn
vrMx93MW14leqrRIs2Kwf+LXg9ThcoIcxF2ctlBhPJ+XudJaa8n9gyIM/N1IJ0YZsYjovh1iKJt4
8bR0Phg/XbrWxAe8sE7HI1BuL/KgnaUM3+sbbb8YRm8OEUnvnlYWqGbfIrwYU+ouP4VBt2msgiPy
CWKB9hy75yw6ocpxBlOfbTFjmyJ1UcojgpV5FxcsPHosvij/zxm0Kpl82nEiWaSPEusthwfeY7cC
bL/PzbfvTqdXFGS9nTqO4ko9ITOuOzEigPKM3W91kATRsSzkx/0/7tovXNNvo2s6ioXNMaMmmy3m
MwRVkF/Yaax7wDdiEWYEcvJEXhMFbwusIK0Xx9ZT4OMEq9JGf1P2teVI0BNVNzX7irRZalXeDNQL
4ZxP8Y1C0MNgUGsUFOBGgrScbBgaI3htkJjY95zw5D2m876VdVvbUvTHxM8gOrIq1QLISHRtzO8i
d72GFyo3C3E8zrEbrgPpWA2UhyXFJm4K43Tj+UQWBXN0mq0KowIcX5FkyY9IsFEhpGKBFPrVYMtp
sTRl6sZnXfLjt1J+OkZ6GaB2vFghU7KorTBrG9O//OEJowqW8lPJt6ssFY6WZr/NubGd6BUQMVDr
AWfTANNJfVrcZ4GJO+/ylBq3qyE/xgL8UF+bVPOnVsqBj6lZ1VMHiZfeRTyINw1VXTrnQpe7vaob
HNCLvs9qyb8r3tgrOPLQq/uBk1KrvcM0r1NJdfjPMlbWLCBufiTvOqQS4+Q+Bvq27eUlhdJcv0Py
p6rjs24fGIQdmTlkx9XBy8D2FxqvlNBQlAzl5OHLw1IrLHYy7Pd9yGlzMdVvkb/n/jrHSFjdBY52
FAD43r/wxizEgV6LYjg3lMCMBx7QPE1BRfe1GTeSX/rTXUO988kzq0tqwzj8IsPlNUG8+1ynqKFk
qg+djCenfWrWWH8gwi4Vs99T+6blJ56ofoDirmKAsBqPCmjHqovOdGskqatkfYTaPNU/C+LfCnb8
ImC2LFUHrsvhrYmmRMXoWZLtMbxOx8F+9c+PvK1V9mJn+2WY2jqYfXQwgoUe7GSMlJugyJen9ZcA
d2SsORRQCHDCQpns1W/GdxsNMOqsZgZp6ZZMJ6Nai8NpP/UDgBPlwBlh2vfx371Ke1eZpUaAb5e5
WpRP5otG2HyCkkO/Kui8u1Z+aQj+RNWT9SOlgixou+NLaHDXf9AyABk2PZ+7XqzD2bOLKY7GLGcP
vJbLfw6ARRH2TdU7hVdjADN0jHg1h0HTb1an846Cy0EjJojHesCZUoEsF9nZrMShjlA+PdvnBv1v
vtCI3G1AHslSixbIa6K460fFX5fhTstHppc4Lr834TU3UvgHKiFqM6bqn5UHpr+6Kd9PkW3RKehO
dpeS1hJr9Bbu8KaiHu9dOIlvpbKQ2jXIEmYrDE+6b6jJo2BDsGHFGNNzv4+abefbb0B6FZ7rMz9f
WzUWcl6ar1Yf81zHAQ9YLwUs+QtkIf0mmKVEGqnrL5HH2R2mqRXlmy1B8nyzH0Zf1FgsXBPw0fuo
Metaj/9q10EqTwCeozqcXHNpj8BeBVYvwsMOWb2HmPTrZ5gym5kbsr4IBQSt4qnd15W7gy8DarSs
IAR9vIZz+SoWSRoxZ9V/SSN6cjPS1yNyRa2ews33Han9fsjw/lR4GAPzapxnnzbIv4UCJb3uXDjY
nGo3rxEEy1m76/L++Mx++/3X/3b6Fa1jFasLEmjMfIpxaTI9RWr4ZGYzbfiNj1aVhx53QSlI8Zcm
jdKIlBEfpgTUfbzzBNql4J5crx4AuXbVA1RfowzIGNz2+s4HYttxJPGh154zFyXVCfy4pdmnxCJp
evy3UQJ9/ekvuKm8CHd4gFBZI94Zb8Ci/rCG1voNYfEjbrAXdip5U2canQ8kGDHLEMqfqcb/DMQX
cT7nRlgQIfoWbYj/aJg4khCC//vo8nA9ZGiiC39Y/Wq0/Fs8z0AcZ+KbKRPJY7g+yzkrhaLNeRu/
GkyIt0kh6ZpzaLAG8i+b+oJGAdNIWoGgvLGwdFODG0DQAvttOrBUYij4lU5wjqgg03Zy0uVrwACW
1P4FlxmQvHO4f2Ry3Soj/6dFc4GZRj2e1oASdREbQRD0NHpIukQ+K9iGi6YnwKPaeU99C8HNBH5G
puUjErEGBI+Os1rF+OgesN8CBjZv4PRMDc/g7WN5UKlKlak6A9VXQ/8PsePgay6CpC9mmCfNKdzq
+N9ss5X4aBkdf9Us9c6bw9s5P7USm53S+9O0AXZ3CXt5qmWc3/dfAIQMVvoEHW3/clzWgepq9rht
lm9zExQxQVjXIJ9iWCtEWwawkJewt/J5irXdazHYOvJfH4q6GZgxTCydLB5IH65jwe3dpi28B2/e
PQjKhsgLbqGt9ZummGeOqZxqEnRfVF7EBTXSxLoKV3lJLadEC7S78HOUqDJ6d92o12XQxRjiMO20
Bax4SeFU2I7rYTX6I2mdwRAM/Ux42vMR8vFxf8cdESxY5mqxTJ5wC/pTUn/mmq+cPLPZBFMNiDia
NXCDRz+dFvpBkiJnJLQAUrhU+Udc5w9zaH8G2tedbB9vW8G1YunEAm2Q6WYIR4Op/jBdSuNaPU/i
sueieFA6ChtfBdkVYJagaSwQbP15WZl0koPizw8ipvTHbDEOBPtOgkZulrQM6iLGjQuqSbvw5bRp
92Zf4B5tFvHgC7jyD65nUi+o24qhi38L6hKQ1FF98aSIUUVk1C2+jb46SfG9/MBT8FsfxGaWzX5m
eQY2Wq3jjws5DBQsYuI4o/WPhuqmWbx3uQ9YQcQSQqphduH4WbeMqmGsdXusN13D3PGG6XA7I1DB
hX/IdYOGrOAYPIVOYFtjgyzOmgchecV4zcxV77UKmPc4Wuk+WXg64gdZbDakW7/h48ERKdXU773P
u2mRUpF9orIDj4yuSCCvSdrW+Mse+sXmUUiuvcHdSbk8JYdCrSwmSzpATWaIEzM9akWXaprYSvWX
jRJh0DE2q86QYk3ozYySudZVLXGBQ4HkvwZM7bgaWnEZ1k3JGexqoLae35xsQLLC6fsG+0uGdlox
PHfDIXJp8TXA0ld1aZFZ71Hubu4/LnaWnymshfCDdcHUcIRfJp7Qy4o+m9+A/4beThurvnKxrZSv
RqW7WR5mRgRzedzNAOsMoDxnLoXMY/Rz+ILkZ/JGxz5TSlq0zgu6UZ7h/xAFvwwAVTTRM+nSBJyx
wYVbVyDK32KMNtS3kvi8MHTKD9SDJf4beiLDbVOoDhAIbLfxEIJKG9HmWwQpdT1PE+VUwCGQ5s0K
/zvXmSEeG0Bhg2iTI3d/m2SjD+S5sRmH7YISEiJ9r/bVEDACBCMY/80i5KlEqDSPRSS3cG178g3U
+rIyCFEmiNARpVafpBJmFoQrGFTtVoSltdCCYNTv6RbpQW0GlIiIoQ00B7jdnp7ni7O4FPUbsy7x
X2D5CuJzp+8CpmcohPNRf/5zlBNY1IBfi5KMEprtuEu7DKrrP1UESmJRsRcrXMicb/nbSMEKAYik
wyBS/3O94GK/X76EJL9JxM4l/hurIzdfRh91Mgzi+nbVk+qvj2O1Jwbo5mwwC35t3R6Gp6Y0Ko7p
SyokKOxR4nls0AAginll4+V/kFRzvem4CnbZCCBAzpflQLSGVaU1ivz8GBa2tNRXqmBkxjfrCYdm
O7B2CV3BtQSSLnvFo/qsGiGhLahW1Btrjsun/onIeNJrvaPV6gpxauJW7lcL6XdV7xWfRqiON2jS
MfM28tVVS81cW03X02KrdbBJBW8FFV5DtKo5FXBKZtz8BslvbOlXq8KXY/ea2cxu4nwNf0VZ3xTc
MguLzkwD14xc7FPc30PTm2hOd0cFHRVDdgKcXOSEvy46nOEl/S3YTV37xvx1BrTIh1zkZwTgV5GS
d8A4+huz7AooplJmIei4mUMIj0bzgJ8AJJ/C6oEeVF6GW0hBc3DZLN/UPF9+VoA5PxUMgkB8uwJN
Syb12LN2Ps93/vgHRhuR9CntZSC30xsY+9X0LJ+DIwdnEreV/+i+CGT/qupDPyd0pn3O8yo604/v
8Np3is0pp8VeE/I3odoiBtvzp3ZmBNaqXGU1TqoXl8uPfr9Vrn87X9hbq+NzYlGU67keWG9eltqV
OGv5SP/5LMnR7fayqIPBpGDPkAZvR+4P1CvmMAuTQVQUwzj8u+6tXUVA5fXs5DYq09cx/irGx265
1LYP3kghblTAGGC0WbfySioR9WLKOXxLaF6pXfMIwtjXq8Opcr17ziiuQ7PwnT6xtMfD0MntRKre
hmNujAiRSbLtJEqoAgClmeRW+x6uxQRHp0ik/OJkMnzir47sLlu1rd1vRlrJbc5T7pvglc4yyv7y
hXCrNTiEHF3/x6wF9Sg4eLvc1rZEpU2Y58iPnGh1+Tq7SbLYDf9e/SS0r0zlL/wkyh9fxCPk/sUm
+rnxmLYFmL6AtW3uIVY4GrywGf1+hE8ABlnbRlgvaWhrS3Imyf3PuwhiZ05LF3wosNZBEVkFUWP1
KUKRQrrt8bLZENc78o2fvfAHiJ5v83O/oIiod/6g/NMdYeshXX8Xpp22jPc276xgVES0dDk2D3rw
m1E5W+DujcWhGg+1xjc9gd9YxiQbv4O5rdltHAKKSU/km5eAV4e5B/O2YCCGMDwzDgIs1AJTFkrh
ErQa88p9FbDwGMUaLF1InHyHaBBSvm74EgUOF7vDgWuOaHf+5CPBqkdRc+AJ+3/EwJRWxe57sjaZ
51UT1XJWUj7ktfilRZAySQ+b8NfH/16hJFQN87TCcfEIOgjt/w6EYRQ7FsfdNjRfegH2pkdZ1ufQ
nnMFtAkiqdyGSoe0xH+m1EiNwl8CALOjOTb/XFSupI6fXpKvkSU5lBrdRBybQ4sJXvFNLsni+aX2
CqpuwT8i54U63DJCZh7QA24PeiPJ11ysVIeyuk/dQcnjiCiqOzdDQMxcHl5TzfE5w/l5QfF/uC3/
q7LWu3I0r9nr/QURCz+o7yAfxxUf2tIlvBjfGw/NePKsTijjHmd9XNm4ECTc4V5s5nsOSCNw1eGK
azd/Q0TulUKe9uuxyvFLnng4BtWXJSf65Z9fsRusxhTa562Y7SBKSOIS0XHim2caVHFUmh5eZJlg
BNiS9KGcdnTQwOl3uQebp2KDDwaoGTZgnPloyydXyYyhdFjeuSq26G3reSW4CNrqFBE39iWwuDY0
W6efBT0e3HWo+sgBX8ndFR6EY1fxgBFKDezgnAFqehSOg6npmMV7mBrbJRKB6fruRkozFa7UIQss
lUmlPud7kYf27FrAjKme7/ooJx5GguCMMjP1sR6lXzR8VPVjGYyXXP7FmPvRqTRfUXYi2ijtBHUh
DbjqTz3on2AJgFPlXedzFUsqmSNc184Q0n8WZTfW9/tWikQneWzfXWps8pxucWhkE0ZpZAwNA4g+
xZb2fxuLHaHXgovRCPneKecHg2qxpHvGG6voGVzqstCrV2ALcgSZrB/cnIXNN/OaRGbbm+zvBsoE
5PG+3BRmGraVx6IK+pQzBYPHLFEdWZHyrejvcL6s1PlFMURU5Q/5AnOFehJ9B8MllBioQlm5ZJ7R
27aA13hhnbFrmMoqnS99XqPiTfuHspXGMRk8iBhPChkZd9E+1Vft/2gYvxe6O6ZyLLGXOFWz/YH2
WsfPr0rOaukShZln0op/l4vni+1Yffvtjdfr0cxwkaJCmIECFBJ071qB9+zKBIIo2sb74ApZpqZ0
PHcGNWZECKwZjccU3jOcNg2fvLjnhzt3ILOLgWWlwl5dHJvX0VKu1DOZ8lbidRyyRLRO5ZF/b++x
kbrGp0l8bUGru2U+K+hv5e0XBZUX9NS2W7eBlT4372RPOgovafdnNEhW34Rw0G37bCbvY4HlmzAC
1SongNCgzD9J8xc/mfpeHuK1JKWZmHcZaSZfm/doGbMJcCuIQLeBIhGYlvnoyGI4nS/QY7bG0ZBo
3PhXe9R9zOTSXrMz9gXbfnBNSFYcmUpdYgxMMPUzutsC8SkCmyJePe3Ypxws1sOmRBhrJl5XsGxu
5X3EX+yqZlDCp5sg/DxIGTtkcCKAtoHjud+VPB68jWCGspHDKtTCni9eaO+y864NRbf/u0//A3wr
wjCaiyF2ycP7DayeQ+E63kZQhqdRXWqyuepLSKpRE8oSkdfscu9GVTFPzfZsNFng4fs9PrrL4yGp
18MiRTnqtvEF1/otlGZtkFOJh/g5mHqPP62KUPy/bJE+Xjem4XoAN7LnzooiUaAuwi4WNUaPZgcS
qPnOW4ktW2D8M3bWRE8ecLJXJYpWp5bcNLeTWVmCV/fgV3wNc1/3PH+SJF6WELHh5x+pq3kuBEi7
3X2timVBTwdck4J7XQ4RVpknj6DKyl9vtAPAwiXOGJK3bNZ3o68ZuXpLzc+qQgljg8ZLFbSQ0xyH
6zd3KHGeXQFgClD4ZuX0de5rVa0vnYVwaRcltRI+Tdb3/4ZI7rb2R3o+edh/7+FBQKM4CCk8YyAq
EBGG0j2SY5N6mZ+vCiorAAsRaF5V/KUHJmfV59KHrnit1Excg7jqSQLZffGTyxf7uPUvlWyv3fSy
Exx+3JsaoSbhBUpTwPdYvs0mnq9wR409V+EzHijRjBndyATM7nP/vAURmyIWK6o4Tvt6cnacGIPH
3sj/YJflTy8mDSrVgZaletsTZlwNrAYZcnTFmBjX3fXMgeuxQwvNw0CvU0EmkyecBCcBsmyN2f45
GBGtClzBaff1k1ldqO6wNmtzVlUEXAZ5g4BBhF8bEtMtwhsyDxnUo0uDJYVc539KqGFC8qXn1e01
1+vqSpjvDf7NDaJTKS8p9YB4kIJmV+JxtrpO2Ua5F0q0lhxoae4e0fNyjek8ai+Hv6EhC+90Hn5x
76klVi3jX5Emmcx1U5PH2lUBcA5Ob6t/dXNi6MdbG/aBmxDtGbsv4E3RDja2T6LXPbVLwka+KzTK
+tm1jev19VaHLOvfaeZAiiklmi1BOHwt44caf/mMXpyX4f2HnVykEekXIbrIrG+Dj3yyLipkVHD1
eFyRUEtowlUjC+IHrmmC7tsuZy713vwLymydyMv+Lyz9ULHX4GmI4zlirz0bBhjdGwO+ReNw8G/5
lLewr+h+39UOYxei4GyRtUfLKzPxIqD04yHhTEwrVIkO20QzJS4D7OoXV1QNNuinjT+TAsajIk1i
zSX63XppPiwmlUTFmekmqRSI4W7phgYu+zsOMB+hVWKeiVzU6H6t9K4F1J130omecq18ejgOBj0+
YCzMPNC94Z2XCp5xxuaUat5fuU3J9F8RevXE/hZXFn7rzq18zUngQrSBsBCmj4h7EBRS3h3DHIMi
4mt1KH6Zkzc+8XAj4Ns+gIJG83L920ZShFiferKE2whcUqsT7DhQMWg4ayUF/fRoVDM5cIZM1avM
RBrSNnKy/1o6NUjFchIgAAGJRdsYqvdO3ArLaP6mX6a6zhQsw3LXcvfFRFtknx6JcIpSqSxXeuBz
hZrpyzu/gG+9QX9t39Mu4+AFLz0lpc0yUNPLeiL+3LHat9OnFzE9k3DlhNJ/+c27mvQwGPMyl6Gl
aawyhWDU+5bv5lH7/T2RDsFNu4CfUhQ439I4iax/Hq2Stx60a6e2RJo3Ro/FkwbD/AQW/T8OdWKv
U5W2+6JnUzsEHxfNiTOpsnWWf/xvip4PLyfS8/0kwY8bzxWWT3ZB2tWiElDGTx9gIoyOAZ+6Ffaf
cykgwFTcELp/a3O2JO8Fx7Uw4XZtNogFXPsEhEbm1VoE3CARa4jR8EDLlJRGsOrK1b1NYX+xKgKI
wLq7rCWf2ku0LQONXVaGAa5/0+I6/XL8cn/qTClTr6ubO5j//xoTW8XQZnBTXsZBXxCalq+0SEWq
iCrb56t01v+lKGmryeoBLQM5HxLDOzOdGpF1uwj1HJbfsUS0sRnUmvj6NnOS7Yy1aS6Axzvhtiot
x/fUUFbHFSJNBwlpqvr03RPTEdiFl0Ac/w5Ry4wE6LVw4lKxADsEx4/nNEyStJ+v4zOSFNm0ZZ8Y
GvIeYcB1lpmJ3IDj2eGnkx51hkWrlKn7P4nZ9DRYZ9a3uO0G+zuLDZhOA8Jg+S4+MVfyhoDFD0Ua
qOjJlhBpsjfT1zMdeZWYBcbrO6uIFWWYcH1ScZnM9NPjqMyZR7CW0vk9erTjnSjjKKggY96Ngrh+
i/vpuSExxNaN8/g0r+xuI8glmjtkQHWSwZR6jLtGERPlU8b30rcMaRT9zVoB5uT0y6C3PmFu/hSE
RkJ1zpIXVfBrRGfmhOWZeO767n9APQjqeEXmVNPgt/jZKZTmQ1IcIAa0VrWIAukVBekIzR8+hgZg
O75lJhwDRccyt1ZIHuFeLiuM2cXqtBZQ7LI0fEDHxtR65lB+/IenguEVyYZhapJwFYoKWy7fGXY8
mIYkTbeJyi8b4iKAXJ6hxUg62p3cv/Qp5c8FGFbZtY8gA2fa+gnmy18tWDpokWleoT5EiBEMFT11
5HPMcCduOSUNYHahX5lIjTURn0T9dpONKOT8SQdBwa47BJr5AsefPUh0JaA4cHODyHS40JMB9fkk
ZV4G3UZUIEFX0cYko6agjQiBM/eq9N3DYfi143qTlG6ycjXaRtasvY9pj+hEl0mDYahaSB//YAAj
o0qEI6KcfRpVmOvw3qqijd+tapsW5pXUHkRzegunww2C50fMzygx+vDA+sNg403Ipoooa8R15HPd
KezdSi2X4UVFAM8AYs+9fZKVqs5JCYlOqs7OxLhWJ8J+JfGRa0/9Cf0VaoM1AwPcWRIpmCNhIE61
lV/MjIa+lpwwVxfefZ09ss9soOXv0e8W3R/lCI0culB2ZoTA8z3gK4RIOOibwfIcuLqAtmdQmTAi
3ngXG3xMOBPb+iWfKOQLPWi697YLSB33OnxrHws/VhUqOlBHiTGHKs7XUPYRFbmFv6lbRL0ah746
MRXasmJAl2HRtiVpFP2R6qhyvPDcC6uWhCfFmIJWpFb+zHtwICQJ01ErIkLuJODEQguTdKrKOYNe
teCQaPzR/x8jcW3MTK3/j0/dZY6yNFIYl3NeD/rZuLxoj+36+uiAGTu+4Q6ZeAXVpINM/D7VhFeA
FWwixFYqWpqM5gH885fQvNQhSfcwEqD0393wLGnxbW6yaUtx/mB7f1vHaAotreYNqmKfc35jP/ub
/uOtKVkblN36cU/RZVYNqxaOpVo3Lj5Ku6WmDvuavEuCjsbyIbtC/PdHG8OCxttKZ8SAQhxOjYoi
nMSebMtDkKYkFNQ6CgYQmke7tRLWheX4EjFpia/jLCCRgjoaOVnstP94O2kzmRUf14Q466nnp5xm
Q775RMnpa7OrTrpoahYVdHceTkg306hrBuXIeekh+5Ra4F530QDVlzxEgCNFT202iydTqMP4bj0A
G1Pcy7UXGt3TAo9hGW5WN9r5gmjbNLH2dPL1Mz5MUuYYIhJJCGnzVwLVV3SHMAd3EwkV0onsNQ3W
OwWiOZKUMjdRUatMF4FnMjL1P23NbcAo+OXZlX0O9id6G06mM3kePnXyf2jiWFLCB1cpN9ATdd+O
qTVCwuLcPjRFz31vraX8mj63dcw2uQnMzpqPZZEAZ/cTomzJJY7cD61OdKVTkusEuH6yWg7jhpCk
2H2RWP+sI2PMCofepcdLxnM6+ThmCQY5Ajw5mQgOgKhPcVho9oPDbgpJC7+Yb2lo8NKpJRI+cVj0
hJVDUc5b+2R/alIf2Kh0C7P0rpPLNF7KIh4RHAp11xNaOVO9806+w7r1RvdPYH/tkEDPn+pA0/5y
vJb1jOpPXVtzX54a82qY1Y71pfG7JmAE16aZvru23fjaboyxn1Dcw1QRJ/qrttOTuTpzk6St4M4d
6wUmlRAvvAl+QWTNa31XAkocfSnidusAuzwWGDMVadcRfOG4kJhU6BWCYlJs7z+EOckrA+v5XJT+
+tQ47COhpkpGdOJIaEVA1koVzF5hNQ1QZfWwhxBlcA4eu77n69cbuZt+T0z2nsKtp942mULcTKs2
ANlhwwjocWqPCd+wICDuRm+1c3vm021IvfT+Ekok+/tTYgF++rh9NtJTd+HxyKJ3Fgqza9ranF2y
f3gqoUmqe20DOzB9/yH9V8yQ77fSCFOoaYECQAfMaGohV0GYVIL/i3kUuZeaMYDTJ33izT5s+fMB
CE28KPj9LLv/gL/d28Xx0UwYTTFaud0W5FA0Q7LQCO8E4mPt66q7md83ndeaxwJXzXBg0ShjHUsa
rVTblif39joMuuewh6Eb79yC0NBTs6JsSlGS18iaMuaqjDRfaKjXWvwIjat+CTuiWwhJys3AIQiu
EgPil9GiHdI/jw8c/tKWE4YSQJriOZ6WCTp6dZ8raF/j36lwY6vkRYswOU39JC6OLSIZ5j5csVGx
xPXJyXK1lhm9KEv3RL5oMKLOQCIekgNO9z/EIiQigVZTmwsW4sNckf+ICxtHQF8shR6xNzV1y36f
SQTEUdUyxpc8CcqUaPze4234VOJRP7hgjUvnlehuMvFstd5fEugAoipYvkQEhflzlhfhxuCSBbKs
BCUs47+uEZcaxjBuUjcT7PMzOgaWgl5rXUQhlSxmXqweJr7OtUp8dwTxsWnaD72k0QArdosDXAcT
331o1qBHsKwlYK4sRAJ9Ei85mD+pYLJB2KVPClvV2hI09WmH5pDjYkeez7bVZksNxFXIDoxeSBer
mmvhllBqolMqNE6pH+1ZzK1iPZN2J7Xp0lVzFL5fG+A7S7/jXF0ieoEegzTA9r4cqFcIlh29cvOn
/1hoHB8vJfO2GIJE07HIxJOXATjS/w20lmAjmAsha/p272ZGY89Un4mVTkapii/+j4loDf7Y6BoD
uAfM2qMmEba9clrBiFo5GtIYQu+Hmh3v2vqajODa6+9O8fINJm8EFrl95m1Z/SEijqIo0gTseTTH
pMMJCD56N9vcaGU6fLxB0nbCjgvLWMkrkIYplqA/rs5JnIGVfypEUzVz2YrBdngFmxXJXEQRHfBh
r+tivqo4lQ8kDo+1xZ0mVTawJptj5Vx2/dJlKbp/xtIB0oxfrhJvXZ/nH2EpO5y2T417qc0rey9T
NSa/gLEIS1gNx8vqoKHeiv2ugkhG0dTP0a9+N5V9jn4T+XerRkkRnauvF19jVD6O+kvxzT7kjjxw
0fPZsi8JVz0wNwkOEZZ+UPRr4RQ9otLw2knGJZt0ODDqUd/KTpf9uCmdp5lDA+n3nO7Q7cV9EuXx
6pk7NONPMG26CKqkO2R+7wroyl9P/a427GPlICARd4zPveoRABsKDG7Ok8P4vIiE9FX0nkMDpWnQ
3TZSgkOcUIGmj7BKFQMRdGtOVedyZwgqKxTebTnGZJ7SOgBBi0geFJDb3CJrQZxFQ58RMn6HhoY6
eaDuqGW0tsDtth+LnFSsQKMOpXXG06e7nG1MmZzpifzYjHfS48tNrSRPWQ0+PUVXwJdDpFPuorY2
yQ2TOro2SGjFZChBFep6aOzXy0v4wG12tenEgHSuf5sXyxh4BaUlLSUOeGLLZa7RZCMnPYh+7XM9
XtDR60Jk8VFIUGvab0foxQaK1zN7hDSTgzpdiMK3QRTml62AAbAeFvB0ojcurgXM9Zj7EE2minSF
pbWS20X9hsSZT1AwqiX742C3L54QQvOwHr1saOq7otrY9NGjbSZy9VHUlT8VrqF7f/Hp63cUNaEO
jEJ1632y+9ILKANkJpgUhx11ZJ5Wc/ypwZIrngosHqCpDjfiv4rs9VxCcE5LIeFn/rC+Sxa2FiUo
dm/21uukBCKmV56Q8ZnAJkog4JfhhRYXs4DTD2Q8S4Frwc2SMkJZhFOOF9LpR5cNvNVeK0cICgOR
tOhzqWFgpH3kUBviE4sWu8q7cdHXejjWWq3NX4u2IIv51z+Gf23Ahml7dhrsID1RU9C27/1DSq5x
p8KizJPRq50547HKhTHbiC7qMoqKvmzBp3DDZ7TcycKFxGaG6OBJY+qkM5cjAjGx6lpT/0dIY1QU
TuBDvZzybp2RWzzW2bAuUV01bgedPIo9yee4B/EU595iDrwiASJK90WisnaA+s3p593nBlJ6nt8v
TjKEpJi8I4t12pD1fmHjgOeiDdXW94OFiqGWIwPV9t9uZ7jR2sI2I6ECitX8ZwlR4fytQynnp3Hl
B651Cl58JjteDMlYQ4VvsNbX8CwvX8D5XgTa9FE6r46/VZajGQJMlOxXkpRi0m9bUG0sEVJiGLzb
WyUnlc8bK+b14NEVCUlec+P9hmff9i3kA4wXGlUSU/K4ZUO8omcf70iIRAfJq9kRnQ7VqK5BmY8V
iqTZ2n5sRUUzw5eCPOAUb0S4Jk6r7tppZMKpk4y9zgzdhSEyxQG+S0yG5twlKQ8bBC1vKtVwauHO
2heqPxI58Ms7o8YBfpwiGBJBCKTtw9zY/14uC3DXymfBYiXXAOxALLCQpGwg90hV3BC5szG4SDb/
y7JOGoKohdnE7dIjxBRhfDd9YWuAeLUGhUKHL7nTdW9oQPE4XXJ3dE8iT7l2rHYEE+Kq3pB3GGj1
dF3oUsftYVawp0kMix2MBB1YENTVukLcUTh8OI5nIL5eysfG00sd0tp5XBAomaeYWBs+tqHZ3NN5
7R6EkwuvaorIKHW6WaOZ9XBCcfMoH9prcE2VbYtjTKhSxG7ks8If+6b7HlH9xse6PrHqI5ECNbOu
pCXGwItpsBRd8KuN58NdDenVsDOY8gnaTSzZ5wRtb/xtlHkNd6R/SPpRJJvAJyMEaolRNAy1HiVm
w5trdt83ykx4+oVtHTOzQ6OdX8x7FmX/TmRHHNZGKql132Hf+57r+Ic1Q2XTSpLRK4icwNCC8Pdd
Ob9p+wQyUnjXHC93EfMMeSaaLd/K6gH4mVXEmW7Uzx+tGliBXCEdCPQ4xa2HcsjLQ7KJAz/On32o
Ze86fpWO5KiZ0Fl+eUiPRPKYxogzmtDSBJyk1ZBLZ3igMCwqrvtfHpteMkG2rzL5f2rF9EI1LjqI
sIF2ZGWM4vOu+ouXKJsk3GVRW6U0p/7Z4eMeX2O/X8yk70/fKnUHd8DKRBtBvJlWt5nJRCWi7gAw
3vIbFgp8IdBOVk81qKBZkH0JAy5XHj2oOC4p3xZ1Z89FstmN6N8y+Jwsd/xddC+wx/vUXgsLASDu
lWsp/vS7WDHUjKKoHra/KkSG1Oc28LpqqPHmQPzso7hQD266OIEOc4IYqE+mXaR9ukyMZCqgRNvE
00xLsNIPA13HdR5kkuOlcKXGE0ZxK/Xu/5DaiNIeo1V5/7LeQGk6M2oOyvbBOYec4e1+VeyZqZpR
oRZ35oWPgmPgZR1rqbHGxxGi47PwUmgOT3H3z9ocrH4CyDDbZEwrJetJZ3SAi49beM1JAaQhwVVq
x5BferPgRa1Dtd+r+xNZAlbkKeLalThfyX6+vC94RVlsmF4RXnyKAL0+oobFthVu7SItbV9KU9XV
LQ3uYYHElfw2RJ8VzWUPxcoH/cm8ciQhZltFxYdEkB4SHpjvEfPr4goZQkx23jqS1ttTYnUDOP2F
FR8OfjfvK2ajQQPKbaW9KDEtzTENyQGIwhmnvoadjJcHws6cziuhEZRB1vJnapX3WkzWEF2PBxHJ
dZsFM6iurKZNhbOuVkS9KcvuN+zElgfAQ7XPlUQIVEKtwUa/WD6LE+NyklaWDaybUpVDyjSn26IM
OOqT5kBvc/N8/ViW4yvwOGc8YXEbD7m8xBSNPd/i3jZgWf9epvKofeEBOJIcSGee9p6HoORZDR/D
40E2IbvqpU1gjPUVqrccgnqWLwMUUAHyWlEq4evkWNN/xiEt20Ck3w9e0h38lMzgMyG377QFkSc0
fOBobnvw0U0IrAoi9fGcQvjfnfst0It65wcQJ3UvnPVylWKRJdLa6pWYkEXpUkPg5PIo1B/Rkakn
8QKdROuhU6da/zcpAPGscBKQPys9XsDAtc3aG0/zNlI4LoF06IA+K/Xaco4wVaTNc98dhfDcC8Sa
8kG1GRYkIupgvKKMn+8teq76+iJ5OsNHcVyB8DljP6hafxxrth0XxOhTO8Riyh5HZoGLWrp/p/tg
TmAEH/aW37xI2vJ40mRqV73Rf+IRClV7dFSZ1vxm09tfestJx1NoOMAxKXpuJ/Txkr2No+BjbwP6
Js3s3HExSX7KhduSXuF023N/50NjTkb+p+09v2kyKkUWXLtQxJGLE0ripXMlM+NUqqket+Zglibk
NJFqo7vfWv76D5fggfWryET5Isw9RBq0WOaSEl++08umKfhW/Gi5fgkeQuZDLqS1xXzPHdN/XTae
ZXkGflxHMV+Rr8rC1GhOlnEQIfe+VFjzCd874aNgXPEqgFKCKjkMpOV7tDo0puhFRh8cNP1x7TIq
pfVbEeaRi2JSVb70oQv2gfXGHNN6ATMMEWgMPAO2Q0gg1wRbzPZJHRVlihNJgf+IOsxNB+Z0LKWO
7t1W3a79GYmh81XcI6t8y+gJKeEX4XxwjvtUGKhqRlta3i2O+A5LsBAOyJKZ9KceiT4nI+xMoCd/
VeQmUxff19jPQ9nw+yrAPOCXbjstVmMOopjKKFHBYaF3qyd5Z6N0YK/y+KBckPwYIaRPwS1RYOqd
DsmoUwNy+meTG0nJxRzj9YDoIYjMWliv7gsmATuFm8CWSMwIlm5NUKfi0L8RwnAWPrMArzGBtsBo
PUUhRUu6vrIyL5USaHSJr4yCKBAZHd0X23i3u+r6Bm4XIqqY2l/+Xyb5qtcFqdsYaa9xu/yvcKcJ
Dr0nvuUES/4gqBP6lxvIifZf9VA6SbX6WK0Qv9Pnbnn4sXyhhJ5s0o6uGM6tOQsWKRkYLrUhPP/8
FH5KL8mGpn/ULbjp99A1ZsPA583m5k2x0bNjzObLp4cleNDr/lCTl6yyjxztLievbbAYheaNhw0V
BomWAAqEtkhBtkP+WpEYMHPiinayFmF86CbB4CCtteLXZepj5neW8GN4nz43SrIJbYLRF6cRokpQ
9bn10w/NU0VHOyIEBur9oZtbPcpi1xfAru5wKJ83WdoGHfEyMpdfCQ3lvtwShuKaQ2H5PIn53cAG
KPkQ5WAKCWEqluq/zs++biSttvsHh8ofBd7l212fqqJfQhLzWmfKaMs+63mG0+m/hhIuwXJpFb8F
CXP5VlUgR9ftMm3STqBPP9t+VjOFAOlEvVonYzEEaQ3YOTmTxdiGiLa5kgz6UWKumn02KeOrJeUS
L1+RThTQ280b6mxXDb6oRUehEceBfGmatFnR0YG4YT3+C+pUpQrZR9YGFKFnGUn9BZskQTkvI5uu
+IjKyEHBXXeh+Z1C/GDgrm9k7jNkKlwtwyW6LIOR157bPFFB/JcTabBaAXd5/mJNe3lL93LnNgqu
qNdWyByb3RZs/KuVod+6JsMNFA9CcW2okxB0hMfAwMqnrNcU/cwYjr0yQrDb4eTgwgrzWJXiQcDc
Yhn/AfpmfWpdvLDPFT8sPJXuWAQdcUysuktb1tOrm79+q/Xdgp4gRPTfob3bmMgmmzqtuGPYbQbD
peep/4PsDa9HLzL/lNJn7qHBnMFWCpN9yibg1GD6LrlqnhG3EZ1bJNqEFHY2O2n44CMJ7IR8lYbD
NspWOYRfvR7oFWRpSQtBJ/fR3raZSj2t2ywmLF5NKXBkzTJnZgTIGUWCmCVME8dJ/mWtsiKlqeD4
tiWeyhQFIdRuxWWsq9gLARlf/1qTwkaNv/rVWCftJ9s5KutQb8VxcafFKLnCqyusHJmcZQYpgc13
sDVYCz0Goo025DjVchYciBBVWK2niun6JvLh+RwGdTAPJOZa4vISAvhODq7bmrMMoaduKWYWLOa6
0ZI9FVEgqSkqQkOhhU4ktop8LGvrVpcW8f+PDts2wJo6FlBUy+7HRtcj3Py1Qs1ljGckdh4XyKO/
8e4Sn++jzbLQfbYlq3LMhzhIhTyhG3aOO1ZwA8jfMokms+ms6xKENK4hndDUnZhO6wa4YffJHMEx
Gs4hCnrcq6SVstigd2vLC5RoRWoJQCw48CXzQSNnIdODhVSR0NwY3Y/VAi2wBo0mhb8NNgxvUxa+
6gkhpTuTef3n315n1YoDIItywaIAIlHSuESAA51DuS9hB6ELnTqrHCCBN6N7PkHRXRR52cT43QmB
SOA7SpcNgAgIcZy3JknV42LpOsDAkULWB651WYWHm6JGsqYtqmXU+hCVt0sWS4krAXcXZM2Kx+cH
qCrfGFn+/1541v/GPvlum8pHj0Ewm202mOv9xHnZa+hzkJ7LASXoC2Dfybrhhxnd2HeluUXF4KoV
Eyg7RX58NZjNMOi/xlmkqtf+dUhBLAnX5ThOxq2A3k6FmPeYjFHcep48SmMNbShPFZj5sYccwTR5
6WcLRWhAL1Cz54GpI3/MiK3dnbEtgmiczAyXZy7SdiRjIwTkDfsIMmUNLydjtfsdZKpow+dkEDyW
rCvpClTD6Fd79Z+Nepklq5iA8bCFwMvfmS/zvG+X6pQb0zy3Hu2hAPky8BpQejfk4EKCMVRp5VJh
9WkZvmLn+4TNpDr5yvAlWVLBQaiJAMQ22U2ziuB+ObKDXicEX5uVX1HcOq3U/IYexbLLovvWCNYH
W+0QUUQhPvYD2tYIkG75P712RxiBHYLDjjK45TEPNdSMkIH6xBZzd2DH46qORVPQX6kcWa3t076K
sik/2jhIRZkeg3R+1PeBVRZROs4jJ33WEcyCVT4FuPmvmPu1GDBHNldZa5zbxuoO2Q5tD9t52465
5sqwTrK2j1OuMpTpLxNNWPeUN+ZkIJhBFcni/ByLIlcQO8P8qEXNVA0HmZWjBGjtiQC23wUGw6r1
DmZ9wivVl9tFHGo+dSVTH/c3nY4UG4cdoh/6OBzDquQwqUR6u5toGqipyFjFV3oGrOaeYS8Ms0wB
mKXp+GOA+rU7BlI1uuU1wO/oNuRs371z0htMpE0FztiBATknRs0/TjLeb+qpNhDmgkwu9iy2c44G
Ls3n0/Fxn8CABo88l4YV/+BVJtLFApy3oqXm5mdMFnLuELUX7N22B5ppGEUEHX7rqSOsxQZJI5MJ
YbGTuTf7uy7FJ2TDlDoI5yUMNKGf0H/FhUgCYtbkdkTvnoMy+I8+DgCltZ9vO3rpMqPDM0jzUOv0
lyScdbJ86Y/InUl8prLyybvyfGnCM02BD9+VCwEjiWYaCEUwUs5lAZ48/b5yfbylEV5xqnb4DXN+
k7slZzTzdFMjmU7FAak+fxfLR1+jADOM3h57PSa0zwrdj5+FQEdV4yk27xnwd5r4rBK+LKPqcFXn
cJVrbyhP0q2jvcydDqfDHkfm0f3u3Kogm8tGrJw6iaDCy/srXsyRZfpKmU5C4Kl7OPen6F9lKgEo
ZTUShWaxCSe7PQcl8P9eZMmcBbJ8gHedtKie/+bgOTPLt422bpUdnPdT07Cax76JKPaub//wwxxu
oQSavcIwbTQYfhHx4+BX7MfyefKKNsKTzPnAwhqvIriX/QC9BDy8Yz7lu4wGGFyEP8CQMYVv+SAI
2vvjU9+XpD27xk81WMy3QoQNSLfayahHwy7YY/tsdiVUX6TLq1TMUtt5vdwELBtn7g69kb+nUvHO
aCn8YGdytGiL7S75KY4vQmrHAXRT5ygJU1vnszrrDJCPWLnewAAdiX7DqV2DN9JkePrqBQA3w1CP
Lda7zatQB73eOHnv4quvCc2HhZevSGlqiFDn9Z4GUTiYUf1g/xcG5rTdMc3/0mpMuHCxz/Itf/vT
qjyaGRCn0cvLYg7jgNibu3wHPuvK9HCmSirwJeWj93bVPpNnWEn4Ki1pAzT0S3zdl2HiCcrgJCVc
lepyus6CMEApXVVGpYxEr3jSjtKgW9ciBNH3jTagV5a/EBVZwUKTz+cCJAOadMoTUrrElMnPxhnS
I0BcpBjydZvrdSSRQA2GS+ejaDMogXolG3CG1d07eJAy9iw8AYqwj5/cGih0bFBhexUzw0a71jK8
AJTR/AI4xN7M+nBmo7zVf4AsANGO3v8oeBJftRo2JWyx2khHbdBpvbiKgdQPuHVnVqOArUIgOYZ0
CkDCiMKkor5jqVdbii5pgZ2K8hP0oIlMn3gR2jYcCyucBhodH9k2YsMIVsk0BGqhn2z95+rmBrMx
NA8zDukbqkldY8UnjXSydT3OqqDiCaoQpPJ+5EpaaGA16piC/FEs9wxKwYj9GUBVzo5IYNNdm0R3
u1+WILJ0dU8kgoNvHPrQWGO0rvxT9Gkq9K9bgnE43zB/V2RVdF5r8TbzLik7H1MS5PZu+J4RR6FA
unj6TbjQaNMHPHd9MZFwkN7ixtFksJn+J1jsdgq29diowzAfc2a3sC/pVV6axqjRZtXWUAt4EEF2
UVRWsQ8ZypBi/KOguTvJIHBfifQLDx2LrsjHiV3e3M6lDmx0twgar8JwcCED2XM98HBJyl9cfdJS
BYA7UbtQLu1xJKkw/ImK7jrse0kT1v7zRf9hnKbPBZQLULt+FKIcSlpVqqw54B9TrjZ3WPWQQG+b
Ws7ydlWTrw9HcxduCsIIX+nL287lWawW5+vg/9lIdtCAV7RmNrhrBzB13fEoBgowPtfOu7jcnovM
NTokTgvTyP1sfyhAq1w0sY0yLnqbV23GzrrOTUqzydQ6fbwi549L/c2d29uOQOPDSQ0AQBn/CZHM
E433IWb7RzcsOzBQkBJWtkt6A2NnAf72Bymb/84sXreXx20ni+bHx1SG7Y/H6hAP51bx/n5LHyUH
UZ63xnKS6Rv+B1qLR5Z3mPSXoTDpqi4EEJoYaA/uJlSphfi5Wh+b9aCkY1MDdAdijoF/CV3PjkpE
jwnO0ULdzdJaIvHVZWxqBGnqbI/jrGJ/RTcYEYZdCThdsbmlesHzSzUjwjs3L5dXmwH7prTMfLKf
sfWuP3f9obVZkx918sNapEaCfhUJzyigg7QluliZT/muJJ6uce91rx6QhBoF/DIeINHLZtQCiTgU
Jx3QNoSg2+qJcNtB/zbMeXSkFE924XTkmUUGroNZ6ocqgOX0e+HjP8Ml/kcMdSOV4aZPi+cFenF0
+sL5iK9a5RWddmwGasBHBHk/SDU6ihPJvgVD+16xVkvWldS+HsrJg8kQyTgZeuieCBywH3indW7K
D//gHVWqA/7uFUDLTrF9LN50M4ifDzKgbdTtPxVEsZiuDcExQz6TBQCWUKRq8PIRKt16KRp/llQB
1qKcB2Of7pjnY8PvhmHWOgKcYKPB6z7jJ+fCpWOodrgMfLsPRYYzBeguL7xPfS8i4ioYb+vYiHLT
99I+GasqbnOM3/FD1vy9u+slhGB8ISTDEHboWr64t3TIRdAE5P/AUG7gIjAnxjYl29kpi/moytDz
viGQ/CNZxvaczoL5fvu+TQolY+CEt4X7naG6/p9uUCGsCkWqEK7V4/jEb0JlsoqhWNsh84LTjveP
mdpXz60eqUCB/sUtq/L1nsr1r6esJXytUmPaSTOoS4bwHSVhWA6MnOi25WdPu370KnczfsFnv03o
eQivZ46YRvCv8VGK5+BP3hwFmmGVZTFLJF8JyFME0OZVVNmTz4oAjzZgHLbqaanQWAh8yzt/tQ66
BYW0lV/n6c51fGynilgry3DBkRicFRdslN71kWjK6Attalc6u5rfe4x2SXW0SaydErHOW2wUZmIo
IIKQt+y4+tnEbkVgG8DwwciRtG0KPCAdJZbTykUfQ7fvquiIKPo/PKcqz/hSYfsGcfbcu84+7vqN
BMeyPFhg3rBRipPfex7AoEEOnlGiotVU2xodXxI76xKF70EENJ1DKHfKQqCe4XoYAxcE5+CIQBPm
HQvKwJF9I7yrQmlnethjmiHHdAsCabog78Be/MVSvtZwZt6DJQDw7D3rDI5ozxzBBNj72JEw47YV
0VzQ6D+MU+/0ZQ4c+YNXMdRTrEDE47ForO9oMvGRXqpX6KqV+PEJKmhiFO5IcShgyEjZSmsVDv39
Onu5qSkYIs/CRlZYL+1n/t1L2jf8VfcvvCXyzUy7R4CIpuNlGQhH+VAXXf5/pQBdxyVwAaLuN8aO
gQjGWhc1Yf1mYOfvo/LnV/Sf7kNmXDkutM8njFT4YBOV+dwWs3nQCsef1xCibCnJeIbcgYhv8mys
Dp1oPAjc1+KWhABzs5XzmrR43U74NFTRkblh2/vQdLC4AHc+QHCrt/tLWCIZttHy7kwNM2cMp5eb
zeFKH9MvYucsFYGFk/mj5/weWrSv8bUOEzwMdoBEqvZuGtX8yBv3HZ5GMdlSTozx1SYt0u2PzwhV
awAHWzpTRiZ34at6tomYFtn67c/Fsqrw9a504tDftihUECxgxb7YRD9gklL/9J/picjECiErpQMR
z4ZSfElZaGudMRd9ml0zRBWlYJvTL0ak7uuGaIcb1dgqvv3Af7/OnsMUnPJWcCMRlERMGsHzX2tI
d/nnXhWvBy2MYZkMKxkRDMOUEl67efT+8QSIVrhe3pcgsvA/s1PL9yKZJpefecIM6NGd1jQFn6Tb
nEZmfgq6FKTCYRpKKcNvwmA3//8ugbhYRkPt3D6vbsVsfehhd0iAoWS/lCqECvL4AW3lOGV+iAaN
wTt2GG9bX/+mXfATE0ozDEVafP9DkIpIex+YrdwBMO64yh0US2iYea80MuucEZ5zxtNCluEzuEyX
xt9+85sFYS09wi2EgdqfVXuXnpLWVavIiRmF/XFnDTszxeeP3fAywS6D5rbAkx5oawUzW8WqDs5h
ldnw+WNSjfHAdxzX73JX8GepUg1mwaXpFJPBECdEQpXhWev4E72G8vwFKItEa/xRdb3Szh3zFalp
ZQ/o0wUTXOmLJ4EPjx2txIGR4a7k2Xa/DL2Y0Ggmu9X/nwSvj1bXrAD71hZhVmtRtLY+GhmrGUs+
5TBbmEiuklpY8c1lVX1ofpqhKqhEIezVSKTUBRPsYdfO/4xGb6nO3sw6+muoo2GLoeBZ+H2MLIVe
K3JuQBGSiAfdW/tpAP2uYgZr2DwK0CX6oPw+FNvkd9SvdGuNe7G+2feeTo2TPCmaGAUu7WwWepOf
WshRXFkvg4CQRfoeboAaYIRrtAIkF66akKudDi2EqdrfrhmoX5FVyeCW1iByokeWjp24cBdgsqHV
IpKwpr+BW+4LgOs9l/HWhs94ZnY7uqazaVGCFvnPL/UYFPEMs3S8CUynX/RM96KO9tFAcZ/w1G84
sZSthF6F8Fps6jNnrxnKeUKZKZ+FJGBAoD8l2CM9t3Mt7pYtLNFT3VaZIMb+X+2GPmEtDysTS63g
TESZR+bFIfJX4hy5WetptiLFks4CvNusmMCLVJ0k6ZWU/ehkwudsShyii0WIysg56qr1UyoRJj+/
j6mROPM7H7DuJfURSlRiPC1xBfH2UqNg9yDXgS6QFfvEei8lxzlyP392JHpgfhN4n6HOHTCyLKcL
zbzr9Wj2Y9nUhYR7KzDNhhNJSHy7Bdx5VhnaJvF2Tzd5ME9l2FKJc/X2/FQBD3XpvgDahbLq9Jyn
PZCPm/s6WjU7lcRGXn8UDxAtI19Tfs7rxL1XdKToiouA5KRA9aSCKo3ofIqurjVsZJi3pb5n+mw6
p442Nn0ABlhvy4zisW5nC3LF8NG5ftVWrmcKvrGv9IaIB4XB3UPtd05/TWHO2YOFZ8n7N6IS7Sdm
QTcRMauVMQ4yuNsrfNhuY4ZX+YilxAVHcyCND+Li0WeJw5+pu0E3PfC8KV/NhfhbG3wRE4r6FWE7
lHJGUWjiKFYr2KmA46tiwmZwRrR2mQKHY5wo8NAoLT7tmnd07pT7ejI+hDmQ95VCRnKvit6rWAbK
I4ulcSMsPyJ1XobiKNw1ChpT8swiFONaUtBSYT4JEEDm5KoVWvjKbwEzqSeNyEmCeBoNtfNH8GwQ
Tt97j+Q4H/34wCve0B5BRLckKfze5bDL2Y0n4QM0KLsuL2N82V6rj3i17sQNsrpdA4/zLCZoVV01
LwZjECJ8JbhWg0e5ij6Qrj1f/Y3/FGy9CfzvG37tJGjQun7pRaO5cTIgt2RXAqns3xK/7I2jom5K
7Br37XGSS/IdJFzfgaM3RpVqnbQUvJhn+ZTkbeeeqA5Ju5cQqgOARY0pvaCjacw0Lc9c154gnch4
8QUqExGmaj+2koZTiYy7c9lNazcNMBS3R/If8bwpm+S1uWX3Et6rpA99OYF0DbXvrUAIegT+i868
zOdSPJtdnmsbBJZ9Y8onD9IdwIoYZTIzjay6SzgmWoRaJwlTRmHmVrCmIcir7QOK1i2Y/WVICr8K
h7LLoCpd8nZruLtT0uKyS6mXKJdOnqLCxrYnVv1DThfHvALUInW4QftemV937XTcT+0uRfqhExom
FV1HbTYd8WPMw302UGwOO16XIg94mouCiyk9of/mdAOTWyPtNNnwml957K8cw6On6G9Uqs7OtTL2
DjVKoEvvUAO4/a7N0cOyj9knxj0ec9WKzldYVHaJF7X9/BsdXwwLFxG7dvr9F3c5Z0ZD4lLXrCEu
HeAwy9YOXzUKLC/owzaA5J5c7nwYjDTPwmPq7IAxrOTpNKWxBCwCgtrHPPIVFzBPv4aU37DmmFUA
36qDAxi0AW8ak+b7x2q6ztgjd1usPwnb8vUx7AfbAbO//Ug5IcYLyDsZVqfMjD7Z1N6/aTYWRsiQ
brG2Fu1ioLjezwWqOF/Wzz60Xy1ewed12wbzlNCWPJwKftk4JVKUmf02pzhEmKZhEQjLRBWoHBgK
LeUjp0IYpjylXTR5woL4U2Z9nORkvm7Q0Jldd7jwsgaXvGIvxlps3siv8VY2GOlR1GhY5tnHw68+
vDarhMcO01ktgC6ayTup1hc0E8wgWS/goGNjejm1OC90g6K2ggGJHHlPwFs81F3nwzBmU/eLohIS
PwOdJHOQGK2WlV8SbqZky4m06SxxvU3ejAXU5C8iRXz7bF4240RxvGmxUPVeg5/TNqZzD5fIEiaO
0e1PnLl+oFkiSSR99UpMeOXCaQG+PbyR8cVLh6eh6f1p36Qaw8XM66Fyl63XNYnkY3wQMase4FvM
VAOCb3iL1L27qEDKM2UQlVWarZuSFlpwonRBj7TicVEDABuawVsbdFvaUkhMeUC4ppACusDK9P0l
RllCUFuVH9LfYLyR48mqWb1TKrscH3QYThbXEj1spSPSfxDLcifpq4m+bnZ94TZ7+R5dVsp3z7hC
QgG97Os+e3XFFEgM+7EOu/OMi09gqPW3KqvW24Zx4pnOR83ERTWfpNSeb3l0khHmqsHji/gi44C5
uJt73AUZqxBT1u6pwpPJeTXx/5XeXIvGPnYKLyAn+//3UA1spDU+UpHdCdz266mQ2s7QMGRo3Ady
HueVemhryaotcC5RKy4YyaVD4IwIPRfXvrxH6Yf8oSb70ASmVof8DjxhG5MtATFer+9GcEVPwNkr
lS9q248uDQfkTPit+Wy9gqiXDHswkpL4EaXnUNpRmYZ8JxTajC1r09vUs2VmJwkXdcFJZWH5IcVM
JqhOdcWw6a9MFDk+Ej1PufuMGEtKbCFnIMvqnMOuR3q0qniGb5nCIeoB/dzVM70kq0eYbC6SkPgO
i1KZoIPU4aUkVL+HW208oeNqtM0xHrG7FXJK1bHv4bsxsUEIQiVPySAWrw8PHio/+lp9w4jaaiMW
MIyi9LWtsJkLv3rlvUOsQ+da3c1wcjFhX7hkuT3DZnMsQT3bRmeS/jx9pqliT1WjY0dftsexZljN
u7ZTC9rpDa5ujWsRf1MILGslrYGwbhRx9crnDhGj3Ct8MNQ2o8Kt3KhiwrXt8HLoQ2sybP5httns
5Vb3QesyuNdhThdViTRBo+Y7sriJgKB/k3rfEQ2RtP5Kv0hjsLmFHjK6two8MauFAXA++64bngJ4
DC9WOmioGB4JidOe6OAXbn386FsRtXuY1tbwOjNrJNiAIN9Iu3H4uw8psOCFPc+CEBt9y8EYF9nx
m+pqUS59t6fBMeoacB4WfDTYxfEUAC0FXDILxGvxFcEELw//lJ+dkBBTK1YcRdn+VlK2C9Y76j8V
30YiWqqnKLZS7Y5svfwHvXf8x88PjY6xOp1TWRggnIlt5+im0IIFpNm/b0IN1DNQtjbVjsIZJFZv
DyPjBWFYk7kyaMHS1/sTHW1cYX0EMXP3Oe5mI8To4kyPX1/Ny4j4dDb7nUMB2Wc74JH4s0cRjBSz
j9ll/2t/2mId0NRFMidcX7OvFHje1UuUf9nZ1VhwLA9/hOe1hArroOm8XQFJRScgAy54Iibuev6S
vcRb73AGx+PILfJHYza4Wy4/ZBtc64qeHK/n6jSPC/PbAyhGj9/yaZMwam818q7hMNqUCWyWeppX
ZnRwHJnV0iYIaOb3bUO2RS2mFKeDtT/5cOoJq+k/BoBfQApYo6+cFnf3vBTKqPKlc9+y4yNqTCib
jS2RkK8yhhSK68ZFUVZenOgocVdoycIsN1VVnwRyga71ctIty3Cps0QDQZsrkzdrW2sbojXgqNt3
orrxAK+Vy7pGGJsHgWGbhHBJHtQsqmAknAkegT96/7XzKpM6E++89u0GdbBmUvrvfzq7+pAGCGSS
GCmtRKJRhyroGXJ55FcR2q6UaeB1L5/lRKjoh7iPqTKULsYSBg2quSeNHTJ0fIG8JW8DShqWQoOk
NwSIWMuMDRICN8/iEBgVQl5NP0eMrkyryqg2oh3uVWtuoP01hcNG4AXgDwbFsYOOAeDV0FmpI+HK
ZNqt+/LFHHK+kiEnc5Wz+69MZ7QMtNc1hrr53XvhR2aR8BXMWns4mlwO/nZ1QmQ65JQGYbNTZ3A5
aTagjZPuSqwz0zAyQMxUOM8rHsFgRVzTkgRMoc0/ejjFsE4LQAVlAJjNgq2R5OfH5OZckZZcgU8T
Ckmlomu8lgrLoDJqcjRJk6sHr1LfMrG57pntb99iU09g2X8T+h05xqrNfrECzr4HPD4be4SxvxFV
A+6OmkqM0yNsUnQ7im+rI5nEhGhcZGIN7oaZc1x41NC7xl2GijUFy7drea0tU6qAAWldI9j7UOqa
JeLfbcJ6firzUwaUYbp2JkUNdFS6lGIlGwjbKKqkonRH1hrTcX0JEfdnosongq8bg1vnAU4DrX/S
gThZcPJjtzsrJDVCUs7vyANTi+bTFsvaHX1Bu2kVdz6lixYOZJWxg9zafPz+dPtRTfdu6gzlGCPk
FGTyXC6gRnTql81WXWFQq1OLNDNeTmOfRKApdy0zybM/Vsy6u/hEU/zbwN7DKndOoEEqx4PYvhSx
Wc2Y55Ej92p+K79TM0YGFxiSr7MhC66oaRJjSv8zjORds4q4hpWNYnS6DrGJ6vGYZEl8sfFF6jxw
uzbNosb2kk5Ie6HUaKLm4u7t+949wu5FnWLA06FoaPdQJ8Y0G4Ox8/eMUAEQ5zME5VJlu4x7tgUy
XQWZA7LU2iD4PoATjxMeOlk8I/hpC2A3AMFHlNEoY80B5RZQwNuQQXJLb7dZr86DL2wP5qWd4Op5
Q//ptwXqvKhydNj4YB9pfJkXvm87+HQZAOk6eh9qcU9eMwO9ZYK4Ys4G+5lCJmwT0+ERx2YwKTSV
wsD29clCDvpAwoWofS60QtxPiyT4RVulnN9OXV1Kd62bXGoIbgNlMtY0liCTFKzKWm56lYQPM3Kc
vSQpo3p6oXhiY3ilP85yFSC70BqcD/VYDKpNfitF5NRNHrz4r6kv+adgelgLrXYR2UpsUKsBRn5v
HJU6OlsN/z8oERYNZwc1AyGlfwwQSIj5jqejUcpOmX9GywbC9tmmz76jZ1NHWx9d6IimkY63qpWk
iozOewTuS+q9ZCosI2/LwOlIiawMHMWqZuYyrQ1SLTr58ePc+SJUX3dfkfCunkZl/NtkJ1p3uE4k
SUqqCQqoknwSoDbgOXB1XZ8UNvMu1nIZWnTxEXRgtbmwP1BJltfKpaTZZktvdL612UqO3iUwMp6u
2n2fboVONxsP+RfrFsDU+OlVqQx7afUDK1YUFziqhSmD3k8LGTEW8RI1wE+7NLaPzL7MnlNY88Q9
KKzRzpa57onHMmt8ugovgAQfLGwV3W6FQDjo8ERBFUXvywdxTZXoyb4RqlVeCJveJd22fgGnXmQi
MgZ2gg0MfGgwE3/aPlIZwS9WLRuanpbKFpwrbkZHvSWxqvhWEaGpYyV3a6WlgbKF+FDaPOpeSs+U
pZ8ZJQwplioHoH7JDBEku650PzSOXRr2WVLtnyv8X7V2msd8+V3W89sgKPsFk4ntGexXvjY9ARa0
xeDR3Tdnx8HQWx2xdbASn0fVMM53D8hrAKleVPn09gfyyxOzPHgtPlLmlqyEtXWacDYWuH/DpK00
Og1mdV/hYjFls0Qg1LpJe2TPLe3Oi8gTO2bhzrzuwiI53bbRnCcH//9pKI4WXN/V2jcgU+wU0myV
35aWAKyHfzC6vpNG1Z9j3Il8NwPrhgZloZhowcBYwB2ROODZZuN/LbUiPmSbJirDK2TlLtTy0ih5
jv3N04yHkCA+dHnKSKVppmTfcsAUcPkZ29WDqxcEhdQ83X5tAlLjQfMYOngrenC44Tv2CnGM30Oy
OkwToiKx6RB2NVWfMqowq9BzX5ya72J6DeBWQ0VOWzvu//Ak/Ytrs9d6F83nsrvcfgGfsc8lQ6KP
6PdoNXxeRqx2UqjdiKQmxUHWYwvbs9ytE+//jyqATcMPrFpMCNLoaNzhGVIh7sFkhRvsjvLyVjYw
46uxvXMz6fNcFC/gVdPDtzb5TdIRHU7f5f9gro/bKSe+M6VDsaqP5WzSqsGBZbJbKQvIeZqfbovV
B9yGdQsq+v1uGfb/LWLz7NgEWWHAhVr6YJUmnnC7uOdW/hx3dBPZenLYeD5T/ug18ZV970RtZDRz
WjGGux7xAOpWFxo7V+I6Th+37GACGAX0ag/hYKz2Wrfhf+pTLIqKt3RnKtBQ0uL5NKiAzZagqG8n
WdVKNRTFoZt0aAdw4Dw3WdM0GfSZJztV/ndEC2vK6EhdeTBEGvRqSeE4jUlKFjUZBywOtg/ixtlJ
Ls0czXYZyDbuCzBFlmvZFKvI4KTZnTSTGFYc62/GcbhY1b3YYtNL0dpPQFsheROVFFWup2PLESoi
KlhtOnKcbSiw9iN1rN4rq3YKGBjuSpsrXxF4ckjnvnbYzjKNMBrUHHcQZor6Br5uY9nVQqfY7e/S
y4OsDM2NZsYfblPsft1ScL2ir55XwIzoHYvKCvn6bimVmpyu17T5YzCO4RgdwraqBlos/m6/5NIA
mw8vzwfFggehjySgDdGcXBRPw3rFzAf40urIol0Ot2JB/JrHdR8B+Z0ZnlGg4rOuw72rjWqiva2e
n7hEcktaYoW7zzzKRM3toB6zZ5joYvo+AV3+2i/yZvx3Hd4KFdO+/Upql9GMlWjgJMWicYgMCojY
2og18lqxArTqFPOMPdNi9WleD1NoNTvlwv59tFj3mccG0/8sPu7ZNCDHRCkEB/I12RQ+gXwV8iVs
aM8ija23WV9lNgSEIXhdXjIRaOPyTaCNBBVBwUgquT/f52B/7NOoO1QxOGy6jPxlhaSYaBTi0c/Y
MXecHgLc6xDXIt7+QuAOrOBEnW4BRHKcA1BjA+VwTUZ0T7F5u3sP1KBuPQmisZQFuMLGKKvdJTKB
y4T/1tN1RhA6RBqlkRWq2nekBrukKJtAxCYcoKMg4fP8YoJIodevfsvFOXgLAqcmp5kdMnD7djPF
Fqi7gj/RHYNweeq9yFtLOoyAkqR7t14UZUuykQJlhe9S++RpNKnWCjFuoZ9MTPEcCHaZupOM2LPc
gu1m/ixII5XZ7BKwsZ+6EEHuAh71oDCvYdzs58FMbXmvlc1W1Tap9GK4s9iLY1gAnMK3NX/Zqy6E
Jz9W5UIbma9V1JIKJGdhzf69ZukiWB5G+cEBNM93AjAebFI5v5nhQZr7XyStVPMdtuRuD7u93d6X
Ezyx5GP2rn/BpR8CiI+OBlt5qyzca3UbEQJATRTMWifYqZFO8EuWeuk/seCfAeJcBHMMh9f+y9h2
bjKDx0hVbp3QTol/QOXC3tUnBn1Uuw+klFeZGriyq+wF0qU+/NpPFqnv3x3baIR0gy1QALx5pVyk
Xrw+DctWlgyaUkxQrtgyfkCJ0Lf7+xjCjqVsJ45wlNdz2GFoFEah77sk9mTWAyWbLtZI6w5VLP4v
WLRHllJa3GA+TqkW7Ml5ewZSbu0QySMbIvqDOAZySBP1Io2i9l4liFufp+g/gtrd91N4AIBgVQt9
7EO+GjKkS2ewM5Va8IIBkb6G6ZtxY/rZccELoF/wGx4E1FkpSwhUw2dnTjBCcgarQiXVui0roar5
Daxk3aplN2UuN3REUSCmxdwJnzWee3Cy0LEieTWr6RHwvzXs/AKQOFC9s9sT1fNX75xGdAQw8piF
PyjqkduYgheDZ+Zv/prb6AGnb5j5NkOMwYGOA5RKg2SuW9jj0u65wHuBFqiE5foaITWzzAEZwDRF
hmG3hNVQaLJzdBAZ7dWBmD+Ymr16NQMu6ZbEozdxbVQn91L+gHkxe2LeN5spd0dSIg+eA0E2g0hl
zV6uFWPVzD1Qsf38csxBZmSE8czAEoPQ090/WXdcdGBfrjH+a149/SBPEsp0qpuaOLuSd2GlJPTQ
ld9TOmHXaUYV9SzuHxuNaDnlek1tIieNe56y/He7SWr3Wfl+1XdlscF6y5D1ebwTZndANuWUvz7m
9Qwm7SprctLc4N3ixfFsVC3B9lzZKSwNq/uX8h3saG3syC38bz7zIAT2aHq4zyN4sbcm22T//XzA
gJM9QYv4VO2+XIxaE9lgKhPTlJJHmhmqYWbtNBs+W0nFtA3Rs4bAMwcdrY6rs+LbJH6JFnk9HWvw
oe3wqsHh094+smPR24d/rnnFgWhC3Fs3O8Iy3Q1r18Sl0SXN6FMKum3oHqNLI8pHEM5JdCeoyly+
AELc7XoGU2bRWHCnbwa/Nky2FJLjtxM85iwQTgfWpZVZF4dXyvAlV3HKHoOW6JASToThXJnhkX7n
yw63dnj9yi7SfTRoBiPJ+w+91YVE0l/bE8GqWksKS0jCk2LebCrKhgGMFA60/R3CBYW6OsBaNFMZ
hboUcfmUsFFCA5v6KGeEFl0PomejK7xJ3S38YmVut2NT0/TD5KX5i35BdxxeWMso1RxFbC/CR9TD
scjZxXd9CGNuVFXb1phqsArNWDHcSCHRhNJDqBVnx6Ti3xUS1nfv7VbkS2VLeN+Lc1799Tt1iIzl
6CRP20MLS7TXEGkTV9mWr+McNCwqkSZxeRaL+NNaYDs4lAOeB+6QKeUvCyfeKLtUXv4YlIHHcuvs
r9ahYJTg5TdhBLEyBhV43j9CR8p6uI0dVecDQBk/9fa01jDD97aFs23zZ9mo8y5BCzw2fFJSne7F
0n342KIk31+x2LuyATqurr+UEPb6li1axs/g9TWm7OKT6x657v6iemRSLtemCt9WcFB0444Hi8eU
lEZEN5pDDnZ7IEEOiuvPdKYU7TNFCpDeYcbaHewcUJQyEpPbPWWWtHm5moDUnuc9Ho7h8ffVNUTb
dfkWerttJRQUGxip71IFt+/RcRdZ2N59ade0R4e1ZyAZ/daHbOq2llNre3w5DhML5EdQh/KPww2U
AiO6bKmuoxvUY6NipJUBjIQ057yoRn/+XuRYDsuYH1yprtib5yX2+A5nzEqeUGAXE8q0Hzb48D7N
XRVF9RFi5NiV1ZwQoogfDk7JT2H6dEpDjbvIhN9CujHmwjHt2jFycJ0lFRqxscylTt4/ByJvqjdf
+bpshj5PrM5g1ftYImNVMVM0kyiHoQNp2lE8J+rR4IPU7b/UvQIttN4TJyQ0saITfYfbhjvlrgqM
wwemouZ9o7E1k1RbFF1VjNiC1IMhhuw9EdO2jEPeX5nhg+fH4Ahu2QdaXQig49p4Xd42xcdZQkZz
0KAmxZYyqfP4hi1te0KrhkI4iYQBaDNODFbWPaPmaN5huloRFGLDp7aAAb0QhLc/a/q8b2cAIERE
3dYlAF5+stiTHrA/lUSK6WvMhQQoF/M/VB3u53FX6k2BG0kqF6+1WkuHCJXWhyKwa8OKrmUrElt+
NSo+0XYFB4cPLDg685qD4b/v4GBkhbLT80eogYX/LaVs+4y5r0UU+IrwICqwFOWaHtgPk1P/BI97
1+vHz7ZJStaYcNAl2q9rljy0uXwIULyE/cFnvt+p17ASEurT/tqIXUauaHdvCyc/ClN9+gUmbMQI
Y25MhmNJr5TtFgkDxZY2Eu9nRwpSQ/42x3INn/WXjteJA+MQYbEE1GNQv/07ADvb6tIQm/WKETwJ
2y6DFrVVbpPO/fWVYWXk9Ix1AvvhHLNdf8beKSLuRzTUfxpD+bPXCymY1SgpEGrIwqWVvGWjC0CO
ZOo+7Fj3SbjGvdHMsafu4aIyBoIPYK87i4flwPAlho/z813qARTXbZFFDyXKrQHjvhTE5IanjDiw
8uWaP4Wp/DzPCMrhYdYb0cYZmiWJUfk1I3y9zsdyg6KZrhuIS6OOCy/pT1mKXFRpWTEd+zI4TlfX
W6+4xwk4UcVbRTEoax0xpwRhnfAr0Dd1uBwIrYT3TgcniwwqaScvMMdk5V1zZXN/jcoxXy8g0p0m
Pjjr9Df95H7SgqioLcPRaH3s9sAwDTggEKvcbkuW2GQ2RjOdCy/vLt1+4vmRDF4Ywxjp2kBiVvVR
cry2CtKxDiB7R750jnrPpVUvyB42+fw2zhyh2ZrfbBeRW0gNhjstDKXfdRTnnpZbxLrG8YUzspDr
ox9TqS9UA8KeubVTIwtZ8BOq+Yq90yOZTdNGyZal724Mewl127COQ2kVaWUyyMmc4+kOKFJ6wgvW
RbOrawNTG/+/Yp4p8PlXszS7Olnf2ejIgq1d88CV4gUOVlcI0ZzhjsBA0ZX1QtWaB0MzY4MyJjN0
qBcNpsye6ddr3H9TR/0/rnPSl/Gag57czlXLWWO68YtlMf7TVXuTBoSnDvVIsPmqR5WORX/Zdzgr
pX+JJNP7h9DVHUZs4X/1HGEDiSTOcs/LwKl1pIRrdHOccQ+nLuJGJgO9oNNQijWsshMbNWhOEW9b
CAWSk4RvD5Bxhkps+XMkcinKUGTLGw2G2LRMELKIbj2YVMyD7JKk6xlg5scoW4IhT2bplEulsYhr
UY1WBCoGL7UbyxLyVqpPn2Oy0ovgpO+VW6sq4bLUm3XBhddzd3uPUmsA68MCbFhLYeF12fkwVGAR
HMieVb/AFLe/d+vZl2exVO6DkwMY5hEAg3NcCjymH69z/zyUm1ruPHn1lpnTMykKjfmemrZz3ls3
jVxoFP7vz6sTzf4F3IKkps8gwzIRmOaweNmJ1CEj0X503znIEhOMZgM8PAbLPrG4wgDgwxPqzjuA
SQSawDdRE2rxW0Bdw9pwdDV6Bnv4xZZheGLi5CyugFiL/EUZfbMhu4QwvoEP+yLuI5NqEKxqWU1c
VX/q0CC5SOShxV1YqLlxQCwLAmhEjhQLSN4LRZPck8LI3dpI5CyyoS2rkksQX0ATiSqfHZ6krOm9
O6mP0AQ6u4linWUtqTds53fynUgANdh3XZb1uet0p6NRq/VE1R46LUPsnM9uroXPnuAxiXU6H70I
mrXuRIQE6fMUE58z/sin9uaMif5djoQOJDhWL8StUMcmmUVoN7uH6qByVV0FbDIjJbek4c29bXvy
oAYPfyNh0+iBGsRn3DXHJFtYABVE0v/gSrQY7D8mQTrzDlhQBd7Igu8JgJyy53fVePf30tXrZ+qu
vX7mS00UaLPk1UQzOV/ZKA5uFFVMbY2MceLFPu9K6Iuej88P6OEPLtdaoi7+P68jFqFUFcCu3bTZ
OKcg6MJ0r6QNsxW/b0dviFncWnSGPTl1MgCiaeiXL+RhMYKU0wiLkhILBeqlp/rHsBvmOczwGGqY
yp60NYTrs3m2QwcDbHc/zsaMJKXG2yOmwdA0gputE/CXCWg60ssqvt/XR9UA50Lh/LfHINjpKr+L
SVLrLPXLoB5jUjNSWfMACJf3x7czbsvOfTp6Qdhd541yaTO2YaM2FmmSJWE5/9cj8Zy/PN54HKrQ
T26pGBzOl0BPBLlKZH7gQ89af8E32SE7wxJs12IDi9w2vU64Xd/JRrOPWHmRT5/bd5VVr3kQYTg4
0RtVpI7PGg2q1kMp7z+Tj+gCl0t/WnJbirhLiParXUTR69/ZS/Igg/L0UOol5q72de+0xh9B4axc
nA+tfyFNk5kl+NlRIgj72Pkab/AxPYsOg1pmL3E4P07r/VD9VOesALNJbjpi/7rActs+v0rrunV8
YTvab1wkYh3Rl6bQLSQYAF9Rw7wuPT7JJNpa2HbS25vaahfzFl/4q0mkweIcRLAZtm3W62W++gIE
4fzIkYyl7Jdgh4iHsci8D0RGsfgtKeGmjE52tSSzoAd00WIFS8KxIXTv0rS319WB6qXqIVri/x5v
1al2+YJym6KMZtgPoHjpVUyLXqygsRRLFO7wdVB0IQ3nEpIFeWpCj1AXThaTnMsRel/CCE9WY7mi
Ntq/s/gFDVdLLjmkdo5fM/Tb+RummlcHgaJcNJN1HfKxJN9HoWYx9dMAAcU7d4HibLH9Q5Oeo+Ml
4qT8W2EeffqTlOIR5QwagndqbO8kjgjfZR/PbHPvPVafEor7hdVk/MTnI/qLz8sUmPJNr4vAj9Qz
Qj99z9xVwIlT+FuMjJXHpPlEx4+JcGz16vsYy8XJGzCnZqbucj9Pt0pPc61MkH0yVX7iNTukVQ3J
8Rw0k3/xGGPGffPeobYe6NMdsh7Tq5R0feQLkg6ibsWNq75n8l8MsN3ilcMkxas6uhnawjvrXLgV
Ag2N8SMkmzJXmm695F2kh9+kVh3ospJBEjMeAKLmfmz1EaLz43hSQY/jbitu2tDCMEInC4+RzxDq
QxBqyb3Zm/FXgeEQh/XNVYN8Cb25s84QLD5XZJ46/da6ZTi8hAt9Sdvnk7vlhYc3wYoZq/ZgcZib
HHPwIa+k0OZggQ4xSKk7uAtbKeagfnz8iCoESFz2Z+Z4O/+UAEZxGNAuUG/1rqEZbN9C9+C5DoVM
8RcWGq6UycblBySZjKP97ZId8J9rjWhZT9HGoMXoFHET1n2D9wShcyK++qseyb1mfZiXATTEq0DR
6veOcxaQactVdYfkZ4O+HoX/7kyMT3suMnjxbnxhj4vVWnhyN6XmbYrkHtxPKfpHflbre2cuS6m3
P1oWoX2k/gyiatCRE5YKAD4SOz+IHXzJlD+X5EBR+p0AfFM5xY/Fvly2wlnGuQcznvjXj0ugnLZP
EoiJy+U2l74JzNbqEbP00TXqUV4ivo3xWrSsTDPIb/qLkJom/Z0dZ2kJfhCL3u1G+ODvCIkxw4Rs
vwArTOmESWUkSFOJWZDlZhcyhnA47ZDIIOUHh27sHhiUeI7V1Yhe0AUFDXKMYro3gfJ6kSrg99XD
63QytnuKGDPZ4gtvnAGhzWPozOqHt4ajYYGgkndfrSUIgEeNhIJps3ImXpR+tPz14AFKNNA9gXCr
L0SCzqQ1ETOCmg8c7JAk3zeuPBGcoLqPvyqfMrsZ48T6j70ITOiIVFLsOZt56XhV6KqXTHR50ZiJ
r6p8l1USCw3Uh5SHPpyI/X4cC0dH/Ry67BWDRZliXj9T6Dy0wVQU8QQP60k4W0ukNtPcnjxBFAND
f+g1FK2YhiUJBsjf5dyING61Hs/ZFJLi4+ev1EPie5sSkjb7dsbo1kaD23x7Ul6cvbQHR3W6jZnE
1imvBcfnLd3vaXOeQQeRuoXeU19WifW0+jwP+ZXZypZrJIo5bYQJ8EO0LhyexY5VLFPw2VUHS6Ra
1v/MeQMxWy3W6ksCV/cYuaQb1dvWL1bKio+z2bXfOLrxA8cnjYOND9TIoYpCWDkooMgQDKImObNt
9roRjnNbMz9bMDsufnQxPh2Zd88h3T+FuPbmD4FUrTFo/lmwPzj0rgZUx0IlZS5pZvYAhYsPfzP0
k2EiDOynMjzk24w87L1eVfRABfrkmjjFo8u8L06K0wVIiRxDoepWqDnzDCXMP7nEmyy6Uc5zW2Ne
MIkNthu2hRayh377M0Sclo+aAbx+ZySS9iemYX9jl6zsptn6wfH9Ldd114GQl2LCHLi7mkoWQPdX
fTzjSKpfjmwnEUbi1S23DujERp7dmhb7EnSnvG5WR/TAXFT98LNmHk9IZAYUoKpb8TnTtbv4fai/
Zyk2cvGIUXgrje3SgUNASAOiOngXPd0oWkfN/aSyRo1Huix+VqiNufXjlf0rKCg8Ypekd8UBJxya
bgJEKGdrmsedrKr86J5mMaPGoWi4afi/A7b8A+qs0sIScKwYO8gs0BJzRKbNFNiS6DsOSuZ+26XB
uYpt986q8cB6EA55DPo+A6l9le2dHSrKxnSCFNdfJiD6Phyc7wGcJ94jxOtM8+AhTkO9MD56pbXS
9VsvVbgsJhJuxSPG1y3gED+OaZ/DQqf+7xOyur1INiUxVM5SKdyR+nRQOaN8wOYlZQm254heXKLP
BvSRN8NuB2ME7TevARrclbtkoOT3hj6E6+IPyAujaRTjg1ii/tDO/CSDw2B3o+QJXNJA5+FvAmov
bbYSUOyMF6awZ5TYPP2BmGjMTA4/npurJiMFF25vnIVvzlgMB1TKZMBbIm52nuGZdSL54lkiT52x
JDVMjwqKJAfpPndr7iRkwmjHsJ7cCON4ij5vNAVoFcky65LpbHC5L16lrC921dlgO7qxipZUHVC1
ugXowY9sQAl+c6wlzIoRoYny9q+XjYtnK9wg+5cIaQzlFknh/A3gt4pNlZx7c9PD34ZS7kE60ZCX
C/DoSQ/2TfRJ6awPkFnNJFdadsGvN1RFp5YmL8bzvHHhqaNPUFNPnUKm1xIKlDhCpxesjfxNqppM
J483mjsBNNTA0kpps44KBRtiaSA92WHUxlpFol4/F1ejCy4C5sBYn+0r0/3cD67XiRj6p99fI3H2
Otp1G6q57XT6rIjXaQoGrPZNTEYCR5DAAlf4Q/p2lDlkOdMXas4sFeNfpUisrzNcjm4/Gwybu7DV
FWmckaX1hpkZUvjlqsYKSPAa4hK5t4kYOXOs9/iSax2xaZpYsRE+jgoTslNjqgDSeLQT71FE6sii
Bds1l+nNqFtuK1CGwjlvIGWnv9K72yXqljlyHo+nClStZk/3ItSZp+krjmBI+9KYLXg35J3W2K5o
R6luMZVyAr3Ji3AtMwvk2sbd0MyaxNulq/tu9iTirI7+EmVN2rDvvrn4QK+Qfb1/17P/W8B3Dar0
JbRGWNqwHXbocbfxtH6yU+g5L+ar9qnmJHndp35zZfvUH31lbUSmR9Sel6trsndmZMM6Hh5DVQXy
QjoeACnAsfgh4zqcigd6jWfIzaJ+55FeAwZUxAFSwGspyYOpxzCGwmac1+WUKr+CLn6Ix/YBMTZ7
361oD/N3Brz0kYBrErbhTzdl0yIiGRu0naPP+KURS2lUrQE8357NF1Z3JbDfVnCTdXiJTaBFGPv0
vDONhoyx2gQ7cGu883z259RmqSjzM3wPTgYjK8Tik/Ly81mKmdykyKc4jaCyFZeBKpgcjCcldQGp
O1EeIe27nmDpfaFjQ+UdEcxQMVQP/3GBcKC6+eBEG9DKBYhnmuxbzsyMxtE0vkEi4gVYxVxCeqC8
hqge3CYwvKqV5N6nAHay2snuugTu9fvYnPjJ8YRMCkjM0nR3uYoo59Z7xeX8ydlXfeUVHfbFrFQR
XuDP64Gt+KLPT2BuEojmI16bU3DAG0TG3aWZb+IfCPsRtfUNLmDmxCWImt8O1CmZMNby2om3QC03
77D0DLGfaYmKjRnTMUg6lnmjcENhWjssDMx8rXSOQ6/NFqfkc7wIh96zAYwYbde1NTTsFafgEsyO
QpZnfDxtjsluI1NRLFUUoyqdXq37ryBNN0dR8SR6Dvv8Vb8B0tgrTN/CVNgosZ6OQKugNN10ALQ7
qgEgu9a3HU7+jy5zO5AFgPR/l/07mRNFyoRbRLSdVBA0/AxXPiegSennG9pTvScVk3oFiPHHAX1L
5Mjf0gkd1L8Dc4sNt4jsJEkpJNOAviw/2EGSDJ5RqUIWyOKL5l/2O92CWnZg+hm/fkf5P9TbO1YA
e1WF1BaEX6PNIZkiAWErZvk8luaeh+CPkX9Q8tNRACoUPmlqP45VDcpnS633N2VNszy9ZCoickOM
Vm92XsoptBHu46eDNbxG9mgurFg7KA6bG7lF01KKYFEXhbCjLRbIbuKkNrEq45scC8VQKEUtZoWm
mWep2Tvu/vJftMAbamWp2QyzR7LyZ/ayG3N1pTxBebYUGNOtTMyrAipOxn1ZSONIK/WHQtwS3nL8
MmeZ1LZ4K+UPIfjIfz4lSxhUqTx9Tnjm+axanT0rVWpLqzuRgLKNV2kCENqVp39m4trYKb05tOCO
skKGIFubfWQVA2BNu4DyYLDdn3Tfu7mJ1J5bLtzO3v+beJixQinBUhyIRIE4BMU1NTzB+GAXEOD0
RL8OrYCBWgqJy7qgIHrzKIVMTs1kD6PqDBxZ+MB2VIczmjMt9ai8C7bC7qUC9JH+pSq9ViNqZuWe
NSG+EqVsSU+LMU6W76DstDOxeEo4smN+yF+aYGEFX6w97o2hK5TQmYWM1Rf28xT4K9px50LZVExo
cz7nHJCiA+Dupix51fZBstDZkRNvwpy2/Xblo+XlvPPmJEdslSf6sLBQkiXXBRB0GOaJlNXKQMBH
VowEH8X65YaGIpLPIG/2IKWCOL3iUb7dSjSSBEikludZwthTnjTmIsNLaFJTUZ3/iJQcdA6d5gDa
5EWSCurQJreH5w/N74ZySWr2KjXEIl4d8DN5BLCvncWXoTZVuPHVpOBGg8HQmVGGhDT8chWjb0GM
LWjOrB3AInowsc5kT/x3GQM+dHxodkHOrwbZGLkhQO4moVrY+hNNaZB/4yTVrAE707nKwrTFwOI6
hxfea0//nO3/v5p+TUXTzHj9FF40CMorwFBs6O7vYDpiOLEaorAN0LIuW2ivd+PP9OW0KuEv1qeQ
/vr0X8/oN6Udv4TmRtj/mj9P5dpXJg1Hi+Fo5KjvPE0Gh9xIseWNrTlgZe/4AuNslq8Y1X8OcE6g
23Pklt5T+Gk+FozVX5oBmbK3aOkO8kzWUBdSuwL5yXPQ4yln+WhMW5MGuqZfoNp5zNt+ZU+f8HXz
6stzmVEj5yx0mr16Jd16IfgpW9wlssW61TA/R3VT/P6vyD5Ah2FBuAxDd2PaC+Vs9SeW4Y1uOv1f
WjGF6E9nNcJtM5gm/z91Zt+b3zOG/l1GAw1tdpaLbVsrAu8YxaMOdEE7kX0wz6WaIV4qNzYb2Zv0
hor84Mc9ii4fu2mO4bbwXscMUX6SVSbnlnd+sPjuXq4jCVgUSxK76DrIfdneeDRj9Ma0yTHet8/Z
gLJD+jtCLEv2EjvpYfuPqhgKQw6eZ6jGsqB9rw/9A2wY6jtYInvg3B+QxVG4kvmi6FHwEoJmEuEw
FM1n8gidY5HKjeNKYwWnywrMQqHPml1imKqRTFsQGoC8UxbWFqYXbKLWbgjLOYP3TcWmcnmtwJJh
LRyoLbYG8YiibG/6N/6JmCaHZlGJ1JX04XWDLnmZGbiQaRyFlKE4ma9ylYgNpYYZdaXmsjanqdg5
ESNL47CtTEGh3EpRnLEhucrRS5Kp9uK+Tp5UejuKqueRiA21/+yi7Tf5WqIQ06ai2wmCdiLfbfsQ
uZ9A1M2DvrFlGqGyBY6WCPZDW6Vm87lbCqqCoi4nSRKt8jJElCY5v2KXEpg976piTNMmGjZYEO90
GBtEQvFs+UHSJveWZCSAPf6UOT3Qy9YB+DVptkUAmMltOjDkT/KBo73crNEvylXQwzd06RXe9Y1I
LkA9f/BfC5uiJh7Ka5c65Prw5kpXBmguJYNZqW12DJbJpqZGUte0aSDqlHCxBKdjfcdGmQMoBKak
4tVF+VMJYHTiNGUQHhLuzjS+87qANA+zqmHQ0gK5xnoBfjcwNdgfUsTDOT7Xb3Cw6N0R7Hb/a8BH
NTiSvw16mdBKxJpvAJUVQdZpV7ZBfcdM5a/qc8EOX7MThIA1WUZH3d9DWMQVlBITK3YlmD5f3opO
BVmm5vPNc0k4FCV22Sz/Y9E05NanEOm3kzTQfJAehCHvdA7LKPGso8KYY38M5+5nTsnnMkfejngB
TK7ormj8ybFYHQfIR1272ka65Upe1Hh7UHQAH3j82Hl9RcKUMmfOrAIQ37Q3/U7vag2VC6dEA1ZH
Xii/RRUzSwU/IvnyWtPlni6YFamnt8afiel1aEB1qGBRe5KAoEo97sffpFhgijuMNBAJm/IfvRkI
YJdS8LGtL/ykwcL49TFDp/VhJ+zyBOtHfTW9Yp+Ana/AY4IaUDqlIKCfRSkzrlPsEc7bIcX9mDrH
IwVoJUMeB9IKnwTrly0fTAUBR5l5PYxRaqerGv36EiEef2qqHEcWJDfqcfFMg1NDn12mi2eyj8fr
eXbrXumDk7BkW0uFQBU5/eWCFvIncUWINVLNBjSBSAfAHfgI7jyXq8yA1KqQS+3aRS4l+PyWR6gG
YQNtEbRHlLtqre8MyR2SxnBD54QX14YoOl6GzxpeUbfFurIyYNwzbloLZEGWfU4eEHvCFHAgR/Jb
MI9eVVLL2JyZ+0Gas9NGgggARgPKc/ymrukgTMVcf/7ArUXtOmePotpNGZK5J+RuEwuobawVlFNH
6whfuUH1ejD2I9gfRhGzWcaYOVzeqFyzlVZJhIGKCCV42bYr7GLYZwo2v2IAOwUx4sg3lbWAkctm
waT4nfxTA9aA+XeMB4oh06VB4tJ2X5alHOJlu1+2lQc+dGNjrwIKPvMCyZJ5Q2SJ5gXn3GRDBt3p
HjwO3fHFSfALcb++icY26fgiV9SOs+Io7oK6Ypb76lsGMiZucC5umqFmFAze4NdWCIZrSAHp7KI8
GeAYoNaRpdznA6wT6PHdaQrp4nbL/MXqoNZd/EXjMHG/rpO0V+dKXehv7GjOdvIpzCiOhomA0Wzz
+V+qoVNJuLKRyjEzMNJMJlwm4EKbPvmZ1jUDUM3D7WMmoow3f4Sv1WOFpYIIRkMMKVF0OJgolfWZ
k+6sitxMQVk5soTHb6i9A1AV7wXoFtN/zsBi1iI/pT3IFv2TKVUx9JgeIMmwYrLkpKUl7UUgz0sl
8h/z+e5qOPTQz9iUG/I8QUuyhznqKT4xz/2hmLXLw3XpbryOomzTD7ejV6chFfXdpsF+VWgkH0H+
AT/tLIs7i4r2hKnHBEQAQ8H1yFVN7J5tjHiFEELcp87U20SNrIxHPF/ovHLylTFJYzSsx71CwOss
Rbm8dR5TR7KvPQ+w22U8pVdaTxEusH/hDVDwry4orHIKPVWuVwV1cHPzUHfg1BvRZOCzb2cnfGmD
5ByPsR7DdeD2d56ENmsBGBUVLpZdO2mspbKrpYlHU1qLk/143ycINE9P/IB+jj11hr539GlE698u
o1gLPE9dh90TFh4puf+ql0rfpVpw4ge/9x1RPaZLl+rCKxqlywDYl4s7d/daCAdqLMMaWGcyab2U
U/Q8g8QbwDl/v5wju2nDqwU2NEIC3MmPI8rDHNAGqzAyJnsMo1z/vqThkK9Au+W42S1hIOgVZNFW
h5Yjkde3JhW7JItaL8eapVA73ZJySFBzIKIUKlBbqy8fU2Fxxgh48bJwj1WbefyRBt77hEmg6/6Q
ukX1XliidSAnuhb7cfLhauhfk7hQaFNshoKx3ujq1N8HWJ8o7WoOYmfqwOJ8qWDUM50wlQfRqoVD
B8SYRHZC6Q+8rCck9k8p5OWwUsS6PWr+bigi+WMhsZ/RX1mwGd3YRsNdVZVgajYt1AeeznV0fVhk
xfcNhUR7mtuWwtNeUFVnLO+spJ8itW4Cpu1rIky2sOm0okPrGK9++JlUduFjTOU9j1FYMpvYP1yj
HqSaVLh1qHbW2Ew089nCEkWdppl9lvP81I5KlYIc6+G9+1jBCJoqCJOQQzXni6kIRaa60rpT9sEp
z4wjI3TDky/21KRvjxcSI0KPFNRfh4bu55Ca4xdNeiilqjFLcJ5oExqxh59nh/ZlwZVEGyPfH0es
ZmIhP6aB2cRcmIB2AQme2rGU+4XpRhFPk21KbCHfPIffGHc76ZQKGssPLU9tvXe48qxFA4bYzoxb
TxkvgsUCjxf8xGEFpfrJbk3tDZNZAGp3KRAl7JXYKCcqfOVcsw9kTXDXBx6SyGa3BCaVVxyzheO8
AfY+fXnXYe3L/WjRm3/A9wEV2rCIs6Pl7pYmClZRJnaxUggOtNwExx48+RQCKn5EWk6K0aBdnSsj
P4oGomRc1u57jJQTv4jcSh/8GaE6X6OkxzEJvKGirKHB8etRS4zUXO9UUYk9ruGrYa8TpI7v++0B
12p1h2jnmKIxYk+nfkmAYQLck8il9ZraP8GYw2iZAlp1yJLh7T754mYZSdMy6mUE9xb8yq4uVAX0
4cEFUrgtNXd6veHOtGLnTYB3qTnwTHLUsyPfgH6D2MMoVGMepIV3Ih+6g+kClnCA32xWIus+40Gh
gjRJAi6OFrkbX7Cp/e+nXwSMeBMIRj+ZBVL7fnSQWplfzqw1xe1VoifSHa1hBEu3Ye9hiatIPejX
2syc7yzrIWeSRHoZ7MxEKa2OfYJoH1xsGfmNPR/JT5dtCnpbdNs4vvQjmI/2Q0/KSPwpGigqljMJ
A6WR1HfT4LZf0gFXBVNeUoK4gJZqs0AS3/zTFPH6BbJKLL+Y+8oA5pZhmagu5fzieCLE/96sOjR/
Vbxm4Hs6yhRt0mIbEU1+yqFUU3poskjaRIwN71CnJEHE47d835QMZZDOOhdsgj1yUukm0tNptLqd
/P32gxGJ7OVBnffBzni5QKUaIYFSycjR/tX/p7fMUY41QD6TVN9NgypDWH8cy41oKd3PiYB9g0IM
cwUgjaSmtt2pD1kjLS5A6P/Hw8khHDHjk9V4hTxXglEjwmao/UScCItmqyjp1bsF6yaywrta4rPa
WFkhT8MmFSCN/gdMeV4nuIlzsb1uC789NmS8naq/1Flz2Tvwlg95T3OaLCy+pPfrhW2Q0N0EMBZK
J0N28ynrV2ynk7L/Zi8Bjecs9qNPnV73fnwCYlgtm12ym0gO/FeQTQo/Tm0tUp3tqkkSKvTgqhkd
e5UJDOgZ0QxJyq20MjSW1lFEKAlu4t0c2LWap2Amvl1q8jvnBaCuP5HKKvs3mk5rAhywTEiIMO7r
yv04Ae11E2164VcL0hmsoBbuHojRdJQgAFnX4JiuYQgizcW0bJVl3wtij8QWe6yAkgxA1UDc4uD1
9ZlIP57SdkyhrBX0vOt9MtOedQPPyncGSgW33uqZ3RkmImdYkmLAWo9LKLem6zFJ0BBPkMoTk9GC
jnMwaRadaXyEhiqxgNdnBm4PIIRR+xQSYNyAJ28Naf62VouSou97sb4W9y2SnQZ00PZ3pb1yk7Jm
V1ux7mrIenmwqUhEOK/iwn1h1NdcLYFpUNLxLozq9fA1FskZ5DEFwt0qoIvrdMlNC7dVieDudjmH
KBbwHYo1D/VCNf1mgZZd/FkhVkTtmDeeow8XGEFEjVg+tWHxVuFVRdGBDUxyg/M1sGFBiMd4rH1T
S+Tv7hkV89AO8/02ftIAuSWqjBjz5tTJd2XgBJmPpFHdcAoGPc9Pd3o1h1WhvURRZ6CYQE9nrbK4
hty6nYjodRYbz1RVX9R5iYJ/4y/KXAznRp1m5nNz8jVMc67IYvZIUFdQ2H6kPFBVGi7tOGV0kfAu
TiTElWbKKVu5VS2rmVlRKbqyIgX0D2Qzle80FkUSS35b/QL7xucSMqFNYijhunchnGqtJMz0sg1K
gl52pILV02SraCgys7zDhMDKW+pn7CB60ah9dUrynB0/gz7zpZnVWTVM+5VGXeGOF+NLbdZITX9J
UXS6yKcXXurBoEj6bARisnEcc2cQ8vjtT/VSHm/Rczm+Q2dNlGpwF+Uj68SGPHribK3eZTQ4WKt7
yUqvL6Ewcgy3wm+K+Jtvhm2zCneesvYmBRu0/pcKEpPZBnyLNzb0AjIcZKznicBDfvE2eCwcS6+5
zhiGQBAfX8pgtV3FqZQ+N/thoxnBUKysCJsdWG7q7GGSmW14QytDzE3YsfGxhalKq50d3vBMk3I3
XXq3RVDq+l4Eetp7ltoYKeCZcWp5NtAZjSURTgvfLkUg6cIKNDzyqoQXS9A4zfG9nTyEL2cNyszR
AL9XS5eSj7aT93OA/ImGh023LRuJGcD6IfiDnr2jfm8Hg5zL+zLRZ6Vc9Bzb5Hwn6JMWisbFiFfx
sST+K5Hr+MyGW+b1dI0e7+vWRsAFtTEIWkEPTp1S0eO20TMrGrVmcPo826ONHarVn3T8zg9HazJ2
1s5u0qC5/9MHfXAirfW2K+fEmvUrhoy/sqC/Gby9dTOlezQpsPdB/m/8HDaMnJWyaHHPU9/q31kH
331HOD19TWIR3G2DV5RdvglHAgQ2yniFWHQ/kkp75235kL8cvGq814j9djFcAkzyqKTmYMtwY3Yo
NQU9/Ohte0WA0hvlm7hY8vPfPTSLCfgThS3WOxPz2At3Bhc400dI4+F0gUaTlEM72+OObHuQ3KG2
dtYqWhajq4ZuNifcvMoZY+/ZJUJKm52gM0bIgtCLrlEsoSvz3VPp6wrMInSHdveiYJ2N5h6EhdPZ
/ljW57QCb2ex9WWb0QxNT7s+xBsETWy1aSq1upiUEXCAJ8xdNaebGExSzLPy5CpaO8UUJzcMlfer
kz7uUkSrDT1qRltvLp8JQyZzL/yzrffD0VyDbQhv9DfHwAPSRoodzeGLwR6TeY3nM7D0AJl2Ddsn
TXigO5ecuBOkDJUzN77cFNbwhHvw8ycsccRDAF39W/qkt2JLADeV10sc9fENU9YrBU7GTT3yKJho
kP67aWZAWGorYEfazaQIPH7Z/wQqnRuBvBE1vtQU4qnA0jgc/RLU6M6QuC4GW8STWGfduISt/0Py
hYtVa6M9glhDSpcSVWgU7rDHbJqGnsDKWFcNc/LI2UGPWyy7P9iTEUAAEynApLBFSnmN6nIj3nBv
8398DXwWkShX1VkOW0Fl1FYzUOT8YJmt/fuK7siefdIL8sIYMLHQFmjsSXRxA0/DSsCM9HFFo3Wm
V9GkrVk24TzJfATWJUTGT2PxBs0FUzdNUt4QGO4mwyzSyhFOTXy4OSqngF7Emk/Ixn73IUz5pjla
DPddFk0kQPrAa0a27U3GmKu7esFdg4nDPfalbasOkk4laLIbMmuunvBgGB+ZSO9X6GrC/uph/Ucc
xIp2L1et3PEHgNSuNPBLhcQ6Gas0DpRfOVrMR6VMlBXf8dId1DWOaWjJamgg9dXAko1m8+X8+O1z
OBkgoL6y+MyvobqEsGk11Tl/Xj7l4d4+2rs+x1QBiqPZrK/TTLKqfkimqPzT+E+IoIndqcf63yj/
iM6cZ9PHzFacQBjltuxbyC1uWPJ52qHap3Rr8oPp+1BVAW0Syoo4Cn7e0ykarcTDVuqO9QUPBGlZ
9Ek2NrcZdP1meYaIGF3Vt94tI4XHC2EkSps42q7elqzpkvOqx3eCuyuFnMuJpoTPoA7oImTeZNWY
NLStbHv+EfDpZg2DEPebu43bLzaWG929t2yMo6rpmrZyDIOS3FKRcQMIwY8qCLFlZryRUNLZlqrl
iV05ORT31TFH6JeSJjz+NO9nz9JkzKsZgoGJ8/hlWc44wsw/4W+0ORRN0VJP8MX+IdKGuKZnFvaq
Ob2SIoGlM66o4OhsewDX+AT63mlyeC9ZRdjzHKdy2HnFaxeIV4vJPQXxLeLJ9JuD4HsJR3Inchw1
zNJ4dyjJDgHLXLFlc6M3E4DvicPG9h9BPA41BpKR3wr+LQ8efvQcatJ6mLG89SObqJcW0uDLhaIM
g7HUA2trpliV7HSSG5j4VUcmrxyELa8Y2GJ23LqUKxwUK6ZbbbWXbzE7AGxmJSi/iBJyrg/r8Uf0
n2Md64B6zPeF0XbsGMhsbyrBQQ47Qm5rE1LYq0e520r71brHc/fl/yXNx0VQ01nlFebHh4rfnCsn
+YYrwyqYF6UlolW9pu5zDygBF79e4XTaCosfa+kHHxlfZWhn628syWmkGhUvUTh/tvjNdO+Fp5UW
vLyCTYWP9Idw0CRu1dghZSCdrSu6wAaskqZ6m+UquILjH4Stlivui2cqg2QAfsJZtoFLug3f1i4X
FWAC/W6+PUjfxOxtW1Y6wLQSs+t12B2Hw+AkQhA1sO9ZRRNtgrrsIqJK1quVPzb5tD5Zxraw1vDi
AEZMkyjIAZApHJdllMJPaHB/XrlgaMCNpLUBF7WDzq9EzBmIW/eO24kK4A1GTYHrSomP3L6xGU1s
Q/6GBtCLcvVjJMdASLEr35DXymMcwlILOTqNQ3DVjThrmZqVK5g97YURndQQnFSauDjV6qqubEa+
JSkijtmIBysWWooIg++KNCIDLcZujgs3vk/0UxfwTyCNTIlIVBueiIlC/4voDU3au+u0NXQWA+MV
On7WrxsLPbhfiA0q6wym6hDZBdINjNrbV/QSGlTYHWHZiLfU63LTLV1J/E40xrUPgeDycuu0fjnN
t7V5bXLa3Q9biM5/5lcDOolHt+6hXWI15z7YHhmPqkyO8jvJF2aWxLHXqvu6iCZCKCN9Ye7BDV8I
c0LbpcNz7TI82f1vbssaigNABqdRnpyaW9sf9VOJLNYQsdy/pXI+OaVvAwRbKBDaRlS32SFTahVL
qAGgUZG0+GA7WEc3BR4g1UcR8w4j+p0YQ5PoWWwr6Xo13oJg/Kqs/2+rSJGZpAvDg5/1D6JpFQNQ
m6/KMek/a2ePS1MjNlkhJoGAquqsM+cezujzTq5sVhydh6F9BT4t81zTqZiQj45zCPokiL/k0jee
eKMrWzRJ4L+V5hltM3SXRopiIx/GikY5tYI8Re6RmU6cNw3GjWE9CUcUMD2CeHO1kk3MdpVBZM/Q
ZPNxGcA1xinFPN0/BQkOAiqwQ8mJYjmdS3G5bmZlsfTgU9HIgroWfq49TI/OOwL0n6WLQ64SVbU6
nVKxFjBx7485MojfRC5v1qNN2jJWOMf/B16QIU85sGi6jSbdgKDPZn9uaN1rSJzwjUxf/8KyUtIf
0f6EYT6+EfvB3K/RTo57lazImYKSdldj60iVKOau4y39NGy/fnfj0nsQm4nfrbKf33C2/2pP2MJ9
ROcMQifRBS71/WMdo6r3tf3AMSiiqY7ePFXfVlW5NPUWrjRHxUeHNR6iTReAEbiL8C46or1UbxQj
zbtR81BFREqpL13lFvJYJKlqzAzoLrBgv8P1O7BDKxwQKj/GH4X5S69u+OMnNmPliop5JRh6NEH1
hCXnAFnc7c5PMLLceeyDK4E2iamKZ5EabJu4C6EDhmmhdDs0RKIRp3A27G0hoGEpkSf+xEyaH5+N
82E4tgqmnwFPuuN72e99PhXfBxhWJjTdbAEaAwoXPYntB/ZNM+ykuEVP1hTAOR82JvFG3gvXduEn
ULeb2NdsHY6EXK7Y+qLpIZs41/W7uO/DTcFYBM7lcvNPCUhr/nKoGU8sABCVaXOdfzMTRbx1i886
32HsQWRCRQRh4C1JzmaHvO1QvH3kigO69txJivAUSqdYtHeV7k+TVS4oL+euawYrT+kjeRLBCzL0
EfzFyPl1AwO3BnU5LdHxQCBEmL0z38RyQ73AMpa1NMSVgtdGOU5ukHsN1JYF5YM1upbE0SAvwvie
eV5AhlDNcKYPjZa55eEzbclAROt8ZfZ/XDZQSuwzaAadoKiq2h9j5Shl8OwGkIk0A+5UIm0pBEtP
uX210srxGFZ6OCAqEL0xeB02obmz/b54U2HDY+BjVENhyjAwW2kTfYgABtT0BtElNOQcg1fYdPMl
5PMmsuY9AbF7zhm505qch+/T0GaChW0aqrHzoAj7c+RSJO9+2SdcqPBms7yGVHxdaVUq8zU9uZNP
pJKmIWKlmKk0fKQfz67sMIitC9bUAEaP5qRBb1/pniCzoTmb4naj3IERKq5+kkcE2uVYiXo0MWPK
DpJjAD0rn3+vgxVqV5+8/E4GguoiX+9krRMPgQn9J+1IUbWL8iY5imuxH2w1BrqX0ahjrm34EmxC
IjN0OXfPQ82L3C1N7fomo2tcOMvJilCJAaNg9mVXanYc5A/4OUkQ7+CdAB9WPN1OLmPeqaL55t5n
kmvrXwdUZvPr+Ib0wZ7LgQuFUfYlqfUbi2mWh7EY7VwTaHFEqc86V1Sq1yZwSy1MgzeZ2k/b+QVq
VL0YdQil94Jw2F2m5HFjfz9Jl7/f//OHA+Mpwc11XAcG0j9gk9OhKATQKfK5n7g4f4X0QN217qaJ
Y4Cz316XdrqHk0FkXzdu9XoMWosOubZA7tZsNtFWsWJPY/nt1KLlAklGt3j8Bhevxaq38BdsA1R5
KUCThWzmf9trF09JsTfplJQd/JURvQKnm5DXXKnOmpn9KBYtZWNUH9zhoEjcrIxKRU4P2qlD3o/G
aUVfGIAc34sLd6yZSShwTJN5z8rYGikTwZkrUzk65z/0m/q3gZaG9SGsbZ1g1SyZOlmN/v1dbxjE
kqHIuYXa4om+6U9k6faAiYHj2SN3QXtNHZpBpglIQwgbXLeWSiZGeSYjtxEZDsiBOwNF3Z2g/CPV
3YbPFijXo6ANHfqEiWL3K2wrRzvqJR60OBVgtba+4umSdcg76FGFyPh7SnxKNFISVpvj0FDup1zW
nXxNOZWmT468WZiEDfYnvRqI4wKlwTyx42wXK+YQWPeujUUW2Yiwr25bJc76RQvOlXyx+0JsIdlD
hALJG1QA4z/9dnVslCxs0OeRdHk4n71c7fu8RlMwsr3dHv1H3vcEtyPZtSo/ebcT7lZINnNIlWP0
lbSr6tZ3vXYwY580UuXs9V2q1oORr0O9hgQSS2UnbIPKet8Hii+LRGzWm2lT1WTRN16fdC2V7AmM
XTJNRYrnrYlMA85c/79ry0Fa0tZPxPXyErDDJYr2+HMESjILhUOOFj8PndFWFAUgoE2t92LTfVd5
laG0B9e10uLP2rfFzd1JRHg3EOpBopYSTd0E5rbD7UaTcNIM7B91tvJ9LDQvGDilc82M6WHpBdkq
xsrcmChLEi2ClbXAfyv0FGUiVj98/Aw4AZGC6ImAoODBmKC2StWGHdusvu7ZvAltNEiuoPqHxWxn
FHGfw4dNYLa/trbjBcg/M5X8jqQiQBJ+hZADsY1rs3kn5WniPDTS8aFm7c8uSoE3Tx+jew3/g13S
9ZWCCO/p5OPeQbUu9QnQNhE+F9vgwGTGgU68L+eTVkNB1ZjqQfUUFMXM+++psGxf4ZNyKuQwCwSF
c8PPSRNa9ZMfya3ITHsAw9mtYB5ymoj+RXDDnqO4/HXxv1P2BFEhgALrV7dgG3gWhX7XgN8tjFvU
z6m1nTYhwyn1kMArDUqYkbA0jt4/aKfL80qeEfqOp+nLtlENS7/jiG/yK/iIx1M+6dx7MgblNDfX
dLdVlGdNZTRWjz9Crhp9mC3giyBOJpyziV2aN7ZKpk8+c2AaSYKly4w6qgenZVcYXTR22fDZVMM5
jlKgg96l5j5BhF8wdqT2fhrf2uD3cktLSQuFZlcP3AqexGmYdkVPBpLF5Wn8rAI8pGV3wXnJ36R/
T2DbGKiM8mtf7RxBjyVudztNAt4H9VUfcnCxNJMl03+VHOsLWT+38Y3QgGLmzlJtOeOaWBj/VJoK
+e43/7p0GhZ5gkukkRdp9l52mtKnvBzYM+NsZgJgyF+/K05Wqx2dLTmfjdVBq35V6MmTz1V9gqH6
FDCnSehjQdsuAoZC09lOC9MCC41Y3HurYL3BgmMJjNOMiNcYsf+kXdw3VrjAONCYwxm8UfKGSKP8
bBMOEZaA9jqDi1J6QYq7yrYygHR1fevbh2QDj1AGuqbG/eqmCmovWuzUCzgjaidcF9waGz3tQdkt
5fb5qP9oIw2IRpVIgU6eiVbA1pB1BUQmNFDdQXTymOtwzmTr7cWXoV2O0DyWv176ud99VIENRdPj
gpK7D8oIv0tYYXIuCa0i6p21wdr3jvztxyDdZO9EUpU3YkwQKvjCCJQulxv/2bd2k3xxFTAScNih
35PbHn+hp9h/a7/+1xa0zTRgTYAhN+STL6PakwH42/Sp+B2X5xLZwiJyYfaxy9jNQAnB83R6cVLG
BvvU1aPi6+u8B+4wVxnWrLNHSixIKwpZ71AoKcqIeKt2iooAEZisdmdJVnuhY7h88DDDi5MeE25w
ixO9PYz/wpRhPGyqYr2dUWNKf0b3hPJCYKCxTNqCxI3pGk8PryyDbrno0x6DCwaLfK218GWRuKhB
e6ThQ/9lzGZpcdYplpSod1+wijXyHuhq0dWLwl3nHxOHGwom6aEf/42l8jtmWa3g6tL+JTMoIF1r
fYUk/I0smP8pJOVDUwonF+Wu1/bmPsxE2mvzqctxNyj2DH7bnSzMH1pUeOj1ReIyJp5qMaqGKVhd
N1um1Xtf6J8afPnsl2exY4dPMo2ArdcU0sq4iJts/0RqKKY9zPhYWnwskRxMwIj7S6fj0phOH0Fn
MqFa9MD0j7Ckpwzj2LMfQb4eqB8J50LW8fftP+syVZlcjBopTG30DD1srblqe7JnesGOlh6XI3Y8
Rv8kD4T8RTr59kyssYaEPt0fFgj9yoa3j5ZC76aWmt+AgeOhkPRPFD86rJ1rbGgwcz2x7DyT+uXY
LA7zBS7yvxAtLCmx8utboq1Z/+LGDGAdu+vn3DhCCHLJw6A8+Dy47ytXlmmVeJyGL+wEga4TQb1I
cUqHMAs8QrEOpLueXXlUh6jsswdf/bcqjwcSYUHHKP9FA9OXbjNQ8QR192jgJiLwSGPmCCh1oj1l
0RZy6wLgy23jrnYBApb+ekkbt9gvinG7fdbcsA55SFmPfHHtOE2u0ufR5cdiOZoYDaFetwwvpMtQ
RBoHdD5oEL8r0OT6+NSC8toCPkfB7JVR6RPM8pVKIG0/v77QSKjUNB5ZotFxxSMEOWoFxRaCNgmp
eLj60cj31J0YSPU+XYGWoq00cagqn8uTa67LGlLT6NVZwNzATx5j/LEJSe7ZFBWcL+5igB7JcecY
S0p149h9WlF3bVmlmd2el27c9icIQIeMjICDlMklFymAdikOBUzZtD7Qc6PtmRsClqiRoZ+S4eL7
3sCpRQniIXsPhDfGbzTgTXRHBbD+N2B+MNaWmpR51CF8s4aYehU3Leaew3xNRjVeweiFr45jzzx9
hYIsInayZZMF+SM/m9SUeAtvCHTl0mUUn+EHBOMdX4E86XdGz/VhPyGdsWrEdRgPEvrWYs+K6A9o
4ckZRNUsgThIMv6LChWWemp2c6rm1DsRliukZ3nXCrOy8EVwnQKcuCiPI75ywxd24p+KCnIjmYjI
Uh2Jatkl9L/MWpvnJ66fxSNgbSht9UvzYfiG01he0+N9tfNraP/GaYTWBbEhVhg7vA7c71inndQa
6gdJ0HCiqnmULybw9sdMjilszvzPPwD1wxcteJn6Si/TO/C9IPnc27H8YwnJeu+Dohp5RwxlSrqe
2mmun7O83+37zc/tWM5Eb4FpdEEM41skCV6tAJzKSW9nn471eQK0zaXdjlNmq+LLiwVxy8kQRDKg
ggDeXlBG7N8Pa3nQO03Mk382fhUXq64QHCkN4P9F4VaCYGVQsvBHDhOnI3jQ9uZhZ5OX7EB47OHL
TH+ZRMgsl3bAmsGLy/GvgH2wR5N+0ELdbrGXK0gljNrWniCX7cnZdhlK4Xo9qXbcIxUoKLoKvFx+
7pbVrGYLiQ/HfInLrlt/ZJWWoImVec6aWtjen+DaJY11AfNxt0RfDWk0BaWTifLMRftdORwUW28G
vvnX9f75HjblfoHlDepI6Y3Z6Bgd+u2SWvLzgMylJqEhfTOL/oHM3lIs1yqWcNUIecatuhD/SLxG
zDWoX2pNV54Fil63dV7qtidL3ZqJG/YxEhj88bQUAWhgw6Y93LYk2qKIZA6GDenp6qQbMEr9Nah4
A7wd6dO4v3MNIXG9ua0Fc4MArVBkxltv7kcbXvWi20q5o+Rme82QvInBq40ZET28QiSj9xxH3st/
vek/Xiz6MUmYCWjYilcagGuBabTF7fEhhday2inhpbJwK+sl1oYhq6K9sR+twvpJqmwaUdKe6fkL
/U5kVhNTgVGyLOSczpl7eXDD/yVTjD67eBb5BTRRieLcFmHRToj4sqrMZpsSMNkauuOP+Dzn+dvx
LyITei1j/E1ZXpCJNPQykHC5t3X/QWXL69icBsIlzuXT5rmBNmo7Pue0gnpT8tPxKQaytwMNRTEP
v8LGS1B0Dz4snBNAf7pN/lwyIioOsJc3FmZNIgFiPOHX0cOLlC9ylESx5/E3Qr7pd+plifdR9noA
anPj3HHge8SCqjRj72qtMwjL5bq1lWPVZEEDaiDu479vty9UAftGPiWgzvwPrj2k/1whHg3clRoN
uZuvTEO25TWUkWibHboTkX3UwaaYIyoNISZgNxQoa5VhGjhDmjkodcp9CXYO7idcRaOi+ITC2vW7
C5cnIFq+AyN+3fP15wo5SGppF87fXUwP2Ko5sotEmKd27OHPYUZATQDtzJ5Ayp3talKgGI9qBLm4
PfVPkfmRWV7BzTbrFucceVQkn2B/viO2UzVgl5kfs+BvBRFn2DPmAGrQcZKkEyDSWADMlgMRKzx9
qZ0LzvIbLxFwWsTurWLfaiLxqOt+pFYOd63JCYHPpjMsyWBsPd8fNkJL6y85CRYKtpqWB6UQe5G9
uEAGlIuwSkBkJXGPAf1j8bpAut9bC7VjW33WM+mUqLfS44iRsBwKKGM1UWINqr89AEznuDp0f03P
qreb21F7k42Q+7JC8ng8t8P/JSVMZiH1m+Ql+I2vo+GKiL7Fxfbwbe+BGjyLH5LReRM2s/owXcL3
iKIBHmRJZ240P/t3YBaz8wwZHQJzNvUKPdegGnWl2ocHGZ9K4eCAVFpqhhAgxBPfEbdCT389iLZH
3Wu2ZTSTQUOTD95mHG5Rkg5DKKLrKYZ7EKRyRbv4NH+Y7bAArxcxXiuEAvaXefFsSfEMtpQJE7yE
2RMDOhnxBaKl90uEoI2+D2oy5YP5K0eL4XRDwx6cpg1PkZlEyTGDWknDe87BbMI0kfhoHbEE49JM
dXhPfIwO+kcg9rKq5OOjwMdCqsv9sGQdQGhP/b0vHo+DZClHm2edmqulHpudB+KTmu30BrIIZKHC
4ypxwKbXzYdiBpdRe7T52ZGpA/uOqi1Pog9/vCUT75sOvzOnlIzJ9ZM1tzOuBBJG79GXg8ssJK6N
LCdJgwBvRS/Z7fxT5uAEJvUa01URhV2DhhnaDL//7r2oRu1zsg1AP9Zr4AgpRm7FyyLE8TDYgW0x
zIb6bqffWsBD1UiYRKYLq2rGbEfCVaD+eZoIdQWL14gr70cvDD58KrfbP3Ey9jqfvVXib4JgOeGD
i9FXepmV1gLlR9xTOP8W0pEJsYQ53/c/v3uTUpEfyt4Nyenb4OduKPcgQHRNDS1KE6sAz5TjWwuo
XxNUY6oHpMq+AgGXGncAY7F1P2zC59uJcnDdqJo2ODLFUQVEGy+kjZ5HHDtD0CnrQdvEdsXm75HI
leEon2BLbj6/kwHvgytXSHmI0dBRP0aMBh67FhomEQ0vuLRHRLSL1Aq9aHKGXPWNy96avOlUMn7x
v1+W/dbkwIS6r9CFr1up98trYrzQ8Drxbr6eRbK4RDks450DAA5VbsNZIzKzoys3n68rz9bBm+sI
ysPOAseOSAhl965cRhmwl3O664wAAncItaV9guYAb865YqiMs6DOCruYFsmrvIj1FjN/S5u96LQi
ss/XReLYm78+gjFhdlcjdFyg3gqfZtGIxVKvnhWttDeQclqq/fgQbyywynV4tTeq/qMSTj5ncfrF
/FeOmzYhfqdSqyWD1eg9RIh1d1C7Wad5/B4LrZFpJq4UckpYJjt5a8tLuMvbsY4h0sIUxvtQCHWS
bKqQU0Fi/jukKn4sxSfoEME4c2WgaYD9QDRqfutE/jrC77D4peEbn4eif8Es5VCQ4azAkLp6T8Je
NiulJKUrxzrfMeVFPhGyGhhs8gXCxYae2YQHB74XWEOqEjUT1Yfw/Hc/dmWAemWPPkgH+BNb1iow
n47b3Fiv9JvKeemYC0LxpR8ME4SkRJ8S4SCzljn7gqVZqk1/2XKDZ0YtsfyROQPULM+8mqEEypj9
yBDY23I41Knm7nlNXmoV0fHJ0f/sBj+QAlCc2I2BpApbIcRvRxof6N/hxTcARUdDZ0XmJYViOjuQ
bzP1pat7DUjzSDjBO4kZqo/IjamNbmZLOGqkHFLKTyuIFu6sK/CJIEJdQEEy3ZjBh0z9wooexW73
3ufJMXSaBJmxZdN5O3sPhRk/SIGK5lFo0WBiLsgi7lRo4Gp9CfxeynrhtocOgDzwZ6nwNC6EQWER
t5/4s/F2QIBV3aUKMdB0YgoqZRIJ+0FAX7ehLsQApKOXxhug8BOtPMOyOnpd4pdmI3kXL3D5xDPF
weq4NQESaPsOlmv2Q2x/yEV5SUiXgKEfNhW7RKwDnKtsxKuMfiKdd/6LykNoMAfihLqgAgI3k4yQ
e98OISfGxnSy5nmDB4naRn7TLxCjzRQ9mTM7PVDJ7me2V+pvKFDGSSEZNZeeaDEM0DWUUC9sZC3l
5LnbK8c4cz+azecdu50hjZJQYm3UoQmZvasUrqhYcvEqnarc/w0cCW4I28NdUC7/g8wlYGYI4qmr
issJyQUk1BSo3ZYE4tgIkEOw4bk3jmJCqBGYForEfPCWuM/ZtLq2yyhuQC4qzj2rN9JmmurkeBc0
3tzUNS3e1grIfG78UiRNteb/MPRpLHEj1M4t1nAK+qkujwZq6Z8uafd9HT8cCZL94YfxliS9Ijjg
Vsrx5lLZe7kbR1mRHBAtj1mRjknWsBXGRRyABhVxXt2rWsqUe24ufYFuduMmTyumyZxuLvOUpCrj
oxTONZK+VL2ouX0medK2abuSwQ33Zt7zPixWswIKcjDaY1kiu7RIGl9cCTvtRn0Zb+MraJDb30lw
4eshR+XFBIQGi1djjxZ/5N2iGQ0iijutpCXQVWQ2JwMdZK6nh2kNXyBoNTQwBvsxXIztAb59G7BU
ScWUpqmoXxNGUfELBm3tfR/NXmVYC3nArmSwz/T+ZfI5Lb+QHli+Z/hBRfeAOn5Njd94fzaU8asS
wMIEWWhOVKTzG24wsKPWMZaTActIp27CrvFGiFVTPDUT6b+tvcCTQZ+6YkIc+gLWbcI1/SxfuIgV
QIQtHd4m6wvOdGH12l+IbGygH6IbmhzOmwxCp/MOv1YKe5XqDT4CZfiWDD722M1sMxJN6LdDZolO
6FZTajhF6KLIZ7N4AgqC41hTD1FLQjUFPFKcGCaI9ihc4/MOtwvSe/WmHBY+2vwVE6S6thoJ/AoX
/HXMaecwT8hA+igyCVhTlvZ9OXz7sV7UTLtJiQ1AqxN0c4IrnMvK1o5ao6bEpJTX7PtBXv5z19dr
9GeFyBBFCo4tUnAn6UD85BTG5w3xitVDcgTlCeAVykuJC8B3yt7hPuXP5PUYGIDecf9q6Po9PDus
0ZEhbAcQ3v2O9SA2H3gogvsXOfhckRb92dfvPU/dmdWKuHlOXNpeWVmKMtuMwF8Tzkh1C8v8GUSc
T2AyqCVlW/FW5qzVhnbBUZNNGN22iRlmJ/wqecxh8fU1EZH1/WXDFtjWWBi6nZFvDPxMQrncOlG8
W+FZdg6OqxL6565eMIE0MjrTg7/VYwfJtzEy5x7DbayQVT1ScAS4quRHIMo2O2IK0vDE7kHY5TV1
AAw20yQrJmC1IBxv6Da+qip39RJUaY0UW+7CU0azK84YARk3pieCz9K+leqxPNQrQwSXf9Izmk5o
z0OzzgrMUXPuqP43w4PWshFIednuBLhnE6uGVyvAUvDc358MEb72Vzd9jmfrWYnYL8SZt5Wb4s8g
kgug/nsJ9PXffeQB5Dkb4mZJTRJ5dRIsgzuQd4OPXkr6h5CffpU2MX6SobHhLKXW7lA6TPtAR/GX
Mp9QvB+IopsSHJub+MGLZ0qD7TCfD+BZeW8QDDqZGkkCePKGoPI914sRPvH3AQaaxawEasLrk1lv
MeCkPmKJxD+PhMaV/V92A/F9i8g1JY2YdNviEfkmL3AX5kDuRSo1l0XhbZdACTUxQWJtwCpWf364
c+R2enztAlTt2JfQtXiEwMzgM61QSGUDorIQmSBpaCd4nEO1agB16sLf8XJ1e/i6QSzhcr/8Zega
h112GT+wBOaIh+jgBp6XCIoqAHoGJDu34IUDlde1D/4DKXER87K/a1P2a/El5EbPPEjMBpKm092X
aP1Noynd2o5UpQG+nbkW3q52tSPPAKBoRQ63RMiIO15j081x3ZNA2z9uAVX4OBFr8RYPPuQdUvM5
eCDYVg9KNzc9NT2nrncZRA8q95GQwsGjChRUViUUkMb6AHtSd3kqTA0QYZwQ1cvlEUV1ulM0PvTB
DnckNoCEfetqa6xWJdPgvdMMeNe2ADF9WQzoGX9/cS6rSi+mCqoqDet91/8cf3bosUu2r8GBPFra
+kcRrcUIxXMkF9bn7RYVsrzAu+IMtx6gIwvaOrK7IydgfW9Xi7T0FIxUXs24QIjT306AQbZURnvK
ffMc1bDKvfkNhIN/sWHHtFl6mWlSZ52kl11gWEurn93WIi3XZxTAsJbfDWPfR0IOBZ2Wn32jbX5N
B3zx4/TkYytNlHHkzrg6rnwsj/FYSJ8sYyOXjcr/7OVzAAfg+3poWvBEpu8eIuwV/l2ZIy6YCuQY
zFEpBWyI1y3yn+KlOSM1kP088sYFkM1D3MkdN61Ydx8f8laucdnGSEhUUdtTpgg0hux6kIeUWQc1
SgNJVNIvavwEy6HiaZ0TNIVUuD0uYr+alTSrEX/c7FmS6+mJ8alkNlxzPa3Y9Q/G00BTKRQAdXzZ
Lp3mWK13ihai03Qhv4GhOXkEUV9HK78WpE8YWO8grkeRM2C0P2Ixm0I1JEIf23BHKo0OiOBaW8BJ
+htCF7CHsdopZbbVPSqUtex6ec6VqFolmP9Son0MtK6mvYk+ZFUDadXSm3nqmnBNbV+9F1uAOTi4
c2+vPFHvmmWU8mWW+EFsNDOMV3nrnywE02ePwyv8ryYR6ixyfh41NyQ0iNxiNEfTmgycKI6mnN1q
C9q4s/yiLkUT7AUsG8RIyZ1ekIiA8iahD7U9pL4uf+GALovN7IYbLhTN8r9OazgDOJcQsZpq7iWb
09f2tJa59i1vYGZqhYY6BB0ibIh8E7GR7t+rP5jwLa93H3nW7Bih4KXvkPHVqNg6UmvgUqbrD8b4
VQGEmat6uY3+yVYsUCU1NB2cSeCJdi0z+nQyQ/YCnTDP31HvYCxfAQmrWLerZP5MB2mcGmYAgsYo
RHoA1TKx0+adTbMfmK3onMC6r7b22E7boqclxXNSX5guL9bVu5Ghy9UMfAxBnoH52huUCqTP39rS
XQS6ZbYR8VZByyovFfb+Sd095V4d52XaKU3M6GaNZfhtwdiK43ftVsXcfxxsy3mcqJw+k9rQ26Qu
YV2tV6j8Lp5RAB3L++7pYPEEZ40iSRhwfyC/ubNg8eXOJWw34LpJeottTcsKL7cl5TEo3FOk8kpX
441mJGQbGb9EOSERgoieAPXm7+e+ZDJM/Sow91WJjeD5Aw1v3E4Mbj+t0JcM5epKILVk2MSvW0IU
ieruVfborYsqscZBSrnI31uf3aOrfqgiwnyAZzr3DMzVsIAhUwQi8pNAs4IzpNXSoshy27ZoS3rF
tSTRv34XFymU3oqNCrIqaibAp60pr8CBXcvYooof3/QMg6N/on+pyrC+z7nlWBXReQOkxoKQ3GwE
k6siU4kIWhYqKIo3Gmh7rlYhTbCbKXGWCTp81ssZ3x9qxb5l4cpPA+8eN814Uv4vDYlQlrBrzH8w
G+jSHODG7XxOsqHzzKQpirSB10NEOhOpolFFxFb4KvbPd/WnRjNA6rCUGXVqT0rkopg5A2Uk05iv
N4Dn9Y6D6HsUli+vcTw9M/Pn9Hbfm5Fl7Ool1jBt/gZeLSenBZLKFD49eU6tJ0BedKdLPnunlLGR
qum2KYB2nM8A5hN31ItY1X/D18pwoZdmMBXrwLb9e5nkZzrKwciAv11SDwrOlVflwsiNUAI9DHdw
ug+C1DyWsJU/ZY1sXt4CB/sc6bztipqiFiWxqx4Q1p0D1hgZcb6/HBXrm6PS9drMFMhznWbYzWH9
NTs6CfobiVcY81yexkFrrdpA7LGgwSpySd2pJHWZmNsD0GicctL6AkCuY/DEp5WocHdHhO0NjyT0
FDC6o8RAo8d+635Eu0GrlXGe5u2qj7lD4vEOl51NAcjzVGK382tf8BXfPbUIFo8KjSQkHga9nzJc
OYpcYo0ZmUB4hAYLSU4T5e0PATQbMYYsqFy3Ja+2sbxZmvomzBA56r6btLU/BuUgdYYO+8IP9cKD
um3vLL3N75CUtj016zdNxfBhkQdGss8HTwPAKieRjEgAP41rAxmm9EQN4vH8zhCsGjVWHobCgIq8
D20mw2+KBcKTUZx25Q0EbL9mGKtL+h/kh+bCxgXqKSfj9psrVNzHS+fPRU3i3CZkirxMpfkZmh2u
TaWnzQARJJOPndAAF7mJihur7letmrDsfxwgI1jDB3KF2CnEVO5GzNHU3ETaqaXru+XjBVDIwcMY
6xP5ptBsVAYkgqZZ5XoC9wv3YE/BK4Ic1+nRhmkseiSstkMiqEkKlSF2oSp7J5ji/7cMhj9OLVMT
j/1vHWFZcOIXGifAo4XR/J0ORZoyjEZTsMxJsOIkrBQ12uibk9sPI0S5hVJCkGo7zzmo1mR/TOMb
jm5OEoZMJrIYK0MOlWZrY/EF/zkgPxHo8DHB/foDqtkG4ynzAj9Iloukt1FdoG2PY36gMUiZZXu1
qPr//J+Myu5Fg1rfuJwmWTLeyHmpXc4S3A5Mu6QoORNbUSoZ9O2LKPQ7VMMxM9dd6ne4EBBvOfRo
Aez3ozTU26VNauk2NDU7L8BHd0sC8k+AyxXm+cXKJi/heOyPahCroULXlKVFimcqH3hXN70P59Wo
9TUOg/cdc3gtCs37IS9PE7eiUfSVj6vohFPhy5qKhmHnRxkPLt/lX84Kb5zZju6KW+ybjP0Ylff4
Hu39BqmwItLsLd5Edv7fppkMR7l9VP8+COcbvHUJov6ABEVNHocYvHBoNAs0MgVRRNdZC9yGh280
RzRQ5SuDgwuznQuWjsGK4rftD6lWIhyIKFYrR0Od3tsl8mdgluDHydUdnZEO+k2kD23xf1iq+GS+
8CqDMAqxdb6ExgcjIUhIVmJpGLvKS72aed9/xl3xwgnyZ4bZpqjEzGt3O7gZICgyzjD1Lx1gw3bH
jb8wBn/WLZpsYU2hr4dAK8NHi2jDybdLdquaUDWEdAX6hufWMY/Ij/ptJ+/0T2YEz4+3droyM6Se
Fe2+5yh3UE/mQl/HNxxzeW3Lo7O1lDVd7MrU3CtluATyTUxgcNG4jID9z2yYmpiYUYW7zk1c3vT0
BGL0Z6g7j2j47wGTw9jILAWvxJ+Et79ZzKXDslCuu0Ee4eNiQ0x0LXmMnT1cd8Kwhh4BrlQfYS2K
NE23EoUbkJBVmRCq4agXIDU/o9RUKwhmPNit0ANYcCLzUGaJQn3RdVCoRUL6TZVrtkMObfhVbiwu
5R4tPiK9wzZaPEuDbulr8URhhH6XNQ2CwDiTEgftzr1DtxakpJQ/MLVDdhFhKaKGsJoH+Q+zPuH0
Lrku+mX7npT6Ky//yQ8/zNquHhnoZXQKsyBQ6p28NUBKNxIdnX1NPlbZbrYZmop6VTsX01T3WnEn
zJVjH12L8r1nGH23XtGR0vE2+bmN+vkdko6gHszIbAvCo3GddEnoSOpQSoA1ddzdCNspjl3dpMcN
t0RZBYBHWwIpR8XqVrRhok37VpKd6RG99/tbi+c9iIDUKQfaaeYbFXpro1wF5ap+xsOHFbuFcR0u
H45vWAO+MNXAFq3vSm2VhCmb0Dg6NldSEV/UX1rQq22/9C7ZCksTF8WdTFDc0TssU/KRjd4QDrKk
zXc6FAPny1fCQbr0IfXQQaoyZnpmZQGb1cdO5eSqr851CRxYV5Hjbu7NqNl1DswPETpuAOS89AA4
si8pHfm2ZmrttyMqN7EIog7EUh2aHGmfu5JGMiNp89rV5Mk14WpSj1byLQvb4STtXq9tHSFR+0kX
JJH4fzVynSczly7Ds2Nj+fPDMeZfq9hGHpQwpVhkcqcJDfYZ4AO5VmN9PioyGkWMu/c2g3NAB7Bf
LOFP5PWpTOZ0PA70lCcVMimeKgZY5h/OSFE0wH7Uvye6+7pqGbsawnrvAgcab5KQiaZcR8+rWjab
QsrQHr1ijqjNE1Fee6fMtIgy/Z6Gwp57JsIIe62eYAhGA7wiOA+Jri9rR45+iRV4EwnvzphsWBpC
LshJfzgCQdWey6cngmYWRvq1XQcB6XtrBy2D64XCgK2fBINd8LTD8omc3Ghmbf/UDL/O3nK8Kngp
RBXAhIB2w1RQBzRvesuMBitXArHM3f+oMQy7EoocMd20ahAUT8cGiONrhyW6TIKlugcU9eTy4avu
YutnIgt8+Rwk4mnNFy2HTSKIKnaTUppYcid6fwQ1uTAhtaBexBZxK+FHjmamCjo228Sv3SLA3Ixh
nIE7ol3eQIfQcYxH27rWzshOBr9raoO1WqQS3MILxdrxo+BDv91y4GDx2UfiOWIUNWmqhXBGcKEv
eZWmr6YpoM4EywZQAGMLfrBT5D73C1uyaG25zE9vOYC+zoz2z5+TWatriya0bD2sflatT+Gx82/e
d92pl85i57qTwEIOOpz+JNcOmF3skqQNz4hvpHTtwAtsUJC6nBpab/AfIXfGOYMleMLqwJMTDwcA
bu6akrDx+/KF+BjmUl6b+hG6VZyeL8toMbtQe+FMh2+DM8sMkv26zwn9loIWtUBhbWDCSzZKjSWQ
VnNljlhOGUY0xMR07q2c0RXVjKXB10kOopz2UCD0HXkqcjWKVBKMuqv7Ngh1HgqHQa2wAiRcsp+i
rMeVD7hO3lTesx1iRxW/eaTtSMDeoWHCfMqBlA6GlFLV6SGHyK0vZRdZWsXcxKxhD12RRIr8YukP
6y5gxV/KArJo4oXT3tC4EAMzyZiEbksPjatapHPpHUkMGf1KFwHxjZ9OsQsW6pbZQdbk7yEHnkzE
sH7Imdmn0YdPCbkIMq7zJwNzMf5JevlLLKOdtdzKYvYyrXA4czx/Tv2apUVG1qceCw9UR+ou9ruv
yCTJGcXN8gWJJATIMyjpm4VkgbGm/Agtp/PVxS7ytrL7RaXKjuBhd/7znWFcx0MuFZzoDCzeiXxY
zBC4k3eubtxxCy1GREMYkR/aKnL/EOeyomZMIUISM8aUwYrV3ilaznWYhz9ol7cgPLSDIgycGc4K
P8dor9+IzcYG0d9/LOnEeHPY1twvexfm3ky79ESUMLpefIPgIouFuGGXOH2oMUC0vzf19s+P0T37
TRJdryB3DFFDRPEWivskS9RoyhVcgTEvsuib601ifPTRA1JJEkGBcUaU+zZD4mWudmmYFeJX9Dg1
Hpa5SfUC6zVUje3bfjWaTRbrdWQjRmcyzUGxL+QB2YOaz5f2lcav+g2twknIMR7z5SyPznQtxvS7
S3FMjbD2/3shODxbr0Gne1hPz1rdFqSMtYMi/qVOTg8K/cavJwuNrvYSQtybA76HDH09v3xp/KC+
6VrVsJldgMFXGs2/mYJotidvoGaHgaHaCmmhFr3jK1xfGgR5fLBCeKqqHzK6Dc6wQGTAokI2mb3S
1BfcXTXhhXj++JXLaNMt1fhreVL/sIW/pROi1Cw3j/pIv7a9jCzl0ghbNMP158qOddUVJMqwmoVN
sxuhkyDdMOKjjnTu3crqsTKurkUxGvHPDwZgajH80w3SjGbKzcDEig6m5QjftbZu+lTV72p/5XtQ
UGklbWIFpbMwaEQ50XdZPGRk4BVXRtly4Z/kndkTIuevJOtAv8+90wRyb/wgiCvKD7KCgCasONmy
1jKUPRLxIbWHzdCE32ojlCEndwYzsWyNJ588rntP2I896l00WdKDX5A8VWjFsfcgE61Hw7/cJtgQ
73s6FxiZFL2abpqXDbVYtdoLsQcLX8/ZLLf9yKBBPQ0Qg0g6bT8UumfbXLwWe7U8lzUP11NxFgV3
luEkddXJdXNozATJPSgA62Kb2J2fHIK5jb0LVkJ7SXL6rFZpUpnifW86ZJFSoNsftYWb+RYN4H7q
s4xNDxPOSo9glYnHmjSBeNs/zVsPyGRwiAx6k/GmW63rvyXIOH/DKxV/otMtxNS5OQdiJSzrGT5j
AE0phbiDoeazWnTAAbJ1UvReKPvmVVtNc77ViwIhLgdgBt3RSosUxK0cp8PahCpLBWrVwD1vfh+B
rTemHQZCwXXWzG1MJWz8un0z1r81s1vy57Inaz+bgEWyjDIBCdlMb8nwt3UdDFtYuKiLAb1xacf8
fUTwO4TN+2QxVPgCF9VW3txhunC366VwldphnFyyTzdB8m5XTEw/A+JhPvEi6ihVZ8F+ex5ZhehS
uT7aYbhBSloj95GZG1RFshFhFsQef3gPkm4oMI9Qu+TJIGaCFkR7jr0YKFHws5S7Seyz2YuuObDy
O9F8wT60DyU8TNub2uGzm/Eb2WuR3hT6A+H5vFcYp0MKpqTzRoMdKWsBGRR4BxsQa/1m7+fcstqx
f/uarZDrpHhqQtjU951ToPN+8FtcnG3b5KdF2XmP8in6oZf2BQxvEmhCYG/aYZSEBUoxpuSQj6JS
MtAoe0pnxLtpMlsPbJnHFjCPW5BXSW7lGPbJIO94TpLiJfebwDfYkUaDv7PAEuXESvLToa8fLZxT
Bl3XFW8uNNoONpLFpGqKV7JreS940nWQxqnG85/PiyJ0IwMz2jhVQK80qcTd8MeEe+Zvt55YuFOZ
RU7uFFIilXLCeHRntVcDasDXZpPAnfCh9ohsAfmNZWQjetkTuPbyHEQB1qoeMYYioSocijrr6B2G
SVX10cd4pZLglyJIRIIFs5nVxkmDOgzWM+CcWMwk0gfXD4/bReTNfbUwUQSbP9AB3oH902m8U6Ou
bzq5+mUTdMrINYrDmu4qkbeqYjYeOtXg+oEy/TLg2LgQ7NHIrIRNrbYU4FTa5045UPXQhaBWulqG
eqO1xeRiBjUjxCZZ+sfH+EEmhRTRp5ipqdKO5J0zZTIbNRmDJny4dlBQsaG4Y0N4QfDQK24KOAyU
MMansDj2XRU4ByEDwC1ui9jlIlMfnlxtNsVF5cDg2u5d3S83MXp0RCEWPWvWMCYZkXCvm6POw2Hp
95LSr+rUwykoVWdVAh1qTB0oJbDzCJmABjVUcgeOczu2HYpaJ1vyuSLzd5r7Z7+7BfiCocVqTFDj
qpEl8lWhX6fb9q9eKikI2iVT9T4yJBhYJyALnHD+rsWz5SQEQIiyHGPNEP0tf/7RpAZnACx5IJJH
a5a6bmVmgb88HumIeOeF2kkyHhkQHXe6vw5ghCcx4ZxGHpmCaBz0W5Sz6h8GkKn8vu/qz25alK1B
P75isJrxVufi/J660N6LmVzgtNKkEMtHIXri6g3XwP21RQUg7kFl9x5WNtV0w7iHIUhT4WllwSma
mub+/pTsFeXR7ST8jAEAwimIw1g/9FVnGyukk1JK2aLvu880WerzPMed/kK/f/62IaBWoj369Y4N
uSam4Vx0yBmHqTonoXZ1ijMYDw2VI+P/ouZXMtQkp7A/5QKaf71mbjz71Epi7x5v0nGZq1Db2V/r
Vlo0Xp8e6jHF90GltlOg8awxZicrsv9obrF1JZgbBXpYUY7X3PAKn3DCWpewtcOixW9ncUN20xD1
NDzkzVE8y08obGxz44g96VnjvS4KOhykeL9sYuaOURFZonJcIz7/bQ/+A3Kc1btucovjB+PSDqzJ
chcuUpME4qpnKV5kDoDlM6kjcvViBJ7gzT7Mh5AvwcxziBiJtXCA+3pv0knqJOZDmgEYkILexcVu
7bWASpGqAs/5JrUMMatUi5CczzUntsF6YCrimmmwM8o10oCIzidYVVcpLzk/Rg5V1wa0vn4kqjqr
aj0Y+4hB2cDoApd9rGXXiCrLRvx/qaj3NvtPwol/GH+mPzrpNCPli3X1kQb1BupPh6lXXGX/n9od
1cmC7YS5yvBREC1ox8evRISYikUyq8W13ty08ESncvJN94buuZMiV0AHc5l2qn4MXzFBAHHmZR9z
SzgW0nbmh28lQ9f7oWSfCqPIUGotLoTqCKBNM05NbzM0fygOIK8UPL+F9PHss0VsFgr4S1J7AfFj
zFM/cem+B8u+LgVXkjaHnJd/aHoSN2wSBl/0xacIOVyZIf3W4pzAMK9h6MvKbAIO7BppukaT86u8
14TBmwuHz7CkEvtBXygWj7nH+/Ik8KtsJwUmDAFv+sBxtQDwpp6nr0qbR/Fzlma1IBKz/Dq88m8z
VYPHSVyoj5APo8qaqCR8Dupph3y6lLLSQ/fAm+iISUsWl1qgXMSqid1z17+lJuGc4mroPTMBG7H8
p4Xntpglok2icK3dMD0oaXSMH5RKkyCKklLRaAbpvcnIjnN9IPhYrddbnFzgM4ZToeIvYor+0Ubf
zTBKFcAwIJM3gw3WB6uPBW18Tsag+tA54WvmuOnwM2FrGhTEsiAbkxm8SalfHCG0k2Px15oxp8Jl
hxmt8kKyZW48XxHf6c5uSKeIDYDAkjm5EpzQ5RgcmCgGybwqy6/YQiWRQs8Z/gP6HH2D4G1sC6jJ
wpHqo0ny4lQHUckmJDtcREwyAVNPDIHWJGkCF5jYPhMozzpOXEj1B3v6XuTuYDJUsw4Uek7xoRto
mzASQQpevI+/VRg5AWeZDnW3DEkexrl/w4NmAC9YzVtAogMCGuLwX2PUtYmnooTG1U9HUAHOjni6
YX5DyxAdvKV2h78DUNEqSpnDxNEut3TJSBSkbzDJFg92qrK3lPA+bjNG1xUdUS3T+H95yZCt49Gh
GG4wBZjolLOGZptewZLYeE0gVAJkswwmrmXhz6XF+KTuraNeCttkqw0/LbNU1o4PWUnXa8LHcjUD
JrrUv2SaTpaGdw3jcKKF1S/XDil7jIeQjlW4aHNn2a1y34IntIzqqHjfKd1XkthiFJdTO3eCLF4M
wyCI1lF5BwIh4YxvHRrLwmSoJNd8ZkRnYb1ob7y3p/x13whYQ54Oeu8dshiUBJnfO6aFaEM5LzNb
ahYV2fBOcMBd3AAMBj/KyEOlldjeax5n//qoUJ1bDyRH8MGBeBi6qRWf1rvU74NODuItJWlo3uck
ToOSeaq/DXtODu0ypLnIjZUDv7l741r2Y5Z5uVcG/8HEJM61fzpQgYuH9pPi3nJfHHiTdbopKhlh
YFxiooM2SdLo1NXYQMIkEnnhs1TDIkx43WBlOVEttuv0yq+jGeUX3gu6ndcw4kBhnOzZWz5AbIKv
gzIl7Ao3f47LQ0y+B5vTRj1b6Z/iRRFPdRELC+i3kFuCQ5zB4KG8/b9La7oArnJcVmUfhDz6+cnx
R7eNAjuEocSCAjKMl0+NHUdvfQ05+ZO7Dfl3bOe8EvvAdtX0gCxOvKBPALxmMwD++Lfjcj62WSeX
bwOrtnIiLNgKqdNInACUEUPDsDgtwy5ozEcjTINa1XuHFIKQN5gVzdFn3aRhYi1o1PXHEhhVGjVx
QFCHpghbcVSfnkr54WLnbJrvA41MVOtnEvoJ82xbXf98LrpHUpNGbuaRLhHmYFdoie0PPcJet8dY
fA6WgPxNmK0YISNnHlmzoNbUnaGgYuIPhf/GpRciwL8KoXEEDrQvUQxfAbcfBJpqB1z19r1ooM0r
rcEJAUFucMk8wfCLS0/MGycYQYi4NfjI7ZiI/4WvtJ/27E40Z52w/dIvxBo+INTG3emhqNMyLqX0
oFEceVUPtJDv1vwhRBl79qKND8xEU47/XtM1wILGtlPzd/GknwQUGi4eHgS9Hi14p95hSD2msX+8
pnNNKJDcJdZnGwtgEiVvyY24M8ge4eiBHR6+dwnE5fNgcrwl2V+FegDxrcWrG5wlH1dyHyYsQ/a+
dUZ43aUfcGWsuJoLsM6AM7FcOeZZUKgdp9hSk4NIWMD6EpqBVBsVJN7rXte5LuaXYj6UN+T2p7ai
CnDGqIF22RyHJEiDiYhi39W6xqKW9J8m9nhJMgqSdT2FV+atTTyXCREpBDWPFiWXd4uDBjvSV22d
meooBQ9m01hLHbu9XgLApJhqJUEADzf93P38dixc+kogQ9Gz79oXQtqt4zpL2oN5aDaIXis7iRCK
wREE3Tt+HOmof3FjxrHj3kgRbLoBxDxfAABq939hnoso+O43MwQYjGl97dmVxdXkAiwLkpTjCerq
rhb5PzAlr7nFN+UYSOAvtt0cMuJ562Ga2s2V8fGASeJEqsTgrSbip5ddIaenb+wwAx7NvYes/26c
YbkjuY5vWDF/hCxAGdfdx5TYhfRZ/sc1RbO2cL37uPTeH7Xlpdo/xdxILJFVrRtS16a66h+yJj+3
4l3p3JPBfL6PRpA+x70Emlq7gSMysMmXoatfw4N1NdI071ZCy3832Gxf7TSsRQDfUe1jeKAoLL1I
93O4fvQK44j1dXbF+bxIDDX4CAjdSpeyaRGcRX3IbkPLFXesXQDhgCZsZzyAKGfRSfi/K6eczkUE
w8XhK8yWYJ6nqynt0HBcDD6i23Cc1S3CmhqFup7Nn282os69NxnHP/oPrsijiv6LJdVafdcxqM9I
ijZugt1oTSAG3W6Es8DXXvOj45ZnqojOojQ3ro7omJdMOhXRVwIHxX0ABro94GnJf6kTLMeIYjIx
vQdQEuVJzDPaSUQ0SECI9iM6E66lRPHOYl6J1O8veMtBDGe1BTh1sKMJR4MDFXLnnr/oWwEofW+g
NL+YerhZE7a46CmVhP17xi8uKs/j58110IRoo3pv8WKNybhllnGnGE/532xIi5kS+5VIOS7dg9bn
yfgsHDn6XAM+EsFiVmSZTBqRQfqZ7gwZoqgjDcOH1dAAkrNmv39+jo+jIKoE18CrxZq3qye/f35e
eRVDRAIYuZktcnho7N8bTlzDVl4AXUjfMM3hC+ogIhx2Rq+NwsmHCQiq6SHUm5WMZaKYWJJE6y4B
xYaOj2tzyv//4EQv/KKlpjWPDLjZK3zUS8w3UOwANIt+HT6vHCharUJDzBk98PwEDrUOUQBAi3gO
bQhrLnRjH1XLv7shbCZlDSgEw+bsc8pde4FMkl5LsxAOo5ukXQ/MXUPoVu0pgzQnWzL/APDwhF4N
8EZAQ/+C5N7XuO+JgAj9gZqUUke04f+M5acKorUJVNOubrZ0QOLLs4KAbcCQcS2HPQQq2BcdNTvt
ASUtO6lt5HjbtCM2xKgsDbDrqMZBZLeo8M7Uxs3xEyN/1/Qykw3H4L1oMalIzrBIyBfDacvld8fW
65xJTAwQlVunsC0wRj+EUG7uttDZfdPMiTW0HcOQhUCDPcbCEKUnl3g/35jOuG0BQr1jS/XhlMN5
liLEh5hBvYyLfZrkI3Rj9bxf0akvSv5y4bTqO5G51qxumxzPNnfW9wiaqrIUey6rSsY3yRnbz/u5
w/plMqYSXj6n3LgvkF+dHwumNA5BOQIwkz4cCAkNYzJjuZ7yCyDGfur2M//0VHQ5MQZdUUwa6w38
Pqb35r40uPLZl6rfu/bWUauOdfB7ED83/89msf6I/VSw1Sa94YFk9pmWZLuK5JPQDBktovw6UevC
hF8oHfVKfZg+NYsQwEJ79Qeo9dMr7qR2ai7EM5zyPwRK5eReFlnI0Gqz/dxZD1bsZHFdZkS+0Omy
r5ZBYerkY6PNThTvcVnLjCvixHSgDxXXjbYR01gDjG7u4UzOQ+QAUjy0tVN//gzfWypb6XD0h9BQ
0K9QrTM9TEfEkRW2HViECodS3nUIsIkPc1ZYf5T5AIWa3RoIiVRdWdUZ1+XUfH4D2TZ9QYvwjSoW
r67hHaqYKSnYneiOJJp5Woet1oK8/Dnp8KbNyDDTlWWiDr/6Ei/NXUmkoz9RnX+F0NrwU4oe9Oul
L0TeZxKQgc4sXfSlGSpsb5xmCW74ejmXUnPiaHF80ogsjxayiiVMfJDpaVjJEh+1pl1hBqR2qHgv
/RK6KxZRXUDSlQbsjWnY4/vZ5E/iwTiXZABQ14BuNDOjIO/2XIZJXKSberL9CQXEsW/6qfoERyGO
AgQqiGom+OIpFy2p6c/KbGzDNmSY0DboqfmCPGSHHpdRYs4J+iohrZREaUywDijVGetERg9lWMwX
xQRelQuvT6BOBgvfOxeNsfnEKOyaid2aLpc/EHsyv0nqiIX7LTInkt+f4Sho5YO8D4GVIgw1rSZW
8o7fPhpr1vPIcgsfBZ2cGnMyUELZo3GwPIujxGUniFM6MTxN+EDnnTi77LA6BrxnA5UryRLucauL
8NCDVfw7ys5lKEF7x0tVLFVKecpnnYF6IMzY8jmHAmHunzvSE6VHYIuTsw+7/RLWLBHd37qExFaV
0CBQTzSemO1Xc4Y8gArLAaxqxf/egFgOT018eXzWuHCeL5qhqVKj3c+FBlKWsj/9rnRpU2js5gP9
/6eDxmPN+jbel5xm4xYU15dLPYmrL+LBAaCN5PSJ6cYHhpffmiN9seyfvPb+o7Tvd/nKCADrUNmh
IrNSeWnep5+yRI/l8UuS46B0sZcqjyhjMbF5qrEg6+4efzwVESsP5jgP7ihUsyH5Hx/9x+LaFbfz
kRKsMz1eV92X6+6axNt8YWy5ddwJ7QnCNiLvJtI0Q2eYfTtPl+9PJ4M1PRK1qqcup3TkRnQA/9Xj
oAz+xC87BUYILdrLMh/EwB01IsLcKynuROoi40y0bEldaebbQQDz5EiTVJRy9bdlBioCv9paCx0w
+gEv2MtjtsjUt48NhG+nW9dD/FfBVleiSdcX6kCAJRbcGV95DtA5BOkHcx64sVZExL5LgrN6bX/N
GVcRCifKdAla51CBg7FUrJInIdw06WFAM7OFacMnIBLkziliMojrwwqu3PrlIqJBhU+NuYIFoXPh
DIE+NKpUpnVbGjc4GUho+0SkUOcFMkdtp4aAN2NixBv9x8BKS4ec5Zk43RdkdAWaz14cxcp4fbUo
5ZU8eJNVHJR2BMwI+vFFhnDdS+iBJVS6WaaFGQvZDAAFxuPToOXiUEaOuoaR/nkRNYQMXymd8fPk
eZMurYa8WWTyNLhCenIBKmxeV3Vocc/yzlpeIqZE5mX3Gb3SYHjK/2V6A+0VQUuy14uiCkzAuiDk
ZNW05PP4eJjs/cO2VTjwidqPMp1AbV4fXVpKi/xe2p2ctQBRNMbVo/y5RHBrcKYe8aamteh/IvU1
bdTnz9vNm5TDTrhF3DTxqrU5+Ddyp9MgTA+qAoKYNhAgqWa9GVdfGrAZ8njuJU9ZKEBLmdUIoB3V
QjQkyWLBZsp86BU2ZcP/D0rihnDK8BmzMGizBiZbAR8m3l34bKXkmA+o8GlPkN2SYBpwHS63Hyh7
jDd+zDrF2oXTiSdF/Ip/Hd2NCWbVqFRk+NReg3DVMTtAIhOaoXglBC9pzXXrEOK/5IJvBTwj2vRK
KYZZELCZ6B4y0abfKZ4l68Cg2pywobGPiWCveFGXKahtIhYKp7bjQA5lQ2UJdBGwNiqsX7OnhYKw
7SGq4LcDVbky8/aeDPzstESJcXWpj++HeF0olU5VO9Khlep+DWGMsm64JREWVF2U+1ZdTRVqM1qT
DjnQNVZ0nFZNvbB43gELrw6o+QVgFNf7GSYgpGAb0CmNgXeOuH1zuVPTXQeLIXV8hbIGQ5qbxDoo
8yXNhwpLqKUaP7zXd47IWTtye5ZmyHgGooKsF5oTbWoMS0gsJoGql2Wj2xcYItj1MhrJRNUpoe5R
KQuEah0/YPT70mDdDJ68b0sW2VTZeZ6+YbClqP60Ctvljtl7LseIN81n4117aW+RafhypSpEsXwo
luj8NJyuxj3vOL/x1XtSXdRqqbRzlheUSszYO5vXBlG0xZTaqz0kpwJTbZdDZCFnQsS1zhmtVebz
LPDdWWfQfd1mtEOdlSVrClvbMHiwYq9Cr51z6xWDVs7aQ2GNkRkOuJpTKpgSS3XID5PFG2bFCMDs
MSPmyhHFTA1D79kFsjUBDt7i7rQLrfHCPqn3VptLvgMsaraKTIn/fN2FnrFgtK4y5lNlotA/wpmX
DauIeQAlo1Q4Yh8SypFkahoxb3FEPenQiZ2h8FtyjeK9PeEahfXzoQ2O9u9M2vWJEnL9SDqYXAVL
bz2T+Ios3sd7LQ7aPmOlNYRo0uEtYAEJW97+E7CCshR5SFtWi9CTEuJB2BbIn2fvbWz14Mjes8rg
GO+AFMN23asA0paYEVqP0WSANSmQOSKh/gyBonTlwtrVG4ErOcBkADt+lqatjwI0j+duM6RnuGfG
QBUnjIC8E7raJWg3CoVUqzCWyuFtGmAehfjqNtD5A2Opjl25w/tXRpQMBW2l0+INZK+PqIqG7T4F
o5Zs76vycdub6mlqWu/mqBhkZFh4ZkfjZLQECyBQr8LOGOwsPq1lBWPH1GuohBPJElOmOCBcvufD
LEehhZtRdn1RTWgn2xi+3iI6DDKJrmDtVl+owfFSyHiv9pknYhwdsDvL4Id2EJJB5Gb5J13EJ0q3
PJ6Pn7PodvSr5TRX+n087h7SWR3dOP78Dsf05PXVSZApCuLRPFgB5gHg1jPMVorljAhER7mIab2/
bZ2XAYoseXo/M9RSEjmirQEMxbQccLb54mLnKgzJdCJscysHYiJCIvdPRTebCPmH5kKuOeo4rvox
ogJAc2V22ZQt6oFk4f1hRGUsIYz5PtVCcAKI+GRA7JiMcUXeV9R/wC6BN3kIAnC/FbJW6y9UQMmF
MKKlh0YiL7gG7X9zDquoXNpxl7mG43Lgz7KlfHxblje25+8UBiL6ByL21lcJs2L2OiR3aOpy5nMB
+i5dN9bV4fOdc9SDigABnwp++1rmKz2vMOUn1OHaQ7fpCqulwMMMeNor2LMVV+AmJkqvH+XrGU91
RY8cD3TA5IgZoowYrheq0FBfjd4/4P6hexoL36Fe4Gvbo8jGHGoNp+bknXQtOANR8sOc6CCK4fjI
Oyr67RYkSZaPO+tf4b3djry3kruq2hbZJ95XRpJ6jD9oyln6ttO4MuQM8mxQ9ETdcgJEb/98piIW
1AOfUxpx49Y8fRwoRQ27o+czAK/U+ZMmtqbA9ii6ZJmKv9vsQNGhThEldz1zsZDeVVbmVl0TZFpj
YeP3xsNMytn3iGF6gYx4WPeIdb5CSajkSjliGkFIYvey56Vgdbm+amekmAUAm0y72emlJD9p2i+B
q8DdagezIZKdChqPujYIzKqLETrJlX7ScLOXQ75slKx2Y8BqlcMB7OInL6ebQNIO+ja2nUc8YVy0
DmLpGFW9gmUqrevpS5dVOabgFfrhIHuR+rKAUMdaGwi0UwuNYdMwsJVmj8ykAyywUWH38qmI1l5b
dbVx4dJQ7dyOVzn+GN5M/ofLMY+3UyVUdBdY9Ne2UsGEbWeYiHcnlqjB65JOoFha68zRjS6Higf/
ug1A+WMutbLNPmFkBM0gbOR+kAiVz7jb0B3vgC44as7s1KQYRm2fMpVcqnTzTt4B/MZCCJ7skO+g
YeK5oH3FyddJFV8B/4eYOQAgVJfssZXAp02ieXQf4qUkkrIk2OIAR1+HKG7hEAgJHbkushFgTCRY
08VEXOJjbxo7Y+V5q0du1+w/N5yx1u4mjWdH4Bz03V45CDnai21d0M3ccWTjs0atunbNYFR1bFOu
mEh/waxCmi/prO1xse/7creBCrsJ1kGDuOZfANLporTUJSa80tg/IwYW1oavz1uHFclthGzKXXBD
MnlJLAFfFqjbJpLZgeosUUJKj99zchjB5HfJ6mpvKeB4atlLTGX4NmoNJLpSYPcpsgDvXUE+jy9S
2/bEBEdp1ef/u1WbLwPm3Uw8gr2RxMuS7OHAHhEbB5gj3QN5chXAwwngd4yzeVvzaWCQwBqOu6MC
3q4GlGpXt7C5tsFaQI6DyCSQveY4YLqlm6LalZwcSHJ4w9krj/73AADODffLUknM1s3NKwIbxGQ8
HYeu45PbizAoS9X+iRGDUHaS6wa5Moxjy1JOBCnSIbuOIK3CKfQu7c9x8tWtav4dJpwb+3yAKdJw
rIDILvXlSRBWz8kg7M5Q/PBrYTFSlaXSHHDxHkreyf67XAekV7efVmd1+EBuGDGx3OYROxmsmgrp
vkNV97Bd5QNsasgZxjRgBKo9HTk4VkSLjY2he5lAm0mpVEwH4J5L172KE78WduQZUsOQc3JuZtyZ
wQdqrfKo5HqKJBk+zu+4qt3ZsDmFPa048HzARCC6fWwUm1lSwZ8Q+1eDwfE3JE8Yt58jaCr+iDxH
NLK92JpCMf0H4C3ZdymZENB/4Hc9niRhocqZHyuVub1LE8eJo/zZfAc1PsQmwIv1mr98JuQ1IxBZ
eRSi5AKOqO66Qx2ViLBFgmvQAtbAP9eH/MM01d3WQrscFaHPfiIczSWHmyHWmZyG+2/v1xumL541
zUv/uPaCaGL1A4UaUFLcNNs80VM1W8oJFGGd+rTJcGJ7JLptCknJP1Kqd+s+633dP4Fpij1sTUYl
GvhDlT607cHRfeGZN10kiCmr5EYkLBjyH0v+eYjTigRNTpc8nPF7syrvMI6rjToih1yTaq6TomJL
ifMql1+6/Hbd/msEn+RsHxJDvt/ku+8CtzTBE3AeTCB/zGFQBBvuDQ2OFMWBSqyXjqn9jcvpmBxW
EpY363tpkAa1P8+i7qrCEE42GPwx+P1gQzqXpQfcZhEQEbsfTzXrUQj7I04ygc9smTjZn+G/sMGj
Y1+rksm6XiHzKCW7Oy6RZbGCnotCYC+n9CBuJytCrBEHK1ElfLsHbovgdVKMFiltLYi7q3tIvmaq
8/nTSc9gUPicMAKPxkkXhj0XBGbFrrKo170RbZt31F7RdZ5hZJZj1iEVapwAbR6Yt0lFBO04qhdk
yQy9wqv3xW/1lN+riT7qBXW8Jv/5+EAfOcp66cI1PrHNCn785S4rfCBOUwttwz7YscOzX94o1CXk
YjPVi7RaIruf65TdMuRQlSEAG03fRpA95iwDviM6iF/0NEF1NVxDGCm5NlzFmOQ8rMuz8y0wOSuw
W2lmkQ4bpr7Nmye/fOA+6YgbL1BfysHsfn3sFvMGOno9Sc/Tej7FPPxgqKMPkURoDzUfXwKXg0Bo
4wPTGFutcVk0i+iJNrtiojVxP3Ln6xgx7OEjKDyIzqO7NeOW0m6C02Zoyc42dE1NxAHF8wzVeT1L
ryxE8atdLmjXmSdVQ8GLlnDGmmO86c7dt5VOZIt08ke0kxKPHMCFW1uLxlIaVJLQCOr18ioH/6JV
Kcw6mr+SpRvPc+gFZfIHc7WY6vAaq80DlepKj7mFNQihJNm4eSOvB74ej7NvFkyB7gTlPnr3wgFG
4eUXSHeyS/NYzxMcsJv2rrdUnVHcZfUTFZ7tlYHSaEe8dlj7Aj82RpF6wZJ5heCU3Osd7FkZESoC
7IJyuhcL3iqtXQhi105gN2MUBdwbk4RB2COU35Tlkjserhur85BPRJb45zijTBvgD1xYeD38ProD
SCdyyWSm9Y+QKae79TvUN8zKF3wcCBvtZ2c/2DWqwvntrrG72kc+GGF/+B9TemoV4//gyw9EnexF
yx/1a9tC+vMjGCbezAJETsdLpmnYezvJcLepNrTFg6SIS4zBXNU2z85qd57FRYy/DDn2IhThG1Vk
mnvWCmi2xdON654WNfgUBDkEBPm5ZGtoDr/Av0/4K5st+Qq18N1MhJltwaZW/ZQiPA2IfSy48tzB
uCUroaLVr/q7fhkEHeLao5w2qAzKUloJkwIgTGw2GyVA0jGKU9G1uoT1gqsI4QolPI4nseEhDSsu
Zw6B6og4DgKAWTQtRv9soKPwCCjakwgir2kKgw+FPLr7HKNIPQ2kWo1rgW1SuS7IsE2owl4JtbSc
/RIqZOhWbOjutD6b2f9/7tVEtygyMjrYqD9rGnhAM5pBXhDFXF2WguhbCP4ify/pUDENqCKyIXKI
ZseK3u/NQtlgc1x7vtEOrSU6oj3aEM4ZAPDhQLsNC5ylBgVWsvr8QHSh1C1apqQmCvYpnOoyqavp
O25dUjan7gWUnA6Lv/RdWKJvPnpHlzb7HsfEDszv2OrqbWmMvk44uvWR+WBIcQ4ZXSsXmMknOJVQ
tRzCY7qaqMzro/S3lmd2OjGzjBOHrJb0S19vtWC/jR0Rds8OjIoWmU94CuYM7zwFz0daByojOQQi
kk+xaf/b6pJTiCh1lf2BfyeQD+VQaQ8v8UbzZ9u39d+lKV6OLqP/1sDta2LgvyKl6A0raOTGzgCz
rSKylNDqKQlG99pAUea7yimKxmyYw4xi/nnbo6zx+e2lxHLuLX3R2jhKiWAzClIePIRQ2sm9RRwe
+sMtscLwTckCZTe3PEv0WKbCRukzpyxq0nbuX8rzdJnjOHu+xhwKe/YB1s+m1/NQUsC4zE92I+YJ
UWxHlnP0nssRyslX+mab+k1Q8pZlfnqwhrvDzJa1b4v6noxgSbgUXN/pFqBO5ojMLMH2oVgya+Sk
yk2xdZhnDv1F149McNjoE2fZRA9DcO5QGiYTUsm5aWSb9ZuXtgrqJMVjQfY5aUl2aVSQGSvaHzrC
Ykr+ke0ftkRL/2OkSvtHEv4ULclLyQkXRvsgA+uPHlrXBPdG1X5NgvnJEpNFB0/A6b7JpsZ0f2pZ
5czXed9YSQlw2qUhO9/jJMsqozS68dwwnlHkZTfr3xsnJSFF1aypwIi0jEabURRIbnPqobNtpA3y
gLhYEI+GN5g9bF5NZNUXSDTIqNOLNNdSqkMGYq3lFBM8dMOCEICU95IVGnOoUfOLmubLab8E/1cA
tn7zZfmr1k1QGzOBF43J6eLMyQmtcPKGursu1q7srSEGIPonX7qWXDn83cz2Ue41i8ktTggmHy8j
5jpJnNsGwZ41A7x4Mm910Fkr5AGCdk5ngRnl2cmiWsYM+KvRR/OaglcZX1+ekTStxl7PI3/kc6v+
R3KnV22mANnx9X88FUDdUKnIZi/xMY1dnuZm8Uq1AGvP/wzU1t9SL8hUy4/KzmMk2iZ/1SwPjH8w
MY+dCL57PS6BGrpL82FFnbec7+N7Acq8SNTQXyInu9mtYRJmrB5TT7+u5FLFL8Ocrg2wyT7HpR2i
vbgwOoNbF1odJSXF4aoYjv1d8IAEfECXd0Qbk6BcogIAa308qh5yZA97hs1hv7uX0yrzpgqZVwDN
f7F7ypxhx96IGurOT6mLRM2+iPsPOVxIMb0GfhvODtKMkCVIzVNq6ZixPMKpE6Q9che+S/dqwAT1
AVd1SfnYKKooPrwqP3Xk61ChbeekIfmqJ+fbgrB3YUnagJ3mELsWftlgwGj27M7F99wKwErWEqQR
RJKtqPSoRpLIIEICFz2nI8AevQ6FtFd210N0+mve9GmKByGIDvMJmf6kcASUNm6V1ujnR5tQtH3v
yfJhvOr+/m6HUn9kjm/zQC6vhT0BMTqZ0/zskU5JlDdiqtsxoescQjGGy9v3W4zWWhXPxNDHLyms
JLie0BcSaTzVhTSgSVcGZC8QRg2eNLRxAAVC1+nmuLmK2Y6Y2HL8a2CTR/ogGVyK2Bo7ozkElurj
jvmiNV7j174jRRRG4XoU1WhbOg0WDfJZCp+Bc8aWonDSrFojtdC4oPixI/+2ul3v0kKDtyoApnw3
RS84IezSf85tUA4BuUfEhl2sOPqOILyZBndGw5QHqsS8dsfmDi186DWwt6cNHRLghEg5jKNwSFaz
S4NvMNu5F3r2Bf/xbUde19nzvy+jhFOmh4uSxPU/LNK1EAWw/eJZByJFFcs/gfJoVQhjbuMGfROY
dxDDI5BdgMqB4KoP1rPFqon1dMYGsz07OcnG4uVzMnokqSHLDub8z0e5/pw3wcSn9uehU3ZMdbvj
lrtI3+HEEL10TeudKrWiwruqmZebJ0OVkacf6pGKyenX7SYpVEniWuhblZFrDDmLjqPWQq27dB/F
QqPTJ5JQDQjB9iCu0fnFJ+PKLHWTRgdQghpDZThQmM7iZD4QbBqQh+x9LnYt8uEnV7VLr+l8NRYn
GgGaI4vh2/EOXovhkYau7CFvtToedOzS6VsQXYGfqWLRtIDvyZEXeYWnvE5VLQb/3J86SSRQnifF
hVGp7gDh3295Sxm0Qmn3oWf35W1wNciX0JWnmuaDsgGx7JHHV+Unpl4q1q/Oa8jdpJSbIzZGXUa/
kAmSiBfXOxF9DxbRQyCYR8wyU7mBvPCPZDQfsqorOu8VUDokiWGJIMOHfa7rX7WXGg5d44JMbVx/
vy3GepHhHBeFAvisPZ6ziY1z7gJSnQue1mi5XSXWzak9+/5DUy5Mq0cz4hyyqvZgi9LTJi21wYtI
qgHW2JzWockDELZlndQDC8zxw7CyzIRNpByF3KMgYlbIfQ3u5meafNd3NAu39a9MJOEOGKL1UhIE
qoymkTfZmAeiQVp+fT+dqM/RevlR1AICGA5zY2ioKn39TNmFGpDzfrYtMufb4Dt1ZEfGonofvpQv
aDkJwGCr5VJtUSnP9DUlnGbvDr/y3vdzKrjGAfm7FjdqFdpXkV7/6EaF54933abEG6t4jItbcIun
dvSI0k7HSzQY6LzDuGQMW9sNIiU2O7sYCO3b1KuTnJGspOqst7JNLXUuD9pf7rVT61NBpocU6S58
gGL7Bax+zBJ6V56yAmTG4wekn7LF0dRFxZnwuxjzhuzgy/yTWPdqMI7eyH+OOfZDwp32NZgTFM5s
XWwR33iaggxixnhnnhjlDSGLyKIa6Rj1DK7K+y4caMT9qDILQsjmh1ITGOkQ7y3YcBYPj7uVLKHE
hC8WrDJPceazZasfCYEr4WU/oaQoIs4fpj323DItT2EL4As7gjZZqwXYli3lRzDPLRJzphG2aZb9
xbrGtwqV7lnAXB7tdeFaC6wqkAfmwTdeM3lOd4cjpiusPNdMSqhoIhbx3Oex3AdqkCHMLLiR5qSo
BCu4jabMjhAgrv3a9OWANpFGdkYiF7qHcamLaZHzjnE29Q7Pd2qnnQHfN1VwenguDmMsMsG6o5F7
m+yi2H4w8zQgblZUJGMQLWWK2vD/6gsRob0qyQ1AfaoTMHOyCavBtFK+LNOw+4nBuXwKN78//hp6
VUIMDI69PfZ+AFxreXfB82vNEkbBrhMnXVsOyLj70+o3dwJw86zZLK/VxjGyTxmKSn6J40UE8Acc
4+nHg7U9fXZ1f7PRfGc6t5q2EzLx8WIsaunOW5uOOrnmsF5myl8AWz+X9np3gph6MzI/V3uVPPVG
Se17S4EMsTTJCL+9yxSg7OVxP/PyGt0Jn2CBAsOO+PnCTjovQBi7kILt7HXvLcvROU6ymdyqmTvO
HFzGFhvuchQYoqDLH+T3pEMyT+jBTDKNE2RDfZiOsbPmpfTpK7UiebX7KQsewVEYGqu6ikj0F8fJ
H7xoHoyiNgDraoMjHPr5/AYw2FaNkPh3xAq86l5oem9YRMKUuJrQA0389+C304J7mhtHnjYRIqHf
xyEH9J3WSJTEgcTZP/STQRx6Z6ZLQzvSQVTV+WGGlMdS+3Y80rYZjyFQs35acXy19SKecpPscMhi
xkRGXzKewoDyNGsZ7K/CxcP9Z2zJNq8Nzo634HNjJLvwCaGxFrCKyEu1DxQk443G/M7ZDiBJL4AI
6tN5ZKuH3TRh1KP6A6fRmUjGyLo9jo/ibYAXM4+YkcNsi+nygiQGlFQG6vMytbkHuZtAFV0893rL
A+CHXtloiZFDjT5MWEb0icSKQdCmD6XaGfc8ChXqoV36sKUsmhvgwPdz39DanjabAJP50BpezSYN
YuN3cfYtgOTfiR3jTBw5MZrBHUmBkWbbwfipG3ZZgcOGuvvE26owxYVWQebQMO9aL/lOkGNHfyTD
ZKsf2e7HALU8uDZtmv2+vvO9nEqeaA9hQBxuXpJnUB+dgrJPQo7+GH+c8Ku91RYWO8FI6JSY0ezN
nkQ1pVfoHiVb+Q5kKz2ki3fHvfqW06fL0WfMsU9ZyuhNrulsQkijr2OczjmKvubsfM9Lc35EKt3u
uluQHW6M8atIyVFKSoyi+JHwRdeY49zSeL5pLlHBN3JrqdvuwxfI4oyWl2WUCcsxmfzdVo9s+a5D
JCG5pzTFuF8xxniFR16nh75RoFlSy64Rz++0F92JAPs/kKYFwFQjTWdVJ0UgkMZtgKvrgqJS0epr
n1+TdbHBAJF06ctrgMqQLolODM+RaHo1pZmOIIT3PAd5y5Py3RQS94pIK6WdStgfmK0DxRj7ROHP
nLl24MyGfpAvCNj16x49zXkV5SAppXB1APNKMaN+PRnsL9wdiwzA0SG6+YukjaiZ6ec3rnxLWk8D
8DUBcYVR3xXSFKo4YdHc0eTcjAWi9q0EkdoAFUqwrbqUJqgUA7v22vGdII/6ZWUu/9fnDVABGLNk
Q5WO8JGsQucFQTc3b0OOSmA72T2YMj0evoEifH0GstuNCy6lgjMj5rqmEZheiUVkUSAJIGGulpsM
KfDNk27dsEkT4SfDQBTySiEti8PBSbQ7Lt5i5qvs+wC89gEepUYyL4P7oGEqhcAsvUKpQgAwVHfq
jbdZNMMko36XqZW/GfoygR8C2ObUlrobRqKvJWgRZn1aad0PG1EYoN/9RWx+MUCfc6LpNEZRMPq5
+wjJTsSoyUeI6vVe0T0WQvCfoSsOUzZ6jfQibkL9dfGApLxyW55sURENFYSJVkREXzmrJN0niKg+
tBWDc0fRaJ3u66a81wgNS2v8JbgOMhWUghKzpMs+Mc7ziKw8+rg8q31u7nXUf5I8nnX8gzGvxqdt
G57UY7qfrH9kKZxK83ELMA/Ml7cP6KvZd5Hazl/eQVm5PR62RtoTpLi3VodNbkYWla6Wm7AaBIL5
YXcEMvMeKHCD0euMtpPXl2Lk54mK6VB4aYazqNfAb6f+UqFM8y7Y1R0b0y/xK0IkxPdYf+WZJZIG
Hh/ILsPyAEcbuWZlX9Dy262snyk4U9Uh3wSFbucXDeHxaVhD8ACPRSty0A0VqQMvs/+BlSaJfSgZ
HFNOZyhJLLzBfleCM1s2BNpxowaECBVKeC7vil3jzh+U34kgFY9fBsFQWzGE26YGwRupTmXUAqMF
kRilazwWgAqLu1onZ/ZMHBRYmLg1vtA9qHzCnsUwZttzRfn1SjswnY5DQcI8WleWmjRzMV3H8Ttl
ZwjRVYBZ/WyiAsntoFsvqpjJ9WfuiF2cxlZU6IiAoXnL2NULpuHz0pThtiIdSU4E29oonom4QrRc
in1dFr9nqxYbyVKZg+2Aw6eTi5s0lEpA7RFLKnQxvcrOi27LGCo1u9okYwHTxi97W8CgcOLTwDWA
J6H5Di656ypzMgoRMPfF87f2qKTwJlkOs6758ygriVKUeX+z4Bv0JUEXwpjmjA+NpMnJlHc0131B
5beuWZdyXS0P4Q3I8tRhBYArbKB4KlRnDO7kYUj8lU8sYg6FqIcZ8fSeIZGvvzivY61ERtVdqIps
qZqcFSIRMaDYPATRAhoBT0FyBsBu9DsJWJjxgXxX9xPXI6yska6S8SFwTBGtejndHacfI+So8/sA
jDQPVR1MJ8iuyzXhw8nIMdVU1L/jueTUOO+Z+ZqEK6mBrkl/GnB3csJaqiDnQsyI2yY/1QiZK/Ta
n8m8AgtfP+R16r21M7oXVeP6iHGp90VkwdG01zwv4GWOy8PP+MtmZmhJfqIl4VIWgBnqDwJW8vc9
XF7asxRJZvlBtO2Id4/JFxDP9ohQqtDf5uekarrXlXuz6ivkojA6enHU0enJuCoHW0+FbnOPAE6c
EGsvygPG6KMFfKeUTm9knpXNFU0B/JgvhRMHeT2H9AvEuFCSpniChGXkOSFzuZMYRUCAVzEZBXjv
EDMg33YvSxCrifWqKawvqVka4k8H3pHwhDxgkQBbtjYaSlPCkKq9/q/Db0ociKUKdsbH+ur1Z3i7
gC6CCuNr/Y5tSk1BgmTmtQ8nSGyTBg6oYmPdBKF96QqkDS3PojVSORRkXZSGE9h2j1nBnGJS5iXe
/5krJtxE1BsqDq6MGPT3Fsvokd+xFNiILtRaxSKmkJIoFXWaP5n+/xcDlgWEL2NnakkBuLQM+Abe
0zxfACNDr2tdE9d0uHqoyC3cMIedi5TpNLSV7ocDD/oEay6wzg45/162hDiAJaiimL52UENsxOI3
mOlBu4rUVLauG+hrzFijm+WPvsgru+glkPEgiUCN1m9yF69Mw9lqe1Mdj4BvvhwDc1X6DPBD7NuH
GygOeYPQ6qt1b6Y4/HZIU0FquBMl8XTntlwiLj8k03FRt/0aqAzVjcT37pgBc5MYope2SO+KqVoT
82SPfy/eF5sv/06ARnoJPjB8kca4VoXSQ6J8GYda5gDkvDg5RdMtw7u296tL3cYUXQuxa4ZxTW0r
+AbOUSyF9Eq8FT7lRFBT1sBBtL4F9AWE0CFadlcwDv0IuGPRaq/z3/5rUBIHP9T0XOdZzBgr6JYV
sGV3UJQSRV+yYS1q+endRrFRWhtT9EYdfhmEGOJMLEWf51/imkUXp0XzH1fVGdYMyNxwrsWpoIWl
igsm/RsFXFsHWTlbhE+CK35YwYSZ22Tu8VP4lefnIddfg/dVnohxvKEnNi18ea0Ew9GGSLUhLg76
sngz82Lh4UM6xJ6pikZrGIFw15i9FbO7+EKa2ndNGu1m33U9W2gPImKE7BGv2q4UGyPLg+uFuB97
5rd8O6RKf24u414iqb/oc1XMtCXJu8EWj3nBa4tZ0YdpGmlG9MFrFr4RhOrcrAxpn+Q92E5PGNpC
XB6zxe0iL9vOj71dWsSSYC2gRjghYLq+0Gp2dXLxFNCrdFXTYGDMjjEmkgzaZMJpuGv017J+2ZYk
EIGc8MqImFOIsRkAafIjrqOmDBZwP9Ji7THU3h2IwbiAAD1Y4xQBdZgeZVi3t1oFfQPKy8TBqM1V
K7/SndpzdkZwlONS++jmRh31L6iMwJNrLWZri0cR1u5SsLj1vRKduIrpuMHFLeKWu7DgOscN3kVk
QQ18FBD3hRvilYBJqJSU5fUmTZmaE2pCp+zz+lBlTTK6OAzcJmxGAf/HVz6bk+xgaKlM/mVHzXWT
jfvFoC0QlPgZv2eRbx8n0I+jdkkKDtbbjmVl7bpaleXOTDdZZV8ATZz8nNWgkdIdt5KjW+GTEap2
necodnx9ZQbEI+IU6L0dxaHP8KFLUWI/YFELOymGmh+YQxlCyjpKyopyX+w20IzAdfrQmUGPAcQ4
IXnS/rhFWz110UW/MUjyi2KnPyvQfXIqxECTAPrpx39nF3p5P56iV7OQTyj7Ik3OWyWJoyi/F8f/
VdDShgUbENTw5r6MANYc/iDD/MuVdnK8MLemHn4NdrRx2sj5yBUohNM9HstnVPT2RsGOCffiQudg
jqDp8gjTbuveVBcCTVWuzgIwtiQE9CzphI1MoFamH4yl2GuVW3bHtQtfxS7aALANG/CX8g9iX2OB
lrCf6OGy2Ek1esi2+jZxKbxxrovAfJuTt+k2aPNDWu4hLAtcFVOieP5aQpa/K8RG8OfyDrLMl5/j
cYTsr+ywEdioBbwoC62cdsPfYMyxTfqeprh3wds7Vvqvle9p+ju5VywYahYmiAEk8aEZGrTgrFVz
005tlDZ0cG1jzydsdFIcLm748IybJq6UrdGO+d+ELmb5e3BTdtl7smCk8pn6HT8CIBi/m4sQEyqF
6aPtPHMtLIGxb3kh71sivj6nTfNXsmEkdGBK/SUR5SU9vmk+7YfZkIO+kfMg5r69Y3H0Bc18n35T
3SH7Hcc+fX5wXIPy9jq62WLawb1YQvhHo4VOXsYXgqoQAQPAjEabAZd3FCiz8GyF+/i8LukeNHTi
RgLukdgALLjw6AcU59N2JtR67izxg9esuKJ0CkDm0L35ntF1nwgzHu+PItgrgnDbfJSRtXpF8v2G
kJBuDLAWGjpPVbpfdlT6fedOt5/g4ThNZ4LruIzC5whx6ktVXse6/OW5k8v1wglJKNf+T1MANa8q
aOPvc8fW1u8eynMBPx1rEkEBHNiPGWQhXb5L+fpzp0Z8Lwl25On35l7gNwNBxS/6iA+SxEK58L0R
+Dn8zjHGKLQqo8SwJxHouTYa7rh2bNpWaRj37PZRKu/FCcpuQ1XuaaL1yRH0YRxl37NEhrVJgiD9
vSNdM9u7CbaTA7onAGJxbVtIWUXm/Z43JaZjF9kLnx72VTr5SLOp9A1RIxYylSgz9wP3cvZX+l8d
v3biCFFKIy1Tg166LefGEbV3CmQo9cICbkrL25HQMGWNSI5G5AmwLfTQrRnNedsUY1y4aJuuIWWA
jsdV536cnRqHwMuXP+2+bToNaiZSG0XAOtLrpxzVWA5Mu0ZZov4BDtAaLD9I5BfaWnVrSSQrbakA
th2jLOrbTtwdhCXYNiNRpcaE16ECd8Mj1zh8UULkfx9m1bLwGubcuLQANtS4PvQggdC+/2LFfGsc
JE0aeuZRFWxj3ytMjc9L7BJbWFSonsdxPtPbXAy6WDPG/UPirRmhHHZ9YhWGs1grq3UTY/jPWwpN
lf9BdN7yQsao3hV+chxVEwQ/sZzyn8w7tHll+gaKOz8nsohJevgSgOLkbzxFI+iM05+JFGksN6E9
eZ6YoRgMglUFDYNIHoDOEjtn6j+6/VF7IQxp/ukPHSpVKv6DPbGa2jbvLgHhMhl2gt2WetRl1uqe
GrObttE6FqYBkmj0VG2yuIS30YCZQwHAhG65LS1/BzWQqudEYmhnNXRMi2AGb+3MDDFldEpMMf9F
dnYipS5AtLmebEQjaBh2+3NYzqNvcrpQ6rAehtXKWouOFkaWbb698pMS/RW+g6tfkx0taao44Dx7
9bCYe/fGXNec/Y90iOgLvcfbL+3cxmucUafeOG6HbLO0EKjnvVyRvX7SwwyY2vUT604TaJaRb1u5
V0AcxLc9r6hcgCmqSOkzuj7NwYil1/PwU+pR0LPGq88dvcOk4tTfjTtlGX+qTL6/o8Z+VglWE6oK
jaJTOBUbk+yR0Fuvk3aLBJ77Fi4+eHv5ZlaTsmttfoehXc989KcSMCOGL5/N9AnLe1DX3GjW1FqZ
ZihMqcG7paYm4bZhfRRtGvR8nMKjmmmGVMAB7RxcifEguXE+lW9mRs/kb5ShjdFbnnMPfSiLcpys
J1a8AkQKtQFAPfWHmQNYNwVKX6HzSBCTSPlFfd+NkrJ/Fn6EryainyHVgj8ydwCcVBD0zhgiV6qA
Duz07TIeNhUkvORr3XYnZFi8/dFciMOAtzc/jQgCtHJMEoHR9nRd3E+69wep2cERB8FvzqjA1aCR
eRyuzMn8wRmzqlxKSndN5ihfgUlp8UY3ztMH3JamzEbqSxLStfCa3fmfbNI+P9ukxxr7O3IZ7HSv
XO1R9UVd3UZuyX3VRFvq26BVeNJbk0J40bijHYYzcD2M9SC9Mjt6K+sh0I5N0vu3khDR9fSd0WlB
/ufb0wElGWJLiAp+OtTaSRfYpm30bb/DYFdx310WYjKnUXGVZchuX0pqmm8iqUCeefCljHnR4AGU
id4UDJnHoiNaqq9J7+ccLiLqsPLIpSGGw/Rz31kFGz3UDKLqh4M9/4JJ52p473Ou/CjJ2aChsajX
LAhB3hrlX632dDfhgDec+4Kzz6TKd53XpGfJG6VMnIsq4OmTT0sOlBV93yHp0wJNcIzXgInrU2/L
CWvH7QPH86RVyhvqdOQfo/Nhb4Ns73UGrsuh10qC3zEvha24IbAhYmnYx1Ah54PToGMfTdwB1o7/
ejAvu5gXH+6XFAZ5AGPwc7bwgEVz2Z6L5vvMkBzg92ejLpLp15kBOBBoPmufHeYpVO8E8ITpYCVe
WJKkpgit6AwB3uqeqIuGPaQyZoNjYtGb/n+MR7ILamNCO/ybX6B6VGN7QC+W8yAoMDnDE99T62SU
7VK7qh4XPiDb4LvUB9FJgSgjZEFuiu4Og4+T0K+bmm7tFqMbiTbFgpI+eAQSHQyjKe5k0zOUH3Bc
3dJjrBPBT9NikKmnPwZtfWaPPKE0wIILGLPgeJtjLzZQ+Yq7k5QfnOJVVI5atgWQJOtgtV1d+nk5
ss6BD5X3KsCs+V99//QQIieFXUDNRpUQn7h3qIYoqyWm/zkmscDM6g3mzfJ8XKB0IbwjBbdkbhWz
U/66/sSbbxfz7Q3AfhGCWHP4kTlrvTFMSpVECKgiseWQdACM6bHyB6UWjX4yFiUM3bSCGpbY8PbD
bx9Ilc2BPgzRF3pS+tb4JBhmZjSM6jfg/rIktBxhrsmZiz/EnQ7vfn4cIZYZ3+CXueTPaxgxnBta
TtotP4CyXiU+eg5HqK+56fpK5xGeOzOb6P3wFFm7WOHEBxpMnkh+DxMa6OdhQW2SVB3SVhynLDa+
Rr9GEuNzxx3YY55NUZPk/YQA/Uh9ZK31c9acaJG8DQsTLeNtAoU3pBZrfVisIxWejuGvzCfH6vmp
dpBMN7p59B1VEX9svevpS2Pnueye7ZFNYTGDoZoZVHz6Mwq0PkRQJisi5/4U+tacOkuR2UIVDhmg
59kKszJNnOys8b3zfyv0fTcM/gFhBJ6665F/3c3BaddKbBF1lpDuc2kj0mLbTCCNsiuXmvChlEgE
z5Z/QC7VpUVh3ND7Ww4CYn3CX5Xpyb2QZ4jXh7oC966t+3s0nMso9LYBy/vHoVGvl1dlhFfeuMfU
INgWSArmzUsVTqxD3OUYJzonKQCC06fgq9lkU5cEz7Lf+bjblzTuNr+OESF03hFc4Bpi1Th4Y1Ho
y242chGkfCHeqhomaHbOUXvtQBHikNrFn6mWjqLl/dsSE9VGATzaq4HSX0DW21qGMdoqxk5Ls2z2
0VzMlWQ54vvQwzFzVL3Xtw7TofaJJnOj79bBLhWOrBKw+HHt7xYreNhBo/+4aIi2/yaLt7RkVw97
zsxWKkTYSyxYeAKtarTFaif0ioiZAM9PkBWPxA8+AM2SZujNnyva/hfZvZCXJXPQgk2i8Am12yiN
vAz3iIMa+2MDcsRjMSKYCWc/nZG3GtouKVqXYZ7DHuX+Rc5HEHbIo7Kr68/OMkqkKyFNohU6gyyB
RIoeZiBeA/sflrrs46v4P3UPZe4R5DdgWvwJ6k5iW458cOt05eKgg0WLk8ESWs9Q3ORFjIovdXad
QYIBt0Lm1dwNKS7iptm7kCnTNTHELNc/ucxUbbM/DB/J9SfuwyiOgOtaXMlxQlda27biIz/RfxjK
7NzyYIiB6shoj4DrplY/Jw2JvLZrVvesmlQNYxOWIh9NQnnjhTHQo6fbnNTYqqHn3uJxhF612Ld0
IyV9RBce8LNu4oOhhoMmKTwY47G3LMsVKKsKMcwu0kRVu87qVUfRZPdXXNlfvEjBXcXgZNiaKGJQ
h4IdWbZ//hy5lzweHKjvNezUT/EAFagH5hAlDFyoDMwoV+GWCP9R+DseMHfXu6JMnpFODAcUaG7H
x844ZY2TYjHgiG2ZZV92jaz9K9MEDlMeKoJGuykk+bwx0XYfQYUqjoj5RODmsDP5kiIGBKBvrvhR
Ct1INVhqlSr3PLGsKEqDdy4aOPi8jAM5xSvPrNcAcEXTCNOqaSDTUkHSbS3qyC4ZsbPRQjqp3AIZ
pXX0bFXV9+49Bw/hBnbUoMPksmGnAMRRJPHilH8Mg6cresgWL5u4tuVuEjdqck07hfM5BxPmd+x8
DoONctXJRmAclMhXv6IPcnpNB1IfJSzR5pSLWbSsfGRi6rIOsRZzIMWkk2HXxhBuXrPIcCWbvkjj
g5DifrWWd2NvLukjIe5VMboFmi636hAlYoGHExONzwo7abv5bHF/lP0HQ/pcowhZX4KHvgLvrj4H
9FVz8rF/U4mwbfumq+m0xgBPwE1zI2G+1QXF/a52iERtTdwhpbFgAC+Tdbf5bslAJOEAI8AQnqBU
fsUWNo+exPwQvL5UAwqo5ndCmApUd9a+C73rs7v7bL3f30CGJREjzez1K7iF5e2q/tTCVrYSaN32
OquTJlTi0ymV1Vxiwdsh8A5Kk/6e8P3Cjq/M1WAdh6/5bS3z4OFHsdYi+AFvrlTTUjixoC2inP7F
k+txoZyjWe2k7BP1F6KWca+o0d+kvCADWux0QdDDO6vizeVKd88UDF3OEBNgt1H+6I4MhlWnU9y7
1aETtQ9vtEQkqE2hBYBzMjUvQzgXPYbu/rnVlfui5gmDm4IVpg2CmFJ2Msqk9rsBnM9sz6reetUc
1ebcbT0KNh/tz+sEM1xhAC+jFuokkkgbsKZ7SFv0OxUI90XnA82C3xVM1K6t/1CDSm8wlwobaoNQ
mpeXYXjmMaupTaPPZtz7QsrivYCfT90VSoI6K6QalWB7rnLUV+YMaXzsJdL7Xlh2K6GayT7hcvvQ
YNkkcu0eIBy/JcbAmhGKGKaYtRYhiAFgp4hlRVnk4NeG5/QoLjox9zndHeY37qW+lbTaEXc2sBIM
mJbRkHc7SOnKVJI0GbGNoqdpU0J8lRU1EpxfY1YZw6qShwXpCQrk2fvTwYAQHdo3IY0a1zEatwkC
CfHppo5Hf4Sp6RKw+1r/l6PPO1bPu3bQ6HCuMesoz56xUbeSMhqYbWWcbMi4cLP/Bn9FYbxa6f9U
aD82lBRBrzLGUKbonZNWLdh96/yESIHTtK5UgcV+0HHV7SJ+ZHLV7RAnmFPR7IXG7lnXJTBtb/15
OLrn0KZr79YDS/agye9NmCfhQa+LuT7WMwdAPaRNHMamDQDT9gY7fklvBF8/WiVIKCGCLl/8C7ee
EA0rwrw8aWxo2qGLWzcwWlIFYinZCmKu/gbiEnqJ2v7BAP2KxrfMy7wc/kCqwBLgeKuejCkdwS0H
QTgvJjOmM3axTDJ2UL9MPvJUiaiFc2hiKSfktHMCzabUNBw1J+5KbenKX/WGlgsEqbmqgk5tvWsv
gfgCFTg9sZiZh9OiziK9D/lReApkt0/nBW4heIjXLRnQe012JaiC9ypDrbJaa2adUYAYK/4RlS3T
xts7pZq/adu/zRc5yPyhyWi5NwHblUnE9m+G7phBlO5RGv6r81nM0/W55Q19a5xc3eM0zLGtOvQ/
7d4bsDbRXZ2RU1Ysx3btzDkhcZDa5CEqiwDq/zsJh/BPFoX56mhbPgZhbf9UCbk7CLSatcyribyH
mvVGSJDCIovepDNp/rUqxQpgTu39o0/tbLpjlK5BBBmH1tjWwTNW5Vlqx3IzDDj1EOddS+TZFNxh
oluwgTSdbD1QkAZv+HJbp8TXRnBxfBoXLfTvlzSV0bg7IqI158WO0QVtzImYqqeQ6MSGxGScmzAY
oB/Cqim9DiGniz8oI5MQGfU381gJOYBLLHVcbO/0bSJXoiukgPduEZbbw42hjNz/A6JbtPsIY1S9
VgIBwuVGukjlHR9EQychHxTKLHYU/YwDgbxZQtvRHf3LsZjRu1Zr1QmCkeVh3v/S4V9HEPfXzF42
JbtTCwVYGoEcCEEU8kkP+dETdoqxqeOFQQeO2/psPVmQ5j2Wz3P6v40eza4ctjEpkxv0p8iI2TN+
ea/vnNHzLQeBm1q11JjS73Q9bVFgcGSYUXHYcN0pt9OqwsTHIAUxL14HVHzT3fl6dj9A2CfUZARm
Wjl6iZWlRWcHO6b1dNuZzbITQ9Ie9vblccU24gEcXiNAb5BxJtG/A4zJO5rmiMgN5Md+SnKt7hcd
Yk7n6UlzlgBep+I8RmSucwKder9Key5oyPf11nGuahrOKNAYQk8gSWqce2OUfr0W35qysnhr/Zmx
lBF+rekdsCbuWf29ZMc6G1m+yXIiCPpnCOaTru4oX1Bxdu8Pm3p3wv5Z/oiOa+cWGMmENOGqYRC/
OtQ4vnziI4E41xgRjrj69TuGnVDQ6lQJ0UCbHBbyuPdMhFUQOc32az1S+Pe0G5WQC5CnPM0eLxZp
ZnddL0aRkPfy/9QMVL7mtH/FYjRobfoTu74eVJlMj4N/zEeAgm2qZMHnWDC46by1QHiZ/lDvOeJK
pOQd7vK5F7ds/EJ49HIgakaBBeZ3OlAVFwnlAnbV9jVQwB8py6LO0GI6HfnuBM7Dq8X+7oyF6gUa
Ox+JIeFNIKsfy9nGJehMPwdoTHrRbmPTVAFa++dTEh1mqFR/QLiXQhrPiw1pNHSurHS6c5J57pb8
EjdOWWEIjrK1YtU3TlQnXP31e29qDBhbeLD8DvQLwIUIAQcbFaSliyXWoTtPkcqacm1tJlAAaB/A
crAUx+3bihfB2lf3i4nrS7MAlA24Zjt18YfqoXXzGNMYUAGsCUahTolXg6VI0scT2hiJaNYGxcCd
GShQQD1JY24wc8TCAestv2F/ptrX/yq8UpJl+LlgLdtoeTjC54aIVFj69pL+niWpaLlj/mXiBdy2
3pGIdUk/6/S8xezoeFqL9oMVoVcLLHO2LOqXT8apPMBX2B41D6Isp2vAz/BLvWTJlUnPTinCD1+u
cnE2/26Q5CB1QFNAxeKkIwXtjWcayvvcZ6Sg+oy2BMo6Sm+VHZTg+Cj49CRbVzwmASg5lHoTpBwJ
0LEMCYdTuyf1eylKxwbPogX1e4nr+4wF4JGHFrtPduW/qvmkXUJWAy7sEV/bob8WQR8TA3rEomYo
bpuhTVUyKr8e0X+taHC2wi82g4QQkec2r/n5yX+NP1F1RdSsWD6Aybc2pU570IbvWql9swFcHMBq
Sb8jmdtsaz5qpvtMRlwqNBxRIETY48OLMa0UNa3Xs4OpeWGeUEPAgtSo0WoipsozJAEcRQ9uCyyx
1d3i4UutWbLuH1OY65CEGnpyJbAt0sOCCCoATuJEzQ5oS3btIvD74s/d4lKBSLUA7choPvK0Jrfa
XRceEP7JRT0FyfjJQAyA7ZujiiGYb0FKsajb52Dk9OU87klY1reH0qrPCg9Z9a/TqBGlY3ICKL6o
LpF7m3aRDf4kKHtbbzUTfEn9GLv6XXJ6uRTL/xZRjz46pW2VKegNHNOZ9mpky/Ta78I2Be3In5ZX
oee6kwBO5J9fA/G5SK9E3BotaCHtmteoaShYaIEZKI9oOTqxrKeXidSEgwByd+UEh5cdPfjXDj9T
j5qd4TuGR4iGOos5ix96zQ05sD7/EBYj7YuEccEd0BBupZ7TK9DGbeoa0XvqjiSkY4pJ4HnZ2O9n
Sp7mpyr3uHU82+UKXLSvHJ+kJZgLENs4bwunzbBOIxCGMOjwAt2PVDvWTdx8/prRBfdLp6XgYtd9
+3Cl9Ox4tA3yjDhdMbjpDVJZmaenJLrMb3B3Hs9/NaPmzUpWcbTIE3DbvQ9pT2qeRPBYhWCkY2zX
pFNlLW7cVHCtFZZLxeFQevAdEDb8FJo9I9R2dl5QtEsWFwz+00mi6p0usZocs4dPyoBTqDGNXknx
C50M4b1WqALN3eSSaTtRCPSXJ3uL6WVTbC1vyF3+dUquk9dAfN3SVCTNy8Ybx9Ogib7xgv58/YMB
ExlHtyaWAOi7z7ID+H111UmkGRCdmYzqW9RK9vNxc+xjTfyv4pCQLrxCqJ7JH5QP69braQgXEZfi
ofUpL4liDdeUeSQdEAwf8OD7g1G4k6HNZiaEm7ZpxiOl/V6mkwgzi9QHVZGzm6PY5gwZs1U21oZg
TYrK+xv7sna7u0qE9WRAZAtBV4cVC3yZglsnRdWODt+H/u1ywzuEHeoeNoc9tYATe3d4IPYSerZl
7q6g//egrfswpl8cptWiVd5AimMJFkykHYpkq96YrnfwNk6yzwbZfexWGVeyGX/x6UUXAEDK11WO
7SvWpjgH7ZqMFzy1Dg3u1LH5uKAqHObFAQIg1XiG8zliO6UfQ08LIYBi+9sHHsrJrNZOgd6pV8ly
Z8UHK8Te5fmuMABEXxoDc2CdpY6qnvtSQ5Mcmb1B8Y0MrqMgscTJRXaqoYH0Cg0koJV1+T8Ws2rD
5QSE9W48nfBm7AiDhsJJg5oHi1WpH/02RGCUVw/gSs/t+92IRY/xGcxjEjUKy/olaSUPeF+/H8KD
tFbsR6G/qNeXeGRtYwpokntgUQNg9oJSTGeHBAKQ/+bUOpqKqxbvIM7xC7BCGZ6IBamoJU5SPdBi
VAQZ2fR/b1z6HgqkBwyWfQ93FrrIn1Mwc4uLX6mj3Wkh9TlsZyj1ygegHBUFnVPWYjJbLj1/LLtK
o498sFVqxyc3KCaC3AnUyerZgvhhjWkuru5/+VAxbHUxMyZxdk0RHlKbhJmIqpKifEMmWHZI2cki
n6eIMKzzu3TwSiNBjkCIlZw7Z9oqXM3bTvxOs7/Vj6NYV8zZHZYNauLeVu+PEc7yxNPDxHLhTJpW
e9wYeL2fqf7dkYmfZt4mjT40NlA84No53qvcDWrVHq79BdNEIVcll+1oHiivWrsm7VEuFr3j/FLN
kk0j79UjHDDuRRqipoSNl+NKgEdl4vL7V5Oy/UVw7S25mAoSK/uUjOeUYV7tyf/6K3BpFWqnx4Is
s0fVqlDf7uW/PsHwaR7MFod58jeiLW9+sWlikDRw0PsMmEVhtlP/TVAL54tT6bChXmaWSme9HquJ
z6SjSDfujlz7ecZo8u2+xDgXPr3oBj6RCnHTGdBzFuMlbfu5kVRuhjkvUpGJC8ZUkHbMUhWjk9Sf
2kfGK+o7zqSJQ7duXZuy+UIummilIFE1p069071+QBPt9TrTSBogj056eAjGYehxfU0dlLKd4vva
jsm0a2uXL/3hNO/ggjh6h4ShPiPLjInpDPNEJgh3tR06sYgJo1zYpM+KIdop51IQ6rdBnDWo90lQ
LntrQYsQZT01AIgBgmBJNcDn1B8KTUym5tlJTTJhIzU3crtD/bPWKa/0w4FaSP885RCUt9pVzcPV
MwpIp4ZwtAizbJTUlxuo86NHb0uOSYtzeAVKU/tlEmdu/Gh4lpDhEnyV+T25TQtyCAypFbYIMAmS
pkVpNOcZ9bbHZZRFUdf8cshpWUxmB3ejEMrTIj1nWOqoiP76si0PjMEKb5UIlBiPIEoxTOJq0TJP
ylmjt+Kj2jTSff/NKrNXQqhHeY3lJ+rU/wwo8jcs8GXISyb2APTD8kR9WlxWzbtLeKbPqk1abCdB
jzkgxszEL4oWS6FlntLbZnA5ABlUex1FJJaYnJmhVSsyevUy4q/C379pq3XXc2ZpW7GGM7ljAoky
PBw5wyZXoBpLhLeAPonnt27jG6QkpmaCFIE16AnnnKRI20whuef4Y/A9gIKXz8LIRlb7UKbDY3HW
e/YxcpOiRiD/IlTFrP5vDTAf6PoGNnmt3Wws9Stl42yxlop/+/cXvOb9CQ9nxSGCTahtdxYbOz8j
gR//iWdOmQ1VBv/8TvX8U67lX2YTjyMbDCdyvYMZ4cFaZz6asNuhdUOsLcQKmiQJf0cSObOxW3S+
7c5HPYMRzYirvwgsjYUnwbAqjDquLh9Af6IN3zY7RrokH8vw76dM/gkkXnOH7Bb1YjEVvVtfMNuj
J/CTMB4c9HvaJNw4VxUu/hWMuxTzTexcAVIVgAr5vBOd6i1hitMjq/IkkjrE9fg1JEKUBTBix0Wr
yQ9avdg+aPMoxsABIlEf0duIRBWRjAmUZAjPHCQMJbqDnhnmSB9B+fwN2hDIipbQQb0Q90ITf4Zo
lgrwx/wiWh2ukmhGwBGuukNeUMxrqdMTxYsy5SYOMT09EXjih/kyL2OHBOmPnt69VWbPoVBljTtg
r2qymjwtMEiG0SQdzUO9GA4FzID5vc3swb/5MCIqWEM0ks/SwfyJtiyzBr8Jk+vGspPVygLoncpM
8473rwUiWd0rFmFKZIUEzBLYqweYNno8Jy/08yL+OeCjhmUyI/KXkjuiTSLFncHIhBEJ/W1GINbs
fHukRQzG5OZkMaRddB7fR6XSpz9q0af7UgQ/MO2j7ed5cI2UXoxUSAcqPqR1RkR212i+hXTs0rE0
ra45gswjQ+r21yURrdH1F+09/1t0ZQ7W/GotqdHpS1DGdapdXMzIiqISR0dkskN4L1PJ1JabiP+w
ZHLRb1QviLI1uDXZwbY+ncv9YfcjWabCYlJw4NQGQaJzR3qWqUMfgiJA3T96DAwkZJKGVbDyI9i/
yCN/Yo12zh5WGXxG4keutvj2lzZZ/u7Qc9aOdsGDJPiTUV/UIrWQGWbc4mZuFJuOt8GMebO5YFfq
3zpevVE5vqS3JhdcN/XsMihPQOzNWVzuvE87nQZAFU1BrrkLGVDwHL8ZJ9+OXT87FqPxail/uyhv
7mhq5DW82wCVJd5PhCCsc6mkcQCqc4P8PQvlz71r+NWGcAorinZt7ubuh3LoQDQlJYHZbHf0RG1l
6nZILX1X23fGUWe4TYT+62xPEpaaEMziHMdR5yl6ZeKFxnLx/pIR5WVfwRDyO24OIcExqJ9w8jP1
tuCeOVm9Xj3qzxIAbj/9xQguOjXI2msgk8+ZjwgiPOwuv8a86SKaMzJtzdcFfLo7zH3oAYFcvNwB
xJu7qZ451f3+lsUKOIRkjcGUK288OvR6BaAOaHJkRFsG5fEX0/bptUQV2YhWv9i1CPGxj3Y3IKMH
fMQ5hOKUrYF38y202CmRiGdURBqSboRqTTJurXHT8wnT++xDCVjj50dNrBFQSBUz6Nhx4f8m9/oL
IzC6TB2r/1qBsmS1zr/qJGzl/oMYyhXtQR6//LGQPEkdIeNxiuctmigidtZft7eztonU7I3oid3f
/eSs6TN3SxSzfTQDVjrxciM4pcMoGfd5JIjkQbSgMvbYS68axtG/Dlu72PCtCJdGaPnuItMO29gM
EisnC+XWGrpxZWYa+v0zJHvKxvZilpIu4fUmY+8njDY+SYkMOj0CyoVp5cDC9xR8ux9MSiUJxDYG
FUuOvdIdeg0IQkXJ5eObBxCiVMeg/tJ2f6FsjseUo4iKcU6ZNj0FuqsNT/wTwIlKRAxzPUia+1/4
K65NqTINKUEiQvk9bkL1LxtBwDwyLy3efKqqP+yWFg9+PIIzDfWqS4gFzGsTgnxrU5DkAxchFo8Z
6nz/9vJYr0PaPk+FYrhjkY61EtHY5yT3S8CRiM58etqkoFMFg9vP2Ue3aC+aIdkc19kraq7Zkm8E
6z53NVOZHy02Y7/TmQD+jKxx2rbC00WPDr4rgoUdkwPn8khny91IBZ4xF43FEKBwDuLmwHB319K7
Cwe92eSoq/nnkcUWcw0qEkw4ZWm+OvGt1Mz/dB5g8FlDhaWtfJ+peqSRSFGqaZ3P4XvCipqcAY2V
KtnbZCIcUy2C5Ok2R3UT7ZfSBopVxdMOfh/w69eS/K0kuYLRaAOJyDAs/xrXQsLIZxlAotQvqCBQ
DDQ97zBB5DVFKcKkEz4qIN1Vy0VN6LF1crv/yBmzFbYOQxIJ9TIRpWHm/l+c6Hl0Hfbs2qdKTvrd
bKa35o6IL5uI42GaK8FOt9gEdHQXji6QDMcG6z+iId0WvN4n9aN4NAlLCQ2q4gzfqgfRrcc+M78s
9In77ZTo+e/MoVrUBZEPJjLHN+A/+0B65WB75tewzJgURZZ3J7jvtY0A+n2skv3WihcQVTjDhSSu
H8ko/a5AOv2c2F9J3D0PHpyT7G4jZtPWrH/VVziSVJYs9NFudSZn+iiKLWVI8e2h3L7Wxwe/ZmHa
RfEd1G6jnCuabZNjUUuLTc26Q7XwefVVoqVKvEZbsheoE+VfBY8hj0o4ZxQixF+85xNUqvOcpXKG
I9iVNHLUfyMfZFGp4SB422cgnnzUwpFrjaCM8VEu2dUSeJVlvC93mxi+vBYtRuhfcNFj6zaAS31Y
Q8/kd+3uB8beqlSOyTH4pvzYYetnXQIAJ2gqGgNOKew7Z45fTKUZas2lyXQHH6fkFbjFKC4Yhiv9
lKs3Ouu/q8GvpEv7Z8P8AOqfmyIuafE6VrA7KykBOrIllRvZ29sZtVuK27yEmiHSlRwFwTPaVjaO
TrfHN4iqYj2gRB2V40Os5I17tixutc8Gb4B73oKRzeQtheuUO3FwkZUB/MgP2zmqtqKfIC+V8vrE
jjHyZNNJEmYZ0W95Oxr9qIWqOuUBWMTvEhKItwX2Dwx4T6dBjHAw0eCg2wK63m8GVgn3zb/n4OZ9
8XTpVanEgWJVQeExks4Ax4ZrGMgxN2QV/0rDoLLlxyVaoQXW1+4DKRiJX+r4gX9M7Rgug9i/hsNM
IgQIQcA9/62wAAvtCJU7lF8DUuxl+CkjEU6PuVIkVaHmaYblnpvxMYXkKBF51TN3g068QANGKEr2
e//djIk4dy+fOn2OSo1uOZlElZCMsvA8MVAxsxSFasIRoYhLtOvac4zoJNc2b2mcLZ0g27QYNv9F
7eft+YVWjh8+R2xLE4VrMKk2Z+BESCm3YsyVkLRIStfBwYao3Jj69nH8kCYbQhXR3TXdYbbejr+i
+xwP/iekwgAJDZRCbRaSMeyuG5v4CW3JME5gKnvdne+7eioXFmxY3oy7BAc0W3WkT4821QuAdVZf
/cMifa/a7AQAVUzdB58YF/6e8Ig3oNmnvTeuFYbtk/w1Iq3Htl/g42rFaDVZrefpDTSn+DSU1qSX
e/qxp8X2zmqSZwJvBtHPyIG/HqlkqM9mXJ2W8SbOZGU878wyEPhX5e8zDQYZ70AFS182tzFQPWZA
E6EZwylIqOIwnRh6kJ1ZRgoQ1L6HOggiGE4pf4dE6LeyMtYcdC+TpBQ9nsAlHq2fQgwKJ3wApWqV
jZlh/mSoGo1koxbY5rDM3Nx45MiV9lOHiredUlfyAFEJDkYfn1Vv9ucqcKNBbc6/sgrPS0eegsS8
kqE85VYTi2ZoCONLPhEWpzdYdj5HzFDqcKnfVQvPk/ixMfohkg/77PtAju0psQ5JVjC0Uu4NBZif
tUc1EZoY0/wZuMiHuUh+hrS5RFcFSbzJJs83H5nm8AoCWrHlOB9hLN/SjBAxXr3nMFkWDTjQkc7r
FRKKZZQsQS7/KNYKmEGPNNOvC+srHfKhSOz14XdN655GNDm4NCvmjncgJBH7t4dicYzeKt2Ue2rG
0sqP/2trHDX+i4P3w4Rm5wat9R6kktRXox+Jrtc9/pMn2PefHv0B5IMFOvHxFBkxaRSdM5AQz6s4
WpbJMXj+2Jw4jgwiJdpfH3QojWUZYMXqR7nKcwNHMllUN2cUIY1bYXdVwlqNQO6iGXt/fxR7WWiM
ObGoaFe1rXfimCc0jNJrVuZzn6tGQyFrLGEM4+6dSa/b6V8vl3/7L0gehV/yu1DMiXLYnCQOjfIs
vIhJPy0H+6V6Atn63udhKuuZDLbCKsacsXfyoWD629ZsVJKVhWF70SYkUyhfq9+eE/v1G2BThmA9
MkX8772AOWSaEF6U1sR8bxesh8M15gKrIa9ojZ97qg85J7kWTgKSZXAdrfVmpFYcargFAijNPtIa
RKGNcEwxs5Ct1OQglE6bZwgd6pZFUfp5dG0Z7gamAAfmkmCGrYmebYyhwNK26wN9h1mEr99V0Mrc
vluSLJBLHgVVLXV/7bgjJpOavPRYtoJ70OJO+zYvrtjGThty2dLgXAKlNeNTAhaS53Qb4TepILyA
m1Nh0sHndgns/gViR0c8Jp6sVpa+UyqnPVEC4XyccZkI1jQjfk8J0uYBMgAEoe2/O6uf2sG7Z5va
V7sLspW+sGE3GwNIHUy1pjdRMfLb/nTHqgkpt5kkoqc1Rzk27a+pK2XN+luLZ4B4i0JfoFjOgzY8
Ibx9Fe2M9e5Jcn8kPHQmowJ0J/YxKBi5MWqova0w+o01wSRYGJwbWdZxxLU2SWDbjY1dsVntFEu4
IF7VkhWqTdqHIW0WE6N8U3lLPXNAZllOgqQnieE2xv4yTgmWf7HKcvMG0RxEUTdOpr5lWfIEcYR3
b8TIo0KR/xvoBfl8mh8XeH+qgvjLWacFV5WKafj5/E7GA1lSHqFHmHDSRJeNWehDhXEO7f5eBnD+
kFRxw9cab7YMn9Od1bTfQDF+VxFpSvn0kZs16LHUirWZhVC4d8+WROEQWdLjG71jleIAo0h9KZmK
o6ntoCKrU0BwcrRQ5Hl0grRTXQEhNVHn/IMYDikJPgkyrgIe6AlD2zTdTHZCOJHocPp/Pr73RfPw
7PXj5Sxo45u0P+Jcbk7xc/c5gdR+bCr+LKWiSaUCudPeq8OUsEtLMPb67uZix+D0+vZGZvbhswgv
Sgqz8brOKL3wfrrJL/CMSCUbkdapMb6kRJAXA0glyUiVI1JxdGh+SD3OgfaXgdslOHD1X8IWKcfT
1G20V4YN0RXb7Wj488SDlagrb1KREdaDlb1YsxJKuXc7l84c5x4BFcEm+EICkv3bCeRhqihKxBAX
6DeGWhD+qYylznXO45cSoVJY5H4MQufAB8/ytByC6qUtmuTaDzkMuQFfMAlbzzWpirBi/wge9hmh
Gxu7iNHWW7eYDfvabMPut9pWYXwVG8zlgo9KTb2lfj/MCs3L7iJ2D4tG48iwfvUlXK6n1m0sm7p/
lEj/9aU+0aWHQB4w839xz9d8guZfCdpeEW4L0fpZlEQ4C1S1pXgZtT4hDfEO9mCuCZLyCyJyfEyn
FlyGiYqmWwG25TYdTmxeTAl754hp2RtUh6KlbSUUaAsYJW033y9Aa84oBtw4+vY4oxLrkWuibxb/
5My3ym9sF7r9/JqAEdxPY3Ho418XpdIIMgjhpZdUuDc8qI8bzjwgexERDEjxL+piFKkzp+Q080o0
mmzznWQF7WHBOEMg0DwPZJz+0QL/LQSx1iZTheIHbW/mEEVNniMvoUr9UukXwCwGOdxQ7uLYObDf
tMp7QqyB48oekqpiZkCVdn30WxLxME8yYZVWRjsEaerdk89hiKrQF+pkeam5rss2vmyIZJEhKZEF
K0kE+66EwdV6o30Duxu5Bh7Tk129DEvWGstEMTRknOCT5r3WQLEbsoGIn92XtVUDIkZA+R9uulaJ
dp5YFrXjNpcHpHubEt4ECGjCBSAW5X6yn0/xoez4BsXaD7jBkRGvJ6dbjRH2KnL/5nh9OLe2Ztgp
hsuiqiE17pfjFofh7ybm+xHD6CySf75jtTvqYCkHFPneCYTLa38dU1xMJMGtNU3mImAdCa5dbHkU
H73ePLkuMcKpwERAO+qSu1lAezlm8W9sK0owb7JZ1L7RpIAtIxrWhh44dAuaY5b4tLFQla+zLZey
bdtir9ZsZzfskaLtnCFNUPbFzvLWFJgk7UI91p/jzWizw6M/uaw+vV7tnifY1MVfM/IxjkVUGB5v
tLOkTsMEL8wDBhcLyx+JE3kcjZ+NOOapg3ieBJUIY8LDycFRVEk+Am58lLi5XvNlduwaByhCfwCP
CbQQvNdHe503uMjXt8Wu+W0KxnmeMN73B0RqjpR0b9mE7SJlqGSPlngTy7JtPZVu7K1dhlXp1aeT
TARY7jV8Yfb7cr7UXUmDC1QeobfURDJ4i69Agq8scLYWdvQxKlmdBAv9qjvoIM+nhgrjEBKFKGdy
djhYzHQHDgNhpnYAOcJfwFLDom/pOxwqNICBlb136138sIy4lAOUBi2dZEgze5rMj5n9ia52VLFe
eUlYiJV54zHHfTH5j9oiBpuyFt6dnVtFmY7+ureBh1aBlzxSldCuObV/X0ILpUFqEwTxrSPJvVfH
EfxZd2+M4dfVHX/1PEJj4jPMQ2vqDpGivXZRbi83V+vY3Fgu58oWgNr1qmAPoZI9U+wxBRkmwY1E
DdIFQbU9x3HoYZoqwY13L7Mh5oUKMLgs9u4IVTtfqTlriteQetetEQPYK9wizLyl5iH2z+aE9zRZ
xCLRP7F84hLam59eq2uTch/peZtCaXGy4nA4XsxsxobreYBNfkfPhqtU3wDYzPHoRNu3Ioz8ae2L
BDjdG09jC+6n3BhnsQ1oTk3gIQYLUL5gJqZwmAIJNgPPa5A7Is4XnwnkQdzwEl1YVddnQB/pX++s
dQPrbSqeA1DG/mlSlpJb1WsrQKL3Rta79GMmvNLmLhdgZl9g6IBPa8ZVTHxcbBLRBt9Ps2IY6Qzq
V/NLgA9/iSj0INDLqSVp4uTGvpFa7v+Pxy4/jKaLG3cmJ6ik+nzbj7oCI9ik+ke5/7GWaZppOKWw
vcZGrzZgFu/Tq2Swz/XOFJtObDXfVu6caPN6NCg1Tep5y+liRz9wQ3TMWyzQEUYrt9HDnD7Bvv04
fkvkG1L2VnUJi8/aN9n7sWUFvnmL6ojVrCqaUlgmAitSGm35eC+0Ec57BorW1gORGmWPqjgGFvZ9
brxg4C8uiUPEVSO26TK3fRVnhH3Aow1+y+5G3VqDmh3oQIvmOFLVmIRgKdo7TUBmxih+9f/x8OSY
MEcy1/l0Xo7D4k5M3etpglqOS0a+zm814tIFXF315n/Vr9iZ7/YOdOFb7kxtFLhhMEduuMUD6zv9
jUZSxLj8M5t+jk7h6jeFArgAE8iWMRrT1PzYWZlgL7NyUCyE6uma2/EpBi94zTLnY34vwVtituXq
5pjtEteu0oXm2cXSM0wXixAblXL/JGM3BBfs7yUlRWRp0Es4EHWHYdWXtZZoq+3N8Ld6WSIrau+E
XlaZ/QveiAntI2IBJ1ERPNh3Rf8YBFdqswoSgEyi+qO2mfctgLE6hJoncOmU1eRj8mpYWZVuB9J/
bde/ncBeIUUdX5em7kSfkesR/Fu39darXxFwCs0lpDeL2uP8HcLf14cH895KlLZQvEKoaXMYWEKv
EzoUV3pxLtYkk3AKJxcNpzl5WlMJPA4xihu4x8Uy7h0/lVPZPd72M2EUSRa/X7e5KxT9P9iXEcBV
j5P3hypanwCPlICdXo+sXlk8zv+bdXCUhs1Sext4BdMw388iG8zBhEesBRyX5xQsBTRPQIZHeWZe
Xv9T4yU6Lr2v2V829QuBGgYji6XHL8ooShxLSTMjEXZsQ9Tugg2Cymdv4Uo27Rg6+PKgTmH4a0TC
XeIfznqV4DLP39pl+IYfIkmiGWURmGkFiVp0SmgXU4F3YYsjSnEMFWGXPzkWZA6cUyLWPMz7TU15
B1688v7wtAnPRnHnVABCgX9fcn6wAu+JkKmw6wSKJaXo8ba6jT4KRi4iadrF7RcqPoGR/qRkPDys
rvHrX/ETI3idHuPjyQE0merLd/TOgLxrwP/vVpa8Q2N+yQvcyF28HibP9vz+lm8n6f8ol/Pjtz+e
RNKpon+MqZEg+6t/UHAKLQl7NgsnOiLRFngKdU3Ok5xzRMnd0NOBNp7z7Kie5eAub+Uy2uthBvI8
dM3PLly026oL/+jW//ZV/VAYTRQLVMRF6FlOJIRtmZYBIY7q8PSfNc4aUqQdP3OC+LEPvNulZPxH
G/PcHTfwlZcq2TmGHFWW+C09nt1HP9bNjiR9BpOEjPvFZv1NY1unOan9IxrmtikBfZsDfllNFScz
g1m63JGNgRw+bkfeZviC+coN2pEaIv3w2ng/OlB/npEgM02z8bAHH4MzpBt3QCqYhmt4rMydSK/G
YaM5ZDcy1fr/yLBA7BPSefSxueGr3VOPCO/ObrAeLoKlR4mD1us1OxQLR1yREk3dJQO33Lo6u0aG
m15QIznzf2GjUytk+eXzOYb28E6ZrxXttpxMIM36ALeVv0XlHjg3FXTFjDPT5Z8tKuegl1bWj9YU
IJNddl8URUgOvvcQK62ByGVwEn210rvZkIKtL22LGMhAsY32f8O9RdQqMhgMq2rQLqekiOmgX2oY
Nue+5B/uSM2imcugsy8yhfxHRTHirQo08yobd2G4953vIMqeYyUeKuFxhbPKNOa8Wx1DqmEuNFL3
t7qBwKanq1saRNcrp6NheR/vHu56Dld5n2ilCxk08PZc/pxTx/2BQtBDvdP0xo7R7+6FGEYxJ9l7
stqCDzGbqwDzDRK2B/P5gaAxhmAikFHWJ20Jw9GmiTI3s/Zj02FmlO59Q+CojC1gmBkfDvWdOPAp
cPlZv03nCkb9Osps9c3HeDfB32/OJc+RCQmR3aj3KTpKENMbXSQL0RnICwck0whcfosES8h0pkxK
anBNLVEbkJ7RokQzI8hSyfiq/En/0dQX/OOOAL3qUIbecKhfHVPHJ2CyBoHPuwz/6gPfhHjZ2DHd
JAAKQZ1EY2qYzMECn9nNFW+inQvyNdvaXvLugoU9jXvCBnPQv2+miHo/4ypCMvG+42bzuucJajWq
Rc9vEHlE8m7CbvbllMy31un4yt29Ts8ZU6ffXGqnYC++MEgYFYVN4RJDcVwXjBtGRTanihVQu4dv
whkodlPIuOOJvosz4fF041SxTzqbnUp/C9aIPRJRkvlaxuaEyy220b7XuZ8b9JWTjVHudIN/coug
ASvS+UrvEUMqpImQhJGJe9VyhoeSA8UvqlGa8543t9rEA+0SvzYIQFN5cPnrkMTofmbaL3Ix1y9U
+FfYwzbnWzlNhVa61N87+AzYbR41nFwo9jNdmbDgK3Jr/0jp0faOZGsm6wpeZvpHsOI87wHH882X
CG2GY03NzhQ4wwsTXETJUif2fh+1+akCkn2cP9tFM4r3JuZa3Ex7ABfkpzlmaBBi9XM5myCB69dP
L+fHSwN+RQLW+sKrUwmIdYfU2Y/u/WFOE1d+qcMxWHR7OT4SgKrH9JjOk3gmUgOK/ObX8tQhsAfC
ayfE/GGcUw2G83Alj4fDDm4r60+b4AopCcPLVAJcZjpdrvCImAGvW99HdbCAQ/O6vW0+WM5Ms1cf
hEUcJG5HC2a2s+Q1aBkkZl/0Rw14fwpAHtMML2xH1c0+u/84hkuhmM+tEszxqdBupGQj0NPfyUr3
BYcbyiNBQqAeoKStTgdG1t3QUeV1vUQ8Ocl+Y1stuytRPc5Ws9brdXxTAKt8/r9gbfQ9p6Lr/+yq
O+yFe1E3tujbJodCjU8NSmc4zTyMr2nareHFxvY/j6I+0wIJaGAj8F3iSy7eW2QJSyyHRSyvzi0L
P3Y5e/8EQR0vkz71V0ph+VZG5fc9vm+ALJdnk2+842HzTsJ9Hpdvrf6edXbTJfjRT6Tuc+gRkUWT
Dd6uqdHhQBnFQbIcfRqlOjXqWsFOoze3o+JTuOI9+GtwtdOGFUdX7pXSDM5jVoJEt5OQjezjynmb
dJWpYDWGz3JiMseUGzGoW38KEtqUARHIK39ASj7JwZiYmIWq0iR3ZCjRehcbp4is08xaypNeKvgv
X6yusjQ85H8aEVj2hvUCtzmTSiuVZ/PDhosaWJ13JnQyGkbFo5JA4LfKYcF2XLs5zTBpx774vm2n
S2vvsuYsyzZvXcKkeijCYDIMYXkISEI/NEYbsLzd6/mcAX/xJutniac5gZTiaKqxSXs5Bt2SGdun
5H0JCHqsJ/XQNtf3xLWeSTreh6HGK6cUOMDx8fTwLwSroSv5RUh2pGBVSwzlNugOa4Bg8OrLxSQJ
IbyNlpc4t96e6plbmKJOaA8sRzMZB/O8SMTnj9V8VRWfob0dwr4Ef+B8CrBdzrsKgQDm4TwnTexD
CwkvpER3fWrTCa9KzDM7gANhyBjdYm7ilyhCarBRIRai4NGZUghbyxsCPokU9Qb/gc9z41FXZqmX
tSPfxm8BrVWdHEKKBp6mi0Cx6mh1CzVm5Vm2Do7pzdMOWWl66DaoVQIywMOho8vmQp5S/pHcpkZD
RPzjTW5TUOzHWOUPYfmL0DOcRoONWhPFqiEGTxK+UAtxE6EB4PxmOQpmeESCuJOMnRNRe7bpwuWP
41ILoetieb7q1xrPn5Gv/vqbL0UfOJ0fR+lRvb0p8uF4yED2MbztblfJ95OzEP5vSnb7+ZXEsSEJ
uoWjhQczBDXpLoC65uq/UNfmlcPipVjACUHNN6WLOEZTKsjlP9eMSmQZZtjde908Zg5ERFS1q2QI
dj6MskZuzYtVCGintCfV8EbD2+54VEU8V5uy3+IPzS+m+NbqdVpJscEX41n5yw+sddYZf9xyT1c5
g3cfLodDQQuZFNUQ29n/bKQtk66cYiTspfyU8BkEBL5gvKcNnIw+Tiioz09gKJrj4EJlgRIPABg6
6YBPSRSRIIam4LCxp/Cux3UiPFspEQmXbyVGVqyZMyFX7fhAQbUZpY5BCZzEYvZzuXgKLFS9F/KI
FZty8OATjNOe7zq0gEi71oyxrEKJeduCrCwi8soUNEjAViryaJ3tnAKCebZv7br8mBhLg1/J+DOn
FwiayylnyNS18x7u16ODFC8l/+2ddib+sa1+OONQFKKCu/Yy9VgoIZRTknjYji8qnFJP7rsSZsQh
FarEplpR5JCTo3EihJFUll4aXwu6cOE+xV9YQxtICK3vQK0u0gruM4GTg9XeL0fpG89B7DgrdnMF
JPTvgD3JfBBQfwKGfsRGbKmoLnyX4hrxTmTj2tYCwjQGav10fnfxHY56j8ldxaq8jztkdaZSp820
9Lh5z9Fj2xKkhikMjNPwVsTO8hMMpv6IqIcXpg+7tktwJF/cTxVIs1vHA+zsUa+iZXje1rnz42ag
WctbUac8UiuPQPirDey4SE1HjbX9oR4ax9uc/8yH5w4OOvqKPbYLT0hK+LubrPEegd1APi7cVADf
g0omn7wUZm5Z3GLimw/8WbIdY4qvQwsQNdG9C8gx2cTLiiZ6PkMDdtONCY0cUFEH7JFdlerq4GPv
nTnUqa1v+KhaKj5XndEpL6iE9d58B34NwZskjZu7jOvBryrVU5wx3xmlDCfS4RCe3QWwL6dFrZ8S
cSF1r6p1ZSih+ML5mDxm7k2/pLdQYJUmaFjYtbRU2Vst6XivAEC0LBURcyRWfkYSjUrx57wVsndU
gqiYoaz2M97pga+wuWyK1lM/0A9HgdpQiQNfVyOlJIkfNvQuED1L0u2XFjbTp3U/DYr+f9PqyIkq
Z8BnFvkz4Oatg4MuJQkEn393nzQLSJBFvuvyZzBPSz714pS7nEQgPw259niWLstoC+ddaCYeSxTb
fGxoCgf6qrNLECOWGI8W7SDCjrc8qagje+g5/Pa4HGLirLZTtUQVi93m8QmjN4SBv0fDrf0mgQmd
HKYMhkILy2OdlcAJo6IiObd0hH+tZ4P/lwTFIUnJ+XrDiPbBCnOwNABJtle3JjuakVU5fLsr2uTV
caw21uoiLFhMUbzdYE+pprqRYApmPU12BehCcNBhYu/zrlvJyKuMgwm5vG3GfKV+Xcknrj30D20N
E7rjxfPozAb76xIOQGphoSNRDbRuTz1z18nNnLifvjlk4IFjNbPwobgXnd2JaMHTeAF2hxY8GKF2
rNlwk0hUtjUh7WEiyf80dTq4vwI1ob32HOV/r6wRaSHZ6HKS+dQbxGFRk7wQxmKhCAMXnqMmZ4Hv
49kStPISuBSuG5s8DNoK9SS4RLBrZmiQKEDgBu/vgK75QNrJx49VxJBc/kEsapeM0PjULq2EMux9
Go3fEdl/8mWSk2Ji+wX+4rknP+UX/KnATQGmZPF6SZlfNShTlSkuguha1dVpfDejV055PrJxBIiA
X3xjUvM9pEoX0YTdCW/UOuyIEmFnkQ0EjeO+BnPdKA8WaLG4mog5d8Ta5vcsk+e9RXN9PJgJG6ea
ih54CZ0mRhxGEFKTVqkIrZwyd01VUkmb7pJO1YAzPtBkSeMP6RZFgvcSevfJ919/Fw/CfQTkcLKL
FIo6DFeG8aE4UyHuzyEcyHLJ9g+eBrNnzCmBi1J2VPy8uuDk2YAbEmIX6YmX0YCfl+xTHMvwKyqh
jn09+W0/3Cx7wYsoYm796k7wOd2s6CJSPgcvpbgK926DuTe4XW8IIqpkJTXiCA3vtlqq+cB+CgDd
LwkvDp84fkvIzIijUtInL1Bh84lwFf1XYjl+l3SoPkwGUUzZRu6I+1q786ocTd4NoQYWJ75EGVOP
HQot0Jo+8YsuXHV0t3Di2Fe+18ZLb4/8kQpIpMLc9xprEtiZr3zVSQka/bCm81HXcJOgHBWq6pjS
vFFj4vXc4s9pQZmEPjjMdctoMEHyUnSHQiVqAFW1muyxF7nvkim4vYgjODpg03P5GAUWfmTlFcJL
1ld1Pt8wVytJ8MOaZ5KihcPqHbDEU3jLSUUYRpxzlWmHCoLjDwxVpf7M5w6SBfGDSKTV0a2pbqGe
EWfCu1V/67RAGhMoeNfhbwUsPNm8gATwDeFKCJD1a+5orPy2z+z7t0GntHwsm2Ba7jvKJzHbzKXY
ZHVCab9x17Wh3NKRrHSaL9553O/C7J4zLiciw+/uZKe+R0WAJX+WXwWe5Ef8M4jR3iQMGvN+Seit
yJ5Xab6cuk0xnaI468Q0+CDmNppMoNKFcn1my55l9FwlFBccPB/BeIiafheT24rQQ/oHGbGY3XmS
P//LkvuzaXYOtCmwBVKQa3pQ7F0f0KbKquO3Smvpq62ilGBgd3IfqfgQohdPSZSVCRp97XtZCbxP
oYFANASV/aqbh9iFSCRXiee3v2B/Hw5gNnj3woDnrhfckskX61sMeYDuWOU6uRmbgzt8Is0bnCFU
xjRWtLB6JEeFXEe5EAyyDUjoVT9Dn36RGn6wc3TXSBxWiRZbBoSQ868OA+Et7iGKeEsQw2YPsOtO
cUJS9ss1/+XfkG+mk51c6YyGU2Hp6OREKXJKRE3V/p0cdoidcjTrD0oj0CKj2N23W2kreNgfCSyq
r8heyne7SshEEKDDZWrfDglwCsoUUyOVcoUPeeJHP0HYImCrslhoIrO+1Crr6txThJiajVzHFHnY
UU8AliMJwODksAqnGvlONlVF28VlwQVn+c2sF5A776DyHtcFN53XOQGvZ7Z8h831NjhOzxRUgIGv
29h2vFMC3wusMGoKmIjP7mHhbJNibrGxaU0JfV+PRuDptUleZOnpwnmZhvOuCRGYA4tmGsNY55vp
d7th0sdreSi17Gntr6SmFS5xPSYIoGJuRy+47pFHsP5imVZp/EUCotRa1ErpfC8EnuCdJmTdim3H
R0oIA0WMqy15rTe2s8nWHuwhOLOCK8XrgFGOTrTg52tz8dCQEnwUfdexvO2coMqkZsXOItdasxZ+
vmGE94y3M1wdnXG1zYMg3useaWMRsI5o0qR+5UJjIzaIEwTd07xbLVD+GVzVZrldGhp96m5qb1yk
spRA9kzZG/uNqPXM7PU/gAoqPuB8JLtFnSOrvHhcyhp3f22iktSNzW+9TxH1cURPxxXEn6lX183A
raAfacV32/WujAqy9dbBWrvTHSCeI4/OiCs0mm8fNCqNfNHk/vJjhqJmiRe8sC1l4WAvV1O5g8ut
5+7zeh+QGS3rNB7UTqjVK7rRNOLBNw/6CCoeFNO3H0sEzftGASbRpxkUOkHkQgsA45QXzNgPJ5Y5
r9kGHJSWfkMI9z2UwWPbyMPshdQZpJnH9lji9tV6K4usT0Go8lSCopEFRVyqIstQ7RdXyN8vCsse
BhQg/zpjt2/YPmC7xXdwBsA2YZX+8GYjxUHVTIhpaBqiSd2Dd/n08YPXwJTghasNDznoor2XcVCl
KRL8AgldDsaamx4q2gfc6+wC8Q0Nnale39j6XblWSCL2hgqmHnxYQnHegwaKnYctIvvg1k8rWWUf
JtV14MOv3BRGvtwdQE0ticASYRxSEE73toNlUP5hTQ8sxfgqTbOtEJfpaBRQdG5bjcWsoZRLZb9A
uKkelGhvpK9Eaup+E7uCifZXH0oMmLzrGD5+niRnQb29/YokV7vX9frOCcLDre3jeuAvwTdOBBIs
lZDfBIh6t7OWAniJv/LJuBW33eTuZByuVtp3d/oWF5/6XyUZIxiTyQlrlKaeCA5njkpKSk79VgC2
qzOGO+eZsuQQHNSvUhbH0isv7Fdt1HzzZnuBXNByBkqkhxgTQlJVyhldVIPxGwvkxrS9D5U5Nc8I
EGhcTXHTNkr06NVKzHS/2Lm2AQrg9z+uBbgBhGiNEexkaGLxn+CoDUYMUJJhE72Ilr+kbGxxMODk
jLi88iZJjpAuFNt5POOfEycKVyNHJW8kYBBKVErIVvqm7d7NdAmTdCf+xQCE/WeDJSJ5tMjfRXKj
5ACDuxsDwNaUhACV0aQ6pFMTXxHTRrKF6TAv1lkiRygRctEq7v+8k/4BGZCNcw3dhlPxfsEKaqx8
eFU6YNUmxFbmddeVa20cXbbWTEHx2yEhWJsuqHmboCMKIJPA82fj2PxddJ7c9SXg3FUQl5BLyirt
hr7veX7RHd8T2d1UI15x5ZW6lUs5AwSbGCjQl4wUrwIxWh+8ysGiXvb8YhC5BBbOYiwRrdBWfU2d
YNWx039fPnyKCEi04SHwowPGxd5NxCxkv8F1UGaSr/koLtvO+SlcBlJUePOmbzC8HmG5ox08yC00
HgyADa3TvUWqNOFRbD3Iws+mlzgqx3EbEQE6n6PwA5yi3oDLWaWOtWwvd0JuDyXtS7knr0R1/Dov
B66A18w8zJgFXZW8b/zAR9cV07owgvVhfDg9Zr5VrsvQ54nD4ouZwTscOGyq4K6oYlV1AisLQwKI
cZSFaNKqvfZofXvAmgsSR6gwj+3WxeUCJPaGM3EhmVrDZjIhSmO692x80CDHahQe2Ku/l/dYfQX7
nJtk2XiNZZOKP4mgcEQipIwiY4gjTRji8OyOXLnQ4iJajM0I7Sa/gT6ddD96MwTftwozFL+JqkYa
5Esm2iLoXokJNuXZPTNWYCfzDMoz/wzu8PitbqxU7DOYoZhjtbslnGMk0qxA5VJJCdMBAFu1BuqB
ZMU8UXYjH4h8d9guComr2TRxoUjA3Vykdv3Y4z5+XyNqgd+ElYSi8K+/esd8F97wK2qrAFzJitgu
7NG429A+4ql5YeodMFs8w1fLjopW9ZEEXbTix/epO3PGI2Qb+fzbz3gMcOI7a47VYnJvS+AOy5yU
6lzzVJNosHGtNz/w5GZOgtNOiVQEXjVm1Ox+VYmqLMG7Iw0uvWWjZTTDWfDRNLWYYk4KB+W1M04/
fPCrCLxGvj/s/j1WR/q1ASYfsAzGVK+GPCDi2pvXG74z+TjtHiTrW/67nwVhlQjt0knaO2qjSc7P
ke7BHb31rBcqLldNJmI+8FwfJ3QSIPtLQp4sI9RVCh7FTfQFSm2w1mtJGoVtWVRWTjds22YCM4ye
yps6dE1yDpFSk0UCg1BzHTBOBHdR3nhStwB6CLPgdQo1VL21mHfNlD1lB5vrTKu0f9YZS083dyaC
owm7hyvH0xb4rCALHOVRZ1hqADQHncOFNf9Lyr1RMt0DfvWscjywvFnySixg1Qr+xZwlDI8YnE+M
mbXfi1uBnCWzaKTZ5JQNj4YsgBrBU7PKU/VQFFWWDl/E125bUfiFb1nQHjtmGH6qI8QfloEi+DCB
NhEnPOEIL+SXF2iJvLsQXmE+TjrCqjmX3mALEKtb+d/8LebL7ahru+slCxSw7Su9A8e4tgCvmh6r
zLPVFJpzdxsZHGruVblYI1r6isYtMnKgTjPPUL1qt7BTniQGPWgl1XZK4v7DcapWgXYX5LHdMQSX
wAK9nVT9RZNnU91xa+TuyHU5wal3O5xk+BDOCF/iwHSAqUFIhaQ4tqVPG68G9xjFinJ/ZPC3lQHP
SQFCbEHHLy6k3/BX0sU5lPNrDmhIyMqjrvfftrXFwpsxhvfBcrY7KhQ7a6OYMkYDGMZoON6gr+Wj
73E7svPhT+P7x6vryIPgNCst5kfHLbdtZUMX52kNqzxey1MtSVPEuznDfHDvyxB87fMnPZi1aiYN
LVgpDC0oyN43wz0Bcj2ZvGOoI+WW/7yACwT9XUYY441x5xgFBR1HV0spo6KYQL4axvhOFNZwzhUJ
E5SYbKjpBxHFpti+IUix4guGLk/f2/Vmk7OncwO3McV9Jb+YRUH+8TkjxD46nB8L+NttD2MDHoTo
tFN6aJYCVT5hY5P8bqs1pGOkH3MbXNpDEo0KLMNedz1LDvtCb3w+nqfi3/ploqdELnuA8q+dxd2S
iq9R3z6TI3FFOsA6/6KiOLY3Ak4+vqU1G3T2LO/b3JBbSvLnot0tYXZaDWNrwziGQyZSy/sHlGGf
irVWRMme+DCaVWMDl38rmsjHRVWBypPH9/QpakuWUfd2KHJOpD17HA6OT+Z8m+9zClnJ6G6Alg6+
d20/a4KBhsjLJO60yYYkL1R89qNewMtvm2NSn5qiIBJ2AFruI7t1UCWq2wzroFXeGl8kLwWtk+oQ
W8HGzUrunhvyJfCjCZVvyhMzODxpWAtUlfo1jv44Kii4I7qmWE2uY4WmVcmcct9dqxuNs1PWCcmd
ATVBKV9rxDK0zLL4f9OeEnZLl1PkpfpOiJvZuDyWBnysyGl7zm8m5QjGIyWZFo+sfFXWtuKY4Ux3
4BWnPqAT0Q57w4QuScyu34avrVHl/vujdoHZjh0FjRxvvYwyorxZi/zNeeCz6B7lFE1INmMpBaqD
AK50BpiO8mR6e3eb9JbgX+iS3GJMRgvK3B/JXVX/I7PQKYVxsbvLbBV2GXlCsocMYKJiWY91WAZ4
kEoQQSKqvqmkeXS0MtQFchZ/ljU814B6rsgzP+JXjriEhP318/CW9Wjjbhc1emerhTZQL45qjdwz
t4Ct/MxPwJB82Fll0eHYjkJBZ5Xfgk0hkFg2ygSnbcI+0QuAmAHUS/vW9rGmlLMiGOiYzo+svl2B
KMLCuYV9LHW7k2y3rqe7KEogh0W6dzJbJ6qH03d30197lfLdOtpOCAEyUmIz3GdFXz32e/yisi7f
J43//ibA1wqnYDE3VPFxysOiqZgrBm6qXEUP+E73SSrS6Du+RtWvsJoD1riPgMTEl45oPAiE+bnj
Rvpb2mNJiKAAOMw53SXmIuLWWImSUAxpmKcUNX3ugD2Nnd3vwRIL888gBMaNdlCKfjykwv7Ad0Vq
oqhRf1JhP6/k8L0MqlJOxvkWX4wP/7B68gVFBdP1QpH7m4+9vwpphoGI5xfs2O/kAvQ9w2HgLUx2
nUVqa3ixRXpsXr20w3HLcscPz/eWQ09LNG+hmZ24bJ7zI8aIcyDqB5JFUsj4qsvwf9aVnTH246Oc
b7QhkIYrGq9jcONDG9/yVY9Tt4q9VqU2sMsdBr1//oUH3GAnAx3ScUZz2OQ9Mf1rctTIbhRx7ujW
PydLINW/z2TVLgj8QGFwQdtj1VeLx2RuV/DKW3znZ5cCOciWUSMKz0BsoZ/BJw1FA4xUXjq531oR
XslFpn8TVzkfWIy2yPZZmpI1hZ2S+yM0VTuzLXAIgMzSDXmbj717qXD6BcVpe8kFbZ434Lf1Kl7k
IYJx1Q/rfl9ZNYtNoy6RQQFTlo6/frdHRIJq8g3xSwaOxYuZMENTRFXJd0XUCtIVxIcCGSfWLhAQ
Xyfzfd9DRljCJXi3ukI13NonfmxFkFMrHepcDaz7JYjaeCZcE8dl3fhRL6SXnqbV4MfoqErYRwtS
nqx0IHueHkhz0szUr3wFJSSY9cSkbNgYq90Z/9+iO2/YwVOTiseE1woa8+Ucl73QBuHGVOmVnV1X
tEd4dt3Ute2HcBhvO15bvvSw92AIi1k6CZL6SpB+EAGD+aaRIYZ4LESBrYHBHwDoFbDKt84AXTT0
RdCC8kqe+wVgs/P7F5dFgs82ztH+hTV8HsX52o4JEiJgIg9X4gfxoy9vY8sJEA7u0kP3a0MoEIy6
LlUUj/85cyO0zaDbmQUoLPUyQrwJB8BWeWZq7M9xIjo+3Uf1XnTuZV0x3vo3j3GhnfUzxRxKVajP
rZyRvj9L4fakZt4aJx7Jf/O5IYNGq+nFCqKvy2vWORkhJ58DyqhQkyCqv60IrhfGMmZMVgpJ31pO
FFQ1LYqm7Ic2PRh0DTB6d7EhtVlGO+Pt2fj90dvdRIDBLqjpXLsU40WsES+phS13/wA8EMZkNJqi
THDjwVHGs02AzoAVZx+kUQVk1EOAzTKnl04l+HmmngAeOlvHHvU4UDfmAyQdcXYdN6jRc3sinm4O
NjJELSFhDQrNtmNYNYldJ86Bv5ATEAIpI7tRwzHg+RAHXuIJ80KPmMFUd9fVYN8U+HY2GUhOqma0
PNuu1g1QSFIbcW4B1zRPiO1RKM3csb5EwXg62MzLgQVufn1WGOFtPF9bM5S3zwDTnNMWRtHJ71z7
cNPj9W4uLW5nYPR8qx9cQNsDEDESamPr39RYRTXyWF2w2JJvYu9hnb/afFPkFBCagbxg2xy/SYWO
Dg0vtbPdlLxN5KJWL9A76TWTu9s25Zp7HVhdWb39bEmgZf3oHM7B32PPaj1SWEnLam+kZMKQpBIP
U7GXFrnypZBE9jjoQhiTO5ZGqp0K4SGWh4QJ2TUwMd0juh4/nakiJxS0MwWXTZ9aQMdP9opo5ZhN
dg380XbJyFF87oLMxr4StmF3VKloEP1QzU+KAKeMLLCwsJtNdQPy0+erbc3+MRuDwZBWqmADELkz
7azddrDXZQ1Lda8IIN359iCa8K60Bm6s98zTKSn4XW9e15xgsFvLUuTT/EDd54zdPdeO97WtIv6w
EzP61vZvFaUNyF3PlRSF5/5/4g9le5xOSiw6mYJL9q47tgmbnQKhRoCm5Qd6H7hFHFDZ/zxkTTOF
XQM9q9Q/PLThrHq+/Zm7v3uVT64OmKqG7wl1NyJl287Kbff/HuZooYOqOfhyYhf/VaOO52Q5qeA5
zrgv3BL3eM/Wl9/Dl58/QA2p1VdKeijrYL/oWtx5QpN++4+YQxEDjhuPfuoECNPYazElFv0ju4fD
998knZwhIHEYbkJFNJ5rgA80t1j7a9PGd1kOYiJGaZ16BE62SyPnT2egaSZxczU/tOeLDWU9gmDe
knJ3oy08uy7Ku75wehHgQn0j9pV6Fe5K0NR5FZEwOvFy6QbbURKbTX1CimijGh9pHXNlLZUHgITe
eqYgC8jQvxHsdA6mDsSXeio8oo0sUTa5SXNH4dZZ8jI6I9uNU5oAQul5v0vvWpRrhPzdYAWoCyR9
3tZ443Fat0XFGncEvSfAZE+boDrgb2ziDK57NMGgsIm1locbnGTF8PyHVAgLHoX0c2MuoaIDmEy/
Z8mI9AG+FCpt/zclC5hr/UyFgCcNG23C7kTZH5FgihHikyrxMefL/YGMQUFDLwMmgxOO60PdUOzO
PY6lspvA4sUMUyRVL3frQ2fXWqe7gMaZ2zWhdqW2zbw5/ZHDACrIWWGrHSuZtNnseJJRHpSZgoZ+
FzMZnPYciLzjhNlrnrMlqhqPFd6TaNM2cLJgjOn8wygbNQhuxieTyic2DwINmjEK5LTjYGT6ggO8
dNHpsgMbaEWz0VIP8imMihfyhxGKOQWI29bHi2A3d9rx0wJfWrWwgzBYfTdbZ46sqfNhRa9w5BAZ
cf+M45LvY5F0gRx/0uL8tPHxOcttXSKmMOWM5CD9xaisVo3BETt6yBzcjBr/PfulmBymCUj2hetM
ognDBhnb2/twOBX8SsOZbQm0D1ontAYrfHfbEQmUSv4qeUbALP0vqjYB49hiKLM/ok8+Mj/xab5m
PLRGF9n7p14QfA9dxGs3p9zt2AScghGivb4xHKVpQ8AsFNG5HK0EzCONaFqfgFRFN06ejJa3LoEM
p0R/MD0B6AETnlRoztKtEBrQxlftl2l+09juRsJZPOsAnySXU2WNlVJB+qJh6DZyO4bSVMRQ00C0
4eOHo6y9aY3c/LqPnh3gh+fhzc/pm7t6L83sS6TMTua3oB1W3mKM59qxo7KeGPjCZxE8NoDwdCOH
MSPHfqTHGP5D0FR7zBBak0QHIRcQNvRusiz782T54gDzgCYFydXkxaMVHcjhY/eT22LUK+z3F2Ap
DPtR96ISebrfKm/4H0HRSs6xw2NtcLAaNn11sWy+YE2+maLM5VYmtp6qPzekahaA+RqTzOVOogPi
sffGry+b+hnurDbUC3wYs34dwFbzyhAHaalVkYj0pJ3/vHB8foMIjCXvHRAKEXQnemjCMxJdPsPa
qHuWZ+q44MYNca17enNE+97zdzoR7nw/RBDKjfqTeZIlGApy4w1wwae+zvjYOdzQys+UU1C06/Ek
WRpyyzhMnP3VSYcTAiCqX5cuqExqayT1aFrmd1RTifYHsvTKHoADCvAmyvJ6DL4j0psMWudksGje
ocrwiDuFmC7OIO3NFU2XU+cv8mWV9RuoQH9OiP7n/0Pu4Nfo5mXModTUEqCYGwfJMKl65RyuYShK
93kD2qysmyp5H4GTXiHcLZkAP8ImgAAEEit4I7jXQSqG9rXGTgcpGcirUH7eZO9yD5AUL42X+bIa
bQinGU2hzjHTQd+ZVsyaMkjzTpE5kc/9JLlBhIAVoAyzTTX2hcJvJSvG7INtcUwr42kQ4SfLeX3u
Hhfvbvz38o3hNjGwiSr3ICEOYZpQ9kjKm8wSoScyyS+MNIGQ2LKGL+txoG5XTMMk0q2iYBSDI0cv
907bsVDPviaNjBfFYX40LHRaXNIg1DH23JOTs3n8cEAR6pVvbd2S1omLVq4bTKGw7wklShzoBbyZ
4MBJ3Gl0OxuRCl0L5Ev2Zgwb5uM3qhyRJJTxi5pH2No7Wf3PgHGV1clZYWWhLAzuXJpyY3ZD5QM5
QiOsNhSYBYko8Vuwnu8l0veSSbBIMCh2RTjxsk0hcz60z7C+iysnW9Og3yjyOqjwASNYx1nrjwW/
r9T0G+/d40ZrclD0EbqJeKyMbOPoHDrS3P0ZGMFLJFK2hIa6VvSin/RyB65cxZ3ECebmkS1IS12o
POKyYV5uZQw8G5ll4yu2JQQ30WojKdhrmkN5EfGBV8vr2cSV1hxmK2g6dqNC+K7+gEuJXCkc7SNF
0xUvBTw627JwLlaA3bpM8EFwIzEdPA7uEEcoO1jsEFXqh34tc0f2FmVRLYY1XFrmTHt/bDpshACO
nP39NOV9m46N9Llv+QhRBE22ZuPyrbcssen6JptFNWIgGoKHTc/OOwCfLCQb6Ba4FHmf7L5dgYfX
6nIYmbyei+aNaEiGlMfHqQrxHV08RUW35UHRWHFujed3+hXwH+8vYBbgE/GkB/rDiSLCq5mivG+/
oNkVh8yc+m4wXDZEVv+DPLPM0u40ZyJFUTyc2GhF0Xc5x/JTEFt2ObPRNggUwnHqeu0LnqLttmhV
vYoJkRp1W07HlxzFW0OZkMQrS2XG36jCTNa47AGNhQdl+4WfUYEokIHwbxJu3z+nsRQS/bGFEZ8k
fSckOYc+nyWbW+jSXC1QIFhaRU5Jf3OjN/LbaJPQKVapOBoqZ35CR9CY9ORZQniw4y712y3rNOLf
AtHTwug0sWLibS9Y/f7+zxDBlhRT99mt+zDFjaYbK0np6jA0+6Dah2ttbMMvx5/UI4DRWnOf2JDj
fxB4u8zvdtp1LtglvBjCXhZV/UJ4cW+N5pU2OeqO6cK40LpJAzkednigNn/188BzBnTlzY17Tcjf
jyPAiIBR/p9LRrp/iizithSiizofo7PjfvAixkj+6flldp7+sXvAdXL5cet9BV5G1bW1OqJWpdej
zPiBWamStQL5Ap0eeOdTyRCKZcqivlq4Uw9TI/oIsKXNzzv5NdArTP552C1iRzVmc9avR40r2+Ck
D1GHI3EVqs42sfFV8pbf2OdhTsTMzzyzKTa1uspctG/dKR3n6rnJNWb9xTBSlK/Iw1bYdjQHMJJD
6uQNONXTKwuGAUvQbO8uLKW5JQCpC/AL4x7fKTpqP74FEgAtWOlRr+N6GVdIskeSw9KzdDIp6nCn
ESFRF4soxhry4b4vD4jS+s5YznYE54DRxNl4lEaKiQJARD/dPyTHGCqMdjSiZrxLqy+1gyJxX6nj
SW7TyS171s9cNpvVx7/7rR5mZzIq3dY7VqGir07RE2iZNLCJqAW8nhqTGSvfsjS1xt7RlGMTo5EG
KzWo30u3pcCVBNGgvVe086uSbkp7RCOkZi/H6vJHmYK0RrIAmOG8TR4YDlZEOTNaeG3tSxZ8VvuA
GOM0u51O5+Atl15fU4YqmviXLJxPhHuanKzf1kboaRXELZtRfBM0A3LJsoyNyMlpYl4pB10GCSUB
/PbsI74fmsRkMcsoJOnsAtdGxYYMX+j8KYXhkn7SR6pi+XwCkJtJRgkaWDYMTK5yJDzQOxSoCX8Q
7cLzBOckJJqAUItsrmGZ5SkxA3vFFS8icw8CLzvynLMOoeF8fJXl/mgu3CgGqHT7RmjSVjDgONc0
fsTGckfFJKar9U47TKd6GWQLM1/OoKJOOchrqBVBTM3uJPwiDemumZfdRfnoDBLXygOCHR+RaOfD
OtlhghfPmh/N6jy5D2k6pn1sVXTF1OpNA5cY2svTIXo9E99EzXeVbDpJypt+rvAyj8eHf3T0pK2P
uhTFLG7Qs3OR770ZAs5Frh793YS3SZbitKoMhvfSPIM62afPJS4PpjmJSsdHNcBRiyv2gu62WXK5
Ytnkv+DeetfRDUJzJiEktwqpPu+6AXoKEWRSvJzRo19Sc94wNwxU11QyFmGO9/Qb/N+1AlU6ujOX
9cRRBwXEC2JdJnADnk2rIayQUAlHiB+o6KdJQeWZ22g7n9MmEltjjqwZmZl/bAN8uCjwioLwNr3Q
JluuG1bp8NMscxS7luiLAcKeSKPNOhqF5um+8DWqF7Y4Nj5lQDUfLijfF3RhRa2ngxujZZIIpcoQ
E+f7XBkgbHJCwoOMOLMjjukF+HDDmzLZLVY7tyGwXibs8qU/wi210kf+z1aSW7uCUnVZbQyisQgb
rLPpbgbZKi8Z6AEmPwGE9W6WvK18mcY/1k8K/g/ICSGxZTjYdtDdi7ydNIO+1TjfEH+6mw71ad7a
6xj9ZYmiPUJnfGzc/BUCDZ56JWmP+O4RO2MhkXAi/OkmcXwG/oB6kA/IrFIsxqq5Wd+eNYrvZGfb
JtbPhsQjgjDWy7yN/pfuUBIjr3af3DU5xNWLnWKeqI+sjBJt60kYtoq5agyXAyORnD+oGevjYXUI
0kLo20evNIO+V9xNn7bDQ1hGPcMl/wC6kax8YAZj/hE20r4YADQePwXvBl+gtdwjj807fDQBUOFt
xYyBejKjF263tu1I+01HomXH9ger2LIYTb5KtvDrhBybZV1pq0dqQYke2giIN8e2svo9KUnvtaw9
lD8SxsMagX1ogAXYN0cUXv5+sozEH5QdF8zQhTwFadGQMcXnbAT5LaAGrOZXJjVOQs/eOhmaiHfN
AmB8H6jD3zsLLhW49Fr/te4yaThbxmDiPhkyv5Xtr9rNBXti9LonrlGkODE+MxOjqXWe8T1/nQ9w
ykLJ1UyqMAuUCN3f3PvCbCr8pfqW71vB/mBpgazUNGiscYix2pkARIdjBIBRW6L3cXxQyvzK++e4
0CLpqqwl08qDv0eH4ugrBe7dh7utm1YRGmpdatY/ySfnCnd0+8R6JFAuEwZhM/QCSIjSDfeELsvb
krnwtgWL0yHeXT/9bW3eVBE8Pc0qO6YGpRI8bTZLPATNFQy4Oj7yQwvmf551nK7UkmZlqsnd4Thc
G0grGdr5A8SNrV/gPD0Mnvg9Egdo4jzIXSUAnZc3FptCN7Nqtr4Ni72GHfb9+/7pG4ThDt5SI272
1fqUPPDMNQkI7NPFcUScHo7VWaGmcx0mCUGtc8rMRXyfPyy28NRyVVP1lcwgMUfidQHFOMC4/wAX
1v0L3xt7OXhv1dM+HUFS8IJ+hc2HqFDmorufKb1d7F5D2R7TtAVczIeHXbtifKac0+Y6aeEJpQtA
DoHOQ+ZvKIGa0J3ZFsXVBWQl+Doa/mnuQ+B4AV0A5f5fy/TtExFZLMFu6SzPggMJKJ0EWYImFpA5
8IUtpYa93UrPqrlXwXRDCjtZoyUvnDZhZNUzXQ7oVa+2N3PwfZVQW6OGOL7W7N08fZe58sJqv2UQ
8tAZJJmbg5En3gmtEsvqRnOJJ7Rs7ndDvBJ8wUCvJRR0e1UE2lwlMI7wLhSvS2iQEVb4YoA2lHUA
vr9fExkPt9tBQAs5c31WiNwltUdEQbDFw3B9uCtR8mef3OhSJtYRrj0+E6JZkNBi+U1xmZHsEkHN
4xzgCb5CIRu66Afme6A8lPUC3Tc/d8Eej9UX81Mc3oRXmtBaZykkLwDfFNsOenuYG14MulTNdTTr
EHwsk6bzAz/AU4nnBr4uNEVkVdQ+4pXlqnbz8hKWmIb4RokhWPCV621Ai7DMp4Kj02BGs/WyHfAJ
SKMFtvD15RS4cprwSYs82oMrLtI8G79zRO9fRcLAeDzYaPbkE3DqbLCs22goze1MuOKmCCsFdDWZ
OSX8qwH8+D60kHNogbbRD6p7kCwu/lCRbxce3jD9qRM9piOoXCJ5CjdyrDG0EUZ7BqjYSoYk7bB/
jYrjWGbAim5TJlmqLV1aLZkP5v/4hC4+q0HxDV/0HaGqj62LAh742azX+q8yO3C+3cNfyMOaBD7d
jPeD0iC5HwVM+kvqX9e52Vj6vhbsrQXT7VvHs/U0r+ZkcsmOYHBInEowNDwdovK7k0q4FkU6xGVK
RPcdZ0KIsA4k1t/g5DYFiGVNmnFj6lPJpSQS8iIp6pUkxSdp3vyPmF45oFmefHgMHYCNpJ213w3B
viwIut96PFlDRYSvFxj7/druy8XT6LI+NHFrUT9Qd+Z9B0Z38/2gGU50mcSKri/RlOacNHM0hFt4
pu7g1gttfne412JW/lEPjyERWOLiNprv1gnnOKAhDb40l8nB+yuDcsA+buR+0geybGQxDSyTQfes
tWpqXuYBlYnpGSuddDXcpP9ZPoAt3V/0mvmEkAJuI8yUcav/sSB4pMMYlFbeNSw+Q7X702/0zS9Z
6Zpe6lJLXElA7IGwpEYFCvBhwpQDPXCbBqy6DNcP8Cpmsx02EuTJJwohp/prK2xStfa1/0BLp0KQ
nvM/6oGW93y9SGmQiUqYgM4g5e4JsKfhI+l9KaN4jhfVbntNoNWHKD94U4cD4OL3w6uqaevUNn6Y
er9BlfeK1foNh+D4iWTKDHncomGSC0htW3rf6u3EB4HqEnPhi+bptRgCq97Nq/7rNG9evsKa6uOU
Z4WuD0K15E7mFHi7AdEA1jnZ051kVBjeHVU0kuYFXWQGAsOqY6mN9Ea+h7wclvduu32Wh8qaKSf1
0H4xt1KnvTAjZcOKb5zpTdZZEZq0BT+vyZe34v3r+821TkWYp/UU03s498Zc4LDsVvvY0SlxwGhG
KCaXEeI5kx/AlCurvsi4TU65NNl4PJ4+U0wyCyxGySeNS5Ng1FGBScttAmNaUxa3h3m28vdcEQbc
/6/585/zCix48yl45R+xlODsYaXGiE7KaeWTU2sOoyqlCvXMbGrUPx0m/p0mekSQVS8PaNkBB27e
mTOResK/AQU9pX9MduGD/7r/Nc+s976j/a1ZGqqUSNEWe/J/N2UQ+UYTD0NSeeTmZijyjoSow89k
Yql6sgIGaHRxadCPuKlzBhivVC7Lr4s2/uTYCHR5B9SzvQrrySdZmJP3tjrnBQlG6LslnF4OiAlu
85mqsbHqahu+qcAx6aOiUFvJck7nxLcTPTsCtfgyJeiVBpSSttfkAVFtOyVV5o0AuBjsjBEdKqGR
DNwF7G0DBnAUD8aHzK4RKLMW0k5WSyORkNiXeEgHcEKtATxGAOCnvj0P2qG4GlhKley96MMeD8M5
cFsviMpyGOI5yemny1vU9dGPLOk81D2slQMjURfqIHSayxHqDUtPcvvR7lwypx643/S+ibyTWFZm
iu9IGqAnxXgUl73RGWh5B5OcnlgLnmA1TSJIiQNmOwDhkxtNZVKNYNwJ+MM4obFkaLOXSReEeGVn
Be1JpD8N2TUFOXYNWIdfpNzkfU0WsG6TgC4TNYnKdFxdUuMov8UMU3DBpVkEtnWvBQDBMMAZmjch
978EjYRq91nTeSl0WKxhnzIUkEnog131Mw3IWavaASV3XDkCNGudpWFtozdSR4LvQEjNcVMJX/Uk
bApvxsSl6pY+OXYImOAIGRjCnDFlLhnxpirW2EAPfpAyzXsmd/vcRQJGPJeOar2GlJkao/a5j5Ik
Tizl/DXAUArBJ69PiVEAXrzHnZAEnildn4/3/otDtRBn/o9C2aQQhKDNt7oTAqTvWfgmAeZdLR7G
9IOfHVAIVrT2bKHNvrtD7SwhU45n5G/Z4Pi79qB7Wq6H7Za85O9o2QG7BxF0KhPPkADLeubYAlrn
DUzT+XRUYKw6wyKXzRjsA7ra3VpLJ8hYBpFu4kvZ0462X73Nkx82NvcxZ1EBQpU2HJd/Fi6qdT2q
Rq4NY2mCPPvOQ/JFyeSQcGfokYBnUSEUSFEuJlPHWCv/9a8QnpOjOAo1E2/CQa0M/67F7i/fVptw
njRiLLKqz/Vi8XkUYvDqmGHNzmw6gQqCJpnF7oK9fVRgz0YFV17nmmKcXOvi14WHPjVr/PxfoK5f
QyulGESfnubWXo3TkFeTIN70/j83MVRAKjj9zYcyI/xb7c73YKFr9n0N3bhf1x0qjamd7DRXZCHZ
JoVEizEdCNmo9ArjyMQIEgQlcyHgyHBZ4/U1iEzTMEtm62AcUe+DXWl7n4DLHh7FIDcfZkc+IZVN
g+4E1+QbsVFGQsaJwczRKDqCRWx0rTmhzgpCU77yT9M7JEc6j5y7EvgJvgrbBKAkaEW+ruYJu5Yl
vpwqHIHSD9puR8Z0kbKzulTkrhjsr4MVKIUfq3tgAJ3xjA8h6K/NZ03GM3BdVDmrsRjYMxRVLAtM
j7yaycmQ3vVa+n/+CbhGjzRuYIHe7Ii7vhOFjCrjIgLg6Olpn3SDgFagBv5l9NmGFuO8GGKZ83mB
eRF2SR2hmw9KcMRuyLtRNSqYkAfx2uE+ypstOXkb+GIg0ye3NBa1Q2RSwLZbCJCj/BUJw1sJ6NfH
C7lDi/OJ3USgp+zPmqyUaxMwmNXSv4MrOS6taG6yjWh5oCSGEfClXKL8i4oXjwOnWYd4IZ/ITytv
MElmZk6yXgLXzJm+QFWG5ImxRRcEfNxQaaa2iXJBfnnCHTbaevoU3uzHfoZsDNcqVcMS/oj+I8EM
UmS8D24DMazVfi2nldrwkJ/cXnO4QeFnub5HaqExYJPbBc8RlwdY+OWHsF0zEVD8TIC9NGdkxsND
9F0FscoE6et/Ntt8OiDMyK5OQouChWggYuRb4GaHOjr1Qk0EpJ+LnYzWhVj+iojPs8GUMcSl5kwA
vThpcuN+NAzc00FFT4etvhGRkfTsOfKgqdRZoi3tLTScEad5cMT1Fc/S5oQc6GS7aaysYl0HqveS
nlUXawhe2WuGX5X6aZZBr3xbeVgUGhpUw8dMRG4xpVzmaZvCLumZ8vVR7pNOAml8WSjDJ7DqcjV2
IQqqdKtCMuQCGSZLFbqwDXcAQnRceX+oQJJi74y05SosEP7rixhn/pyf8ERoPbBxl81muA8QRiSb
qAFOCsyAT1ZSetDVAuvMK+VLi89sG4kr/9zCUQKkePr7E5DjUgwMKibJIPp/XDDpDPKVUQG9Y5Q0
jWbpuyQKsqR7UeXL37XDBUQbyrd+ubQgXqhj72NXz2cNp2QLBIbvmU+Vi2DL/EzJZw3p+ZMUj0QV
GNym4SDjRD5Bk/C/cwL8YpaY7NTS2AOb7ANbdGd7E7Lnmb0+RUP3OtlTfL2AggywjOiBnznH2R0w
NPXhjCc1LSWEs39MZ8nJdVxiYgF9Tozc/THPZVei+BSWJWHQ0DSdyQ0FgQ6jvF5n864UvZuxyaKH
nNmNjkSOqRXBbFQsjnnGX/QWzWUu2Ucr/p09Tj09RrPHztf2qt14vacQHM0iHFF2wYWbt3HuLbhJ
62vZ1RKFOufLICMLPeg8NURJ3zVyLiwkwJMYWcN9FDmjpIqRQivQ957xGKQgg42TtnDs6vgdOMZq
22e8Usnvm3WJ+erhoVrWn4badDKrQcu7GnYlNZUflFbyjcPIO593FI08i73Dh8IwQ7ui7/tUkepx
INvyzWabVV5enNXtT0FJ4DpQPylmP9ZB2vGmwK7nPWSvSQRpWsFhLMdrs4Lx0lNCxVZwTTEd+kRT
HusfFXR73UWNtbI4mk1G7G1M8sFq8zmd1HCsu/UDYtY/ZdQoyGTC+qvY6DmUzriclH2xaZgDA1wK
Qsslugg5yMCFFcOyuUktq1dsFnMU7VAs8LrAjfN1JpD1+73ybYZiLggH1Cg4rEbjns9g7Qt7HD6H
U4TYT7OBOO37oJK7sNAUc2CCulyjWmLcS3aatBZD3VwevmpU+Q8lwO8LJNSr2zPK6ECNSiEawspv
6Z5jqXTRj3UX4EwbdWV2DQXpbuQhYhkJa8jXOcgBjnyCYepDb6VFckhXFtlPRNgMjDCwz2ceNMGw
rzXNkf0ULeOEFNCbXZHWGhlGr3rR/uQQW5tCVzigOy9ObrZfImB/ZDYG7+nOzeFWJeFQG6IzDHwv
UfRHRxR0TbizuwbtXc624Cd6gkKxpxTfvmvooDBRa84m1hUd0Kl5BQTxezBDTMKY5T8e2YpasG4b
QSeZFWBuPt7wf8wHeLGglQi2sPX2WgSvrdn8gxgYJu3gj0fhMl6Wn83kpDScWQn6LSxH7X2aeDjX
Zv5q4Bn4wrjoPeuZHVAJ9POzJUsP9wKK33Vj8k4mRYkLrtXH7dMeV+sPWCJBOt1ZaEq4aLnvrrM2
uAcU9lGydf6TAcceNaTq2kBO9ukg3hX3UlWa72dibyrty7bf9lgWaNTU3/fym6yH78SSrdXx5qip
P4yOCOFl+XlSe/f2Ag2n0OgWsR7Tti3PNrRF2nssClkYSVRrQnnrRihccrstUEf+VTR3vMVgWZWP
fkLjiipNk5aBXiaicgHaA/tTx15TPt5eJvmY3Ah2c/L5g8JUOrxdLTOg+9F/2/8sYuH6GHtA4Z3K
nbrTo5rVjVHurKmgsV6XLNLYLw0a1/ylJcTmk2g/KeHRmmZT09THegf+bZal590QtqdpRkSSpRrV
2lMrluEiinhWYmLZGhHg+ZB5NX0vuFcDjaxM8rAI6pvzFoGCvPRckP0bNWXzzIWJlKsi6ciao+Yz
VYwnMf+6g9DzeBccFeZYYNDWP0dxKwib73IK+G/aXRn9+KUYYNLUtLpCKltKwPQN7SLtewMnMDT2
U9/0kuVOaAME5blVJJJpod0qVTkC3FM+bgPRhL/cAPp+jUHRyEo7uBoNMMmkXYh2ZNh4NsmF/zBv
OvYrbr+6pPxCr1Wxh/eHTOGGb5eQ99DXddlXYVHWxGkHqEX+ZVakdlYWnr7BtFSESK1J/Xtn7emt
Kya/fLwJi+fUM35n+iuDge72N0/Rmx8SZoptyNzJtq7SumQPwMVQmDVaWBj9A76FAVjwm2aTeWqv
PfpH21XzAYxYyBEHoceWKe9nQ5cY2p17vYxO1RLya17eIhsidCLYqEP+5RIRv/aZ1b4f80+yOps4
c3Dx1hIIqK0dkHeFMtooDLXIXVJv0w52A+LBIzNt+4+oiw3zQYSLdoixU9gXTU+2F1EuZlEYbCr1
cuVcd9NS59lwo0chIySmfgQ38Yvb07QWjfmJWUJiqqbatRFp5amvG61jVvvCyby+z0FZFa96G/Wm
4BF3CEhCndRTkEAI31hoJSEivErCsO5Ohh+vktYN908nBE631wTu+Alq1uB5X7ihjCOcJ+BybEpE
QOxkUQWOTFfPgOf/oF9UhB6PEncvRFw9kJFHwZXzvpvsP20Jd3a3+602JTT9jAVD+SLVlshiSG0g
Iaa7iFL5/LTIWXG+iOmaoxZ1ETkV91FHh6mliQ3Ta1YzueZ6qMKO6lXuWowTCJgeRZ/X/ScSb/U7
uaPR0vXZwQ0Wn6Xfor0h6vlKT1jGkfemu4fpio8amgvRt1xynXzETrRMtXHT3I1CHKvKxRihCNB1
CsliuA6YKvD1hKwQRF1PF5BrCbI3eBblNuEuln32VoXre1Et+8RXgSVmcLrlpqTOBuuzvyvDxM9C
bEqKo2UJOQ4ph4CG6uPu4kVLjdgahOWob5pgWX4NoLkmGAQYhNNm3mKkUE1/5kLTCF36emoa9QsI
tQSntAxGSaxUixNkUUEwBJ0C+SAfiwnQ4oBd0DHT0CixhjqZ531ZA5FJM6PABO2oiu8KSzgtgX78
91dwXeMlaI3m+Vfd06vFIaAMcUUiUltHC2fPCE1hlsTmW+tnHK4U531oKmbFZzaBAVfbIovGnPX1
SsfJQpQHQR7BHiKyrsuO0MhNioUANW++/s1dzlx+2BJ1ABSUHNM0POfeL/Woh1JAx+EpKG60zsaP
lnEDz8Wx5ABj3pdy5GHfOclE45Az70f4DfEyj+jOzxvwzUx9n4BakWWf35/MQx7hqU3D0jz04u8u
jOsLpUIsqzRP+iK+F4ZQB9Z5mzaqBNv1PXD0dNI+mVChOlv9I3DFXxrzbC1DYHGYtrW8CweNMd2m
tpuTuI51t70Ai/37GY1Xfa5soL5MghE6TTq3x0dSN5L393fGEOHNPp4RpwJIlV1dx8sLfTuUg9uM
nmEn6a8I88Z70hot16WNHWCgTVbjPZ+yI3Cut7ZTUl9GtpKxZyncAvuZW6mfkn/mif7BJYW2rUTV
jDHVO5hxUu0+f9cFErhDoY9vCSN1mBMTwxsxwHADvfolW1LY7fXpoDtLgzXBD+AoLXLAl+v4hXBJ
UpZSEUWoVZDrwFYT0gK+3eHm39YdPIAbsa3CV+i8tYHzBhHaT4okuTOr2nSnPlDo2cQr7LW6+xvO
amhmQtcjslzq0+7yB23qWMWlId2MqHxkmYOccscBnZ+rj2JbSh/OqKievkAUyXyaGOxSZETep1kb
BCWjmnjJYjzA9VS2TCAHE7nJmoKpRgI9eZOSag/aIe95re2YTTQ8jCW/oI66EHWemwfKNwmzNERR
Hm6Ypx4cFgHzHfdTBJ95ojFZE6ZV4jQ45eYUelmmpCcHCNxRyZDUFgFpJ0DpCMg94Og0oRC7YLwy
bN6EqD3C7SfcWA2NLJWZFT1gYzCU680YsL5qmGHj/3Ax7dhTrijW5hLYj8R7UPWX+svx/kIHLdZO
Hep33ohbhMdiMriAxGmIdLGUhhPxqecB48YldnNozLvdZ/7leX5zntl6vOaEXVvV9TDYwmV2KdBJ
dsOkvAdNrHYca30o1Akaq74oFisY+7G4I8GGbO1cq86pCojqb0GlsRCyQkTR1C4l2mEIkmp7w5/A
wqdv52eisptiX+yxGxPTpb7TneLzFv0s+5ZKB6W1qG361Fqh/t8yacqwAzBHHzCeNs2hraAsy1gy
ixzEYcKfrdoHQ/nSM9VZkyBK/cMVAKKJQUnIWv8kARSWAv5sYvlfTN2EjL+wfmEU5vOgJS6JVwKC
4rtIR4wyUt+LEEVD5+bweBu9z/JTH+a27y11Bbh4oS0u/5nS8DJAXfNtv/P2UropOEAwZL1mlwW7
DFFUMDp69xnV2BLWsTR5fy8DQjgpmZsoX5IY+IYzXzYY7DinVd5SrhAIxe2qvXM/Dzfn5dMkZjzI
FNEuK1eBzOeHXMje++66SE0jAKZfZ2vGBFzBrxS9sJ2Qm9sV2esmpLBFua9yV+MR71i27PX4aLI0
nfy0wwejq9eVvCABMhI9C1lRON/qLBMZibF8MPDEJvaNMVyhWRprjNxUZ26Moch/3C5vYHMOCdrJ
yWaP5vYvfQokJG6tDLvC70fpIve0ZRBH/v+aaJ/9xbdQCJqSybq8qPUj/Vv8QqW1DgDhTG1sFNJL
62SMX0lnkakYdP1Mln0GmLJK5Mud/SNk7kMyZhaKjAM6LSAeIP0CwEB0FSPdc0ZVdkD6WRboI9gC
X72HpBYROVZ5kjXUDK7OZJUb7Bar+frmUDbeQJod9oZtIcJtIJfA1ApjLuP0zwWxS7Gco2JMAsHk
quL/exnuNQyfKUwALQwq6w5xnNc5P1z/2fStCR6MhNPvutGgVU+zjvTXsrwVoKVBmZzi5DesPNDI
VqxUSxgz1SnGXZaEvsecX7gimRKe2HtVvQiHUdpuwtl88RjjhA2k2H4EOniZ2XzY2VeD/ACe5w7r
PPllntvwvtDP8bv8LNy4K5vlmxgjJGDGo7978KRO+6YP7Fh5jpOHN5anS4D3N1uATtm8HUml/PG1
DxiM5cvvYfv2xc8zFCG9i7CWykfW8+cfi4PoIs0V4snA8KohzPJDnq6Jd5mafb9JgZItNZhhpMXm
++6yFZGJUx1tYlORgxSH2qo0eAwkLxWRUT7/ezgO1zWDo+2i1t6Rn2EinPfiRr4rXauSVmhpqRfM
+lJWYirmgzlI5BNqE1u+oVVT1zuzmDzYgXJxWriNrn9ReHKqOhLrPXhPAVpiWBFvv7fnBMKPyDFw
6KH5sOd77ZhehEgWUmzx2x46jTrD0zvfpINi8YX9FKOfdGSDFkAK4noZ0ygP1J/ijQGdufTdUsry
1juRdoBNq04nk5tSBuTGGkBAB5pzdjZiRNIzVryADJllUKVTav5mC/f0OpGj2MnMuA27UX/I73Ua
QwSL04MLVduF5sNDTo52utIFzEGX61WpI/P/bh8l3T5dWi7I5W5j9IBWW+xGcuehUlQDu8H29Mk6
O5gl79/h1Ey61zo8mgRF8hDWN+EwcCBEDHxLHMIPXOklS7IBPUqKo53357roDdyTXgkA7/6umFeX
W7GCzV0RMcZVmBIk1OQxWatDyTCazgJOyuHTQSLDN1kpqPlFngUOnf7Bg4qthmzL1QVeH0akn7CO
7w5BfThGYWP6EHSvXZ9pzCTN3il+4HYkwVPyOKVxY5EfOMvBiADeB/uYFn1fRHI0ZxkCDjOq1Pfe
OZiQfuB+Udkv96p5qvxQqlkV+zYRYB9hh1ua+t3kTHi3FQB6BsOUxcqMDwIOxApCvF6OTSJE8LJW
1+CSsH+Wi4QErVqrmlOerbdusFPNRD0800defzBlZOLxY+ecwpQ9Z92RXMYCnrJk+JkJmT7zktFT
io1+bWrCqGyzbT/iO0G0/UR7XFXtWxqaUs2xswLBhB/1PStNBraN7xr1PSeilPShtQYgRlHFCBLX
m/2+/ss/hmHP6MBZ7+XS2yG/DcBBPq+84L/M8dW2IhNoIvOyq71W5zDr0rx6zJL6kmW8pG7JHwGs
WIQUAQKCd/CBkmAk2BWPCxjvJ+OGpmfVjw5QYWZqbD0u0FVaKxiUot2o73KjNcG0ozGYnLtgvMJt
4spU1FSZTnyysX9ihnLxjYT18Uy2TZ3wT7qwfUt4kzANFzytUJUAbJPzgnW+CJx+UOAPCdSBi8e4
lE3qtFXz+qHRdcF+01Uj913zOMvcCyJ91QqXQrvhyuCXrd6RuobhxzyQM7s3p5zfJid60kXo3TFZ
0tUFzbJiVvyijXLd2tjzEo+aX3Gxc61F2oUqC37mGXeB/lYQf4JwZWkA6al7DyBqY17L2NSxi7YQ
x37CL1ne7HDj0pAeZVSj8FKROIfNusp1glaSRNM49AagDvg6eh8L+IIBqIZNggqqhNODGZ1sU7aI
guL9mHQ2SizNMuyH/p2IGvhx8HYtrP8huh6VnvO72z25wnNLB4AG4HW1Vb5QHeRBqF2ubajrGRET
tjvbgfr3e0vJwont14RVhFz5oK/xSPL/NMLvQFWloF0Z5Z8Gh9J94Z2ug1rFSA1nTPDLO5Lf4VjR
tufcqokJBWctMyJGZl4KRES/55BjwOqhmYEL/t3CDmj0U0ilPI4PFBPUTKZv9C7So1Lb21tlZ271
w+3oHOrQj3mulwT2pf8VIuFmkPfB41c4T3U54xHldqqug6eJTPgznU0GcygAkF3Jwx7WYFiQOnIl
l2uUDeI1yUvXCnNXpuN+yVu8MI8cqTVQDcFv4RXXaaJZftjYqI6enVmie1uxA79yshee/8H8Vz77
TwLVkcThDWyMDTNAhIKK0VWMR5s4GlOrwDbabO+8ymyBFLjF1YAIg4h6p8FGcKH6PFl8KGoTlrwo
SjIeckewgQ5wPmM8/VSh0OvJFbPAHMGOGOYvlYITv6T/5x7h2ZQniP+MUpsixl+v7Sbawtn+sHoW
puVAxV4+T39rp1ioY0SdMkKjaBRbS4QY2vr60hFCH2vj8sBhrbDHPjUoXfOM6pjzVZ6ZATGVvfsv
f0lG7Gm/CxCsEfmAXz6ViMsap9GA+lAwWs2jd0Z4kmV6EQ2Z+e75i6UfvYabq04sh9dhf/YIo9XK
1M9kPFbx2R3GAUSNSdOOBbYKS8Klq4012CdO0RLzpBOdpZsayGS0nXTxFMRbqx9JdfmIUZKK7iMG
6r49xN4W+sa6KZORt+EMTA47Cmoj3lCTNXBa1YUy9bIcEQ8urS5i+3uNqaBMzE7jRkN/doRuvrle
uUIPSmDZB2eOnRnX0OXhSjq4DlWhUw7QIy8clGJTVKvej/DFgSAcQ7Yup6F681Gs84NOwtd1jedm
KA5TAYtVKpiav2CeCNG/MrweSvTQKQaLHIa7KNBHn566op1mF8jrokNj7fshxqPuHtS/40ci7jWY
uENuyG1P2F3VDXaI8FcJ/jsLJJUq/nSv4i1/RIKDwmc85QRPEryHiBYCmV3TebsoZ3m8cb+nVtUO
EwMlcCpcC3WUkVY1OYrTxP4RKXRpv0NnO/0e0Rb9eWXPs/f7mTM5MvS/3lXDmPXXvBUaUwfz5MOw
N37ssMdNXIuww4kgtCdZijTGOYfskawBwSie29oJUYi1TDbEG8D96T7fdiGLW8MevXsEhVdYbFjO
cjCJhFCJ29iHK35nFnViJvNtMhtxClEgtqaCU12WTaL0wOeOqLkFCcKQOPQcjgwmMJC0lKz9mZTU
n94w+B/fHU+XPXiccEdqgUpU8rmafJvdiqzt8lgjTpKdlAMnm8LAosp1WSqOPydpplORue6YmazT
ASi4m2ObSdV28r8fJEstJqx7y9eMWrIxu58EXEiCAFV0NiPh923HbvngeZcHBny0Cfyx7oMr1onY
+Do8Fgo1fiCFDsSag16ucRjHNh5uC1+LaK1dNC6rCQKq8ztuC3a8mzObV/THEt5+XMeuXfD1zFr8
mqZJSKZz2soZIjROnKy5HZOqiGzIFuaouH/3rRtmi/VkCXoK67g61Z1ZX1Nfl/n9IL9gPC+PSR6D
wiX7T6TF8hgAhVqmmaUz1CVC2YEif9Jp/Gs0+REpa2nkBCELgxK92Y4rnauQdvGYNGp3ve/f7l76
/4llDBb4Jr3O18rGahiy0ZWrSbxhD/MSFirOMm0Si2iS8FIYenF1q19IOY8ZUT0L+zPpbnj30ITd
xDmBypxJpQ6M/bMlpHtISZ78krfA0W+1+ppUD0lqMyInlnJ3KYsIDaajIFOP4mXaoxMqqpOZTst0
OLd22J2mgEVjssBTYe1nhul9HIMrmtvppO6LAa58MIPQAm8s9y0OdsVVbxN0roZIwjgtvzjI09Jg
FbBppqAMYewXkZUwdfrm6UGJ62d+hXBSqOR69dhvoXxPWGjHRLd1II/qY1EgzOgDqasyoOgv2eHm
MbSjlhh2CYwtjnUAhjznoveVcZMrsMRacKJzzHwDO/ikkiU86DrVmVuJhv77S33UQy7NOKwkOr5k
M2quF5qAkOYU4AfE9K2TZbS2+KNOah4ZbHpIZt/ZwBUcwfql+26lgGxHkXKArOPKnnoAFifXQTmu
ChtpJzMswvOVLNZVm9VjXMdHl/3ZptM+e4QmDxClr4cLO9gi/xM0JOu9cXeex2MDoUt+FB2f979w
ilB9KY2cXrJskU75zvj8V2OqO38HH4JdYV5iASVT5hSuEKic33qirq5RTuB+YHmmTJktG2UmDD2P
u8BvNMH1uUwBvNo5JwjmT3Cx/pFzXXdXV1XGqAB6uW4CXoEbEJjRa2w4sPTbYLZzG/JV0uxVdhmK
jM2cr1JQpnGVD3Tck+0v3CDCmWsRs2gwndJVi5kN/ruL9Ad4N5i8W3mc4b3nH/91wGqvD5d+hiN7
vJNReyF7cKVAAcbrAHtLgNcbU47GY0mCA073+K/4H8dQ1mrUE1NY3xNuYK4FzvgGqumbHDB3x9n8
SwC0/ks1Y0B6ZstflgmIrzPdoBD+nLVKYNA6eOSPvMZ7O/8NatwVI5YMAOhhUAfc1hLnQ9NPVdgh
FBFv9ofO/cEDBvp6GNWgcAeM8HT+OPnvmvjjTov4gTdUU3Gpwa0ADgn/azyiEsDtq3/Gs6rUiLII
SuHEb1yQzxTIUnjNhugW/Eg3s3R59vuGSC6q04hQDpysLjxYdE7Ws7hNM5p6PqwT7kP2ZzbHdse/
UgahN/g10cn2usgsWeHrSX7n/Po5V7v9C29yWv0CwakHzfaJKzeMV51BIrl7N50qQ7+G03eK8s/x
Mlfrvg8oqvhWjcZ31fqaYJ1Zlzl2NVCRKnAJG6NFlPIvyk+UZlWT601LaQYMWaAozGDvNWrhZrn2
C74CPOCblW2Z+UJ0MvvsviINZyc+t+xpk255bunzO4SAiIiClxLmSLZBNO+OTQ/pWUr/qQ+4AIny
wbA3Fj3pa/Oaq5uV6fBJcl1bWTUHddjwNnnWZCF9aMlFNZThBfZiSCEvbPjLhcIyt/Oe3CP5/3Gn
iri+x64074ir9jF/fO4buxqAxteiXlXVfz2zSRMpulnAfDhDOsvRnmCF7ACNHPg9fnpn4shh9z6K
12wS4eExbaQ2yWD58F+URKuvNCtUN8aDjQOKVFsaMaYbhLZoLKzgpXyYvbskMOCXxoQR3fW/OYcQ
Ci0CITqdOj/sivXbuyahZvAg2JuAnRDt3bCITea+BiL0JFsPyAoK4zVXBiQlQn/Hzoaimqx5tCE6
nW4R3iWVyQY7MuN5nKlTia4mlRHSL2K8x6qANr2Yyp1KLaYcp0vGzat3LOxe1y3dWaOeg4xqFUOX
tENXzdx4p82b7fobLwJrzSsF1aD1becE3RPKFlTCCqnz+jQ8C4FxCitoybTr++9Y1BuNma7EkSZ1
jZGzlXDCASphTZfh5YxxbREXeLQm6c4snkxeXHmd3YrwdeF/g5S9a9SaJ0PljDtHI4rEcpk0DiLE
kB3KE1ME+xoUeXN2It7MPap21M/liHAoxAYXNA+CYMYT3Dh//egx3EXhYU3Y67I8HXivIFKOTpcw
npUfGFcq7QbpdgVUgV6I7ho+/ChFPLM62C85/dYgabda1StCjoEC3SYYEJkV5Cs08Y5TyZfIye7z
n30j5DJsDxwDnDBtkilIKrh98RWIKQt4kr8oLHkn/etP8iJWVm+ayvbQbRkJ65UpfNE4KiGc4fT6
43VuEAOsv9i7nuq1ZoonI+qbAwK5/Dzu8yKC+wO4V4Lxi0+WMGmyvCfFrObaO92VaLcaN0UrbN12
k89aIjtoECIWkZWo/Wt943sblVYam04ouqhaPRH8nekS9r3Piu6c0dNMULB23cwhPWuoIAYOm0XC
LoQDKdQUeG+mkN1rw4dVkvuNISW0nLtYTY1GsucMf07mARmXTVFAgMABCpTMQTtjSe1DzjOFmjYO
ffOo+eztzLa/8SvSdihuIZgb93SrUjDpDSU8tn1fxdnw8WPwfZokcQxf0+kogysxD9GPihOT0kAg
KNSC7E4Sh104ZNqnZAI2ZW2wWhIGRkGO7JwyEtD9TLGbYGmwJxj6Y3N5TptzHFiEna39Y4BhJl+T
3HhhCoCz1nCfPICFftUPwCTrSOBjzywXRfykaXsgl5Z2xBW71dwoFrHEIPa19FrF8EHjCpx8xGsj
/y4LVqLel4rG75LHud5tyy2egih9erOfqVzMuGYW0vb7Ue+EJqCvmo5VXc7Uuk3VKGUpI/TEtNnr
xFpCxvjkNv7WOUo9vHbj01HkW9yQU7308OzgOUMuwdR7s9i4N4DEs2+ARpQksnSdepPMYnQBPywb
H+jsyQjmVwxbq6n1VZFBTa+5KlwNA7Wt7/LzswqX3LKc7gXPUdk9iieTNWPOBzRPkRbcKvSfk+TO
/ElzSCeXbC16LS6S0kfx4D+idJLYlQcxi7mEXd1P1zMxD9M0no3OiF0bXWE2hfnbduGz45y8mrOx
o9gRDm+1qcl99rXQYWR2qD1Axixmo6ggdYfrTi9bVJNme3GSdeG6Z5C4Q+iliCx6/1cSlvqsnuCK
Xj6xLQz8GRax+DMLE58qJMmEhD4tCWCC01zePHESnp3wWeSNV6WRrpefDJ6SATCHrz06OoGsQsy/
Za+mipbws+lUxvNpt/9tbuhBHqygvgo7Ovbh9eUVNpqauGEEycPReXrG5JOlG0psXfJn06+aE+zc
i1nbiW2b7I4YCZE+nZbGGY6uKTZggq0onylEymAuIDRwHDdrYO9fMlPLgojR3pSUnEK/2UO6dFr7
sWODl/WY3jVhTbXTlPJcMTz5G7yF6EUrc3S3IV/5An6IdBOg8+jT5ZpYZCqITy1V3AfqrUGK5jVK
wSkFK6y+JFcRxMG61f3kkZ5fJMMi3fxGevzMQWwnj1g/yEJyvCCdulcFzOb1LOVZRiHImhW8Uowa
D6Kl8KlmwbVexs1vYoCT59VVqfROUoIsNk298WgdmOlugECXMq7D1yM0IMOQGDJ+9kEFmiNyw0aZ
LZWZ8ZLNtOTyzPLzO2EuS3Ok3uBc6cYCNEUnPc6nhAb6UYpk9unMKktPYceXsauaT9m9x6yswreA
iZLevLvJK/HuWdWY84pp/wnUA6lrwrtHX6he+XnKAWungaLcuWZVPJfowpO3yBiTgl4lV7HWcILL
KZ6sIhruz+btDjMO/N7lKR5CurREG8yLijYHoNTKbT0f1LZYkFlwzwXee6g3ZqX82S6cEkGhltZ8
0vuURsu5pzy361HKwAy+hjUG2/WDzuWpktAEFYs3opwrKLt4pIG9KF115G7pF7G4mTqvk7n5RxMW
EtfFjN1NKvRCR/vbRa4QcrupA7z0fd3K5WWiNS69M0Un0oHEBDoThIeX6ldk583hq8Yt/ZPVT9HO
TyUuappNqnGysgazAulBnRiYij1aMhJo23aCbDL/LZusxnNNwgkxjYfpx76pezPfcv2Y8Z3mzXTT
89nhsYF0nIzY8sZZQAUz+VJ4leG72LMsSSERl7MIXnopYytk5Cd2fzrrUBkKBf16MkJrA5q/d6Jf
+5Rai+h56kKy+5XM3DDtZ51hTg8nuzHsEXA+s3hGt2wO+daaO5K4EglygydY/uNB23YJE5Y/u5Z1
xie2co390kBuNT6IfZS+OTdD0TR80JnXjpkaAuhd1K/77lGnzjWcJYZ+g2+7TkgEfbaI4u6qoMcp
hjX4fN135E0xFExGpoj5VQpF5EpG+wSnMzbB9yzRbiy7SCqlgW/uo5n2BfhezBRPnopI7ZUNSFj7
WSWL964sw8semXD2iEiIl0NX6meVJ5IZIBL+vLpMABLmQWOvqQC2tObmDHy4BOrzOwwg7NwN+/Es
+7jVeDAU/ooggyFub1r/ydJuuKfPs3jVgp7YSfxNDap0GVOpqsbEskc2w9l1uYVr7JjZ00pyWHwe
LQNfSJ8tCc+wcJXPTbB4kP4mp19Salf+QSdOae6TTPZDsTwcuL5e8NYz02Z1uxUqqlz9FQlC4jdO
2enoevEzBJcTRle0B/PyxA0j0dfLRPc5iXSMO4JoCHdR36F6i5+L/RcPTb90GKJLGeXgv1MYqHvH
cwXfOC66H0g+BacFo4v99wJLhhP5x8EHD8+m9toMD83WO1SLgArn5pItGID566TG2P6TPcRG1MF8
ApuvCEyubl7qEPM9vyhhx48BYhPano/QZftdH5NZZZVpxOwbevPXvZVhMAUHqdlNHiDlp43eYfZC
0CaWnV1f8djKYgyBN+GiVGqoc0z1DYSnD6X4PutEjF8z+vM7CZ5l0lA1YcIutg3X9pP9tBNDWBMV
kW4RRadDblMGQZ2L+jVNTJScmHP9lBHYApqDpOjBh1Utb6lfmOa6/uJX3DuJCIUAmaWZQfZMUkP0
Db6RRBr1wAio8cvNkwodlbRVLtQE6ABNkveT1LeaYDfoCprGhFenOl515cMdWzSNk1uWMcdustVJ
ezku70EYty8qJyLBLgf4xOQgzkV800MIhvdGdhSPrjdaiusZbweR7xyiX0YfxJ2D/z19cA3C3Zzq
JtWEVqpXxyG55M7AG8mjdhSwHy2UhGwj1QQsweOE0QymnfZlwJNmhR0hITy5WaJbhwAoctQLfw1a
NAqcFHYYFM/ST9T2afFiDS6/96ACpXbGXXPq7kqpObCGHZovHw0yhKz+NnYXTrE6gTSn4HUijHiX
FDZYBZrigUURJR2f4D/9rLr2PhLRWE0u5jSvxcKrPP2sKzRG90IQvcf5XQBzYAoHH0W2ovYgXWpS
zbepQvxoobTrR1afM9S0LXJhBkkqg7/MeKA5cejw7t3fhj+rhT+QRauuWMPG5hdh/4HKyKeZAMI6
XscDaND1Ugv5R499rKA2CePWcSu7nR2Ag0fBG+aSyKm94zo4KiGZtdC/wfhKpvxXVpPUri9blSTI
ztuU54dgRlJxl7JgPxLjBzn1jrUcbfYmy5HSYJQSa+1wwiQMcUX0Vmxq5AKGq4mIqGtwJNtOPxq5
V2DuyDorHIeGIuWN+dpRUEWa6TUpxnRc+WvsRIbgKPxY69xTMWQmQCaAdTu1rDJOvwTPB1MMZvBD
y2a7u2H4JIkRpc54VBpn5XKlmv8iJW8WHfQK/eJyOGRxLC1vzQ6+zBK16FCws5x40YVICW9nxicT
lV9pd0dOQW5JJROrCUu6os298AvC5Sc1PX85cttG1QnG5WW/OLysqOuIM4XK1wsAUJJM4RGVOWNG
q/bWstEie6fDK77siSFiF9nedqgvevgrFnABJQaf89wRT+5PVXIG4p2DXtordpYnehjAV8rH34h7
rFumWDG9b+zYugC+zb6j70KcPLMWWygoTv7s1/gpnvhtgDVLQjuj7PgADyUlpriCa9/gK7+yz489
Hhm9bQlS1Y3DBLRx80qI0UxJlFjUCQRj3bbITQnQDBw1lrKobWotzEZooZRvgPEyL/1hkVAWgPoX
+tE0gh3MSi63F8Yw+qs5XaEOCjcyAmuSYziEV3OnJFpUUFPKACGAEvrVFAEnzY0MEwU614YLNSu8
sCbsu78Tmno4+OsaDMR2rq4AqqqNAUpRtEnyFm3prvuvers51wwOtDQMqTphN6naXGsS5YTHIiEG
q8tJxgjPV2uI1TFWOPrjiMwBOqgE2YYE3LySC6FGQXL1sBpvOMJ9Se9LDsZSD/0r8Sdu9fdNvuNb
/S/gaqzFzUSEsuh4jF6bhTuF2T+9jgcfL9t6Za7ldlDiRSpPISZqP6J3afnqQ0Cg4CtyBkA2Npzn
wLgcX0i/5q1ixhB2LPBJX1w9AVBxj1qEc2eVeNnm6oS1pTB8nH+lIor9RBU9cw9DKSBsP+wTeEbn
9lharXwhk6kpBc5yfn6RUCSjquduM+J9fgZcqYshowuMzjUvBFjmsdxx03w/b8YQ/DniPmlD2rJH
On3y+OZK9m0AVFVRQNdQGTfwDVPSphI7q8DF9vScg5cAiCGJ3mqS7EMQhAfUgnod+NbJzkewj0gR
nMz/skrRx2BITFRFmMMED2E0dVqdzbDlVLwsZ97fOvsOh/Um4N4yZ0D70nltLgOM5TpoIwDTHpDo
uydo5FnoQzu9CdDRAg0LwaUuKSQ5C2LtxfXBgRlSy8UM/7pWG74cu03AG8ND6Qc7IwdPHthJLkOs
zCjAGANYJn3OLfLDkEWdTbS+7Tsn1PNSjrozm8dZ46qb8KUgQVunBuuu/hakxr6ajHP/DsHSaQiF
jCsAj6N6Oj1ygYkXZSKJDRwakZV7io97BYfdS8NbxI3R5PitQwibtQTEVwjURZGKtSgoQcQxWHSF
U7Mra0dbocVYm1odtosW4u+aD6mEYz8lg1lJYg7AO61DpTy8QTRml9psBRynnNxBddz+4wENag5w
G+xUpM/RjAvCJsLDoqirbLMbBEWQ6USBCAox0iV4OyEGLftI43/c0ybjHsFMiWn8OaScg+eVJnVp
7UKH4XXUotzSlyBtS2J/avO1x3ibrvSh5QJ5aPRhmfgu9rc8QpOZ9yjALCLHC9QKNGOyIU9A15hQ
Z9L+Lrx3Crt6n9/cKKqVXyLcZt2U7Hx9v5baSJ/XBS3jJowG2tt05XjngoFwLp9RMNdRA9nvK75i
SnuSO2SIInaIelrhqBlHlcn5ncAzWwVDnoK7s6Se6tF9+/46ps8rqEBIJ6dJk8zU2Ty2CDKVcxMe
hVeuokJAy2uf48/dQ51PjV+zsXMkyfSHVTc5SeNILMvZUH4UuIiDk2qCf4ADDHzmFw6rVGUSGXdC
QBZAan663SCsGaiSl2nxMDvZ/pidhJWE4us24jiw27tN3cP+VIIvDouZXMz28ujy4IsvAGgeivpa
ACwSpnSqxacAMlQUnsG/GLjnSnzBK/T+mNhy5HuFlynbfJaQJLWcbYOS7ABdYBxpOn2CStBiNhIl
PM9tXIZJDN+njb75Z63yamjQhEyuvo565js0rCXfG3Zow0940xBzf9fDSn9o+HecdtOkETWsfu5Y
MXuXtJIGacwhVFUTtIIPewuDgGqmkcaUolzvadGemyShY6sRx4GPpakYYVpBC5hXMu4XFBj9Y40c
RfnVI2+Cz86eWX80CFvoabZOMgYKaulH4fwJy66k/CoQZUHvWoBS+kZ/TdGQcGujmPdWuuMt+GlE
TasaQo11w9e8blkvyyI87803HoDuApeQ7MVQuD+3QOKakmOTm3avdqoNEOdh1isSwuq2zjq3GqUw
5lwtUN4epppEfyZcuXu8of08P2UzklVrT676g1H1fNix/av8nSA6ViNPJ6ljqFRGNNLuI40umvVK
B5s8r+QKOU56uO+llcVWzpTB4IGmdQbQyWZeOooy2/kJrPyATp4jfBVSt3jsOwUctIzGU6VdVyn8
nw3rqWwDJBPXYPt7sw9t3VHa5p9iLjbpdNWCL9jp0K8ZE0n2SkBOFI1dVxQEvzjxaY2po6SKeqwe
uZgwrfp5KupXUfxG9UQ4h7xfJEL7APsoxL4MAYwSAqdtWLpwUIrbAHpOCNLCKxV8vHG/zJaLmeG8
GLCK8MP29Z0uwZw6G7KbNekR+z9ieiDQiQOLA5IVuak4nf3sy3ERNXrjYL3wiI5uHZgLf5Dv5GAZ
b6Ru6LJhpabUta9LP8xoTql4GRdU8Jn1HdZQkOkNTAKF9KgbP0Ih4cd/UYq+UP6Ap6iBe1R0HDAb
Cs1wZ557V17MXEd+kCl3WxZEl5KJ7gCDAtD4dlup4ktjD5p2+oFJVe9ZZPidZRRRcsGjDejaLO+0
aGRW/T1aAzyEdO1JkgLI4wzhBBsO6Y8R7Nc/cxQojWJib6lINEpHlyTTYNivvfHaBtZyqIDXzMDK
DPDuknr0dOugBIvUWJtuGfapr+8gkb02zkB5P7guMFGC1DptDowxEg0VYF44UowWvVKMyVtztTNO
z+aK0Z9VQIEd3lMVyQui+goJxXJbsuLpzgPCUp4iqR7bFOb4V1FLqZFSmUz8X3UOo8lVnYXnhjRq
HLJYmj96u3VM5IbUq+vHgvI12VCnIFzh9bsY5591FMQaLwNtjkVh06gkH5eooSvZKBFfe/lFYBl0
GBpN/FeCBc7FK0/6/UhYlecxHUvzCiusHD446/YGkTn0Ar0kl2z0Axu8TXMZ0YynFT+FoyjZuAPT
yiDIFVFQknl3taH0e/P2Y2+EyY2T3Q9ApLgoVYL4yqdvvNlfq6ScSEpB1uc2barlnlL+DAEy0EHz
hXmtMj/a+EBx5T83ABNKlV+RS3qujLKfoZ+UZlmd8Q8fJTjbtKqTR6x1hNObeMKnwEpcY/KFMADv
YqBtolKKSlvGdj6KczqqrWWhaw2Bl7j9uVlbnQIyWf+x+6l0TKIlZ0M/07twkDHV+m6r3llzE/aZ
c/LDL+o/lt0KnO4vpp1s6kWMToAPaKAzTRyZM764eASbHYs3fSCscvb9HWdCtJA+tEVYkz77ybh7
n3AV6W8mdFr2zHsjp5HwDJPzwXFvPzKtCckRXSyWKy1/23zp8iUkC0qRhjY5mPJPXby+tCm0rHw0
jRl5JXwbaKKs0Y+YpsT12P5GcRXP2nBQzp8vXo5s34wnQ3rLLeBPxrb0RBNSpiEgP1Kzvb9tVB21
dpyUKtfPgufsmzrPswNLVP72ZrVsejxkPil0lzke4ESERcC8QXFk7A/Zfh2lTOGopHCJ72MseZmj
OdmHcuih+woN5diSIbBf/V6GryBrQYJ2+ksCt04bzy0w7fjT2VbzIUDr7J0FW8+4ZjWZIYUmomJi
Kb68kEKhn5n1xEJq0QdfounxvMtu9kd6TAsBp7aqsccM7/nPRsxPlyTlXBkx4nPaTYbwIlModS/1
f4QAJmbRwYfwVUdKyXkFtCGXgPG+a3MRHMOQd2z/7SK+yHMEfYCwonRE/hN16UqGag3r1OW8Truv
zZjD6EjuCnEKqRHwF6VQglbyDASvk5+zEKddXKhre/8DNXC4U6w84RqxpWX/xO5JvY7Rg7AUyv+6
Ie1tgPxdQfqkxRWabkuOhlk1G+TllhvoZBRbuKpZJ1aLWxOHjxiPgLe1gyFVi+0eXe3mlgNeXQkW
Vc2/Fs34fAPpxZ5e2UqXyD14UtIMwLp7gunU1tJw8urXuoiBZXwDZCITQJp1WIDYDUmdhMCZY3if
3k73CQNIpLMzoKvLR8U5eT455+XLiUQQumJA4cqMKtDhk7dGq9FyKjNFlOB9G0Zz1/HkxzbziYMM
3v1pci+VTOk5z0wbMa6vfteUrgZHdnjcMkktuTBD3xRlJJdS9X0CiqJlYArxs1WK3vhXkuHhNsiO
2VPURRw8/h74v3aRbCihS1U3PP6ZB7VcPKXzq6ajSEqRClPNa156SqrimP4+zbvPWDsKqKdwj7DP
uVJBc6KLkSbwVl8hrrGubmxFEPg7YwTH0L49KUhcbZBWxxmZxH/9YGKoZPGIGnJUMdFkh31bfXOv
iATu1PnrfAd/LvOT+lClP8Urkp7uuS9H45nKuLpopWoker5pToMXHiMr008G2mDkCBzwO5Jr8JN9
N9ydF9REYzsi7y/3Tr9czJhD93hG56S+BcZnWxKEkLIbkOWclG8idSzGEVQgjjJn2c/yKpmxih/H
IA98x14PQ09boYnYmEupZcVSCOHmtIevIqeVAtjFyQEbXGfefUp+jGLv4EdiK7OZUHO8Ox7tdcH+
bn7GqOGn/6HUU7JjSqTSQeb1EnECtvGx255Ijzyx298Ifs5ZJCLf9hPHg5+jMo9etpKfbRFjqpDw
4hwEf9NmAv3sFbphw4NtREEGRw7ii3O+Lxf3onwp8qKBebfRtLk/dMgUbZYV9ELXn46h3kz2SxSQ
qxJj3rLnmr18lprpI+rLD8CRoNgRGl7Uwh5Sf4bcc3zfgpF3+30k7rS+5gYRY7+7vqNv+PKRROUl
3WC3cJr8A7f/uHb0OcBRG1d5TrJMNc/ym/NmWS24z5l2BYYEfig3rhTUGnf/kjwrKHFLShyFdrJs
vys51OoRntcDF3AcC8jkvo4SbKXKJYYSBHrLgsZuDBf5pZbiugHzG8uxl4eDRUZ62g+3I2EnrgOc
clrW021N+4zvaelwe/6njBQAeHwPNTUkPNy9vdkKiREQKY/uxGEWEWA62cF+glUAVr0Kh8piKiI6
LStYWh4nrQChqBthDTnFxkXYES0Auhhk8IOShzw8d1MlFVFN6d9Z8Vm6Z2seq0XRIvH6BiCCyT1h
eQl2ZUq9y82raTOmN5tmhrPgPlzPCtJqTDoRryen3BAirNF1r6GSHkJIHHNN1pu8SP1lHEP6KEPB
E3ZUFgcFH6z/FolV65FlUN3q6tlBUdvKAAD/Hq4vxQIPeNqiuKrdCanbFxxxdrIVmuEZOc4Lw6C9
uuPKJ87Yow+YeSK7lFuU+YaYqjDx3pLJ2D5jIvsvhTC84XncKZFCYj9uxWf+DzUs0td0ed6Tt+en
7bGDgOQpSlDt0CiNM+6znEqGcqRI0zwGr/ejYnj49hThG40UwUPVaGlGAa0TK0v+vURtECYUEMs1
2uKbfind6Tlye714qPd8AWNHieFAUgWOf3s5WytFKvvn8eM/j/ZYoNSGqek67+oiCPX78fFpkjGA
SCFUv9ywrkME0guwqb2MsPrAlRXnf4DGH2Wur2YOWu8FUKanfCuwFVDxuINPYXM5+ftquglKZEhX
rc6mvh+CJVT3pJv/95v13yuN8tVb4XuyyZvehirJVO9qGwcfagINma/byBkKsH+37VF/TCYvg3Xp
3w9ag0ksbY14RsxFnq+WpXZ2/0Hrm1TwaPgPbyXEhgqrChyJJOunGq6gmN7gWuufk/CoR25qkRPs
XO4fqBtB/8oCj5Tren+C0RclnoCOhlrh4K8d4GZBoRtsuBJJBgs+0BuEjO7hQwfdP1b4Djw/Lizr
OXDUz5137xfMmAKhQo8SsEFrbBVDdvbX97QU1vZcVc6YMoXFWyFWBXv8pyKP46wvNayHTxTf3SXG
MGPjOeTegPUZ+7pZYpIeP/vh/ADeLgIIjU4jrbvVW0Gdqzzg4zPyBHrJnjF+S3Wgx04OMihGvrHc
S/p/dPQMDAHj9lrMDJL3a8nTrLcA23B4FQ8IOvP72cvcY64gNuncGHTgcHJ8q4oYIoC0jUTyB7SK
gID9kDkPXkVLHcUvTAKtn1lstE3yyxtO3nueSUFU3CrKq0CtXU2egImtbYQdJSRRLf33s6v7JAxk
aFkeZpU5g5mj2H4yFgUIEvWXtElCJTJqyvJ6+WB7UXZ3oC775TszK9SRxKmPgamFfsD4HF16nMLQ
ibrVCkj8ri3o9cyEtG1afLlAzEJagRxUCUwrmNnoyDLcDn+cCv+uv6NpdOj3ZdG3ZZgqPgx8QGMp
1lBrLQZq7KFMOmA12/CTQYWOufZzuPh6HeV3eF7rNt/Ls/lRqVx9JYb4Hqm4sYu9bclttTVM0G6B
2ggX2HPVnZux1wddw+K6/oyWglhvBNODGVVH5QEXjlWBKe7H9M3veGwBNlCbXNuxow1n7nDGwilG
OZrzIIMsDNqTDqephQxfr/kaWncmEYfipSr9FjCc2CxWg6Wm/pOH3Y1W5UHxagX+xvazo+C4yIOV
S/+q05VgBQA7Z+I/jhoWhxV3SMRmtbRDziJoUzM/yabq8CLkKUkMDgf3qEr/BbguQLAXu2qIxXv0
vnzisVmvOhb4tYxh/i23zHzoTEVRc83ANNwjRQ9OXzWrSHsoNJpha+mDyLzYrYQUq5iXezrz0zLy
4Jdh/TBN/5iHSnAJgNtWmUrUALzRl5QRnsS4iFviG6dFBQ6b4f+DVqWvoxo54of1+or6JWvqEFtj
x+9QOWLng1nSHKkFTPvIO8WdLpf9l1AOOs2zQnt9eReirxRBx6AYrgwBF9GItOdYkUeSoIYUiSQO
ZW5G7k7OGG67mwar2qi9aMW1qFbNRcpM0R0yxmc0U+w8/03rrVvdl4p/BDqI5uWFaIfOPy3UCWF8
4JgmJv5nhhOgxayO680ZuF9ldbg3ZAo8zxMtluqK/5NX6GnSwiccyckBX0XCdCUGDAesjq30pm87
hK0cDTh/15JN4ta0X8TRJ++2cD9h79sRZvCEdABZXpasEbkWgeJ/I9/CSE1syXoKuz/+dNtd5Xfn
qdm3WnJ9vVwX+mknQcPtL+bHwSFI1fRI1ZIphO9xSzFkq9K4PBrzHVoLBo9YfD3BXlwLigdJLSj7
Q/hoUDi7Zug3ujPWbWd6I4rdjBjqakr9yhP/D23H95K99f/E9C3eVfBZDIBN1C31OGa4Q6b0bDfW
S4WVTgjYg3fUbZeek6gkXE88RfDuQmzFENt3MYrPDpn6+eT9rNvkJPX0PWW4Mah/RDchbMq0G8xs
aAvKR8nTSVFSafk8rDRolws1u9A+FP68C511N4woQjNTPdv1Nb27rvYsp5AxcCZLUan9BA92jMLQ
mtI+lZ6dMxjlRZ6k6kxNDb5KlrDjoU7U4cy9rvZVsPSuw28SgIkX/PRROcNZBln63O0JKpcNiJAD
liZ9Ft1ECumUSi4Z/2bsmigKdlPqMiKLdvsqzga4xp/4K3ZUEjpmGtFmoTvvgrorzL5c9Bkg0HYy
3iXrD67Bp+crly0fgDtZYL7JsLwtq/S8KIVUdyCSukivfbvlyP06G671pwRrkgbm3o/XWmY+ju4d
FH/XYPiK5rbVk8UnUhOk7tJyIdRbPhR6yVn75tAfVTRumxEIn502MCvfU/0CH8pooI7NPHxgROVD
RyZvfwmK0T1bo4MSFPLGRHQMy9wu52QPJThD8VQaAG4uAm1Al358JgI5Hd9mrbdvViUeR5sFYmZn
dmt2Icr9k79AnzUWkKEK2d9jKHSNhXbLwCmE5IJNooThCKtgUIjDY9ZsPF5mozm5vvijXF85wBLq
jvWIvdi9YZXPAuk6GVyMonYgzOoXIq9+CHv+Fu47avzsp10uArUCPCuD3q5S/ykvLcRXTY2gmBtk
tj3Q0PozskgJJW4LMi4QLMrtDQjmdORGWgXbrHbZuYW0Qe9uS5UWCJobcdGoqofOZY3VTCppmQxN
T+q48OEdOm82U2UVXxuVXJLUeEPX0D7ydgHkFx07XisV6eo58fqQeo5e9vADSMuVqkKEwbGxYvkj
tSZPlmut59TxaGU4TeVyQAkTb4lHkrn5fWTFCzmmxOlh/ISkjvwm0FCEjsXBrT08UVC9hG/cUFJh
N8XGJEEgn0kpI6pTuj8to2uq99CHtChqvLxLyzAp4/9i8i1rM/JH3A/TbzeTBEKwiEgU8qrWkizq
fOa3zwoekPOOqRa+brZfgTrlS8QQ7sHvs+HM0PicsCnv40m1eleDgcy0f+8gQQs8V+ZsohwYzTV8
dvnhX3MmGfsNyDWwgWpjANS0ohI8LFvwLfuL8W8JSfZxX+IvPj7eviKv7EpxSu0C0Ga8wQ3vIu1P
DahAH7Qj0EHFM0bDX3xKFeq7JLflDmG1+bUUPH6pmCIc7/izUP2ciWrFHTaZdjmQOiiNpRJAjJbU
FGWoZjdOfCtSR26AyepMyNG1KAAEvm1Fh6+fS+oeWcoJLp899RjupLkt815LML+4JcCEafUCtxVc
ysFoFgwkNO2p36hKIyrtdQFqJJqs+5V8KTRtN5CsZOri9DmrUhzTV4ihn9OVr4tDOmgPswpwVfHv
e5qmE+cMG1NA+aeookyrBoii0jDYzlI7jx8aYyQdoLBeC9Fn5CG12UyuZSxhcy75JlDvtcX4tcBN
AjuXPdN0gdBpfnE17J0v96BC65S/oUZ3w3R+WwJueD7LuHEkfXnNzZwsMkLqApELMQ7SUnd239Lz
aDSMnJXRuecIMk7h7SrcHV3L4IcWAE9ruDx+xXt6HCBtsBOa3+y2nH2ejUtDJxF1fq0km4YRT4Y3
WKW1JqlXHoY8IcKItkC+BUQKVnhGm7bXE9UBE3RcfIFFEpAlQjH8mreXdUMAieqSR0TpAz8dChde
jkvyBye6gc7r6G90OM5g9/t8QMlwS9E+XuXsu9Aul8ZdYQ1D59Q9a8kIFn5WP90lsc7vDU/SUKo0
OKAUqefPv+5WZx00RhKb9+PisvpIiHaAmtDXh9GaEcmClTyebOMoCpNBE82fGFiJEuSgTO+K7nvK
JM0cKpieDJJlKbroL6gREknfZvYwUfWM4Vyhs8UGr4Rjab0XeytkZtBe7/ay7lppBWteRDk0wc0M
SfCzRvDzbVwme/F4ZZOSgRojPLzXmU2PWQKbW/oy1y/MuNSNi1l38kFIQRWcMZii+deS85DhRLFZ
QR/5lt+oUbDP+UBfRLVyMPUkTdFWZJZEXP6dtyrxhbK9fVDGffVPIktwOtI+yJKnQm0mMY141mHf
tXKgO5hKmX+4Lwpq+T/fZAXM/KVzdlq7YfYHd2j42DIwebFVzpJm7O686OJRMR2uyUbOD3icc6p5
qpxmG1UPKM8vRr7hlfvlfWMGtAEXOallNP7oTiTEb5/OOiq/y+7qLMx/5NKaTq8zMHDtaapkWmrw
TAJXth+0u3tgV3xIXtQ1j83oxVc3yMNZcAkR7Hq4miW88NqpndZCassmPoaJi9nB4by1vYmUdlrG
d/WrM2XWW96bmrvnCAHE24ZyrsRaVreiuRSMCGvjC84xCKlpfawx+Jbj3mv/du0eld0RWvLNcrZc
CtxepI1yGkY/9quV7HNDH4JvrSz0BgMUb/YkD3PfA3OcdxnO+/u1eS76mkj4kVe8ZmkArZsrduGt
zA5b+JC+/iDA0NVyJ+srK7GQ1UGzDA0VXMcKAEmRVYVK0FrJCxL6xn41mPZs0gH1mNyFov+J6Zo7
pPNDIKv9i7ymWqkCP8qzdx0T5urDhCsVA44H1oz+FEt9+kHlBho9Fm3WwJpDCz/kS2n26J1Rns3v
2hMh84IV10AjvDJIG+LOIjSutufOcMb93XqW9x7l2uDASUegMZR+g5GOevZuo0thcsPH3dyBsjSc
X9h5wLsnVn7SpAMiLyKqSNWliDp17H6n//s/71H0wdrIf5YntBbbMpm0opEQp87mglqut7RYpuQ6
NOA80cXax1Wtw6XZqs1sA0y5dc77cV6yf/QDtSQ87m4OvZeufjN//aLW7yY3Z//QY7YHiFG4DyZz
0R2B4Qhan/gSuNkkoIvfqwpH3BGPGSUqddHM1NjrjW4JvC3W83Tjd3CshtyRaOs6MjSU1AworHxN
JABsLa9QDRt0ruQri9nIwkS8+aWuLaATTDqmbBJSspDB7e3ukQWRtAJxWjybZXhbCwF6ne4chAfq
inhHv1zn8KwNAVKsfnEZOBchf+teT630g3H6CgiFDwsDgtG3GKi3AngzHzASOxnSUfF7mmfDjN99
dSAZskh5My928cSIAQCCIz8KFGWa8b5fkjNi2RKtcKgrNOy1F3q7WjPLWQWHZTGbcCx4XBNF3kBG
cRKQEuH5kyIaNhnJPBJvG/65iWiujnE/oncszD3rZSExZd812qz+1cida0XlHKWpYsFv993YBeeq
TzUe6UEjz9OI/0zy19c6WiTlavw9vs9kFFmxP9hYN5yDQfy+oimq2Ltuk6uY7lodyI9zR0Jlndhp
jBRVkbTBglsPPjFv4tF3Hn6Tx2PFOmtPrudDMqoCUTuv5pc73PIK6ucaWVL0y209hGST4AOcHg8/
ewf9o8SpZYHkhGqGDghtb9I16LUa4Or9HGA0+jL/MJISBinO/32Z6Mbx24vOuO+B/AhUgppZC2lk
/qWZzvMhriuqPX4kNVySBQaupcQZA/DsWxgqw0I5TZuQPT80hhDmQh2p/3V8/IS1HSIloBPs0xgD
5r20ZDDCIj/xPg2K57E1LZW3pnPsljHX5Wcovg+1j7jZjm8hXSKRvVKk1f+8AUfFPxRb/PIpZpTm
2hHTAvDWcMDrBc3wr5mRo0SFHmecTLuO+reWCZy8tizBcb05C+XCQtw2iVAWvF4/asUE15goglup
q0/hXybVz3HalnH5vpkzyvD6QQAH4AnpFT7lSStb0HjzcStsVRYV+xOJVLN55UykvVmkb1s9Czvr
ahxsLKk6m1d4UpFkMZIJdP+wDOq34xRJlsHmWB0aAzL7yiU1uKl8TSr+P2q0YU1zKyYt1ucHaJZc
2YsU3ttab21T4MIaazDOEH/j+TuLxmvtd2qMHzxuccJE8mc5WTJlk3oCfRy3N49CFDV6HtkIFvNQ
28E3JyvVYdvSg5Ka+2YtA1sK0PO16Kk61Wd/MfoPoe+2+uJeAZqxgOxf7uTDpS4iLC+qB0+56IgM
A7ybjmxobMrsMu+opTKo/ohi4HAgYRXn8BItJDTqGng6dj9p5ea4imNUgl/mYfn+dQmSeKxH/aOJ
n1ckIOhnQdc925jYJC7biAEs7bp/gT8/y66iW01tkM/yCfGAOTdKHDXF0YH4QoDnTZYKjrna51EF
pfr2SDTG9B5vuWw/IiWhzauP8ZtqzjdTz0q/nKLfKluu2Enn5UsD8sUVVIMnOAWhEcLVF3Dyn2ib
Zx8hw0c45HQykabFU+ThthDRNA2wZ5EJemAc0G0NenAQeEXczWRCFiS/L7jeoYu49pvbw/yDYyR9
lrFHqfHEWddZDtozqtZGsA7VOJVxNN0jm52e6V2LFNittDVxiRYF9CeDM9G+GP+Y3BTnEO2n0DAy
AopMbGVqvCKG30S7+jtCGiC8ajcdTGPt2r84oCvcwVXsC2CLCdtIS6krjcDvV/ztS08NdbwEHZOL
eutg6mN4rpuf2hXrUnFgrUaDTPLLh/FJm80XfALHt6U6a30AgskNltu0uuRlQC5F1D1xcs0fnzbz
7/JC+Suwxe49P2Xig783yu/yjxivWTepoBak1egx7fH4eF8K3QtxhK3HbiuGePapPu4L7S1xyCPE
3NfiBfdj7WsTiO7QyGjqx1M62F3uJaB3leo+GcPFAYvvfW6zeaxroGhebd44bFuZyt/u7HxMlI2K
wgdzAyCwSZoG5go8N7XrQtW2Udg/qP2VFiHbWFFCEJUWxvZM9gY3EyUzr2ZPCxqw3E5Cr0WcCZwO
hGCI2vzIoToR002J83AmLlfVzHOEQdg9+0J5LSOr8OuDcpkkEkrC2WZU5+PPM5cmcBVVxLAwltyw
prPVpMuoImGEYq9mb1cBm/jhXiXt+/ZtgalnDoLIKmatoaDn0jZGd+Rs1vbkecXudUr9vEJqGxj0
D4VuMdAfCbQhUc3GE2MQtCqAUOP57wTZpC8CLPAwL1XeHhA1ppbnTrH9w1guHkTm1ra4890XjSzk
wQYwKFm+ItXK2hvUpoxWpedGWKAsncAYQ31Cenynku0cJaJj6Ao82xri0EzTQn0iY8oNn4CGowYM
ivKXEIFkoLWLa55xsOmPQ/JNVY3er+Z//iDc41AjqRqybCzCK2zQ35nsD7RxDli+BkHwhSgpol6+
utMX6a4EW356XdeHKvKbMpKGyluZ0ImW2H/SQT4I0WNSeB+yLCh/wNBvYSWoX3GuQ8f9B+soXaSz
w1PQK6GsOk325k0fciLiJwljNLA6J6k+7LwAvd/14knyPbQJDkpChuAq7qy0bSwKxqGVsec4poHc
YI7vD+t5DOlUicPHVuYORxhn303seVi2S/3oPayXxbL7mR/QJwW+U9mOUqBHEOCXo+xEtrE5P+Ix
EIhStcen4jQTkfPF/lp8f3mI7TQvBvQb0kGPm+D/KHsO825J6UjRWEtFSV4EKEottQ1iUFzUA5jA
ZudPd/F1zZ8L0JJV/zss1GTMe78nzD92JfBPQaNYBYenjWElXHifQJ+ZwJjFYMN0V1VA7uV+S7lF
D/RbIoubIEbtewrxbY2IIbeS/YAexiT1PyTy2WZdMPL6vFKD1OdpTUYxvZyBudLJd12RNHzAJvZx
FQYgQGXZFeih869YrkMFPwq0TIartBhq7qpGalpJE8jh7xSElKQBL+UfpxeMxnoEQzqv3EWQMtRs
F21W7jNq+FT+SGeIv/676RgPma6Rpb53Sx1cbB8Q5CikyLdgKTh+3XmI6aTh0J3v3AzRJVk816N3
GH9shPpS0h1dM9WXZAIvprXBrBUCDOSI6xERjVE6V18nxVGM2O+1aT6H8mF2VWEuHgkDWOnZwoRt
EaI0ta7fb0zhN5A6f/0qP0Nfq8AKxFsDLz4R7h3GbltbuGKxlkLZb6yuj1KbNR/E+y0CRaRUnMOX
8/sMv/lcWSnIpJqn8GWYO63WgWT7MHcZeNAnGBSOuSXHOTraHL1T/RvP9zfMz7ys12X0HJ1Xic2w
8R51234BzqlQUPye0fRhhPH2cPM4Vrqm2Dsm1pXSzpFaORzJXp3c2bMas5xtcTOYVN23unvIruzu
kWnyk8Tigqa8ddCenrdX125Odn1FfLJpRhetj1urIsUutJfcbZ/pX9dRyt7sJ+LAOLr+HpeLgs2W
8ZS/UK1lHxqR1hLzZ5GC8e21BhshDl5cfEYRkAcHWW0Kx7kDlDGCyrdEfYXkOUvOcn7cNPSIXTLI
HvCReKJYFyFq7c632KeJujzT+7yN5A09Tl7JQzOyukjlXSqcxdTyC4UrT+lVr2WVZnvM+79pqZQg
7AVGJRQ4Ac3ucsWx79y4MG+DK98A4L8IVbU1HMuidGnYHk8hxSIjgzRfZP1CDNVBbraA2/IYM8bl
vI+hEcPpeyayRqdF+x6CEAwudwaF7lsz0lf4h1B0dwOCQXgHHfKHtuBqdn0X9v8WPmqpQ249/nZY
ido392IL7SpKwqp4CMUl0F8tyYhhJDtA5LBQ+L8cRXcDNdNwDt7oRFUVjJa3r18HQmaaq/PZjc12
zC0u1OUwOXuvbzkdcTuqSwgQKoEdWVLqKLAgw5vYtxdmdw4j6KEKZZ49+TDLFzkUyfmOClgTuqCe
b9oaloLFoblcmg8tfKd6tS/l4masxWGdIt2C4fyF/AymdBRW9Q3jDn1xvUDuOgt0syEyj2aPdlJp
Gw0m4dziuu/MR2gXRpjfH39cBTfAyWWM6ajuZvxTeyCazBzFmulR60F+Zo8yIkI0Lv5H4cfDpbbO
eG5y7dQaDe6LPisqI7ki2JLJT28DR1rTsEOYgrLSDrRMY+mBopTJ4xbNWqEs5MQsxosjgWcT43ec
GKpAACA5X5Uytztiw9/z+GcKCJ8jPFP603Qj3akW1C5kly0LH7mzDlDGUHBhew3gOu5vFF/sfLq6
QzwvCF+2HSq24+7V1lWos4li2r6UIhlneqFU5RxxWQ7s7KoedY24YPT9iPwO01w2sAqKb14aliwn
V9eOTRM2Agj9MWbE8DjXml4dIIOtjzi4SYbmlbmoRsCEPJ13QgEuKyd0JYsPJU0KjzP8UHI6vx6l
PIxQ/zLpkspd0F6c5muxKheuNEpv83UErmJgBo6nyGONceRRiDnrch5cKgeHnw/vKkJ/5Ptr4VRT
mneb2BohUJI0Rnwk+soWkyGDOuQoJaZ0U5eTFHslEqCbQWpgvSqRQBLrYtENZ55P5XWq9a+MVBqJ
DGbOk6T5V4nkv9eW3LL0G6MmvLUFLhhUUNZnqItA8CG0vg7nBSh/eWiuw9j2bH3VsWS8DWhYeOPJ
FYGSpJksKMPDiEdykEA46O1zHbSAVMwPtcRx8k11Bk6SgwWmPS0aBeCN+RC0KlH1qoc6Fzijy/yd
8tMZffBlzWybEFFAEuRqpwKRpNsGH6FeF2m1ic1UzgBQS3visFmXcM4uhXDt3DiPSZ5pI24uhxXU
SY3tXC9a0qf5lzjWyUZnfHP4uATzqF83ppsKqTlu5vC12zPqixwO4IYpq4httcoqptKKHb9RYBo6
gbZRP5rydp69tJy49SiXAKbPoqE0bpYpVlGZpdGeLOzPwhUPL4Lb904dmb2rklkNIYXl43pTMHEx
Zb41bv2/gk1ZjKBRIJMuqB4KjpoPpPxLZkRL6dUjZMNLYSLoawkaNvGs1LbGd7KtZMWwQbrVtC/L
/9zeQ67vZUvH+2FSbEe7sr5M33DhPHFRpWQFAqVc9BW0ayTc8QJJ1mAGwuRd+iiRpxXIvHIUHeKE
kK/fUDBgfKO03QZhnnuD3eiYoyd6gwRljK+WRAO3jhr7eAGTg0bx04iVxhPUiE58Sso0vRcsPXUR
9kcJRQld7F3JIh2sCt/mG4UsPGidOgtQ6NT/fTTXoeeoCjCT1801gMOIc5egLEBkKW9yxUoeG7n9
rEM9Baj+0c8LXGPTJvEj0MbfCSDs8GKJv/JmCkTB1NgComngt6rt+VcCuOlQtDzyg65C3qgLrJzM
iOyS85gpVpwIlrdGCSfI9nNJRMPhYpAH122xjBSBMd22q9W+19RZe6tVsgFrHqll3VVIEEFITEv5
dioUbKLVsEyX0EhGtz4wOmb6pXmn2t/r/Fa/kLpnaoY2/q1IBvqzC4iGpXYr6ZBMO1mcPfNTJyEv
Dm+dLvZ/941SN7ZTXIVjzot+kRlstwGmWg1Ro8ANUI1iQEo+1d5DvVH3B9+MHHzdTD7VlxvL/wcJ
Ff1JGmjiKWWlOY5B62wgzvmZGh3OY7kr5XJkTnUh7uIJG9daE/heU5AQB3YFgDV9kv+pCWuuSMMC
I2lm9UaoR9cnD/7RavXWoy8jf2ZB/CkNvI3h++sFjaPwNGhddPxXM+wwkQiFSYK22DCHt1lNzWMP
FGhHQ4QsVuPlaag9+Dw3nJ2U3/UaHGPKfs2g6tK5wz1cbjrssUhsE49KZ3KMOBJmNGCBkvsGI1R2
M4qNSTaQ/8RWa61RL+Z+MVdz/BNQMyAtTME9LatOtYEplRqfw7cYZRnJZtqzZ0ZOWxoAE3AEwuyt
2uCZELAkWekGdr4E2bCng1AkQn5sGp1GKnm/1e7tn7JHFCHChnNG+QuJaWQAM4z/IzbfWsC3TuFn
uHTThD74ajvGKbaCNu65bpxTmAtrE4KZMqpC4UNyCGhIm1CZ4tRpivFVe0BmeYRx633u7gh5m3d7
4kMkiB2Qe9Owj5l+st3P4VnOhmgTPan6hcfOTzuS0W/41CEjRCg3aZLxAXTDenRguKivuT2mLLLo
fU6jIMGRNIgC5yWty/MyUOC+wrxSR7V8U+YB7CMFWnBckl0sK5sMSzFL7cSxXdawPzqZXsm7M+pf
tO1e4SOaXZ6MLDyaFjprAlaEBFoupmN75WX+AgEA5NMs6JJ0cXvLR4MVzDa9mxJCNBhg7e7wfKUZ
mdSsM26lhOJrvNve/W4AR/46OhkQPvia/oSBMeiHDRh/RlODaLY86RYGoJKpxOSOGfE3q3ULgwS3
MZv76i2nTjSCXSu/h3r2AZT0U8EBemTd/MCIlLASeuV0CDyfOt+1vvP3UwZRou6DRQNQUh1fvu7t
/35znNQrDb8XvURm8ahTwdKl7IReSyTxknW+GEtV5SwyaBKa2hHmvEYTLQIW3es5zI77qWJuUZeq
qq3r82NP4lZR1olChHeZtzlV5E0aWliFVBBQ4n7ccsErAYOF+lvwsW5SmYxKh+y+x7o94z6oN3yT
xKlAMCcIF8LNjFw4qXkoGW7dTsdh9/z3CCDhBgAF8U0F1w8X809jc3y3Ntg2tYFP9N+3ittGncEl
WVo28dZKTCT8YjsMCy0J/JWukO0ZQmmgeF9wVjCGMJomV7Ez/gJ8FqCMFUz8ecyqoMAMfm+skjOL
oKrQ0RGjKgk99vUp6ePrwhnC7jOyNDWdPp8/mOJwPnmrwwS/oYHd8/MEDweQhjE19zNo7bbXysa9
UKxlQ5AUsqBg6gNCDYIu4N4w5bXFX59P+RJApn0YrgcXwzuZe/1zZgpqgbikexvCneshPMQxk7IM
IMMQ8YB6bR0O//4Nzj9Ig1Zrxwhxdbpx6tDIczR9C8Lhh7dKy5VJTF3isNLNzUdY+BkatpP9mkAp
AS7xxOMLWDxnc11gc/MDhnfI6gBbBn5ZtjNPFE9sJYxoVNmoDcd66tYv/MkYuh1gZK2uo6cD7FcQ
AaAbfbXggXVh0xug/7h4eQGBp6B+gYuPUC3x/aE7RjsW50FcIaffxWYBZDDTwxnqhhud6RGh4nvG
wCTWjm6wERtzTheRVFoJkMY5cQmqcjJbxLfBndF5cN7U0fXkrL/uFeDt9DfAU1caoIf6g2VrK0pX
Q4zlWsWRYtaZNddPkjTLLixTR1/8UC6lHBi2kwVPwYbOKrbZk0fSfMjwR8k9lVxMak+QeXVYTt4w
oba+hyAISZFMxO+bJVP+z7nHUnTfBANcvj/7DrEOrRTcyVyTf8/sC3bJwUWZj1Vfy8Znpk5T4J1t
MrDbjKhjQL1ukAqF0ExtY+Eguw0VocoP7EyUOltbZ6b2G8qX3MSlfvGJGgEmdi9ZutT4pGvSYUv5
oVqtlar0+2FUTci5yKnJwhXdGP+R/7kLseD06Su1LI2+gFhyumYRl2+MgN0PVRv6klJDPI5JPl3e
Gk8QGEGQ01YO/0pp2eumtSjFbJQpfFpbgmTFhjq+rR1ygsLt+F4uRl/lh4z8gQrA2OalU4pxh0Av
UV3fooiX+Bxfk1T37SP7YwJjXjG5sJMiFXZ4gP6kHv3GTZN4/Y5Vb9B/r3Ht55yc7siLlMDjmIcs
jIepRwEkoPk2/OcgLCdqV5TS6wYnYEr0jkbXcyjxtyb5FDgIwo1u6RCgDPVPop39e6SvpM6dEMcu
4ZlWERPFjArX9Sj4O83x8XY1viCMgSDdB239gJ06d+cuJ5Kn/tJ6X87yUWCV/IJl3Ywp8VANttXZ
n2/UsRIMKkkipRTTJsg4VEt2RMF1bAqM57VrAXKaHb8iK1bRg+u5e4OEuAZKsXqaQw9d5cLHFnih
BI63z08yLcA/h+Ahiwzkugr+z+OR9vGFrYBNtGvrf7eBcjsMD+HhN4x7mW0j2UkzHgn0tP1nmk/f
dg15/Uq3s/fID7XjKamvhLrWKkIUMnR9ScFP0e6Np9iuu7FzDjd88CxxfvllaRuUi8p5h4Z2+4gT
kQ9/w3PLHCoBqW+K2/RNlT/3X7F+6495JPPnn1R9zWlmpXjOGcwhWRIRJ/lTLBv4dcm4OZWx59bq
+tUmorttVucmN9u9YgmXK06ji4pn/Vgye3e0E7rZG5EAZrQaQIeQOVu8wg9nVLy66yXYCF627BoO
tBe3goi/NYR5UYINFjVXQ3+WrvXeMFXk8DtqAl+AB27ewtOQwqXzSRCPqMYVWVDPmt01J+E7lAKu
B0dgqpcC599vFAkoO9nvYLIlR5RsXwa4Gt/ULjI0EIuJEB/TZeY8UoDW7Xw2901zdSFFZq1egvcN
Amv+UR4/dcnI/2CqxYX5tmBDoObUoS5Udq9eVYCGSuQ0MxFiiODfjMM0fz4PZZjjl7KFI+X7gsDl
+n4cOXK8d/JxMXw4SuV+4tE7ojYKJD82VVIDSR7koyTs4JFbILAVJbrwMewS5uWt1avLvgTi68zL
U29FZlVumpexpge6L/BsPZ04U3lmCBe/DlGk2aEhgQTHsxYtc9A2hYnszt5D0/A2G6an2PqHIvaE
CKkO9nIpwk5YoNBGxps+ORXyIVDuZOvKv44AvyYojZCzcD322TEAV5rXaoZRU+bDgPaPzYAzCZxL
/v10L2DFAUnS+OVli6WequOi6lRRPWcXoxkghXzLnNfpJVlyFc8CxTHd+25C9Mppg0AwsP4w2cj4
90hhWPnenNSzAndymi53SBO0VtaCo6e0yEhJwEQYG1JbIRpci/iaTFzZbDHpkuti3vwDbAm6Mg4N
3up2usaDm5pFoWClV2YpDVNzncSUA9zuXSf0CDk7yjNLNKU0i1Gl7htuPUmQyVVqlj7vAO9vAn3F
1QbCm3J6qAXwmT1al0sT2Q9yNaID5Il/IXDbxUCFIizbgMGiLKHZIkgVmIVkntXlDKOrBKjZGRQH
iMDPhxWJkeI6JCHJ2WjzWWJbB/5wQLV0eXtltFiS2nEJG451kGlV8EHezj4aN/PSq0qHsqMX62Fo
v1wJXR+6SzZ5ZKP3/M+gCQ5wmW/VUhFkyfahQd+yRSzT9JEFy/rmLLZ9kzJrW0qKpzppSitefBgC
LXUtVmLGtDCw9Oax6RCT6jJ5CVGHRs/UgDg6T+CQbAe0PWaXlLqojKU5ENNmNbz2mWf6gXMcMv0S
7tPnEwI8QjcYyqxUYdDIiEYN1+dQ8BMxebv4SQf+AgExUv4gTElnK2djtK8/fLXyZ40V7ZBwQPzl
YStpA87mYgAm8st2SlGgqc4pWxVZa3oAATyZMife77UypxbR8QzoY7A9ZopL7wrEJbzxcIhdgr0V
AuI65hKeIgn8eTzSoScElQANDT9D2Nz5aLsoe9L/BSR5DYPhQYNn0zEk1YA/L4+86f6PeKvHXO8t
dPoH93zdXXEwzS11Xh7XVGPiNY9Z4MDuxlRx/pwPJtBpLQjZ5+YhAVQujO3U1Gc+GScMUQeXU3/b
BN7GFcKJqOg/l/YFf/sgMP9pkxTEj0/lfGyyDUMM2D1tNwAKkNXaxHdPRmJJrsGdiw2fA/XCSunM
3PYcNEy7EU/lkb0S0lMkipAOkrn5SEmdtq2sbk+4tP8VPDbSpk0EGx7MfhodxEGkCNlQyNjqzu0B
RUX1btEZv3lpm8u+uZ3DJxtZ2AFDlJgTVWVMiSjIoUdP/QeTfN3YH0NEt26TolZfNfcsZoj2OAgC
xyNTuV/PXM1dnnCOZBWWaTg/eJ7XuLZOLrAdz8zYwIskukPnWeTOgr8XNxvBy56uoMp9GLNMhLM0
ku2SvZr8E2M8pKcQUvcqmyyewRtv3tC/0ouDQewhyAjfF2/cI32Y8O35owrgZj8bBBRTLuuwEoNh
hWsNV7/3XSp4N6Jiu3QvZn18slcJCk5A0FOSvgETVpe59anNjbx7CKb/Ouz6Eo0lKVlL7c5WM1kY
+LKKhvQJ07QItjC7VyOW40sfw/1XTf/wds5gSLYemSW4Ob70A1ep6RMeZ+ruZCpvPz7L6+nVveSa
qYukCmxOzzfEi2r0ZG+jQZFQmDXretI/zo3MvH02Gd0zcjd8vjR5oTBtU1yVR3GFr9kOpk6R+9O3
OL3HEiSbzp15+vyVtcnCWN5fADKjvQ5dKOBDL3iCvxTUQJpfHagR3uYc/TMaJrI9ILNla1ejaHEx
IBoGZ1zKNswxxXWfIfqb8pF23Bmvj2W3/lnRevSV54YOiEJZ7t1ES0AohK6yzY32nBZvdjJKj0cl
U1976on4yJluxJ0NYT5vMVPp5RjuBVi5FzpPVzk4CbsM/KOpYIPSYhmHC0Edv94K1sfBsZ9jHvLL
+15aj8MmtApNwcBkpEJ+ntk2DLGQyzjSSZqYY3Haaq3R1+hB2bej6cpop0iS9R/tYMLwjSeCUna+
v1V5VeLyU56xfHeQeDpHmhTs2gxVBU/kB68zLogjDnl7L5u1ygVNdrtTzDqXVclqSn28l6AS7ofh
2y3fltVvJjA8uxE2IYNuvcyv72WRD75vFg9UqMdizVrkXB0q0A96I5A6pdCBFJbTNguRx5Er7EjD
cnn2Io+ZdKuEqOKkW1EtwOD+/zlzBRtnO6DzgK3s8HgVhr38UTeniChDFhscHjiXzJ8xblVlteGN
23ORlAMFsGt1EGNqScgAclYUXg6QmJ+52gh5XymjR/e5L/2rc2foc0hRptKZOSfvambBNifm//1q
5nVprfslY/DEuWgfT+lv4Q7nn+jf9PxuYmVDYp7qxvLecBAe+0akdAA+weGi+4v1TFl6uQT2AURm
X65u+GQ7j2Z/2tvTiLWb5lNKZeyF8IyHGtX+UgEY7dshiW4tfwUpnxXIyzsQQLmQDL16NVW/Ciyz
h3gXwoD3UvMiklXvtSXzAYhbdjoJhnuViyZEW328ALVbT5URebOlSVyGDvfRZK06PDHxNpAN/srV
0xOkAk5C4CSual8PuS0fA9lABfKr6lpy7KnqzOfwiMEQOFpWGgoAcAJ6m+3kd9dsD4Q6RTzS52pX
iLBXshxoPCUi4N+g50UT/zaTaJIUOK8yidda7X7OIC2b1qsmN72wU7XD+yMx06996vWPwDRQsjTK
0bG/rV4TbbJEd7rbNgDKfYQpRDveWalpM7ePBKxsnSEQAHQYUAGywj0jbL+FoiKQiJKic7Rd9cS4
yaSKEeCgkpG/M+NCf1T4mM3pk7JvRq0Ze2Mmjh44tFVNzyWzmAL9ww4BhXH1Yy0GMYVFhVLDy58P
lC6H+ck5VuHva9aizsezmTpCPZXYKULU/dnXcY6BdF862XRzwZ6z6U9d0oMf2MhrEJyFyUWxKT8b
HF7rIjhYAjyp8yQS3E7endc5MzSJcLOG7GSUXove+NWRZLfcaLkz3z/N2QOqcUsiWcuuls5NwcVZ
h+rFCFodQdGoGLsCo0VY8STI6FUSLfNdXobQK+h6AIXQJB+LkRK0GPkqp/KzRCoqxzIv+1QVDgnr
BxqVyk2sApsyLdQXmCHIlXRelBP0yo4M9y78fZGuA+NYrPPTXrMGZswAhGS2gPzZ/0AgQ9TE8EkI
7XZMxS4KdImxrAARI46tpo7xIm85LMwMQdwH8wtqw97YKnkSt7aEkVUbfTHuS2pDNiLO3cbxs08V
BBtCufiG7jVTChz1Y8vmQvU/3tFGSUI/RBRVljl0vC9fxm0d+lfj2iOwxFzARyOJ+N52yVlRep1V
0y4o3yNFb5qw73y6853Nw3/RpbotiPbJJIaTmSPYvrxboauqeVwKwTZRP+1NafhUDkg8C84h363F
b/as2LG0mRVcG1Yk/XpAU0cFUOCauWEKKEaRYIE2Gu/0zkfkYDyeZYbNiFNs2bZCfBddiZyD1Ubz
OUMOYdzOWF94owPufVMStIdgiPTKrlqAiPu/3SlOU8Aww7pZPOw2gUt1vnBTgGdaK9bUcssigRVl
fu65wFxjXUn+HMwUr5uH7pt6PsxguCwXJA5Kth5mw4O7YYMxIW4xwBwimMWbgOTWtXF5JckKBP8M
l9wFdibvFQRtjucUBkN4/GQrNC7de7Xs0IRCrFJ7k6MaP5RHsv05IYihRc8X2VlP/1cQKNe0hFwL
6YEe+AYYePhL+KkijsI7+VnppYi39i2UQ0VZRflpzGxlvZo5dMIJMJIbNXssx6sPJVXLZ2OUmWYd
Usw/2zPw2KeNh0K+JJ+Kqvrdj9gFpNujPvrzSKv2RKtF6Dnp1/ZKm+OwYNh2jq2Nl0NNd1PIPwEh
dqED4hh9TfdQD1zrOid9ldhtB6hdr3WmoecSY73DN+tReiXg9C8DD0uJQBQtiyVrEHJw/abe3v5x
zd3/Lp0Ng55N7yJr15izRedqMnURoHMGoF71v6cUVnGwEeyOphnxIt70S8m9NK5Wv5vnnU6GvDw3
S1Y2VUPbKHdl8y+q/gRR0LrZal0xiDDqU8ewxJavJzT2/ex5ACONxZY4EsJE5+WrKOjsVN05DhmN
5MzPMdB7+U5pqfm7Ed9ISDku4QIAqkt756O03PtVerpxk0ETii0nECZh37kNGSduwRsNp4tayyXW
XgPEeNvo0deINMExsql/GUhQBUg4vrg5wHiQuXgfvIJrUTP7OOTz00T3n2utUIK48QAd2AkAVUnz
aHZM5qZyJhc4A2WIaQv/tMfjfuBImjeztlwvOUrhWgAvdCC5sNXKQwF0MgXCbF58a8mr0VO5WTVO
cjMY8bkgz9mbR3W54fRekQu9svQvanMsJ+yUgeM+qQYTeKZtDgNnNmyiyJ4pEgFNZgBePi5QF7w5
/kKdO+qNVKAqbefNssH9sVYzUs+BxfYnp0pXP7/L5on+sOzhVbjdc1ABiGpfS1GdwASNIEaMwTRe
HW9zrOMqfJXxlhsjBip6rlZeFEUA06rsO3ozuPscPF6Xro4Pq82VjnyPn0y1t2BjjJvLJHYdtEUJ
rlivzasPku6axlM+4oyEWqnTpidhBF+txm4j5ZiNncsjyJLPAU1Vq4910nBs6U1JPwwMekeHkueQ
e5kMtIH2f7mPKKRJ2GP/enNkhNevPkbj6uWleJ19yian/0souiRFPCHFGS+1ecFetA7CYok4np7P
bg0P8RSmFVKY2Q57xR0uhvCUhLYjJD4b3bEQUhbQQusz0kQl1SIvIO7hLGJEybKkHFPL5uSRh4kh
HnUp4MwJLtwritRN/m2GQ3/abvSpw/d7nMW/+sNgDxLnhYK6Wv2fw/LzwoIiFpf5DulQ9E/QrUVj
1V1j+ui64zzLkffVRsW0fPzX0zgo5KDg5DFZ2SXt5ruMHOgwTqbq/uvNEAJFeZNy/plabA6/N7Vc
TXusM9EffWkrxQJTPZmrhwHGwAlAHHCsQl1h3ydM+EcMwN4q7bkjz8BcJt5spje/qaNS9xhu1i3R
PETeUbkQ1VHKjk2/+GD3/EYueNstbeNVdd94mNWjoEVzoeVuLnNOxlhxQ5gMwSkuawNow5QtDo0H
kcxAhcgf6iwbKyumWpKdsD9Z10yz1gb8mdzQd2ooqMr8yZ5V6yxhyF0RL/Wmala4KfxQDy+fMU3A
AiPU8Hivhv4/dUsOZskKhBcHqRe+WQQNY35lHez5XgA2ioFwqGfvRBuN3KV8fWpXxRIdrtApWTRy
fvHhE+uBXIKOy8yTaTXRnBUAoWAj/OIHtomVhp7kLOLRfwPB94q61a6W8vS2plvMJs153HALzlm/
9RCVxEOfd+M3S9uWqQtwrEV2GhD6WOILOvyCg+4SaJCwvI4Uc/1inBBYzoAPdh1K70/tROGwwdDc
om+UBgdoHQLR/D8cGUQTIbr+N5X0j6XcFOhz55GZzDQ8fSvLFoAXfYisBzic+tM5+qzlYhh3ZS52
83VE+89x4bInlp8bs4av/h2oxnIN6IHIKT9gNgtqk95u5ILzoT5FWKdZM/cml9Rey1ln+uSryXqF
OcKECNnHw/cXB8ENqMBHQVohXaIT7ws/RUS4MLhucC/d93d49a0DogShoMwy5QUczlvnMDQQMCao
tCNxTJHov5PrO0ZDaWmfdCi5LKTqCE4ppggnpsKYyS31GIvrXzvRCXTl/whloT17Mi8dEaZOIEz7
xp4ZgF6IQXi98PgTFSd8jmhyB/mKTRknFumnsvOysoD9dqBtp0SHi5VdqEKH/zrrtJVxFQ8s4YkL
fCC3AowfWMgmog9MIfGNWdmas8Xputa33XWn7b3kibcHAy/XzwqDAadOd0MsibHs3/GR92OkLHmw
r1rvbxKulnQ7gmk0IDRThI7CkvHee6VAsFZRfaEpdfAoGIcxGryTNPVAAdAfhX8/UHodG6PL66y6
5rokC2CdIJC5y7V2hpsxSTORNtJMOy1fakkGy1LDQD9SUBS7ZQoQAyImKrG45A5Ql6QMSS02uqI7
sGiJVPgjZgLdCQyXxfGiLYQoXQJoxW0+uqzCynrrfAI8cRJ+zrKLQtqygjpm2YkCxtxQbHOKp23X
e/nu2vkhpuHcffMd3tLSGO4v40s8xOqjO+X/BZ5JjOdhqieq/bbAXiK81CylaKKL+/5Pze0yziNU
fCaM2VLmC23jgxPIqbEug3wQmClxFCxjx7cn8rhuQDWtYkHs6jM1GWB0tG8pIw2bJ2TS3EZJSoRI
XKHL629a7Xu5VpogvNYJEX3o7LF2RJ4uRQSNNw5JI31ObAJLPHy7FPuXkCK5vStLdVH78Ndkwiyp
xEi0S1SCyoHRV9DDHRfBh8uWe8PnUZ5yHmYz1EgQ1TIn0WhHBhRzOuWq6WjupdFreqMa4XYzROWP
oGwQrHeWDqTcg7WcPYXf0oULT+iNFJtxnRdG7CPEX7Zbn0NHbzW60mDPgzLxcgiKzC+EHzDQtH2A
u+Z14d/82mV0nqi6YUvzk0PHW9TBEUamO3KybfZlkEaSABJ0g9vwdX3rwnQrCAMgV4dVthxqLViX
pEraMpR8AnqtuKPr0/6E32fAY/FtJLJ+gJUvJ7mYqyzAHFBADoIFgV7niSRhSm/9e5XVNR6nRQ+q
71iKEME4V6/+jeTngKL2FoYbDQR8dQg6v5Mj6ZXgB2D+GPKqL/8B5kVdQy+Nd6w9yHa3mRdCcNlz
DJX3wz+N52KzICqgNBqoHdvUoPan0u2A6EvK7BcZzzQ3G1Jxc2HNir74cSIBJ9uXc1B60G+nZHJj
aRFw3lNjWKTtMyHBxwtbGfehQox+4tK91yOVtPKtMeRjyX9XuhFIQI4lX++DLs1PQBS2L434Bk/I
s4++xSDlEiqe5HwjQ7Z8aXSZpA0ReQfqm8IvK8VHBYBZm7av1Kg2PAnvOk54ljQ3MKZxC3JD7Ben
wwqoMKoUpat9zbbdac1mAiut4akzu50W1ukXjQZViKBRTw0FjYSQzPr04MlK1FyWqynswMS1IRJ1
jOop90b+yj2HS5yt/N+8AnsMv8cCHiFmJ9h2HFAqDNIeueFfpsXPAZgPqt4q3VwH/w4KVJO4bWx2
4vu3ZVaFp+F/EKFC6cj+eJoaR2ezO55LXttn2G1FfWx4O0locKqfJNQssPMcZqux4XC0hOZ10c5d
QR86eRDtXJQapIM6/EMVU5VHA2NjnsH6HXtB3MkQcMsruEqJQE2No7EqwERhRu9RNaunmRah4sWf
iXe+ftdRokoJ3FnOSlBJp4SHGRUWvQ8jHr8u2FEFNW1ZCJDdorHEXR7Pl8eL4i7WEiAsISMPCA4G
p6up9CBmBWmffx6jXcp7km5wRJJNwI5fiIeB6zPLWo5I5lmFa6AwUwuUFUTCTiNI28saSjooBXH0
7zBOmGla3+B9/5Y8htVh4dFCPk+xTRt1+unNR5U//bTnjE9IaZ9oJ9IeSf+LVzIFEjQ0kEDmrd8u
s9tBFW4JfCZ6Ow14eppmYLoN/xNRWW6n3A7SioRGuVikKZLC/juPi/+vUZYAdh5u1NFaWAmb9NDa
t5h7N0xMTz/Z9C+vc9s9zXuxsmdD6DfoopFM6nwsmbIGX2LRN8oMffilpWXYC0E/cEjItKFCtFQb
DlvY8Ig0VJsO4Y1x2M9ajfc8wDgUXUBK1AucVbx4OJJACoa2WxOCDgiMm8BeZ2mB29eVaLe3ijYL
BKUSYT82OS6OYX2kEqLfRxGXAJC5Z9ytzHts12mFTx0ZKSGKeQhmobzOQMXIlp/kmiyR5tO7flW8
/KA0gpsv18GEn4h/RRflzA8/5aQm5VNNdEFwTMVKf7yIOjtqlM17rFwdpUC5gj9DpgyuTZsQTsci
tJIsWaHwplVBXlvfhmL6ilZGpAVKSruBZfX/34igBYAqOAdY3+PL6hInNnU/i9VCa8YtbfYMTH8y
TZYWD5nG7aemU4WW5H0soRiRdGZDFUW0ae14B2aEuyGqdDyzwnvzljQ0WJT22fCLeGkfcH7dtdH/
28ZJSl+Uyfn6dJat016jtEMSnI1+VZXuC5lTLseVEzq7n8vrFjfViHjhJNgbplw2ScyJ7MKtrwV/
H2W+lAJDfH1llo1Y/KGnVG6tOsAELVPGFpBzzGX3boyR7868YPK+WXtjEsxyjZNbJ86boAbAXUPk
77KiPDYi4s3QhYkQKTEZukeGBpuJ4YjD68Zff/Mv7QgzjTDAjUXNnNFxKOwFxbeEAEYoGpWtZLQq
0XUYJK2qbrVr5qSZfYSAFo7xAu2pBCGWLP65rmIU6JnwiuoU+b9CB7XHTjgdSA4hrSPGOKW9LsSz
MuieckmjBxU/FYqd7sct3BHYhPMClM8ZwQBitlDGrW6X/5BPNSeMTDrRBW/cEDuqeQEYq+Wu5APv
NnBpw+LvZMHX9K+SLMDcQhayKocg7K43bAnZYnZ7BmzV6BHvrIk1nYWezPxxOOX2qahyFShOF5JP
GSBDf/2TyVL2HJFCww3GxRbvroWFt4xRUdk0z3IoTzum1KnYp25+WWIbfmxNavNWD++v2nGrvN6N
yVlln7JugriOlRh5xlGkJ7sMg/Ac/zsT+KQh5xji5KAO+pPirK/Hwyxii+7IEf9K7OWz8TZvKN0n
AFQwMIyIbz6EYpWJF8xIhRMJZqDixcM0iAhhfLxIb0qRVATKq4QK5bFZVB6n5EsrQaw9APFAF4Dm
IXyVkMBHZFesD2q4+8wNBNiXRdVf2gI/wBJcZb2631dqu5V6THHWSqqgWsKkN/K3mVxNxvH1ugm+
R3/hS90xl3F0IwDwaTmifn5tPIR6vVbl0x+GlvDfOo1gjLClsxBguFzIvEUmX+T2C+9ZfYvPzj1t
mUFv1Ns5BS4NAgp2oBnkMs/B7Rq63LcOfdMxUcc3TZ9skkDsCTh3h3gELNlSKBlltjl9ricbxyVM
Evh2SVTmSRUpykL8kbmgvjXtWdgxhtMj1X8FsuNGq3TsEPDC+ah1duUjBznAln2q5b37uIWq+6vh
JasKf6HXW1wJgUa0/XjhGwP1HV/YqyrUOy31QkaiASwHldmIsY13PBCtEiykH469rYvElHkXzOt3
9r6ZiJM2tCkHt2RruUQZNjYsLcim1WFeTBTGgNpclD7bKbZYS9znvWfQwVZMez+/pwV6DRElLaTn
KN9CkNyA19Z7Lm3cHg1Cy7hgU2A/pz3/4T1g3XAklODsxcOLTJpcP2GRcGW9gvKj8sDSmYT5X3yK
6KsdSpcmBsTXfJeg68jBbSk6lIaNJxaUc578JZATLLTGwtBVnPCtcBV3GBoaD+GEqlRBd2UbBAHs
/sWwVnD13XE/h718x1HEjG/8GIuZwjMQbQCPinO8LCVWNQuNYEdZVxFHj3+N14MOBFFRAFUBpIMV
5TwoJHUoZIs3P6OG9KmXILcJPBL2q0+V+LW5WZcR2XQJdJ+/mobXBqIXUnMswZK+2JX0slpt7sY8
SQHsmvexFXZH1OxK9NqA79IH6hxmYp2gMknWlARBISVmATORk1C+dT5buz55D56h8dSHAz3NMzxk
uDE6eJxR3CTCu8J9P6Gks+8xWxYQqPMqs86X0qRfiQ85XyWpxIt48SKGYz37Cgsy1W7LZW27hiaj
5N0m8MK/tLOdckiGD0Z92ranDuyKKpLF+s+n6F42EHGWbyi/w48i5PYRuDmBcS8c1dDiCE1YUxYT
YOGVfgAnlKcJzH7LqGzZBhCB4KUHcXTO8ORaedJy1434OIBUo34sBFXdxLRbsCRaLItMMg4yfi54
rR0REuMeqBlwpZqn7LdUrRUH9tbGXQFSOx40nKWxrL0QVGx7UkVhQsrXHZwwOFoBfCSrg2+tFYKM
Zg6dURiLfgohu2kOv2LmhaXBL3w9xHgc/BBwj/FnAlBLeMwb6hh11ablqsNU5SreuRwdGxwKAIDw
INLQaYL5rgF24lyk3cy1wq7K3u46RnNddCyYPBoTl0OzulG7fUVgv5Bx2PuTSlwM/1M0N9qxNpp6
R0QxeNhniSu1weuhvIn/QqeAc4N/uElU/fIjRaHARc6Xod57xJeMTXBSSopHU1kjm8eFUhxUS8ou
LMWa/Z6wfjJfHShkS07vU9q5dVNAW/ra5q5ePpHAk/xNzDb1WCA9/4rJzDYt29kgUXc1CkOeK2v5
mFXrRz7Pa3FfT36yAkCXI33DNfSNCDJowyY/rmeb0FmWtcoFJRXIID14r1ejO8dW1Z4zoG1Ia54D
XUlenQPCK3A8c2G073ce8bgsaz+ZWM/P8cx7ML1EeWA2733Bfaiizo1nYcrA49Q5vj/CRA8HxWEL
SOit7JncL3CvonYeoW4ImaiEqzRTya3kFiztymBISgDrdw8t8dTtsc/Pd/cMI2UYUQPljhJCcmJg
npnXnmL1AMmJxx5bv3Yp/VZh6Fd0/86HuzIFKs6P0IEstnu7/Q3ppZVpRm7h0awNLMFlABkiQSvp
3Cndmk5/PMeWrERQQHLiFLZqOF5w+bil9mfmC7Jc01pgtVbrYLICgA2cI8ngDCXc2lfNsGishP4H
6x97Va6SiGY7CGp7Psc2LmVaCjkvdHWX3vYlF0InXGhwqh/KW0ui6wCRqpZ4hfolQCr9CjXLUW2w
+CK54EjfxahMP7QDqClq3ZvsMJUHEV9YB0HvRfpge6uI7NZaQBfbsPMoZnEPSL0X1/adzw/DfQPi
w9pYLNH8HLe4tnYFdR4u4Y8J+8frfQIz/NCbrbSUSZCUgv8NFmANwgeuCEcML4Khwxo+95XeVxkI
aG/vQCLKqvPNv/6t3qU4jLOCLb6fC2HgoET9Er+kUVLVvUEpLb+4onI3OlwH1JA5JznChlPjKvlE
wvIDGdX1iFTOlBopYAk4a1dETIteOusFBwsziUMedoQuiaGEOlVTHJlMjdy0OkkpAdZrKCFDvzta
aJE0WIqF9IWK1Gr0/W2I6s1C2gN+xDHPwAKTqp4tEDwsAqT8AV3B6TavG7381xOHjfWqGvXKkEWB
LiVwUcvm6ideVgpHk5ccj31ZtLMKIWlh8Hy38xqHg5XyAoVOktbA90eh+zclmn+E0dYju65SnjCG
EOrXvYeugoGzC19DDqgdBAKzx3kGFcYydl/gKnOhqqKbHSmwgc2CveEf6+KV6TYI7y91pFsXRWVO
/NqvBfDkQMx7SqAp2OKhH6+wZkOjkPXWUQAqSyxMwV6nzIZBqCEU9RqE1Lb36pT/nYqxfjKTpuCm
9BKGq/uZnkuEV+2C4pOP+pfo4nctIZPXHFR/EzUWxKj8yBzkOuS3MUPZkhgBcT28RaUWhI1Xkwzs
2VUAb/OF2MNLiQbZXtxbbJCHCAgbOPZ2ll7+B0mwwuvGN5Y4QS9qSxDQc2tCzSWwb9QEQm5mVWQB
7tZ0S2Bbg2olQr1KaHn3lZ244AwfMYiLnQ81gOnN+ahuL++TEVD7juShFJIgtTe3VKBsU557yuUU
3Ak8vbVbjrzS5+OceZJNOKAjN+9CqdKsrYwiJwNY6VsXF1zF2LrLyFMEaUQrsc/gHxrr6JK39UwQ
GcXtyaV5nRroGa4KFZ88AWI+QZ07SBEAXADEjM5avB4zb96fvmrtRIWADmV4tWnLxONNZ0nSGxAo
ozo3dnRY2bQtlP9PJkbB8nT9FrHw6A+FnnqzmZL4041UtwaZLE6LFkuu043i2wYnM+WzYtbcZIOR
v/9nLXkOG7P464xzw5B/jyn1I3sWZ7QW2g2QxH2wZ4sxubJ+AFNJ9fDUnyoAFhklukEhrmYdOQ1I
35hSg4V1ps6i1ukLyYgeGlBj7dlJ5fULhVM+EC8S1u5ap8n2iMrg37rVlxrpXt+/3rw/aIhyWniS
O7QbEE5r5TwLZ0cUHTB7a03OUXdmkhmBOsqMwii5XU5VILv2y2yee5asCKXpUJLaaCqB3/iW0IiB
RQlalHHNnwbrXZEoNdXZwobn6S8U1tr6HU45KINd5fkUCMOVuppyBxRijm0zMck64TpC/RyE2HeX
PXAx5mrm1w2vvjOLleyfNuxNlSIY7oIleel07QSDUKLZP7ZNzT+kJDz8NKx+pgnZflCIw0KkSWq6
xxf5360wggEpQ4e5tjmSCQ4qc4KCjaYK1N7vqELKqHBlwu4HiTiouppuov0axDhmwtfbGqrRyjEf
ZP9UJYIA7M+6JQyhciW28HKg2C73QRM3UfiU3Vwra1qPbSlJVzJkmUTcg5ow9ZqNAoKMwqu2RBpL
uGJ1qGmPfzbU31PVdOtxi0aGQboemj7SYL6Ef1IWGQ9amVGIk9ebNLVWl+ZK6ylTNKzUS2aPnuRl
zGi2P/zizQtrvx125hQFUv7kGP1DRtRRpO/m6w1K3n+OtPsPt6iceFKti5II9NT8ZJbv0SY39a+l
ZSJqanqBQSeeR/G08ko4MIoNou7PpqvLoLY1KOn+X8DJP7JIaKYIHq9HlQCVjRUAQqrWNajppjua
u+mrvx86cUOVpuKbGC99HACTumfFfcnZ6klCMr2oK6dwUy7Ub92SKo7pL/EvjqkZQ4wMV6hwAB35
ttOlD6ODURGadnDP7aQPFghfN/L9aieODXWlJWM75UeSfKeocbEin4RjI4ZT4isv0rWI01r0dyp5
YSQMPoJXgJ2mwNaCfdJRfe/HSJnW+pnj+kRyTF/1ZCc2z90uftl8YMfFpYD7j+Fj9NRE4S9UUUFD
B92bGendanKICb0p0LeNuQIWZfrpCYzr3RgxlNU+MIYtU9US8JsuWQBM6hoWiGzPcqeScgmcBBQH
DrUiGreCrvan9b7NvaTYzrNq2wHYBuiwM+QBtZeSzMd+G27pRHGZwF1lfDoMGKfvQqjqpc0TzNHB
c2Li07Y/VA2xOsr1S1GkF5SGW2ovrAu/6lqpNSZLsH6OCIRhd1IhZrZo7CinYtYV51KV+8IWvHOh
O23i2+3eoQpbPJqmJ3hHCm9nPZGT6ulr7ZMGXqib3rDoPGAMbvx4OQTBuQ+O4qCAfCg54DDsUUPN
il4UrfK9E9wAXFSHlxUHZqNiz3gAareNW/wmfj4hCr0gFmEXc0WyrFvV5pzMTv0c8jtlgpvjK8CH
tIxGM8AkIJi+mUpcuiJexGtrYlnMkWQ3Hi6xxM6wo/FG9Om7/Vj+7GDMKh2+B47hST71e/2kkcM4
TqCfQsmUPmL9u3zzLWGvBSKiBHBC1lIsud7Sk7cK8q0crw8s+OnHDc17OFHFlzDs2N3o7dtHm2As
de9aY9J8yNyaJNB/HcQRTyx2HwkmF+W5m4YmAeCA6Lw888rLcW6dPLtxtovgwlzhRmvH+F286KFP
sqYzz780Nb+m4I3kcVQNIKOwqAW4GIyagfbnlZNINxX9MVUrxfcbwC+3YXsIx7im5eES33suyYrG
bzI/N2pgJGognD0UGnYz2BWT6Pmgj32F/Qs7+F2gUYGFQ+wAFCtO8xMXAkVeMOEEW2M/bU4P3npA
bRQHlTUDgMDUOp4kvLjzR3HzPX4IoTtSMAQRSkbt6BS+asX+PDpqZJ/uhiKYx+vdP14F7JEcg/HA
T/ZyMA5mUlEZAzQ6VOu9+Anl2/FVOOOUWMnsx4i336N9ItvYlKdePjkZwO4i+BLfZqbSnk+NCNpa
hrcEYssm35EkQ+F2X6GzjOTQkCP5Zxyq+g2VR3aRBl7UbXXRTStoJ2sEQUfr3HwO3WA4NazOwcyq
mqae2g2XTrJ+LDilRZCPe090XVCaVF2hFVGnM+N2j/g+7ilYw8WsQEIMYvadANOIf1NMglJWxBSn
9cDbGQ2zsSWz7+NyFbuVIYBDkJLnJ/22F3bjnpDHemNKtLrWp4bJQUwKNMMF4zcJto7BtsRrtPLY
UOda6WGV3t2p9t9krpjzQOrjmED0oNGOMXdLQqnGU5M6MMl7SXiShGZ/BBjDONgJFUMnIraVHcx2
DyOBaWKO/vynTXKKvKd6yhgpk5SPMQ3ytbeucXH6+C4PpLo+0Kjv1514haprAnoMbEQzSjiBTrrJ
pZDFDQp1/a4iFz2fMK8AmTxDh/wok4jkkZAkbl/uZYfH9y8eYFBy2qqFbRIWfpqnZ3cmNW2Ctj+6
wmNrohQBSm710pF5grE2ktuNEtZTpA8dkMSX+quGgZRcZXfHZT0QyA+d1wFxXp0H8vqPpgm6v2D2
OK5cW7o7KQ4TAQrrBZr6KqoS9I6hBXTwEd0EtiF/+rXWV5j6/LrGEfLkG6wunW//Zc8gGTKtCIvE
keTud2SwWDa4PFCxJk3+HWNtfm71QvbilZUIcTRwpoyfHsYztqZ98xYnYcBOxARAY41pwC0LisJo
/jXT1GjmEYTuUDHWp7zRn+w7DvEDp7sA2xaaIRxyEVuz5CCGw3bo9p3qj9BUhrcPBtFGLLk/UvFZ
XEdahhNw3T7rpv2TcZ0DdVHIwUPrqcRXc+jBzIU3CYWcUBWWtUz4E55ROaE0QK3PwEsvAz8nCs/A
G3JtRf9pgwS1x/OOijj0p0gOPZgl9oCxxNibbyqKhs105Hu1kqe532zsVqS/0381wAYFoKVjIw8L
xm9HwGo350b7p9A1E8gMaEleYiwlJjkByKJIYMzpCVGq81imRgz2lU2iKJ0TJcb3oXDqhspYuH7+
sZroK0sJfZ9btOLku/05zoEHqc0L9/pJgO8HzjXFyqE9L57+RJMoIjZBbML9pls+hnVKY2wKhrIS
FhLQnmeB7TdOC4x6JwRcXLWicKoU8dbAFFFzKL+rSpNlZl7X2vECbCqOdqbhxW6nFMMYEuhz6rjT
mTSPp6HAmfmDgSBLKp0VoPE6rGgX9x00HZ6UPc5pXMXsqjNfjZisl00vFgFWr01Are8S1kpNaQdz
voZBVvbob6Ooa2O9Ub4lzQyYn4FGrJfDT5z9hQ+K/tfC2Y1LK7THESkjrDepUMHHI9q0AxgJSyYL
vVpniPDX0Y+ggq57oRT3jM1cg2H4eocGsvEtOos1a30HYsa5yOD7GkF27wZlCgmPAVwjgolj4fTE
spS1a04xruadu9Esg7C8U8DdXxUDQwc5vNK5A9ihh5eXTkt416ViVfzw0rWVsFHJ0dfQ6FvdOcGK
nrIgSkUQVjzJ9JaOI5yS4bjE6MvKYXuWF8GdGI5GEKgAgXAa3U5flHVz/udr0ZL02SEeYkcp46yK
DKaXQWU8eUt2rl5eD5H4wyVxoL81tePJucL/K6r9M8e820h/SqgrdYmNI1uniAgrWi1F0+E4eIea
FTDLG2cyFLC97ect6HoAWOrjtzQPcvkz4y0EUX310WMvc4hIAEe9rq4IMtS8CjfGvfWxXWLDy8qA
qeZrIlKG4ImFsOCbHRT6OrRWDuS46QKKX2YwaNphCV2lm7Ay6ApSXcMjnBIW5oNFwiSo130TSXRD
ZH7ivr1LDkOlRPguHMolz3To081ElMeSQvs4levO/Ruum+Z+bhbV6UhZpmtyDp6+QyL4mrhrDqY7
vu21/XNfmzyYVzax9K2EzJ8lqLjuXwWsAZaHi7QC44ua5uHtLsrBDkHH8DYvxLYvuFDn3A4I3S7L
eLFiHJbge05fAYSkVYRKtfqkNJmysnOBzMMms1PXlkIeQm+V2LP337hZqK0VbIt1FMpjqcwnDqua
GkTdk7S/EglYHZ9hqAcEOm2L37pdtnAR03uakA4Q8cD4Rzzf7O9YtoJ9+6884Z3jB2dkfs/nZBNO
CvCu56z4Kt+ghnEdb80uqWExrCnkKBjEQZPoeQT5dWfW5iv4xlVMR5f+F2gHFq5jk4KNpKZbUbyg
iftO6JfWneSGe61uwWh2VyAGdy5Q99Kag4KwyyFnZ2HC7n/8q23S1nMhpgIUl6WZZ29elMn1xaE2
Q0JzkFp+Ub5ZIKR6/ywTY00OVIqMNGpThohoeKqx1H/coMNUCq9mHYleh36mhgkDwHuNwkU0Y8/5
ALZ4x6G5fsE+d3+s8QbgrPl5E4FYHSL56WpXmnUma6wI0q51UVfPG03gDspMkCqZqdVK/91IGxmg
LrvTFwFDCT4g7nQBvPNDfMzwgnvlRc3lgLIaQmP9BU5A2Msn5a/lBceR+HRPd6NQjC99k3zAocfq
w/X+RQJF2ar4bcBF9Zs3NixtKdX4NEto7PFtKCngl8IPgwF301ASku91YJEGgT9seQBafCaLpSd6
TMLtyxc4yfqki2MvuGqc+AW4dBFkdxQslCc+GyftNDFxuC2Gk9SkJlImsjp5BV4t8KmAmdxgkTs8
eACqeSx2aqluklqpNd3x4nR7vI4igE9oYpWnB2AHH/mV4NZLFFwEUsgRi3B+YTlQl1NxnqYiRWwP
FrXwzrBkPDvG15pLnrtb5qIYHEjFfnWGRauFzOE66jBOSYqRMCpC8QNJ6za1V7ck3lyLTF1oYYaU
Bm1USdOJyfk1haTNebLUggzd/7mvoHdkI236OsVexgD0crQZenjghx4qJH5N50YmDkOCnPD2BERO
/Oqq2eezCxByc9g0oqcwrvldsyd8UhkfikvSgfnkEmjd4fhEPcd6A/KTXW9Z/91te2Hd8E70j31y
+H7WELVongmPCerK8k+9aZu1cnsGEsAh2iyswj/oDc8bsHJ2BrvymqmTOT4puVZVh2ucsuOR6vx8
5AL2okhTz9tYpiYftunmlvsi+8r9AjYl7f9BdgSsyMMZYS+a4iZA77Ahms+pzj1lJsxcz5R+pZx9
XbUVYFFPUN9h5t+v8KALAIpQse3GAj39oQU4McTBvGz2cCukdE8N1+TApRw2FApbQkxbSlR6R/l1
PzoOryfHE2jbLjrCHVJwTUrqGyULey+q2KpCm/14NVZi9ni32XTweREvjNcX1MXjQdXGTqkuEXW4
GCkwh5DFgwretFpDA0PFN17XR2dkSQCMYlP4QuHVYeaJvClsenC0Oc0AsKE7iCJWDwJeQVExS/Nm
5pA+vsTaiH22E2nfkDTBaxN8F033OhRJXWcmzhlB1bPm/CCXcjG6nnGWAO92wB74NFSD/knm41fG
K6tljAmWSD7kb95wpoO2yv48GuUWhu3G9mm5LmM2eK6bf5VorJzjBvVt9eXwCoffSa4Upi1iVSnP
1fst64xoGMI+7RtkqF0ydJiVIAtRGNEroymFDRM1ivacYXWWAWUp6/j2zMFLSTTElZNdhhRkmXBx
Og9n0Aq460ZEVPcbpNQ6q1ORu2rRl+SWo4cR3dx1Efhv6JIu+kiruPyuu2XkXqBCg4Eck2fJvxD1
E25X9UPMYjTnQiKykdtWZnDGnl+hsyJs/F5L6ShFt4JcDbocNp9WA8CTEeZfcKeE3QiB61GDvWin
DYS2XU5ChQPBScHeHDGMq1NxNjVlbJBP3oGWdfgJMEOb9muMUTqjK4xEE9Z0CpTWI7Gxn005g/s2
9m5HQG+gLL+3IzwZWtt6YyNW9qDv9lWD8Rro1IeBcswBtftvYdrOKbv8zknsYXPy4X6waiBU6wYi
UpESMQkHUwqebMqs3FJlOU26I5K/dboJ0UD+HWnJExJ+pIqCK/DtodDO0vahujiBcKOU2JLCUz3g
5nShgKPwDMGUCwue985YVpfwrdtEEgtgFoBnKjrwhPAsETwSIDY5Ywzif2lyexciMJ0thOdAabGI
p/JO5VJ7ozFyqKTuowexZmTav2ssLz8IMfTrzUILl3FKSBn4BsKRWMm8qUyJcSjTMYztWqBQFWDg
qVVEX25vqwMWThaZJOLnerSGgmUx3ALGePOL9mdOVmbIVGxbsJE0kC/4T8hLn4L5hwk6JViK7UsR
T7aHzX9JHBHAQfnJWrNzDqWKg8n22mS5N+pGWs8CoiIyhFDLZ+SOLfW7Ztu7UGdK+VtJ6DbxhBbb
dWmmbPLm00HAO3bTJhjLs2Np15l72aXFFoOgyzdgdKE1ioCCobozc2zjzHXdCT7nayXxBEUZjJsN
iOc4uer6UbgZ7p2LxaC5jtaqJfeKm+wmMj/jDZm31QRhA5qXyYzFSScsWXGSl/tSsEvDPEBhDg6Y
HGJwVhQYD9LPX29c1D/e/Hiqx72bDUpWgB5GJuPzTETHA/MtqTTvRVLf2Z9MP0FT5iKUirQ3JmSC
WLifZpg6mmy2LTLS9HT0t6nAc4kqDcH4jkbutGPrrBphjq9HS0Ug48xYwCNn1iFKGLj2WkU+7e9u
rjOZKPxXyv+zlOOIVq927azlgC/waaiaa9pvH/QAKg1pvS2CSsJpgWHuyHO6f3l+2k5FkHblABYV
lI9d7X21wdOeFsZubIpAG1SW4DWWXrvMP5iuJf6W3qZNPrfqkcoHN1L9N3gSP0zisS/edZRp1CSg
w4qZ37sXQy337uBltG1D5C217za1xS13MZ2HHT+p5U97sYUxbon2KPtE+qW7FvMQ+sXWM3gwki3V
k7lAeXi4RJY+qtfNAnp4+RSJn+WeHJHJ7v9fuhH4+jstUpgJMZbD+xWFLsr2yXv/2wn23TD8aZN7
K/ZPgcOaIGQtEn7ql049d0d1pTPp2fKHhDkSL9C5A/32T45Ad2H6/1o6cizmsyflyn5lMUBuFuui
ZbQIHOXcQVaihm2iLGJGXJnsLywK3sKZd/IXt2Wom/6s5e7IPIu9/LhuK7HdYS+eVXgQQl+xoILR
wSO+8S9ysKqYYC96Zt0o7KONvOskHM5aiGjRZDBi03AccBdpWtFCV03CJTeFjCSAEsEVwLXTXSeB
5QelMBBfJQbVlhRYAkwKU5Yswr/jUQvrj/x/ykb5pMZdRm39wbk5W5EnfengcyrNKCH3r2q2x2J6
po9uYHS3+mBW0x8XL2bv8R105y6sXzj4Dw/UuSF2YbIhpERWK1R+fsfzPdEuC/y7fH6VW36Dmccl
DO3abcCw58raK4/wBK/qxeeNvhkjYNoEBgtjdSv12jufcpTHN7GTzNNljeWWiDDiZmCOeTRKXb+z
PeXKhyvjLV/1JZO19zC2p+h+fYhUOGUoZwUcY6EoqLKhdxHiuvNkXUBHUuXkderk7RjAO7sdin6S
b2+DPozwZf13grX5PS0Pivb2yZJlrf/cexkPQ3nIouguEvlcnvN1IBbjukOckLtdvWRQj88zlXUj
w6cATrPTzL1Mji5FqIYnr4NJmr7HIuxolLyJjLWO0tGovg8ePBI/ni5Dqcw5LsJQKY750ZhRMAQp
0lD73L9yUWyCfG7tHukfrbbevRNfpflaYSpVafblhhdrJZwbmMEKc2oz67EJ9IMHT4JWcuWqzjyg
P2lDKzNTb4lvKhUsqGYlFBBQqSxhslhzou5MiYE+6L1uwlIFDkplify8G6WoSHnAdXEmc4Feae1y
QadmluijcrAJgCx+nKzI64Yje9NV2c5zRmRHCN3LLHidtu36ltk22fdx2OiBolIwD0OdRNVN8rdf
HPdR814+UCOJnD6O+aV/TiMIXwQWPMqA9QxpSbuf6d3tq+UZZy0QFEx2q6ctnMFJDceIn7h16SDV
0FQI3saJdhr0qAph1Ez7fbdD8ArkA0nVNgDqIOHgTf0dclzF5FABBGvm5BbwLTW3jLWAKQ3+JsRN
iIcWr0kQK7OUXpg+2xEwHYvOIab5y+sz28AqhypGNMg6YT+cYHEVNE5/MP6MEpuA+g/ABol3zVov
tCCJCxjTsyalhzIukMHPdawbkFkjXgD84pAH4joruBTZX3qQKOoAgMXj9sNzj1QkRihNIP0LMKUd
xPptyx8zvl5lJnSeTHSBvQC8DYwSz9mrjPIrhVop7UznY9NgLt/2XkXd5JR2pU26AxwXMTEMsL4O
e2pt48NIieGzmnvR69js8nfDbuXFnYEycM+sBg5uN+gQEV3ztFziVvbo74ZYV0S8pKP5CRGDDpxv
dvtQSOPtlt+m39rcoSQo+VGTIOOdfUCH07SM96pWiF8lkWafJxCbguEeSj+l6OHh9WTsXz9BTLyo
bD72+seHpxWqkoaxoQJmRhUqo9vcoRJdTooqS38spRRVnc8gKaZU6zn6U6PUOih9FSVDTWqejq8h
42g33erOP7IaKGiE0d/ja4K8mwH03HgBWleVxMWf2hc1iWeLQXAwjnaK5pfGAAbP1xf3JXFtUD7W
ea0e5LzhuD+c/w2+LR1q5jP+SIqvzh1gyQ7zSmf8jxkqJ4+rNSc9HPluWrxe9FIsbnx143GMagTu
rKuGWkpTzbmae1tYDop7vCSo7pkveXQHtEu+qkfIkEcx8X4SBpQeC0sMbOjeiP/kqb78KTY/kQpt
7apqAOiycTmDNY5Ph0cb5DDHPm4T4ouyJXkekBJXFK0pkZ0Of4bzRupcxCGIVg7u1wAfi+F4Zc/D
gGka4ngCImNMDUM1BAHuXLp2NxnazR11rq6r365lcfPrbPwefg+8kB0DlE/mkJRvFLufw3Q8w15I
xma9Ylv9wEe5wAnGRwh0shawh8SSEkjzKAAGJOOr6LrtJ4nXS7VA0V8NNjU3j1koAe1ZvHninEIT
W9mbJcGc+wxtSSCOvbUpQ2HyVJWll5G6inJQDkaf5076wsRNJh9Gy788FR5MIyRmDnw7h8WyDVzh
fB/Ghy0kPkw4NQ2u8ReECewAXaEKIwdGPIbyM2I9gQfIwEBJlfViStcdlGckmEKjxo9udYfMrCvj
oNJOAwbqCxyPHzHk+N5dpWRE9CVm3M5o4RrPgRB9TS6GU9u78aS8xvJQhtn6CXyjUhAYeLir5Ja+
2kwbQxHwkP/dHh9Iq5Zcejox98eb80lpZRJ/jEL5gG/9VbWHwKCbQCjqaUdjd08DM0rH44B1/zU6
cdsWcTEn5eUwvohYbi+siP0BK5KBBn9xaAauJG6jVD1I8kC55erCh7RIvnfmc5yEreY9QSLMJUSD
S/rAGbJpqhWD4pqaY1L+SIv5nj4ZBil8hHNjOdwQLlivGmzj4O9WqHkifYO92QoRVxsHUFNB5dsE
r4lwF9elwEAWrlZv21utRZQK6/8LQEIxHbR4k1PQ1gEitODk5o0ZvNJlB/stqjF7cZudmAU+bhPo
1O2jGLin6ofU6O6CseyGCjUU1SH3f6tCVGPUAdZUyqIqMpSuee/ekJBfq8DyRE9Fj8y718sv1BtL
o8v1Vos0y2+zlq1SlxSzHFGBoDd3AxcGXSnWkOGuztb9VRR+2uhYBTwzdSF2VrQhinWmDJethCS3
FlgSy3drdS+f4ySV7KYmlma8BdeiDZbgWgek4faoF/2PWtnL1F/1qDE51io6tc9XTvMghrakKHg7
FlN7UKxhHUFv3YupKwtG1G+q4B0WSLXms3u8PgcFBl5WleXYtHB9E8QDMCLJqVdrJMderKGwZyfE
CRVMHiNV7Th5Ch+C9szDhCFUZXZTWpUn/kVw+9vTQijNZdEJ0tysMgZ8TfbPMw4s4WsxUnYHKLS1
tBqzEuZxZjP/jCxtk4NNRlyWnJcWaO9y1AqoZPKZC/yHyMHvTsHvQtHU9Y9tAEgvBy6kTMEccaSr
kwVh60/+NPuW2bwno9VzBJwEL3iU1lMW+2hXwCU9xXVvMjVKCfsITWRnGRG/WniWW3Kl2gf/URdY
C89apO20H0Z20wDw5Vnj+zgwYp2VWqQDASVEhVn9fqIP1wklKojos+wA+3h0T+5HhyOu20OgSfkh
cTQHyabygaUyQUnarUhCY8yPrbICl7uY/u5f3dIciDT9ik3pdLhLCbXMROimKZMkwkrwxbu39utw
t5nkQx6BsWKn6q7hd4EADVzSd3T1+6/Xenvh6S/9ZGlu6o4ldl4kqlN/LSp/KG21bsDx2Qj8FeA6
xnG6hJWGj/miL1cWP/ijAKhYCrn9NZz2J7QJnipkvDd3RMoZYjJ/mxWknpH1M+XU62jDZI91T6vp
r+QY6s85R1YMIrA/qCNe/MBTJmjcd5lJ/k/Mf2DRCVHmmMCatMXq5vNandyGOPa74TOzqQIxviaV
iHkr8kt4blH5x7ZcEU0KU+yrK5eF7hg8ewWkyuWoyOJ35+VbXeoXnMHu8xSWbINPkDPTfwbmyPNF
KZkvsC+WQB0VZ5+c1Rt1GKuTUe0Eub15LzHXmx0JmRzPbH6FBUmIbf1TIMZdW7jRXa3Tm4hqzfK2
Sg35HCxuL74+LSrqAtk7jkn47Bjid68az82dS/cITtYRjDd/mJNkwBvFcO224gzpocgFAM6ZKgqa
ymh+PpW1dP5Y+fE01QMVLV75CVLSCbdGmas3kmcwGnGlb7FNM6EKOOIw2Wl/Jj9gU9vw5nP2W9NH
1EPZ9TMgHeqLqZze7gabCnuBwjTJLfXVldQf4vgBRb/B1QTl8B0f3U/DPEgKWcV66U2HNLyLhnBg
alUgBmOBarvHgOYP3EOb/U5ay1fLz6doUIAUYQ9R5FuHNeCP1rwfNSgPOBTPw9JgI1EVSadnsfFD
r7bDa6fmwZhd3Ts3ScC1wzYRourYfCvC1f8yVmy+IXmvf6yBtMcmH8MsF0PVfpPwSLLKk2N5vEDH
ZMjjzuZnsBMGqBa5QarKEDIm4mXKf81HuPJxW3jR8sOyzgkeVsh1ssTFTCdxjss0sVovVMj8U542
twhVeblH/epaiyL0LUfwZg5c/tp5BwP1Dg+EF+wAUHD9rZ7cG6fY49e1DpKI51Nukwte7HmQiTcA
GBcySFznVNIENpJqw/pZeHDrI0Osc7ieDBov0SSfA4Ch62DVm+UK7tVeTMt9EYb6lHa6KCv7lvW0
wnZzkh1sm1ycIfgdLwzwrLf+b0WDKV3uy0EYVGmWQKTyIsPnR2hRUL5yGvZ9LAZeavhPaTJPgBmq
39yRUNfIkwnhBD9hE03hIz4QdSbKsmSIplnRRlJj+CczLCEMxON2eS5++BV6h6VGYe69asJjqBDJ
qJq5Llsi3ryl7vZPnTR1gQIkfbW1CpQZa6z3LQVMrMAvpCXdXjFP2PXp2uqqhflEu72Om2fgf8Bz
6XdOyr9lHzQNoSIkRBA22bMNmAuAQDTfEozWc2AsTxrZEI/xrIP85dRGAaP20buMNhnAWmsqMtTH
4yIjLi4mSACx13y6DcnQGOoktUyA7ioC68K1z1kwp2Uq+1EO0u+XB4QL15No8vPIG8R5Z6ckZcF6
G0BoAKUDFZ8LIrnr/wmhxytOozMAG6r1gQCe2PVvvEoeg1cXZtCx+2N8Y9bo4Uevbqr46IL96QVD
YohbTMx1PNtoK0t/gGplORdFLJBa3DUvXqVecgmEUAWQgT3GVTqv+ZXrC27P7fjmhzv64n+nj/aA
JEU7WXllqIWMtO4TUUK+ZNCAmRUl97y3wJXpLxNMO5W9Tc3kl1sZly00SvsitCogfhqlcesLarrW
OPtJpyfODLwQCVV8MCq8WjYP3LUARTKJu9cJWZiILmiuASk09wiJwYQCJT5xpVVWiftWA2a7H/3l
i9esJM5TTV05Q1QYkXVd/8FKebrMHmJNuc5i+By65Bc6WOJg07HyrEGjifSR/GjC+4mMUdTsiwXL
G8s91HWYW9dH7UK9uBF43Aj/P+1CTzR/cCPNi6Kr55YkxJ5jR+re9guIii9K43MDloLuEpY+xxaQ
9A7NTIStgdEDl4Rk1zNLDGB3OejabuIhL1GeK+aS2hGybUWPIiTDcoYR6Nfx0lL59rybgrBKFjX2
avSnR2EKYWmQYpD6pqFm0Snic4ccjkYsQtdbAu7wlY4CGb3hL+mcAB6LF9iJuxdAd5MqRk2+7H31
MB+tVyTWbelVaAo/XHYaMwE/haXKQOWxSbHubNMGwJRiXQlbcpM3p/nf9VQD4MlEBf+gp+F8eO1H
3Jrphlvsmec9PWd4YnkFda6/J4m7jlPqd+p/UO9rHIUcuJ1/BMA7/mMpI3To85bRwVR+4vy14PKB
E9VstnU8D6/i9sIPAVQJsXuVY6dPhpTWEPPEBR8yQrA18NKYJkPOsHKGLI0ZwlWFZPSUpzVKR7XM
vQoOhctr5B1bm3Mj8XSTaWCcNYJJKLrnlapPOPvr37cxexgDe3LqcwWocAP8q6/1s5y2nWjaKCES
8CVKmAYPw05Gmwu0hjzq3iNZX+6A2quL7vejfZ2GXtvjdsmQ200U0yli8fzuCKHbw2fegWoCl+mk
A1Gf5Z3EeOkwWWsn0X/9rB8jDgXcahKnTpulZtK9QEMQWf4EIDnLQ9j4hGMSh3HRDXBT3izbOIIk
dAOCZkx/LjT2pnOADRJv5vnYvcZ+xdh2AUUKLsrWJRl0+7maLrQ86Y0qJ+JuJF/Ydrb/Lw1SwWI7
om4MnwzihH63C+z5NfHatBisnlCycOkAR3JIJmAmb7vcMK2dfb/Jr/9vrdSA4Nu0pntMHif6gzTL
95bILTBox4n70rqr71TsWnfjJcr4O4dqRTmA1nW3v94912nKK2SYnWwEIETdSbX7VE9secJQ/7nq
6K07+f8qW6acPSIGCc1TbGt+Ike6ADiSv6yOcUwVIXH+2W2pCR9sLFwuvWx1gHkVny+aQkpFGdYh
gJMpZaI6VHWuCEZLmmlhek4n7jSP+Ptq5cyIcR90YkdcQsbf5a6H+5BvvcwVNMwphTuMrU6WVEe+
mn6Z0PnZUF0YOrz8CUWXL9vj6YQdv+OnE5jlXNAIiHgF5VL40EQahpPFKXnGesqi2pGis1/de1+E
HhpKRlQfE8XWdzf/3RfHi3DJYj3e2igTPii73es6vPbyFjIfcUIIuA57RUcKIuYZUDQmdEhqnT0V
m3r4LooNOxnE05BtWed1SooPzW3LfrAAN5nuZjoFUnbFAysZw7kdmOyTbw3MmF+TxP9IksDzQHGg
0r0QapNwy7FT71InXfMpGOrihAdPmh0e9l5g4iaZHskJZlzzbcZBndG5bT2n+CUbMU4+x0zSIgyX
gRSu+gs7faZpsIzUWplrj1pGlfamg1BoxGJZEmvK8x+kdoAFr2I8arXYRcgCHa6InmeFkp41kOhC
K/igDQrkJqsaULQX9lIaq0DU1gMdqzOhQikLE5w/sr8dBb0VXP8PlH0G7AD2PTzrkGATQ4mtpfdA
6ZtnmtY+a3nj+t5IrKzOkkVtMS7wBvzSshlBWDxSVA4AdzKKesZPqsNMxk2K5h8A4C9IojYBPQY3
+0nqLfzXjGJ9qn9PMO1k45aAxEVnvhpMhFGwlkCdBTqb+Vs477Qsa4pkKAzpvrMvpdgIqdZppYv/
DzZXfCzbCYJIARjE6pX9FZH2XEon2wPeVMGpV5ESTqBLY78FqwvWdJ2FqfKmuDT1zFnxs2VDWmQH
muYqy5LZ58k1nMWkvychEHpIRZ/lNVlIG8yMS6b7Sat+Sga8J+t6wWa3JEvkDIbOOtFA22OEHsZf
zhHjhIN5nD7YvwPhvieagHyn8A4s+xkxAsUfQ1yHLlM26SJne29Sr5bTbq6y8AHkoZt17fqiyBZz
ikNn7c0Q+39k9/dKBITrzalSIvC0BVLAs/CgM0pGFgk/kxH3oz14wdGtXeBzfO2xQWvGbeZPUyzL
ZRlclXejnjv6yAwx+wSDNASZB2lvv9DtxvZXKzETBJINObMGvNQmJaCa6MBwJ8+lR9vdyEdTFGf0
Cp1yE7Tjde6LuhhkK84+CPjnGvQ1PE2CNt1qCryr1j95TZNOpkMrAuQJfJjTuHezWfmCUqwa4Pbx
V6kQ+wVI/b7tgtWG5zKGRqp0Y53YkPuk97/AcmV92v799rV7iaSWXUNOJ+pbf+Me6nh1gKJBP/fC
AysX0VkQCFqQj7Vf7EeNUw1yrE2hiqJ+nG4dSZWYZcED6VMomanYdY0mP68ZWlajJV7E9qhoBjn7
ZdfOR+vK5rdb2wJURnWJ/xmbqMuC8s/7s59/I1tupiCreWX3eQ1BTklLuthk5xUvJ2xu+vb2rlAd
vX+hBqgxsU+g47NWaomQmpMAG5mbfbPnlsUUM1IaS7liOUnyKW/y+ODal1GCoEhBMBuPcmnWE2PO
N+EznlGGDxgVh6CtXC/LkKeRA6evEnAefu1ZoaAQ8owk0kgMSaCVAWJ7ToIUbDuEkwYHe1WtvjuU
hQfn/3Fqn+0l+MJ9iLET6YDjxbnZW6AH5Cka6BioWDTXGEuUw4OMrWOzriOFNKAZ39pWlIz4rDfu
OkejIOQf9qWRFdsLz6YUdtxGo5XFZxQO/wezBh94kbCLr2KPYMGi3qStkdLhZTkY6waXPjMF4kEK
QFcQLxyNaiw76wZfHjVi/sB3efeiPCeSfiAtm1JH6oMDx4rY7ljYShzWlc4hVgt3UlYyEmrjePOB
sp7V3XJydxSGM3VeC78UjsQ0HTUVYAj6jKoNK8CcmdAgRiHwyShlmrFFehSMWJ8LDPdCi4jz2gZf
E2Z4RVe5n1N6sgvu1RlSd3YXNtc07Gwxp1GSqcySndR+cGvkO5Ph0Le9QMugQhv7/u3G9ubnz3m0
8eMGn/ql4Y8BTADxyKDnT13dqm3nOfvAUdslJxu1oh6bZigHALt+pP9z1JgWjfFzZ5+5FByG5bCo
NSdNOIG4+QDvYBN7ToEx4UlRNOxmCQ5AFNr4fB1ooK3vK6/Quadtm+fwgeqGK5BQtKx6OS6G3FgS
vQbSuip5JHLehRG6SfZsVO37PREqvQp5BmTXFko+wng7vJE3fpyI6qEca+klY4RRwwOmrTnabwPy
tGvl6WHhz8yNoIA6hQDq3/ACaE0f2G1jchLG8FSGs1eajwelDPM2bescXaDI+I5tdZmILsR839Kt
kzVAi93LEH3fo1g6FtSir4zYxa+FlWP+sSOOWrDOTsfRG4nP0o4sqzsJFdPG9cGLeYRiKc/aKdYj
OHRbBOd1qVtlxeDqSaHbJmbZKqed9o/e9e85cvp7G7LRzXkpWKkAueFDSzP0G1AXGqrPWO5qYodQ
GUX1NbMFsuv53Ldy4OfwvgH5KJlMODJlwrP86G6eBkWAwj39p238FSvp3Sm84mETuAzJyLmrU2vc
FlKf17EIit7M6TGVKWK+zWeD4hU5FMA/fJ02kno/15VQLmDS3pcfOf6CFuF/IJDypH07RuZj/Dl4
xfwLoCCxvQGQFZRBOPpf74f8Mkrc8mUON6SEVx8/LT3uz1hDHmRrYpQ+AdIopLGrZdJr8wlDVCtY
2jmyETlgJLOIqcZGPvDLjeJGaPfMVhBgj5XWiPBfEiBS8fVpOGxSt8sT2i1LYgSVfdNNyHx61KqY
r2BghedLcbHfW4XJIh+1rZpuGvTHAoq/1wfGGRQZ56dxXIV0Tp2gwK1ilTeAEFyhSIdwq4bYKjpY
HZBAZH3oaWb/VJrlWifNTE/H7SlOt1AokjnzeNI5uxcILtkVhYszqeT6QalS5lhBXFIE+OV7y5F2
cK0nSKj7yqnGyVWbmML5wTXK0Knxg3iwwh4mB1lBKQ9oCFcY6XOR47aieI4Kmrc/rRG5MJZjuoZh
2W3lXf2xq3Hyd/5NRnwYsiNwkpj2gSaQVOfXPcqTWzbp3I8BObtla1zfFjBopP4Qe7mU/etYexli
yWMurN0x/6AincqLjixRnP6/sjXCTUMKd+KrmHMnMCI3w+f2PyRU0yIu3Dpx/zqB9BJxbDJCeL2P
M5LMkm17dM+8csIgXwkIJ9IgYqZo+V6bRGlwHmVtdP/N8B/EiaX/Z8CpnLZeuAOb2Nb4t45wkrZr
rcKDw93YW+cXFqHwxRYRmkl1P3HOZz+iqGYvy01q8QMYcWZrGVH/S1Shybqah3KUOclRKgjxNZ7h
bc2OI3BJyctu49IHd7nMBnt2BFVVR7uF5tQwabi3YVleBtvGjdQ2MypKFM6Ix+bRt3R2/hWXSJAB
ByGO3tcz7l+Es1bQPeB6lx+fmUfoxR2wMdujSQe4NpD+WPjR+tdv200XKApG+KRB60c73wLh+1uG
1WMKEFd1lc5DIGHu9G/A6cOdxHqGy58JNb8fcjIj1kUtNS3vv1zDUpyqoPuSCxIeTKvZnh09arju
r97C23dtlVNMC/bBvob5LszidIlXiGHQykdpI8PS8FA/MkgRWTbaiHFuLRW0tdnSQ9kc1grDDo7X
4jht4nfY5khHrIa5tQtdDU+WlKS2/6kvx3v4vdGOoSDkTdxx5Yt1z+kiN4KsnA03mmtF3a88Ls6A
1N2t5zieyx3+yt0sOKB/boc2/CMAefGfG2jlxksFiBL5qSRDGhhFcjLWllaIA7QknhwG/ivwbYAC
eEYUoT16fb7rPaCLHdP3LQ31pVVs6uI81YkI6spK9dgBZNCGdskFZrn5U82xMV/GRSY3cqiXSX0j
sT/aa8KqbsHYPJRXUm5z7ijgG6+o+WzEl/xR8T5X5QEljLFSr5BKAeBdc+nxrM7/mQHQe2i8RWvx
NEkWaPN7QyUV6jSundVNjYCOHkb/KER5xHPxf7FpNbqusZQWBYvYj8hNRHW1XprM7negOT5readF
Ud8q2jb7lz7ntrCKKLhqzMOjbV8ObCdIyt6CGTWi0E4InDoW5HXLzgPdS4jmlzpnzvdxMbCQKyDa
jiYK0tkmmuwYZIGBuRMvCTTXHVPFUCZvX+cXA6mdhHp0zjVQvIvA/3iRtJpPFC+TiNKADU9akbre
ZLF9bbwICkL+OChnuTltolkA7RUPxfZgsyL26hOw4gUiDztCLnJukPj0ID8omMbA77ihY9a6QkW8
tNRKV6tgF+zIucanuhkgxhNwG5yPmjYRYLU30OfAr+qkvn1u5OXzbn+TXEvCLDLoJ7uxjnS9Gexn
vLz7Z3UDxOfKgFXNoYX3gE4jj++qFH5xFcRPdreaJP8oYO5vWYM2UnGmet/1+VDk3s3O96Ph0FUr
twnxuQr+V6KiMgkUiG65I8VNVj3QThRa9uTbkWpd1OUB8bFFE3ScPFYtI8nNhPmkm4pvoKkRBJ9v
95wGSaXhn0rhgQyRsUx/oVpNxhDleKO6ibsIZXGCa4P//Bnxbg40mUJUkSJzKQ9ZDxZejD1NT/O3
h/MkGjllarfvDDrNX3RG4X2ie+FPE6SHE2vExKbl98UR8yVwC4yfmxbIaWN4PgnXDPSOOJ1CyqBP
T0D+x07AzrwQ++jK9vftXRGoKY3Bm27ihrDdG0oHOemWM/6NaAYRZxK5LTvAZ5fn6oyLwb1Fel+F
kA2rDbIviJcBBPejQQkrlMXtW3B39XUF+9dqzSvgi4hRRstV/BLMoMbSirncdLqCZmR+eFgskBzA
fx+v6txTycXpa+c4dDY/rGOP/3h3VIRmDviSNvvF9RX7iMClqtVNIi1fnoExlwV/nXtAHTQucAXV
GMmPvPQvMfuSx1a2HheGh0VcBDeWsxKdIlml0KT+tp0JJBXJE37nti/xuiNs6vGlNyE3m8V5feby
o9lGQws6McEaKmP2V5/wQKUHp/yWKFtRFntMstCH1o1gyVkU2mgF7ME4gV2zwfJLIFwPzDiSTmX1
3flTrKZB0yu2DpEiPB8qXtzk7ar4cvd+iZ+UXssZ0MJhBSnhBNChMQ8kJFEk/SDikS1FR+ywS9/p
1+eqFG6s7RogR0dK+L+mnKu0agkwQAa0PkD8hivBGSw5HOt7l7cE0emINu1JW6xKl0ER2m/IgprF
5/hrnnv0+xAk/qJjcHBkyU07ZZykk1J/HuPYZvbS52wMY0iAFOZgpSYvbYX64LfxkRiK3ols6BHo
V5OlCHtY7kAZusKdOsYlEYi6Ce8B+UVaaKi/m7XxprcswcUvqBPs9nhfmenTx/9yAmPvHT5XcQz4
ML3ccRuGGFTme5mQxiOrumQy5ks9DOHe+JRnIKsZrqfzDCzfhv11vnPJssRImoGKVl7DoyhBpJQQ
vwYMxYVrCjwxAw/QBUfiyaKIfOOnty9+Y9Cbz6hL2WcwWGBI3ZQvPWtRpqaAI3YtwwPnm5FGTNAh
2dZEooEqpDChPXk+H1w8z4Lhz04ueiOj2Czv3E9y/B7p/dQrbmFTBySgr+d5mDcdhXMolc4gfwvu
szJRxS7lYq/gFiWGMMHyR9AVXkvjKVxbXcDtuZMFse2Ot2fsEKFqyFV1j1at3b5PVFAPrnykp179
SrQwzvpYjDRiky39527rKD5KMdg+bC0TpFMadi2mN01CHrU6u1l3zoI0oEIt+0g/Kxw1Dmc/vfLf
wQolrsn9KeuyAXmeGJsniAdhoCWXT5k299YX5CUhBTTmyJFj7Y1V+4HpiJw3oMhcilGAmOPsbNpp
eCTtuIP+Sp/Woy1ZS7BKYokSmLS1SrneGuHZzxY+THsRiqUATLWrC7LPQ64EtuiCE48Zst4lORT7
00/kvVHS9wCbkcdeo7cCMx8PNCXugtDMzCJeuh0+mz428e1r8E0bS90YW97oW5GH54SejSBQdk3P
WuIMWlJhWizZKFKTwt0Rdb8wGWjmecrFbdR07aZHwxnVNoPDPyTDXsgh4SQzhese5ECPvD0w8k59
z5fZnsWF0p7zI/kDfacCNF0yFr3BqU4Zg+m/oDgwDm0oAGFFqeCxTnqMa9Q15cXIM/ylnPP6J4I6
UJmN4oyYUOSe9RekufErqF+5bKSExYitdQITzTVsxK5WZ3QjxiCKoOLOCKtNMLk9xeUzeZt4vZuT
M2VtrFktel61jJ7euEerrfXAII8WpN72uy6LXUn07TcHBrY+Y4ah60J/50njh/9eZAAgTw+MOd8N
gUqDpQMKJG/XKcw/vXMZODMK0ElBD/6ptv6yP+Mb4x0aCFDuGrpYXmzBTHm9O2VQDRR+Rct4lacN
d0e/QjlB7l2F3uNzg3pXelwcAhTYMXZAbg4hjZwR2u2ZnaVG5hxA92FbozVlaxIRFnGMfXyUHvXn
vPzkvA75HaV7+I2kSpJ/b0L1gOV8KjWfPmawXCcHPjo5W7ct4ZXUDIkdhX7+OcgON8lcm7AtCkRP
44GRcQqOxFCIMUa2kvt8u1BVZcfN/10t9fxRcB7Q0KVMHN1+XEuK6Shlly37R8dNswrpnmT8W+OW
12sZxdFcAJJHzwiGW6oZMv2i3LI3tRQ574c/WNv25qotyS/480b9F2zje0Dvp788WBLQDrXVqDRt
Mi2ds1XnHRyul5F0yIkE0tVaq/i5Z4YjU3sjUCfthGfeXipRteq5+iSH/hELsPPDl9tww9r/3/sL
2uAeBU2PSFBf+OlcWOgL4kW7+gno51Zg/A068oRH1VXOfuzTcUg7C/FanW8BVxPz6Z+Wi9WgO7Ih
ZzJCeJRwi90UWHUGHnSJ0xK5KjceB+8mTV8S4pUROPBXqFNGcNu9hw23g32lGSuh2iHhMJBy0u7a
iqmxEpNeWUnbkPUzsq1HYIOw3QnimSYQkUjOu7FFCBRgb3PbdEE3UKJo1un0lh4DUaKk+erV7szs
vXvu4MbIItrKwJqe7rQrfoua1PGDv9gDN4GUslyLaEvxpHemVPtt32Cve9tmaNvxpBr5w81qwjUE
BdVtDG5uERi9SvqRW54cfBuIyJ90NYJ7n1Y+vYcxR837KSN0cJeGbR9D+zZlvI8HqgF9a0kNU7Uw
HGrSjQ3UY2QKBhM6w8CTCFXeWhUU739Mmmf2E9Bq5LiWBNGZUuVclFCHFxeXLHO8RnzgC2c1qq5H
ze0UMkj4FDJfQAY0GLvIA/1AKipFgVfbza+cDYq6erY9YrHdYgEONxq0egDexr2kmbS7vhvrErO3
sdXoAyDJU88nTLWonjkYmFWj4J3Hhy/V3OICUupQdukLL5Jzg/wDYbe3dguF0FQInoyuq9EyzrXv
73TD/pEcdu5ShwyEbXrqIC8zpJKr+0t5eJpT5ycg6RP3IFCiKrtpkDEGonDYk+oEOGBmT+9F62qq
e2j0DjOJopUTbziwE9YUu5RRBVvMahr1DeerU4cBQI4idnPvnxSxGIjaW+uCghoRimFtdoveHIrX
Pf135HN/reGWpbUM9GcxdRPO896toURHvsyWwPNIOEApFHrJBSlN7oJ5n0WgDbZye/deUj9iGwvd
+93iRlSerKiYMgn12pZS68Tgu0FAzQ30bLi2vKhliPcoUzGGdu7GDnuqI79ietMTVi+ulk9EEjwp
OhTSAcfjIva4tJMWR1XQ4R+eiYxutVQG08s+nT9CVqvagY8hLg8zNAJMfSD+tC3I/UEUZzmBJNz4
snvacC0VFaj/2zlxfuKQU/Ea3zSsKWNGhBTCRYo6SXTuurpsxRzf748d1/Jc2mopxAGrrfBPMR8/
ESlKxf72ZYoRqMVS8EocFfvPDHo7Rvt9DjDgFU+TEyGz6xbgpYTC7fUAsmG3WL28E04E3SWKuKjY
LHRQz40oYvDoKTS0qpifq1ITzn3XdFvIXLE4fG0P6hT13G1YyCWKtvxYl9y/0lwsHvkj89CqlQZN
EbvZFxNNfmXF7zGjQ9KfZEQJRrRfZAPD6bk2Gx0xDHPXHx/P4mDGzHs3i0hzrxO94mRX3pGcRZ0V
aN3geW8mJcUdLNrqcRIgJqSmU13n7wHfKjewh+zjxomAZ7DSTo8rAqQKczozC8wswutV082Kzvjk
AVWg0k+tddCSveCQxeB0TxWiDFAxFgRSFvWk+vxalxZtJMZXoeENSjJHiAo0jZ37w/PsJvb2ZKkC
PG6Z+n883u8kRU5cjvm2ibSU2x1hY4JnzJOWxf1Ym4S32UaBu0s5kscMXSXJnQW/I+r/g5rADcz+
YfESMnR1HqccqZ9Fb09TFVa/SBlGuNgeV6hwcK+1pTVBcyGlP6c/VEXU0gRiJR5TiamMiOZNyRkb
bqiiiGEzNmxWJRT3OFuyKMBAXc17rvb+vUz5sqCp/psLKWR1p6U4271uxhtBno8YYZwZeRyuoCN5
WcPRoGtnh544mitK9L+PPmAeIAVTfn/b8MMMEmknznfAffmE9lVlF9F48K/ByZy6rb5r0DdHsAXp
oFnYWduT74gdIAutgIBFg0ylZfjv+aAmGhMAsDszHj0awkvnc30IhSiLYIMPIWRJoEWFH4/fbvVT
TUiA6rBrChaRSA13fpxQmJFeJGat6fqqLF4A420jeYmBIW1cE91MLd7v84D4JLUsGsN2XITp12gc
OHXYQsNvEruLpjkZqgDyhP47cYKdYAa9boUC46krARgr2824liaD++CP+25lDW3vboFPGG0p1wpP
ktTb526tLZ5Dr9KA05Y3HmDA2AeunQQKrBoujUpOs6HdJ1eYNMoJugKFuFNV5Svtbn2ghCTC1vFB
ay+GY/PrqNlZ6vUPGR0xla/bjsjbl4KcaKKiJ6AUyUZ+cwqVVTxGF/4rnsGBlQJYfbRrBjgOk9oC
cQspx4msvdfIuLj45DZhrWxK19RhhsYaQAj4DBa0qMl+7NgLuMu4HDb8rUJstbaOLmwgGKWxwYdp
XrS0elSnG4QLGldZw0GEqPl4GO8VeUGms/qnySGYM3MNJvaz5vPMbNtVpVo6Hquoi7v11R8QRkhV
aw+ZPkCD0V6xR7HSasfOunKYVJ6j/WjxtcSiWntBmKV9biy0RLTHFVxDNzo6S4aeNVPojtUHLAaK
/WxqbJzPasyqGct2E9UR/kdAO9JV7M1jQm2LBrsOPitCqkN8fYUKGWo3LHeys9XkI602GvVgyIA7
QpTpW7KpLA9eKziHzyNdAUoP2Kj3DfU4sXbcMhVuid1rF6yVvAZjL00l0jIt1ds/gKRhKG1cczOc
MJPa39MUhMVMdfoykDs1cB7bBeqObTVujTd71dfmZa4HZxeUVfMuJEKRmQv2/ginuh7mNF33r1nQ
YJuIJwHGNoxysnPuaDb5oWV+VuUEmPD7kRb2z3Q0+SzhcVmqPwxTk6CJly5qkhEcBEqj+LKoPk1/
ifyFDkNgPHpEIpchSijH/IDvu1W5IpJUijAutPVV4TOtjigYSwo0QkJRhBbefBcMi2RTYtELCQPd
p+nU5kOi69uGvLJppFpWmX7jF+kUWeGXn2iFqAIR+OIdf/TNmFkLHKsbKi4nLKPoZafeSLs9D/Tm
orqmeQoz53J1f5mUt6I2QkHnFVVtVqGuE7j6eAc7r0tdBSCte4p1RlaJxkKaomE3JVGV21DeoOWM
1eFYyj1yJ0ZnVizqGXIhGGEh0jBagW5b+HbgonGvg/Opmrd6T1RH/RNW9v0gzjBnOt64ikGG/3O+
rAEqZD1HR5pLCX00IlBiK+vugU0FpK7hFl42MVLwFvTlAZfUwuUYiTCL7Jq2BSyiHs1/YijVqO+M
CqfnByT4eDzuW3ufkvpkaW2qM9mFywBPwx/7ZFj9sxh/GAaP1/7vRZCS6Pukf4Q4f+TmKjbLzoUF
3ys/WevM3W/4JlIeLS0dWQOkbSYAFsgDdu9ZRcpgn4RCeHYZd8C0StKbj0yHMK6Xv+re78IBsoiC
OBOVxzCBL53DjcxKqpY7yz7S1cd8DQj+cC+ZthddHW/SRgfeMdjwut3emiYajWuABoKXlk6zSdCL
uLWaXA+NAMJ/3zwOlNJqO/qXV576krDguWISulWalvY4f2nAX9iz0kzNahcYu+1aHQ6Mg73wWjlE
6N3JCHayxyJ6B+oe45laiOmJoeMLdG+rjh5H8w4f0wGjS260elz/WooEWxMcbCtgqMgngLtZaEST
99g2+iZx25/EaHHvUD4nvZWIEDyVKzUMLwSFwCce8ZeXcT3ilu8hm0sdPUPEloqxP8f6uhE46EvM
YE9ataLH9qMakTg+EJgxJbSv94sXdfeVAAcHf8Sa0cIU8IP5sq9vdqp8SV+ufJHbFaT44IrhwUo9
SXLcTT+rCaX6PkWmuHlei2F0eczu7XkUpQvCd3k6RHOMp+PetNGfgfTFZllh7LRyzkYhZK7SGLnC
8TPtiNjPj836iko5xU2QRdP4eDpz2EtzYVopl90kugxfV1GBaVgKT+jmuKBex6ruTHCuMSj7zPRR
AbR2X4y6vyrL+DDDSDP2q6275L5E/4oGZsS5nH4kM/NGJVeJq7EbfUObQZCU/hWYEvZDZ1XWXdqA
yrCgPBVsVp47Fw5lOK1a/RZUO/U7334TbCQjw+v2SqPgiQ1ts33h771KYg5ehJwcC2h92Tt7xlz4
aNH+7oiEupY1M+JWzrWv9444XHkgFxGu23HZqPX1bEN3tlRrqL0X4maPfAsRbf7mL9AkmLtJodtf
Qdh99UkWdUjKdcCgCCpQd9UHl9fapDDg4EeSQrAcvGKHqbucQY9BzcJyWs3WmP0qa4RtmUsfbKZi
UqZm0+DbK7EypOa0P1/WLy3EWs+tCX5ohqJ3mrBIOjehh6PwFKtqCkTjmoGnV+huru8Ul/Ciey2V
oGh+9wiOSo2gYr6r+Ivyeq3txL3C67B1/gkRd3dYNxOdqZrsXIL0JQr26EjQicftHvw20jHdbqV3
/jTayVGygFEls3snro4H26Nym55Z0Nc8Hmiun9lZ8GoAPxEHcax9rM5lc03N7fUvPxJNUzgJWinY
IrdW2hV6mIurvCgq2q4JjnS5mq0CFfpDZTuCRCEeDJv6gMy3bxKPoS+NcfXFsYQLGRr+nsabA29l
RH8iHXkLohRaGqapXb0llEOskqvOZCk0MFYP7JwhHtfWlBgSi15jGtkpSFr8weXLPcWjZNaH+x+N
bATzWxjpprRWQ8gyc+bYZ/FP7N3HVTnveliZyoVERMWPAlf482ummnKxXVo5qFjcBkqn0kA81uXj
nhwKJJw1OP6UyQ4nRmdz8/ZKtD9cDhz1wTt2XM79ozdvQqyRavTvI627y+KmH9kYPoNS7x4H9lwM
yHa9WOGZydL/QSqDu1S45EHVsp/99GQiUWyxv0k+dYB+M1KDxWnoI3Wa2LX8RdRKdyoUTRceKdG2
cmipL3EAYnFdlxQ7AEZ1YS0xxHIJBB2gZ7uyrNoJ4R7d/OdbSxSalC4Bt5ANWlbwXS+pWOEmtn0f
cfqDgBMg8ZphITrUYLr5+vQ7IYYi0s/l5xL7G1u1ACmgKRwxkLDf3CVV8IN8ebESnbWq2i/rk7FO
PRvSz74WzkY5SigXomASAOKwB+3fo0BQb9fNSbb6G8MMhguu/aGQlS2FI0S3vXHvfD0dp9/dotS+
mt5Wa1ENRm63C/PY3dSVabScWGHmFNB5sYTVpXLurQNVsNfFFz0bYcUZNa37wWeBtsnayLqcSxq6
wyMr7c10QTa+odAePSLjEJm2nrzX5boQRTUImMdexrU50wWCMfphZKgJa2qoMG0OMNbdi+b7XRUF
cc+m1UdnT+z8COu5Ua/9hknC1xqxjlOeZZeUEZc3+XUkZ1nlzVTGRtxNKhghZj+9lRlUNMwFHGSH
DQvhSikP/p/yPVRtxCSsdGZ7I3S1DJM7Y0pk1lOOLWM1zg76UrrJKrdhU3tbZ1CiSI0t8irirpSW
etiBJ3tOg/2Q5t9/YA0Z1C9OobGsvzSBlvHccDZ72amXmgcIx+ZAVoBDbWX66uy4/hX2uu7yNaTz
z/7kN4Lln1VfIEogZHLHsLKXnYIiA0797IZquIFxrrLSIeNgnzG+hEt46MLv9EgIL2DtRYtCBZEf
St8pYtR2oTun1C4E2HGJWO8KxIiO49aADl5X//FXm8LB7LPzTQnOz4u1E6JgbXVkaJ6Sbrlkjv0f
rN4Ay5/l1aR9AFHA534QOnUGOPsItM8dZrSYtFp4f+ezc86yb022HS33GCFERz+Al6qOViOq/oYl
x+hC+ZZ9szLhZkOTARHVlb5Q1KsAmna8TanMGGkH8dLrHtEC6t5CJSVnd33/Z/kmOqqGW6lZCj4k
dfickS5cr1VHbttH0XPfuljM1yzmq8bPPYhIrNcX8HsxP5UKvZ2PbbZMJgOB8O6CG1vpuriIGCAc
Kc+B4mwC1NZOo2gkASixbXyfzTdP5R4noxGYVaOOs9nPCdLxsKLiUuOvSOdJyCGvWJkDsBU02UQT
Ei/s15lHQRFKVx7Vjhtr1zdk1QyHTbuW3Ij5D/rbKFdVQxnz1jwTIulsM8/0WQD3n3mCtUnx9+Mc
krzyUeMDJoPLy+KPphnCVOj5lcLYHim0XetrhUElinjN35ZaRSAufhW1fysM5zN9znGqGPd+j6Ud
tKVyg+1l+OzVOSC4ckmui29yMCXFcCwJGEkE0Eff4ts+rxaSF8sjg15OT45+Ej3iyAUZx+hEXBNC
7Xza1BS5IwHvLc1tcGNRzQ72ueYTbm4jePZUcaWzZtTg18lLm0vZ5EIAeDIlRbFBBrVbkzqo1fUQ
k+Mfa+jDlSeI72/dUlBhVpPLF5fnFEq5bU2ro2Z/ED9DDNJjXytchtTL7xM+5Z0aaS2iVvbrQY/u
aEaKGvt8lrN/P20y0+4Z1btDqOqgZXMdgd5PgD3afOlI/zRv/vzziYtepauQbshFYGMENnYO1a8r
4dGvUrOLdXZys45lerW95Zb87IAFu/PX+U/zdJruJ/yIUawVGmFKFzzZdTNGha8+NvF79qSuEezI
fIc0NskbabfHkm8GcCUJTtCRIdDN/XJg2bb9i9HXSs3lZeRqg2vxjPPK8pGTjj3C6+O5qZ0hi6GZ
gUmSK0lPPTNVFTEnYSwOjbSNYQhy4pj26MUxjRP4VEyQUXOc7URutcJUIn/ze0oDtve2liumeT/t
sx3JzFXWxdqgY3GVe+pu4Kdkir2cGMTXeTftf0wVE9RK4+x8lyox1aTSzpw+zB7GD0yvVzfWgvqj
SENFc2gktqUCmKGRgVCLHAeYPZL6UiLfgOpKGdQvTkPUzoGg7HW2WXGnR7QVdx2zXrqMgRUZfxzE
ZL8M10xKBF4kCa1RzMw8E4v0MwMGT+7OjYs/AVSGj4mxUJZ291ROU1Ldc5XlWV4a98d1TYdJMiD9
EX4+c35tRRdyTG+VOCPXw0fxM0GFs1xKcbbYInBJGFgLN3NqpUNB0z6gjGPR3VTd5NzbWfPoOQ/x
6cgyCP7RDek9r3bIbeYYOzjmL8sGHZbfHVDwpsa7JMYtu7K+5j+sZITlfTbD3A/wyIUAHC3tGZxO
zwlrEH/VkH+gVhfwwWJLloK9mPmiVjjOsc8sW2d/XZDAO3Y7soM2SUSS2CahcC+Y/36SCIBLgpjr
oLlG5u3O9gQ+jiJ3cSWinxPp9Qyz7WNuNQz2zlwMhyU/m8K6jGSZyBU0Sj2G8aYMIMfjzgjQt9MT
4tu1eJsSvYepZwORz+sxjhXGEmyDz6hlWrpyYC/8MkgXyexgKKm0DYm3iBXWroxYU2CtgP52QSnC
uhfCwwFcIlt7/n1d0piyiBZ4QLvFiitkF6ZLQAbskP1H1/GI/0MUtFxDt+3ROGEXuwF/wSadgUmQ
amJbN3I0SA9UhsLynd9NXkguSxz2jX887y+j1MUQAEMi6tE8cqpfRmipvubkfKNlY751AmZEXKLt
xqCX6t4cMe/gkDIoDZzRpy1ORN1UNn6a4S8GdHVgkEHf9zzAcuOk8ZdtN34OrH5dGjUry68hR+O3
uilAhwqz+SMroJ6JZaxk8NTzRs8ghF4wVjBvGGKSgwAJDmoNqb5bCTqQzbv+hN3WAc//HLT89Z+u
SKGsOruC4U6VAMTc7eXR/irgc/xoSCTBESmu/cVvcywxVk8vzbPQSu+6ruekQwxxAUaFkCzwBPzg
k3c06I1OKECnevDibAgGvy3nKGRqHb0kgORYvze0pu23W/niljZ8HeJPAz7Wkqml8E3KK/gofqWP
HqyHbBFVVBUKhg1+HJLRGvkXdiIgpAbZld8Na2n+yjpos6MIKz5+iTts35wX8S12EYN9/r7LvCVZ
80hE9VGuTaMq7JIcMinJTa85meW60syv37Bi02UdUEURiAUTmLQzg4M54yojq2nk7iOQkJQMnx0M
qvZZuWMfOtbg13QsSyX7C/noLRrXaSGCWDJPeY5XqCfE1Jm0qxv8/uy8xbssjLBr/0NfvKNSJVx4
06vThajf6gSGO+0U5fDNfBEBad6XbA3aU22tfVJ3Cq6RgR09YMgml3JnYmHZInSaMfYCVuZ3hAZ9
zmTiFAWmc8SyTb4BJUvW/JU144awNF3zOMEd49In9dhhh4quE16RR+6dA+F8vLHQaDTwU3XElGdj
9Qd1w4D/jMFA3MFgEIaYu2gRlvA5DProYaEYNuXNOjuPgExLz3LmpS9slcpCWote7xTHCuFF5NtR
sSVu9xMkiQd8QxXPGK9PFeG/0q5iWxzJ/gBFQJg2OApxYo841Yw88SoHQAOsSpSECy6sCIN+pI1w
c2VNfiGUbzcwzvGsGTnLKZ8lGtzZJi/ASt8kTMAXbIbIfBA2ZfFF5TVcEvsW2YUZR4+DiSls32iH
O+0/ALJQMk4xe4S6fHGubwg3HMMuqYIfXcoNAKzjzopU+FnQcsvjbnp660SAnXQqmZrVvbXhZPDv
UyLnmo5XcP2HSFbrcDz3aKUvH7Kk4gc/cDbJlul+Np0MNshUMos622YwmzDr5ZCGrUnEoRnaeB+c
cDQk3nsH8vbBRTY8Oy1TyE2KGNHZZ0rqMwCDObPoRe3vXkfHu8DSd/0OPrex3wSC4+c1K++Feeiq
mE6W0EM4NKnZEj3gaPa7IZ98djEbnu9sOybEK28Qxws6w4bM0JWLnhafcC6Odc7JcBcWnw3s5L3W
A818O3bn4ZEdKKLE/TXrjMP1xz86W8PsfBmFmCGFCzbJyeHCFVA6yIc8N4f+0jS424cyOOpfTPMi
X+Um7Vn6QcRmKpZLx9m8fjidJeMZqhnd9NREvZFPI4wQq2YDYmgaVMn/i1GlYpDKuUKq4CvJGpNi
I/ygvLlV5VxaMi/eVdxIuvkz3F+B4guofE/oZ7XcGO9zfzBz31150tD4UfCINnSJbWab6D+DnbzR
0xQqH5yJvGoWyT+U5zjsryaU7nHyM/4kuj39P2+585GyCB2/zXylcYzV8qeiwOjmUGuX2ieaV2c0
+O0xY30bZO+4PGqjhlFboJVJPG8pywiEHvjyjaEVgixkfBajOAl50fdCcfg913KA1cM/MO6um8N0
wnWy82feaa4LnAqZ73svpTIMEAhPfL1Vu2XoY3EK7RUBXGaewVaQcUf+rT7aiggK4mpqWedgY4l1
31eqwX5DpJVTzFyXWyjkpJBmes7O+VT+uak5ldf2KabJb2cmjRVtidd2qUXjLtRegx8WBYh2dU27
1r62aG8VU9U7KcMvuAdY0kRROwpDzWm6l/yvgjYp7zK4psyT/j4KL2BLHTRCzGIQtOgWlTJWtmhX
iE3oxwlXRApfa4mpdXUe7iNBicEw82IKEb6Gn0FWHQTVxLaTvZIa1IpvXlC0btq1cGmNnN4mHe5I
oCI3UuTTcfXr8KoZxi7XJY6SumCU+2zrvX91z7XaE5oaWx0he1QgpfCe8epCEvBll++gRqsmH4Gn
hZgOpPdHi1p7ufUlwR/oR+tKd7Mp9g14mR6+8kQLcbj3jCncmKoUiJ0Pbtd9NwT+rF8fwTI+ZYkn
yVx7ywExEo4Xsn28RMu7jZbzpXwXhI9K6Sy88KD4YiZV2FdwtLTA4idhGSxc9iRcsMUP596B1jkE
J2bEEJL0y3/xlwsBkxb7chzSIq+vjrO/31Wwii7QbMG44HA7sgi/bPrq9Q9+NzhDiTTsmQpdu6bI
FgtWL7zLzImzJ31hNqmK3sb3AuAsdfAW2Tl1YxiCkm2N5/XiG9huHldaC7gfAH17lf5jOA0Q7Uvi
ORKYC+BSmY3Yd9N1Zu/erCNO+VPgsT3tsqo0ZpZocII5CJL0QRp3KNCxEU8zqmI19wLlZp5c4h9S
S++6sg4AMmHz6SVvFec8NGA/F0++1I9SqKL9a0QNpoZltJPGCELCSHSUw35ACnohrBO8+cmjheAH
/vkOL4Wdg0LMPmBbQzvX6+XpcDz9uzViDqFrrS2ezNH59qWqIhxCj9yl6m7Ye9sVNPkbKQjXh6nW
110gsJIh9PUktq/VG0CNmDrpxWeX77YIiCPoDGkqmOXnUC6xWsgLb+qrxN65Rx+pBJRhBl8AETUt
j+Ud8MtAotbwakHoX6CBJOCzeYwcDWdqcaEIlO09eIgJgPMAFp89RjO5Rk8JjChsP9ZT56mhTpyB
/60C+KpA/jnamtH/fruWPmEbdmpb4+CM2UqRTHNUUmXXjZf9a/mZfB7gQ/Mgf2xJ0tMDd+qSgYTv
qyU/9FSfaljrzFm4rLf8oI4UbQvKXxSuDwLlMFpmNdCWDidfcLlymDeSdkQ/35De7JMcyJepllQR
WOQE4NBKfHRC4HRn/taVD2Gt09k+f8tBufA0FnVo+VVecqOQWsCsH8dfFWOg+nAwDAtBiT8gqNxu
9GMu7qlqPtsviY5blKJwuGn327RFllF+ziB53WGGNjirlSgT64hNbSUv2dj1aIH21RuybsdfoWRf
oKYcc/8sLROMnslMZQ2W+Zg0m9e5XcFYqHtgS8mxpeO02jwHr7Jt6DMlVHpC/M19IZLOzM685JkH
LeBbQ2K7dZKZUs8xAtg4pRB09GErKF5JYRhk+EKXUQgFVJrN6jCKZrm8rApWHPBSP0VRV5ozdBXo
08tHqx2Pd28HPEMRtvN9vkUa3JjobBduKupJ4fKpgdi/D0EN+sm7EdEP1q0zMC9lRQ8Ro9AQmo2L
5hgoRLYrGU5k9sOZmEell68X+LzzBBS6nNi754XAccOVhE2pN2hDBtwn9bGII0wuPu3kD0nVzx8U
UfbD2K1aioO2NY999KsBdDUOHmI0O4qnZNPtF06758kSaJM6anFA9CyuSSrITdpyT/4uA+G6Ep8T
itQxfYUoeCr3dG+bElPk0Ilqk/tyNZ/KUokOTjw3c3cZ06CzA5YOt9onC1irkcRURr6+Ug+fZJps
ACCRXxDN+IbVAqSTuA1UX9xKapeAjbPJIn8pkjmdJ6MOp+DWlQJlmyBLXHrsEZwApcTIRkrC3ATF
AmPk4/erZRaE5xnTeNcOT9MHjvZcT0S1lhmEA1h38keoIuhgwWBz4g2EdBgAXhCu8KArKAxePggf
CUeMUi518l3uxVbE5wg2ZsZu21bN3N/wN39TIG71dSrnMYsc/k8ZguEg17v6ujSfw1lWySPu4v5I
36Fjo2y7UaHmMf9l+5GJ5PBlYsMHgNA3yQob9fsSJJXtRiTVHKINrGYbZKfOTPEDzESRVQ3DkY8F
gLdTWpj86WeidUstG/EczCBMOLqbW9Iv4hFMX6tiAk39eUXdfinuF2bzMrJN843Z0Ca1Q62FIqPS
+04Iau/CxpUGG4Mvxy7vCN9gvLpxm3dVY4x/Uz6lM3P/7dKd961yvFiMQAttg02dtJbCsm8collO
Drl6lHt2Bs+Mco7eDIsGUl69b7KtOOsKj94fdTbMRHx3st5FN26ThRFFHy7Cmm05mQud86UwDPyB
3+XFe9vS6XKbG18BPxOB76xI0aDHZWOGZZXYM+X9GekUUQUfpRmguzdMjZO/T/ZE0Gld16Z4cgpY
AKg0qqDp88iExXLMhjpSI1LoW9n5dZE1L9EBoVKULR4coYkJA6S7Qu0YKpM+AJbAX9WW9KeaS/9q
HdY9eHyewsbN2dxNMKyK5sToMMiL456vLUmVX0MFXER9lY6pC2ZSiZ4qDcoLg18dyVhBvyX78Rvh
S+DNutaWwyhE4XNmDYuJkc1Dac8If39wUzjJfUCkDYVWSrC961MDKsAk908wTdwp94OlTMvOMlqv
ftzq+r+ZLqCjRdZPMf45fkv19tuyScYtPqG6ACQ7/qeinlk4LZRmrVMlYnmaOBMPVu2ULLY6erRu
Tia85VkhqAsHna3GQcVoXFodKxACdWCgOOtq9nwowddqmNYrqp4ab2fc6ycN58QY0eVf9UxzsDZ5
EwavZcLA8ZRxkEj0QPTCYXMMHMub/zSOSlmOUPaFs0KZIMSF4c9HR9+xK6vNt/X0pLsPIHqJx3fX
WkxwT+3NSrauycsiAsdoy7icYatoYcrfKQ/2unP+FeVSxncATJ0CxvS/m9V5XecUVcqWRGzyGJeG
bB3EsiYxhBLiXRN6Ogk9wbokc6+5w1Q9+7fnfsi+P3HNRZueKoaibFBIwNBQcfWZXPvZ5+8WlJb8
eK9l/x3GOFCQ/i6NGcvWkWFyd7a4XB2jpXM2W93w/8rsQL5gb8K9YEDLp4utI6k4svpqthdrgEJE
kKrKBpBEHotEgkp7pt9B1pYocYdSbysZ/hDEohWymVMx/dka+AnaqNRGenAKiRMI3bdT7pcONrXP
BFmiLNK4o7hsg/QWSOJ4aABKszK05icGBFj+sCoXv5gNNKiYFI9/p6GdBQE4DwO72nIrsTJP0+i4
RToE44KVVDPQidIqEoEp0x0c9fbTNdrYMj/CVpGoYvhAqMDV4lDY7/EYDlWm+xEjLl6KikJEaFv2
dON8IudBjSJlctCITdTo6ClRSDsCbzYcnxJQgV7i93LavPdiWKUISs0LcBA3wZ8AI9fVtg8TFGxW
LYkhJGAqbsI45SE7JwrqPm9gZ9a6pVlEy2IxpA3rf8brMTH2pB2nfbSY3Q9yJqRBhsO3barmPIte
h0NwlJDw9KeZOZy+VyaFzepIUUG6EDEjBYRl21uDw3dcLcG5vJkXeVdTtHJWnpM2MZx7r7l2Ev61
FuiKziLzOXkgiopk6BGvVWlNKbiCqB5/9Ogr0uVvcCZiwo4H02Qg6zdU9ykiENGmykeT2Inibhgr
4b4mF/AIypY/EplqgGCS9cMtasRovwVftiqyGfsj3+Aq4dSZy3DyQqJAIvFCrrrzTfwLKznI6t0M
NhjT6lZ+UXQ+TlZfv1GM5B+IrOC+ELVCQki0gJpedg2npuj0l/FRQkj1kAiHTJ13wTRLCK0vaOpL
78rWlDRss51vy/oIVIcSDmXeKeSmGXf9UPSOUXMwpe2jAYHyjFm+pWdO/eJ8UoDryufYOkuHZow+
kIzpWsolnsjMTLCb74lGR55ki2AOHScPs3ydnncEgNQybjQYfkQLBVd/uHSfrxCMzMdhTYFeuzZY
E1v3Ri1qeKPD4CrwoXon8vwROD5k4WIcwmWBObb9fy6bN0z/hicAR7gWiIB7Bhgo0FdAmIEk+pej
994S/KsIGLkFEQUl6mrJnCmINgfjlgK6w501Z704WvUtUMdQdCyugbJk74/EvP90/l38uPNofSXY
hUy5umSbcoA7g7A5JsrReTuAXeWtgJkEK+86zizNYql5iqXTwHfFp/SrJ6dUsoZUb2XsSKpdMzWI
O1QMNpCubV7Z4E2Jh9CDEqW6z+hP0GBWiW9haRDXpCWsc0CU3oyQ7DmJZw4DO10VJDmXAMPQiaDb
Dv2JRmmfTmfjYQkYZzLfNB71cHskBWhav+3fm5Q8kYECSsu0BoCeVGA9LLyQt0R3pcCiIllGPvTv
2+VzgHBIsUnrr1JjEVr80SlXnm7ZUhpZQ6m63JYRQwhzShVPk37usWy/zyp4omLP6tfaMpyTz/2D
pB0vsTGTNioVNJCP8baJL8Bg4iQPGMupoM3Cf3mbuHBndLOa0kLBs7AOpTBLDTzW1zcf0gxK281z
6zpO8ENLwCFBrBI1Q35S8h29Dz/8TrzlIUj4nL4an5zffY1GncRb+UMU2DGy60eDZTcY0G5XkoVl
8gfVABMNMbplo8aNd00IB0vZYbueeatg9+zTD3g6ME+0RIfzTqIejTO45ojgHNykLudG4abscAY2
CsZIB41HD30uEm6bpZPnIL8NTvPYMRPxKwi5xoNmcBK67ZsqROW3X56ViybN5Ow90HXTOx8bLAqZ
ZtQcZes0wzegB38B9OK6kcRSRrH27g2HdVn6YHRYzLUDihH5+7eTTRWLJUbqtSFp0OObQrGpSr8J
dnCs2sP0vRh2GONKmZ0V+3tyL4nZ8P/K979jfLbWvOfYgb0IoTtg/ILTa/maUxaXQW0AyXshS52L
yFvD/zsr/tUp9YVpyQBasZqg1ioKLWFa8rrpuDfUjv5yQfGRH2eEUMIeqp6X1PCjb3qgkPPZ2Rk/
hnT46loWhRm44LG4zrfAqd0mt2iGa5LNLmGhAKFy9dP3t52o3Cij21J5RAaDqMx9QeMtROqZPqZW
qOArP5N5TWsu8SxJ2D+3UZSJHzaNxdZWhwgJcY0zbmvtgdF6RJLph+GdP3drPokXWSU/AzZHyvMK
julEMlfKU6JWsny77xzs3dR3lNwKCWRzubjhvapWnlIwvjzSB2H1POsKqEZdF+lKvZ9Kyc/WGvAs
aEXGsytKizqk2UmMLNeCrdpIGuc/dfC0N8pgQJMTuyMoTzNfcvOcO276uMTUNck7A3y6rXI5KG6T
+afFn6/MiusPGlZrTeR29aZu5gFed3AeIUGB2zfAOoMB5mcrtDTRpbiqAcr+g9Vas8wTo3LMXFg6
ueABguUEYmKreVEtr0CuHzw1Y+O5PIaTMFgdMue8OPWayZwMmB33Q6lxNLvnRxAZFWztzNTZ+28F
gsgiCIShQXLTePKoQ+hmg7xUVXiqmUJd5vwXZALG9FCbGI+hehCYj1c6LsHJ72bfoMxbQjgz3nCk
AiAfjE6rw0Hv7z+xuoquuV66qUflmuwjRe9Yq07Xo/BqFMunc+IG7krMdJJjR1Zpr/g0HFW7AaaR
LTaoM1UFn579cWlT4PmLDoM+A8ofRLsxEGbSI4jxgRtA/l6NTYZVeoSboxkqAa7ksm11zzSq+3CJ
K9YsSLhhXwWIVBBZepsex0pNaXkPsmO4tirDaSh6MxU4E2qxcgGUZ6PLN8NFGqZFCz6hvamFNkwQ
9XZDHWDc4dungMkqOscDwrvq1pi+zv7NJh5snFge/4XjYUYwUiYxRsayqsOKVPF2rSnK6am/ZQVp
srd2v/txguEcBs/kOkAwVHP1SgyxfAXdY0ytb1vvBbnRpLiv9hk8lreDrS/MQRzVmm2NegKmTveX
qJJj1Oy2WPHjh7vkxEze3Rmsdfphm+nmx4lCsd2DvvDfobjsfLlounJ53XIisKc69b6O1lWQkjwf
Zas4zec5UUKa61KC4FN1E7uPUKZiFVHmBf8nTHYInbBZfTbSRGnQl7tmtBx6hlZY7wQH8YHdLQTU
yWhxaBDg5E4AmPZl5Vomef3uaD/HBzPVcYSA6jYu9XwpWRc6IFIRD/Wp+JuLkWnvw1+W7+A45i71
poNo1gSSdcsUK3hbSGJWHC4hwwnwBbWcZcOEgLLPBtUQhCMfw9ggcdMFmho98Ktqw93N+9fyEgD3
XK8iYZ7rXBl8drx0LV9x6+Xkok9OOmIjfyO0GGLo7c6nWw33r+8tsNxWpXTee5CRNwDBht8NUbi0
S3vk4Oowgm58pbjZQRmdeMcOm/x7tSsz8wNBBz+GaICMQnpqLOcD2YkschbJcyHT9L4dwVE3enj7
ZS80rxEypNeHdXzanUtX1oJEXBgEgr0Jl17Aq+ai1ZBATPoFHwmyCjgUr/XpsE9SkChuuBhV8yDP
u8M3Mdmz3NnPyCS2Kc/1p1U4AT5iswUj5cZqY1icoOpwjso2UF0r0mUkaNlIEDtjkD6A5mxOLccs
4xIMRMQW0FP7tm7bZGJ5jwHuz946glHuPPSNn33Eti0BzRv/KXd6D4O12x9X36iLT2Io+7iaTWY3
RG8Pfq/xpoLEciWwEnxeoEYzWsoLwTxOji1XH8yXbzmECxWHjjLEoNamgOnKzZ0eKSEuedqC5e8H
E3ohuLlQMWB1hXjaeqg1YQRZ9a+n2bMi+ptp8f7ldJnZm2AgvC8l1rtQfDE36YgZOHmAYwfMSRZQ
A1rc7L4lecRJMuJvVjvS5twXJ3/CHTggoKFseXMxDvRKeiZgx+eHNGt3FCZL8UPAe5BGqfzc4z4Z
ryYW/Ael0IYLRiAwfW6I2JQfuXt9PVv+106Ov76WFogq8neig+u6TpDQPalezYq2flCUMmDYKkyO
L3GCaL4tLxJWYfU2ZKK32B6lhncxEd75aLNWjL4XrLJGQZxdfv2S88Hscxq5ZyZxpmucWCk1DeFM
3oClp3RjPo39msk2drF9B5nPObEc3+EO+Pvwnxe8SefxMxt3Xsb1IIpINg1ZyN8X3XKnNEvq3VrS
R9FklMrdZoL19+bgyW/7wvGuDLprK8utNeFqRgw0FEOzXmnsL1bhAW2kaHKEFw72/q0In60mVVM1
0p+pyvAUL1Pj9cgkksY948tb0MRURcqvbybwp2LtXvKNcdsVzWJ4HlU9QVDqxBI0cX3efEACAUUX
L8uVLHt1egOGl4zfg0XDINbTXbzZgWvSHQyz4cKDA2WMiwaEn2UGzogunvrw55RPUE212HGVdt6h
rbTDyI1DWDSonvUwKwS7RsESbXcmiHGarZYOlEzi/tmj6oJQU1t7HTal5xirYbUD2tLvNEZhtPo0
NV7LkLhmwgJR+T3vGheaUfmkR31T6L4m6WpXF1aG/QDMiqUyUAZreQd2NiARB5wWuHNp2OaC/s9w
kXv0y6Gi2ZQjkcK5NtQ8DY8+9e0WyXuymnC6N5PdpuSRYwORCZOavgq4FEvcHQ0UzdCvwUEv3SPP
YS/dNo/IYMH1IY6o5arEC5R3wFbYafJn0RsDzcDPfHiy9vogGVNRfThDD4n/Jyquud2gsBEJnWFe
I6z5zCm8sU9kgxyoDo2y9ZNLGg1Kp585Re+8PWsLMMfLtmlkTuSLbyyAE3bKspVeK5lWVTolp/qL
BLY2AWDmOxqpTdj75/kFWbdmo8EiLOTuVUKaQDjdqoRUXMpB2bWAMVS1IdRGigD2Rmwbof4vRPCM
7yFA+vTZ44Ljb0w5D8PurXBElaB0/ONE0DI/22lNwS3X+pVtSkd3W+iS53R0lYDqY9S8uTzyvOWg
x4Gx8FywQiM0Xns1F6jXb1AbVG047P4keTXIcW8RVK9R04KMdz1L4hqgRTdD3XnUoDb+LbcOfGG7
EaDSsvCmExpBwdsxUPRCYo6Eg0MhjskrMBXA3uJwrm1fNWi9op/5/zVTeiAVSNJzF4qz8OlGvA+x
b1c60K8SpluD00TrxuVC8KeEyXm1sNoq1vzM9UDaqJmFmE48SmIbRDgRbbeS0bUglG/Tg/hmiMMC
WB4D1oLBBRvz9zBaRlRRjgoShuix1rSD23hAR9qKpNkooa3ugGLimkus00LUusprbScf3X5jUnj7
QjnXqEgWgKQUTyVY5MbqDwUYNt4fcnb1Uu91WsxSf1jl4/mnVgqpzXNZK+V/lBAxmj4r8fTBN+Mg
c2vXx4dAAjcYpqv9rufPAgaMLFmK8Gj/1H8HZ75HfbBqKhZ3dI4qCVtsn7RiQQ7BVD+q2UGsY6q0
m21uFwyT8EqKCKUngEnozLtNqijuZedaGG5FbH+zeZFQzsNCWCK1/iBsmuQVkFWskAHGuNX4UTVg
UC3LQG8tSExLHcx1zVBRtUbSIGdoR4yQjqfdJc99CDfxrh8d1ev7jInOwtJzyIOb5Vq74MxWrj7E
d+ZT2sYKJ4EKUtFQofV3KoOay1cmnIp2+ipE2GstJZe0EhUqsezjWKm+CsWnKCnUBCvID7N1/5el
0FKqoM1N5fnQ+0CSSC+IeyrT78LVKIEx+X917JvzDPiBW2WMVL9WatPmYtWqhyqbZaEBKPufoHk4
MQO+Z/hMt12eZ4yHFKGRtc+SxU8KH/I+PvHu5UxsAK+2UrtDkeE8UkUmWN+l86isxeqMzaTePc7w
tiuw7zxz8qCNnRimVqwPkDZUxUksdqP5Zvs2B75Tz3QmPSnpLBMHElygECeCXmF0iU2xzvt4P2/A
deWTvM522XcJ9oll2MrfVXf1lJlUdyFBwFzdaGIqUkSt9CRYJZU9yHUsTgN4Nx5yDJ0oBZyd88QQ
gQiALAE/JKdYZkVsa353I39eZljk83wZ7xLklbcvauxOTDcI9GHJMJ36uD7+GdwIYqXWGJ3BQhEg
k9kxj/fLCTSFC31X60Ep5WYocG3IIITwVY2hDDNa8A3+p0pkx1njDNAIM8N1eGG7YnaymRiz6XZE
9zKvv5rrun2O/PG4g0ngcBeEWo0dRCLnLSk0XHKx1j/jcjZLBsWG8Hjq1dn37bLZUBkOv1+nai37
5VpX2v9we0b+8U2kxtw41Qt4mknrKYQNajqCxWx89x8JS54atb8SdfXTscDtU5hfQtbFzbbtdc6P
BEv+NfsKbvi/h3B+MmzyE9LRKeEY6I6Luu43Q5N1ZzfCh/rcOGP1LCf1DBHdEbQpU+/pMxOj1Q7G
G3wzVNqu6OesI+Zwrxx07FIGfh+1yDj5e+gUsILWdqGLzFuUrClRDveoMGrJq794uhXMryCGguqE
l7BfwwlYqF4hC4Cx8iHhjGCM8rIvSZt/NTmeac0lCk+v8B8PFf67scanFqq2Vnhb5Vn/ZMWxwLf6
S+TDvkCFT/wLqYPqlK2p3y+PQIuoTX+31IcNS9t9k9XhT92CSYAa1Amr4zESDq6gC/jlJ6YQDNXh
/8irkeX3Z+SVXICFgRdWPi065lpmd3ywyG9tTFD4YyndK+Q9PoS8vE4FnE0zEsBBS8tyKsdVIOZD
kTYfjhS1KRvst+ZJPK2bCSdGtagPn1GAl/cPMI8EsKQqAivCeyvpR0EHuSkV/bTP+z5cL24xCQoo
HAew1oLfnI886vcV//iPEBrUyJyocdxoglusVXUI9TSrJmoDrh+LdV6dp8sfym/2fiU51ZqYzHvC
9yepSqRg/5K7Z0NB5rX0FrL+lT8gHgDqnYzPCmVQhK6kUqQ4cQ2o5W2w4T53tnyy941RsQ5nIli/
ZAjTJoTX/IoYMfoFEYffPQz0ldZWpZrs0KKFxLLSMM6448iHRBUQaoUazDW0JOSQjgZ3pknCIYuq
WN8JGsRppJK5Vp4fX1YbNQMUf0PLzYuLIUsAXpE78lvx3Zv250KStERRUT1EB9XdNfNNDmhMU3IO
MoJk4ySwH+lo+rcv+NcaVZRImJz+zxxNOx9XPYdTPEWVGn25a1BbxbNkhRXXN3Pv8RMopA5pO3sN
PCVLJcvnip799k4gtyM1OO2/BHARHl8OZES+ASx8XfCTn96u/NIPRChNVTE6SbB4XDlMj1EdbZOa
TQ1DGsw/bHXxRi2LHW0OqLaaPct562S7VAR6evzkz8nS0udyuh+MPx1zrW22GID+LB5fV3uyj4Hv
vRZlhaRmfOrYA1DaalgVri6myI58Qv1tA9hODEj4MjagpegSxoNvWavFaeoNcc8MFLZQ3P+AdM70
BYuZdtzuSrFaYhxT3jExm1YfVo0MIRGsZ+4/Ds/a9Zfayx/g2yqCBGsCG6I9RDOF7f6MjH6Rh3nG
qjijY5IpbZQTb7dan2mFFHfD3cAtzZVILRaYkXCAMUmhEw5hGnuPcRixbifzIo3ge5EeEj8WORob
7P6sefXEUSGtJMTB6rWc0h095mEkIT1aF9zuoEefWJU8HThNkDRmQwmGxVXWC/Aym821sA/m7Ptz
MOWFeJCXM1H9zyNoMLlOewhBvhvpDVCdfUBGnC5Bh5fjiYoX3dsjP4FLjyO5u0+XgzlWe2IqQH9B
WdPVhjMxYz+T4EzVUVuOnZplUdEPeBXtmU58ZiT7CEMsH2W1uxIF6wwtEwQGxEJ94lhJkH4oMDqB
RQ/9qcyeV2VZJ6X55lnIj/kG08Y0bzwJkXE9XrnHl2pIRRDEDDEWahfhUvaYXbDldr3kP1lsuNsx
BhZBocLasXRnaWYzK97TY6H4yRd2Kq7ZAyFbaIemPb/pqayXrlw6nCKiMLx+SDOlQMvpWJ+BicyK
wIy22QIvi+qdDWLzYDC41YGFA/yHIpQrP5ZxSLLFfu8F8JSwyKS2cc+4Z63z2w2sy4BUleUIfWPC
OnFvIm3PK/+OztSAb9O64fz+D5RtHt8celosRc03x2Y1KYliS+ceQZeK3A9rzDh8rHBJWDhxUngZ
g+3kT0marcS6wigVXaMYYDF7eLMs1ZcyWAj9/0srYiAE7E/05aDcnErCMUqla6QcdcTenfW+hV4V
YFyLoHYj6ZwJlC+RvH1OukuWFUlySd2ZmGo4XCkNlFiMyrMr5vpMMqNHVVbQltmzmQJNL1JJ8E5R
hJTz93Qo8cjLfC/TbOpSHvssXoTWwiteH3DDw9feR5pvzRk5PF9rVd1L5YGqMPHQQczRSzwt8Y1x
QGW0lZ/ERuvbXAv3RSB7eonmbMvCzCpKzwJnkP9gsgKksFBBB0mZfvHe9ulbjb35UCKEq/dh/5Tf
+R8RiePn5DXKESDXzt844JoNNqiuCuaoKdoF7rgzV0FlWypwa1tOtd8cUxsmd8B0hhQNThgMiWq5
VyRsWJtZveUz0ps4YYlz5MbXfteyiPkhBV4/5MdkbfJEQ0Iu0tGQp7zohWtzbl4oHKGVXtgU1uDj
rZgkBaXoi/RA/WO0hR5caxYrVdwxMVFXSfgaHuBE0DQocsvem2E7COn0LzTQqZQRBhh+rpEGib3v
iHOwJnydEPN9dBFPuykvUX5y47MtD+C6mWPxIC0QTj5s+cumfGHnd508o8Ld+vFFM35efL9Y11Zn
EAzcfjduC7nOBTu8HLnDkUHUagspOPRg5IzBWYnY0qzaiRkNEY5iZ9unNLUwpk9dSBhp1s8+XzEc
Me7/oDjLxiHNHzuxYcpavYB4tE5LlfeisoaUEK4I+asBhyCJJbv3YY9vXX3FJJbYJ5gRwxqbnVOp
A+YZyvLdwviBigvj3LlCo68XrUYLAoD5DZCdxb/P295tkEvDBwbaN4vrtEKWy11PyXDO+ILPFZx6
+OJTtKJ24wWDSLQ1jqfWpyD3AozMEZ+TLwfjWKaUYKvhzmIvZo60cXD0GJN/W01XYKljqg+slKtA
hn1iJLo2RBzp91E/DfF1mGrHSalQFJG3vYXPA7n9jmwUiUnLnIuUXSJdWagsQcIJ+3IeslYOYWcY
hs3Y1r8F3HVL/BpoW3foMUo0aAGUAh0EuBJbYM6HylJwjQG3pSnTfASsxJnvJUfuxi+svTk1K+Vh
h0dHaKBppts0Jjh10l5Baf/PC3pezBsaREcNmA4dlnEzqHYUeuZ1id41FAjYvUnFz8zO0dcy2aAr
W89q64MKsJlDuig2fkO9OqlJw9qmxlWFcHx3ZJy0QqcH6KGIWeJKf4guMFLWmY7v7g08MalPBE62
voAqh1/kvij51UjxukpbqxSvktoJEmk35TpjtX7zWRrr1iWYF921NH3HgRAJa5y+78xsOlsSX94a
uE4jKf8PB2VDySxur97b1QgVsEbQ0Ym0Zm9y+N06brxzFbltEcxL6Z5PYobdNjsXLamcRfgFDhF9
Xy6eDaeQlmNdLsFA9Yh8IjBACTdRDne2pW2Ouuqc9XcboWooENMRKySRW8wQmwBzA5TtYAVJPdyi
l13NgSEaPhsD5VFHvZX589xIrONDYK7tD70mAdjzba8GpFHBJGW2rrUkWBuv6M1os5MQdqKbfptd
0Vfp2R45l6AMujcqjB9d5tHGfDA2TMLsthE3rKanPvEUjSn3KSXRiITsBW6myW+Z5vo0XJpCyIwU
e61xNeJD226CfB6lJbxaN/WuoBZ6NJQcXJi0LhDwSLO/pBvkCfoidjkbuXIIfU911M1NASjYLAWJ
tM0aOMBJncMLugU2OQHgC4ULUId8lBZ07tKjEcy3yNqXw5PTHCBVADf73yGHFTwBzKFt/fFJn3Ge
IGmidPRg6zwf9DenWyn+g2gR80cCkR+1Jl2boAzgq3oc5Qu9ZuFNQMXmiPDAsr5r58ybblzLnTVR
0NEMI9Rp8pTr2EeM2WHrlM9Jh9Ehw6kYSOvo8h48s1Wqd06LUjH5qJvdv23I56LKteaXGgmQnAc0
qzzC4wQZ0Djg20teBHVX1tIQkjSDFxHqLmgQZ7noDJtH7LhUOTTtOo168fXiR9kHTkNv2pBOPVVC
hgJCfgI7Bugz3WYxmjFI7mycchBHKfPr62vONfSP1YvYvPtVeoM+a8LFNcn29e04IlM0MNIlDNVQ
i4OSOjclDMbYfAg+5XOyrvbsKN2hkCnIPpMmdvdG5WQXIw3qzJvnbpLVXrrLLJfJeG4eUKcuVEu8
F14VD5CYQJEE6DoezM7oI7MawrtnNxmPJlb5T8nIQolBvBmTxzeLnDZ6QS9Uleyg5cy2gKqYSrBY
14MEDF2n5epEwezjBVY9XG1mvEmUGkJXdjpyvpJzOuStzPak7npXvUj9VvYRTn8VxgnkYJ14aatg
3AZ45A2ZcxIzvYsa46M3e/XlJVDBvJ9ABsaEjnAWoCnewKQKQil2ySocbNAS2xaMGSDphxZW8WWm
/rKVfqtnzqRPXiv+moI573n5WXfjIJZRGRyDGeydKtFhouCydJUfWVUkc0lWG2fRdm/oKYnxNlzY
VD1IYMd3bpN46KaHQkH3+Qfr4+oQ3e+PCu0QPAW6TCyUibIhS9s/ClmK6Gcbga3kJ9wGO7zVJHy1
S/qkZTEbJZSsFfBVJ+ry/21i/MDmygb18d9l31ku1IOZHg24xxoo+8BCe7mdBwzOH6pG+vCU9kBA
fJUnDyCl6TFwsyREnYwLV9/AcG/fvLl3crwixc0CHcd3ONMx/aFbjYLxB0vY0CqJuMKXaN/R4/RL
aFuoCRYLdf3VMgE8SzAXYjQa1lAGkC3ySWbiLLAY/VYWkvfO3KdtKtHs4qTd0U6RIrz3MY/PEYbt
NPcNt3xB5rsGRxZTOOT/L+0W6/Mofr5xXv7HzdqPbJe6IvCMIXLiFfbnk8sHJqHs1oObBKxsviu0
CRyecEFWGFzXp10kdhWCcS7fcLbIRIx+T3/S8iUwg2cbkFIZI3UCL6aL4xnR/As7PcKKdrFKiFaM
cgFfndiB4mdkkOiO79SD6jDnyvvTjUpWVRF0rmdMoKtknSiE9e7wFcqbR+sxRI/utN/W+mwsZiCx
nCvo5Mv+2LOMzveND73dKh+e+SdmthxFvjzeKAaf+wzWA32ABkYUKQF+Jo2DL6HxaUpBjLD7Guy8
iHloqtSATjaauCfmUvCONnZCFP8n2Vz56XULKKwfdcRlFXVOORq3N1slxOIKAznQMRrbUK3iioYp
6TT1TZuiNuy6M6HuJMDvo90LZqGoUoe1V8rcRoCy55QIhklZb9oZZCiXn4ZUu8HJewUQgP6y09Sj
7qWE5rNtsNaxJL6DIIJfmxd8O5ZfbDnJNQ9lLi07iJOdsdnj8mf1NEn9Uj24JuWA6eWG+9346LP7
noQx7wnsm672zQTbv6NWz1IkU79ELpxkd/5arom8vRX6eWhBSLwccT8K7ICdZwt0i82EwpZTFfR/
cCzODVromr14Qxk2zMiDDdNGIkp9WGpxK8O+TgskWl4a+uGZ3UtLCgBFQnBeolnJH3zOgJYaZHmQ
Ih3KTrX1XPsewJIYb/5hfEpLXMgFMSNekZ3xWfLkDdgev2Ho9iBDwI8PCsVpeLVeMSeNQ6VLuPTs
yGx8/0PVT2aLBxuWEfabfLo9ssqCJ2n0ZG9g+b7alAaNbWRemtwFe1geMVRuOcJt228kFdE8TUQ4
sa6ov39fsQWe50jPsMIDpldO+3sL5scCcvzx43YyRrYlE2O9WnL6UuyD4IR9XOHu8bL9pxnbAHUY
FGezIn12wP6Ag6WPrDlZSjPb5IFtVBTiqVbuSzypUFF+qRr/p6HmsJHFHCBLRYh0Ydv9Vz1SWZHC
rehxDM1mQKOZ1MclSvrZb8n+NnQq/eTj+1tWEd3xZPcnZ5i5ddSm918TXqphhyoeBIceWTnkYCKK
lxXfYlex5JTPo3UUJeQQq0WuMb2/xXGOqCXB3cEVF1H79RO8KxwZ9kRZ6wE1TTd+TgM4ih2DncZ8
76BDXrGlXI+PC2C3/LpEQsaW9I7EbZeC2lGWeSVZw1CadIH4t8iBv7EkltDUaQ7v2uB9ev+Tk4DA
TpC0n29na4U2+xowywCysqtxY9njoWzYOT7j0Tn4bgnad9NwmXhts/EskZ56BCeQZqrx030cGiNr
IouMLLzTWY/A+CIMiJM6bRD+ur2I4//h2QxPavB3B0ifNDE/bCfBEFv4hQXFWBvmiBYmDzsQNY+Z
ivZtG6X5cmhpMQd39EwLJ9/foii3qZYZdFJRH4afG/lCIECgZ7v6sbkQA+NOgpNE1HwwV2I4KMCU
1XQp+CfUEZBzL9T0WnrQRUDILjhKgQdrH3AJTOQB8XhNES3MB9+SDJqDA1TbyHRHtklUEUdgOYAV
cypMyfEdf4gvyW6XHh8+I478lHAX+kOss4TgJCr2tM4G56oxGWBup12JSQOGHOmYeRqueOTiXr/h
IGasZIF9/W3Ln/cF8+oteI3F2NIMOjicnJ4ELLx8mq1FLDcZI/FqKDKaFFBnBmIHHYOYWrJgxaaM
jXLLqOkRZgqSoWAUmVQ1gdu4+EaEckTafbF1xtZyYb/0wFdeglKdLu3d1TA/tL4nYjbK1sfmWocW
01ipfjvkyzR9/LpTooN8Tni7xaxPqUYR7FR8MKmxqmzfYmaf24tNg0dZOfRSfax9Ft14siwQkCpz
eZcELHmX4FVBiq1aIjC7q3wn5eKTgvJ4SSFxc4DtqoPsxqe+DSAmtgOCzAEs7UcDRkuyieqzryI9
dj3GaL8OBw95B//QiVUPtZ9dQZGbP+u/bB2GYsDGZkC6WSV52WzAWW3Uyq/Kdkw0XZ4WuoB2ufvm
VtA3P/r4ibyU2OTM7GUaXi0dVhL0JFineiJ8ilUmYy/0RbLRRd0X9oOB/6X3TpItgTHdVi7LFB7c
xJvEY/4TNH92h/XQqoPqEnZXW8KGjBtQ4kzcLddybtIDHj6unrASohFa7mQAjWeSSmXg906he4dJ
ic5bl5f2PnGzLk8V4epy+wXG8pcqKbcQLLPA3mfAivdADgEQsBCvkuT7ep4i/eQ+d4PKaK+aOzoO
P1DnfY+ep8BuoAqROBQbos2GzVNIRQF7+rfw7bOvddvcfk2KB+GkVdMdMZJShHFwXmarGQqQhSv9
aRP7WzBL9Dp4Oc6dIwh813aNtjrQsSPDyNAxNR2pfDV9ZxVRhOnKlOqLpEzPtPTXkkiWr1w77byI
McnEKI5DuSygXH6/iUfiGKc3oPnVMkzp9crzABB+Zew/GxZjfFmNh50wWYRYFS7NYOfv5v4FViUV
w/xUwE/GdCm/2q4gaCt4KZRBMtCcsb+18YLhNSpmERdlqxm7UM2EqyeHMLNo7ZcuU7xK4wr6Afyf
Txi4mUw6A4d73y3nwniQOWNlL1DXp20jV9XiDDLjLwHrY/R3ov1ibWpOZO3rdLVR/qkV+oaUlchh
V47pJMWVRBvO5i/YrZLBbo7pw9ot5SIucJ3ts2cIsVfPgrIk7Z6Y0y5uxIsExv23oW0nShdZN9zG
viOoTpGKene2scnjrlyKccmitjNTiCuLUyIKBaSrky74dTewr/TtMsNH/K3y/XbNnN4unwXmIoCd
D1ay3RD78Xmrma/MMO+UGMALZb3S4la+suKMopCzfo5YoLaPddlL2xugda2Bp5fG+GgLxTwiAk9K
CvPsz3geFkXDtPgTGY8XlT9Dv4JJU572nGWarx5pANfePwhKvr99tdWZS2DIN1jo18nnq4JdgdmG
4njsL139Yylk7y2Xmly302dvbF2UxgoCIbhDBoNuJ1vB0tA7s2/JEPphmP7UcoGUFSD24AcOAC4n
udcMNxze1yZ31SDruhOPL7GOZA1P6qyFfpZ4J7+PNFsdLwe0lXuoH8vkfWPCD/QycnL7+peB4e9e
7AHA+9G6fJUpfY91uE1aSW7p5e7RSOD22xnuIO/cadNaWo0Bwn7lRChiJNdyPDkoLvPzmF1uUwiH
8Scx5BuYInMYlZCt6wLPqQDmRlzThlSjnCv5xXXGNr1eBTXxAo3GEhkpWnXC2IApocNSRuJEDuul
6S1wKP5lcA9xuanFkclF+dyPo1jpkaEGCWWd8RvZyrbHfPDGNOq9vhO5m3BfbkFjC4jeGDgnUm52
tuxIgfHqi7GrMck20Wk11wrmghDlKMR6oMD/pjOSO4l/tbcnOWvScELNAkCT3xmUHieXcE2XiJA5
poFHVtfr5nGErda7i6BLJnmfijbAbHQExlAilJw9e58tDulX7nfSC79ZfoeQBrnuCxMfj6WphrH/
WCxoRczqRj+E1UXk9ozH1eMeMdtePMqj280s+RPxRRJ8suHLvWpDzLuNgMbmVb6TL672hahiOdt5
4HX+PGHp137fbLNl7VmXOOT0IZYJTqKian1zoNWf3Mgg69AEvP/CcMq0wP+TuTNijWtbcZVgo+FA
6x98QN6JgJDg6Fo3JwwXljqVzyff9U0gcl2G56cEQPCN82zVxrmcOqmDRXYkJa9xSbiOPW8EIV0Y
JK29LP8PlZnTq6eaYOx0Dyik73dq9Lsi0Bg9kjNEPQnL2w/3hjOGpPLdwBE/V5jXlpgIbEVFWwXd
an447gf8CAIYYWCMR7dz/IyrZOnX90mb2CL3DTCzRcSe03nJqgT3PAeBoidqgBPnRdiUHomtI1Z8
JcXFk0smGHBj4ALuohtGBPbCx1vpfsLlGFc7l2A1g9LrJlfsgG+mNilO99uZy/CC+9XarMbR4p3u
1IqEItJj/lclhJeV3IiWpMJO48oBkLywHQy5tDJyfkk0jvBFaIJShHwsnvPypPNyJ+1WVwVvd453
GhQ3clPVE2QxAJR7hiHURofYUuyyc1d1St9GQmJDPbmYOYQFyH4jiErRFxYDfqXyWIjyxzojeEx+
5CO6NnTOraBccsEX8zdTIs6eRq8OsGG5GyC5R01IZHyDXDo/09bbmlzKgfRfuY+kTS0LgXrf9pgF
z/ctGnfq0DD8abGzjvNYNpg+CL/h9XHBUusiO7QOY24H9xarXZFyLKEK7r8vO0wRAmvgOpzL54e3
WneG67WTKjhK3K8gYKCp6XLr0KNw7U/i7z7395KxQ6sLBqWBLSiBMJDeblr/RjFwYOA98s+5/NcD
hRH9bqUrc6YbGnwlF+c/3wpB+Ac9QO6c46XbBhp1QibiCqtxxJsL9EXQ4aOzH2quIIpNzruJe7g8
17eZvMBjTv0Oeq74JUls5BBue1PLADgZ4omod8l0hajpofEMBnTq65WRHNPiwO+NODliYY7oayxk
E96CQX+TmBrCgSHF/zF26F6nolGtNJgmecyJV6VYW5HJuzKx2UY4pVjSSpCORs5N9PGvzPtFGSQt
ElznDen2fVcAvMETVIVGiXiYiqkSnbGwL5aWR1Gq6r5prIF+NB8zFxOt5UWxOfGlr8CeP0h36rsc
3XtcFARqZ03nc+u14ErOqZD64gpjsN9AtVDvh0Y5EABhr1XzeYz7U4tDFvdJWKF66BKWOfj+JZmr
4aMbQ4cUemI2VwwZEu8FmgSS37MbApaA9THsGpv+z/VNHo6iAMCFtEmElTEojtBokKZkzqyu5TaM
61RBHgUHhOKxOTtzxjJpaanQ+apQmwwoS9r58CxaS2OZKoRvHxw7kmK+wwjBIAhsevM/IpOjZ+uQ
9KV8IEFtJRGOHTWD2TXzEFa7VA/l3OoNNZFDEGAqUHAi+380OtyvVvmKYIVVHxlsToYNViZ9h5KC
vqPOpMkYR+hc7g47A/O7va4Kbg2NkKjxuYlOw7LvFU3e1S8SZ1EFo2bEFiH/78xL9g5aQJdIEb77
g61XiNZp64L3DCqvQwy8nSl8s4Vh+6b6PVo4E1MUgRd1gIF1tOMCaF8acogAZYWVcCj2/H6Lm96N
I0Tsisw/lWFvnvif2kuegOL1aErEWb26julb3Z6Kcf0HbFXwP/I2yN7TfNymuLF6BQRXJz8S7Uzf
nFDRhZVPPhsvpSwlDWpniPufq5jX1bYmPA2RHvIYgT6I2DP1Soo6Hta4QmMZ+ODFnBzEFCfl8iP6
MKfzb/EOp6jp4OsaTtEJTcbNYVwbRZ6mjbGp74BbnFzrKrLdh1pYcD7o+wzxatywwZ+xImSWAY2P
JqXD1opowJ7fx8M3CFaI4U4B0MYr45WdlDmJNCB1Ce75qnulm7Ynwm816acpuB0Te8nST5lJ/2yr
9B4UFk2emhVXo9ZWnC2fS/IYNfGHjEc9CWVnsbDlR+CSsCdfQ0CvNhIopXDu/JUvmlwHzgu8tDDo
ozE18oUw3YNN2qTbD+PsTzjcfBIrgunX2StVd8R45XVdcQ7NZMqt1tvt8w1RV25nGTzLVDXvzz4M
GXnLZC9T/utyfKzK1aVOI22FUeFm/QBpU+DGamVEwqFegEnm4vJ2qI2u4rnHSE5V33vfUSsleNmK
GSYc2HuJEfLhb3tWg9e8WKsAarXDSk0x4G1ttwutfocxXtwZ/Hv7TzfKnlhmYVKyQcAm4BEOXvaR
HTil1xRrQfS5Mhg7UIXzGAvOYWxCvEHmL5Lyk6aCsehLKXKh8iFv0kKUI0qvHPDZOZr7yVc6EqM0
g8zBN0/H1ZasJq+bSWIzVpjexPzSE9dOyjPy3cPYWBI8V0MpBZZY9xKc9UT/SKISCJO6gYbBvKQ1
LlyMHfQzwuDGTyxbwieI1zFqEVcuzRf7JOpA+4srocfkOARg8tDZAzSetjX5xteQjDn4nElNH3+A
3bcuujH1Y4nJ6r186ma3mYlWGeKo2bbce4sSAwKiSfEerdDkO1HdeOi8p/wbJRhMfcRhcHIo1+n/
9YlYsuXjRGoxCtC64MK5CrH/H3Td6plETZ8dA0si9mQt4U+bJvvD/qt9rIU4IVe5w0GvslKlPiwF
SvGJP1cfJmJtPEoYCzpEwqT1S1HZgBM2ZzZJgfNInn9gKOwadqymRpFKQZsymCwXOo5j4gDolv67
P+9Qw9OFkjB6ukS5Tp7ua+pPvTV2/0JKJxqOT0Dp4QRYWfQydb9akJimcqd2AIOA6U3zXfNdLGkJ
wbg6KOjKvh9sK1Bj6KAThQf37kaVNGjfrV9gFec+dh+PC109TIYmbBHSfROzbxuN17cQwCWqeL+I
ZijWJcCfHfOvoZM/kYnPAKEmFgkl/TvXqp5BUzXkJqe+vfvRzdxQHHuCb7zkthFR7KiZm76QhqTp
YEpZMlYsuPCKUNKKMjnxAmb4borVh0tq2Qm4d+KzNNRjHKr5ZJvepNo2WvAgHFNI5gyqOaku6CKG
23dVlVUWpbL3L3kBlq04nrPyEfY6XIX+lwLg272qrbNorX6VrNLMNTiOLw9AqNjCJ+tR1NSRTqFu
qYNanZXW2menAIUKQLY0+GgLRgxO+j+2KTtRW0Bv1Ui/v9rvbk0XFZhfumQfUdSmsgLMFo6VNxZ2
x/FKiJES2qBIJH6zMNg+l6hTVexsd7bM9sktNIvgC17qEourpT1F1fDVJ3cG/AuXuL3bGUCGL8Ox
tTgRurpMxXGJ8h49tlrmKW/5v41xMcqbhXCUFlEEtiFAupgxVzoHYMotPc82lQ1Fx1jw48HntdM0
mJLm4BoI/MlL60rvzH2+3EbUD2n52w0+W5FQLMizgBdn5ZWBB5WRmaCUczys3F/LNk9rBNWPILFp
063iwLlVzJT9VZ89dtKHV2DXUV+bWR6t2I0ZCYel9fmEngNH6Vgo8EL3Y2OkUqFAgu1Y35V3Rxf7
xh+Pp9FliMmrpFw9gkds2dh+CU50VyPa3C1RICOtXX2EFI476IY6ZCP6xFh89121DbR/ilYqg+kD
YFO91NsGLdder8cjyZhZBsGu1UFxT3ffJ4OB5G+ZHmlMb4lXtiyVvPJ8A4/THw4c6g9Y4/Au+mur
csuu/SNJMY61Mvkz+5I1A4KnNC/MVtlS/wD0uLnxxYqVb3FA6J9E16fNeLj0HGsJYu27xBMZE1bV
Rh395fiHQ7ju3Qkt8fhWOLg6r5AlCHs5HNtRz0KAfDxS5pkubSYN///tcYBG0K2OhBfdwiGNyqFY
YuYd/Don5zzCwhV1p/Yk/ntzu44ExfhqIphFgZ9o71MgOOiMtZ0jUsXs6aAduRdPe/s0qGeR3rHW
m4m8S3eJV8+0ab1gzwwjh9wzO2C8RVtwdc4wgscagRR+ycBkRtx/kuX0inHUwhpC1TbrBkuU9pxB
j8ROuY76MYfW4eOkxLD3FsiDngM9FlIhupz9VxcSU9ku3guYw/BlXZXrVxecZpUlcTKrfcSjGa+W
RraRzJmlorBrv3C6ktrN4uUMrZc76MPPtdJDD/pNtXpEsfVYtv8+lu6Nuu7ZGK3c1RVKdyXJoW6L
3HT19mwJ3XL/Xi6DN2wpY5F7ApoANjNewzQz9I9s1i+UhCP/O5ui0bX2VDbhTkWM6NH1mqZoKR++
WJ/JsNvah1BNyy5/tXK213xy4rln2ISEnMYuQAGnWAUky+5jKl2r1zCWt+gWveqiuydsckXGDAif
zD/Nf6uGFpakqRnTUcbOG5AssJ+fqSOcWUeVVSTjDpm6JUONIqLC+aZNkYEbA0ZpX02AcADUBFAK
96as/aubNxesMhaSa7vv4V2oL9FrdwT2KrLJmzg0h5+nSWa/mWQTl4dVTduGUdVTURbLCnz/4ddM
j6n3vXpNUdUiSNLk+Ehy6r+X0yqOoOCgupDQYo2bdvdK1gpJpTvDR2ABjoynRXk9pYu0o0XTKihT
bFcRhQuDoEBmHEwDRnQOnyxLOFDV5cLdIzlrX6wxdf1j8E2sr2XJn+yASpMUXrewwQen1CeGHvAp
p0nXi3d+AwYJ3NmKmxTws8leqbBf1ertbKEhx6Fgo8eYZl3WCKdFOFGCNFXZ/ruwhg3cG1YjyuZg
Wk1+tRm1hEmZJTIuev9mvUpI2HmF3OBbJ6gbfRGG/S/61Zehr0ceh6FYC3d4uw6/Afzu0D/YRHrq
x3SMizmZZ0ZVZRx89VygsWHGLZlQ1yVuMJFfCXj7D9naWKAxYOjb2leA+XmksuIs5XSHdOsin6lq
y/nfLaciI2nfJ99L3hOVfeJ3W2lHCrInuafoERJPt4TfBMQ6HAzW+EG56EIebm7y7J2cBecj+6cP
IfU6bFq/9qmF1VobhwJaSMo8Gt3xcfmo/q0Bytb4MX3cyEp8A+jYaSiCHPbQ4NyVfE4iLriGl9pE
mXPMU4JHRXslSvwCg70mGwTdWqhKQGLoXs3rcETsbb6nSdjzJsI1AjB0gk8QssJacmKj49OSLvDs
g/bIvHzvUn/ZPRce4LP/mPjIqqnYDZM4Dr2OfD+CFgNGeh7v2aqtGjHwYM20w1L1E0hUVJdeKZm1
c5T68L+n1lZXwjBb/YTQbylMNhwcCKYuqJpX/fPOoDDZ42K4hSVyFL1b/zGFvaFKfDoLQ2ZEMEBv
OQjE7oaAia6syW+VFhzzLj+u4oAyAGfSqaU/tzNjPTNi2fkNbzcIyQASzlYu9O55YQCV5aUr3hlv
Jb8uNXf85dR+A3dhprl1smQWVpT6EWubph/t5IpcTepDBJ/p5Ij7l7BNs6bybLe4yIcP954mZVkB
azhVoeud0Uz7sO+IykkMq3PSqTo5hqByJyP6Ps8rpgZF+f4kKzbav7JDrhWWao61mEsfK8jc3ib0
mqkcR6YphPHiBrVBHXF0enwSq76rRXku2shm3zklicxGCRK/BXgPVlsN6l+7CNp/OF4bVwREG4vm
/Qvu+C6m8z+I9donWZG76VvJSr8eBQHbLRzzgonWjEkYFAkC6oBkyyrp837P5jD2iEtEjx7F8GRI
qKmv333hETX3zrHIrMGdnx2ctOwoQO9lA7GxJiKWu7B1fBJLwSxlQifo5vA6OCmlHV9DhbpfWHi4
vxpgVHbj85fBBH7f3X5yyay0ew7Mn+l7oATqGTzue99OoDwYtXX7lIP9kwb+NweMPhMJMX1g7/5m
kAS1ZKv4ALjYsppJ760mIVpJjkGojtd0vdFCq/Je5i2tcN0Tj2cvQbqDlO0KmyD38D3kvvXsAWev
G7sjerirj3GZbzOTYl9UF2Hzy1HuGo6qO2p18ZRl8qWPLsEZgxKeOZ9QlVWgm5FJPNgqfQcQEIDG
IchBHyjKuUf77gmGvoWr6QPQiiKl21CGS8mrStXMGCwsscMkLfWO/yztGXVlR2GasljPwnWrbMoF
eh2JC+gZClPeS+oPYiwi5o+rHH6635TmiznI9gqwXWg7czSG2liqmL1S/gn+KLHak+l1tmyM+iRe
pWxQGnrTIQNUsa1kvaknQfSfDb0H1RyvLgTpj/YdCC6ej7wDG1pS6GbpV1GECVpozGSKWn9L/I9x
aA6xvTcMwcGQZJ2d4bRcHQHf7AtC/l+jbEZjhxjV/UubULjkI/OP96pU0tU/E3U1UBa4CVPqwXem
v3nMK1e4kMyH/FZ5Q5g1X2hs/OEOkaBw5/Rvg1LaBrKrUZT+ksocpzWXjJc5uEpK9mk4SxQ7vppQ
1mCgkW+OWrBuX01feZaqr1fza9wQK+JyKoFCCK5sEK7t9D0Xi/g0OLFfZK6CVEWiVp5/zsy5NfWi
+qedHOXDlxxo4z1jF+2vnOamr5yD5WPc0r0LrgtFsvGm8dZhxKA0PwU41PJCk73rBDghN7YI2U2M
/KUE4bV+y+Wkxv4Ascge3o9xFOzLLpErWKK+ErqD/CUJ1vS2e76sw+87m/Gu5db071HIvd//s0Yq
cQzNAZVGKwB6/oDu6HRyP4vFcR+3Qbe3mfUTA2VpY+gMtTCJh38LWuJxl2uAPS76lHak0IKlnYkr
Q6YOAekltmX7p63q/Mtlj4ZMctitikZmVOu1M7YAq9M52CgB2hiAp6aBz8uCujDj5lFEc8I/Z14q
zFTiTU4imH9zq8106BF48QeAF0/N7WbcLLOh7pFMBbASvlQykRgn42RkQiJceUfDAWfz0aUEJjC2
NSCtoJf5FTzeAraVq2L9/CnCDlNBZJGNhZxcTv2LQrJ29tGeWokuI98nfqjdCbVYaA8YtcHSRs80
erin1vpicjemOPCrmhnbFenrwKl2aq4j8wnIniWpVymaXEyf+0RwSMvUQ1iRBC3pgHAW4s3MnJr9
oOsHtokQsczXEBG2MdNy3iHMn5TUBpZhYe3KIpX4hhFgPkmTPZoehlBLdiQ6dRg2al3AbBoB/8y7
/NPrg1ZnsiU6I5tp/1MZLhKL0VUX0ajQ9JN5cCMWekBP28VwEqExtCUZpZ7g1P2YvH7sTIdVAM2g
OWl+olWlfLnuH4WNno3TtQYbBH6oGDXQqvcEnKt49JLCwqfx7MtstnZ9MtiW3AsruQPMCNMG5VFc
YTS0y9ajggWJl647kIeJqrsGEerErgowjF7ywe4M+7mBZTqvxzqmvU3wx1obfZmwkw37rLtkSXGp
FHVeUFaJPdIdFynCpuoD6dajmtG8t5el1BfS/B21B7GIZ0osPtwGb6A6h38iDrfH8E8wE7e3jxAy
iD1Yb8GsgRZJCIeu4z8EsgAa3Fs3Q7TbN9+sWX0LbCwGAkBZvOJ2d7Q4WRRMeDfR8OjkEQIt+43G
biVI2pKwfIuZenjyx/bhjhXkigGB3Lf8ZYvfYjSo76vebjTqwBG30U3bcqUz6Knmcqby+qjd8yr7
QkkaGdRhDkQuquhn0OEt3if0qB8A0pCiKik0m0bPx2PNUT2y2+92n5IdBkTFFCc0vSEILdcijfuj
KMWaGKm6rR82OfX0EtiEZ5euO9A7CcupDzER/pSylMN00PJzblc9OguXVYwLpYWK8X0P2aDOVhqy
deB/jnGexd2B6Em83coQSeN3omrsuT572XBWE7S4qx7DOZu6oobhbkJwS0HEIkCqHiTHZvW7E6/F
OTwIoY3MD9UkRkQb67M51bxJVkz2D2d6mECPlJ8ICp1pej+HGWLRDc0GW5IN/VaG8zQjMDpyIbhr
FrDuncLP4WiTxW5A8VGbFJig7QBhLMiy9ZP7EtrEXNdA7aIeQQr7xhkIL4FxYiTFtxSr3I+AeqkD
WQGpTpMf7sgwB78TVK18RqVXMUn+5snup/YRl2ERn+ZZneGDLFyAJEmnUELePRj+JMcgIy9Imknc
GlVUMR2OLWech/iaisFKZr5K9Eo2f4mcmn/yzk9FxcFMan2T9sAB4np5/Bs362oulRB3EnNYjT7U
of02QUwr+UXUbXJcw/uUxakIliBTOoWxZnfMYgiza1UQwkOzNGLjiAizjZ+3gBzJTm0t1ofwrdhy
P3VpTLAA5UuQRatOaRa4LD+7c7wUSrX96k7XF5p05zQz76Y6/bbZhoS3++6AQ78/vXPcU49Gb+pL
FGTQQcMg7Zd/XKi30RCS9X2MfM0ZrrMp2jYcqbZl2YsJPsx64MWXDyMUnp6uqQRg0sDKZV+o7BUR
RbuvKKePXQ1tRYO95z507FTe101/e4EYCA9ljaiMC5eHgWu5fdN93flZ/zP7tpS2fnsxz5KYb1/N
je9tprBPREvx7YyJ9GHXkIsDZx0Po7MLI2BDKsCjYlcILHY3Kaxi/cXtG5Km736odTui/N3zDV5M
fv6h86x1xr3f6zN6di/lIw1uK0oe1JJ/DwrLU4EPONz+poPBlX1A2Qg+kIs4TIOh0c0RqZeszwVh
yZGsutsvxs2fOLKfnh5CUaGxwF3aHNz8dMozUeDXqlTnoXq4uAtF09mOHY8XBRx+skIJu1jDrLRQ
lSXJZkrK3pI9PiZ/BU1Mo8gctW2KXx4GlNfrfpEubUctbnrS5u4ame+DJvzLE+kgASZnm0wlgQXm
fBzzfuaVt1bEdyjXN7bhJJCGgzvV82Jmklj8xi/OxwQEHeDY2DMpBxz/0FjPTrAFJFtw+O/g6dpQ
4dp5KPMmzGqbqfCuMnxJmC79WZTAqiFZ2MR5bZTbpqJG/C3rD3D+vKpyENMrTpyxI7U+XIXD4oqj
Vs4xmz1wzw8uXSN9wjQEt7Qrpt8ldEsD5lLNCIbPqFArorwa7KbyDQ7TNlUO+sG2EM5/UZvqmrYS
yyygmhzV5U/9I0hBVbQoqc/jViA4zwOz4gjpiDY4wp/7G1DtTW1SnwPUN/btnFtc5Ujw/ZFfQs/u
U+hGQIAuII3Cs8uE1fkobWs3PrhaZAPule2cWVVSVC6YtTYZwupE/jQbhsEEKas+2jK3YRQuewUU
x0Jp/v+iu9xs1I+AjYO9Ix3ZaF1a8Mz7jRnhGmQCAalrTgvsg+gmayAqV1/akeo8OjEPDg8L/ckD
Mlook6de8nl9psnrVENMiWi5SSgqBvfqQyC+y6Z7W4JH+QS/tE8uif0g2R6cXvBKCVsi9EmJpsua
MYb+4NSu1UKVgwsNerWL/hs0hGa52zFnY0CTFcwb4YK+6BN1ulMGPA5/lUQLYD3sC9ouUJelHGSs
2hySujri+SJA7eAJHnh81YkITeMj7ugxbtRdxhgQEOq9fMzipZ/mFYYqzle3g6XXOateZsRmuJCE
4Woa2+YWUPH69VCKfukKwGrnjN+fyI1jlun9J5SV+q+oiMKErQgQWdXMrUivqUNjNCM7/TTv2v1u
xCw2LSBAA0gDvM+WwqkkBREFLuCn4bd5JSbeRtRHnY8/5Z7aM5VhHVTNhUnmxuf+K6kBc+OnEovr
Ghg0lnTr4k0/diokav+90ftrBj1NYInhwRenVFsJS9CbR6o3+G7spIjdQKBwyjIhASqXVKvxpLko
LQNcz4Wex1ZDmF1RGEL5yimjEeXNr248AxPqgmhyGUqEORoCJT2Up0+xANFnWNk6NXZbxbDTr6qM
x8XtwTEBLBAN6sendsDt6HTEXzTTFQ7Sozx+bAweaZla6utBkCAkNOGR8KAIk9wPlAu5qG2ZjKeK
q8wO/Zy136VbS8P+pdrxMCYV66f4H6pzTSRZ1LIKVDX/hfycY1ZpP0b6DTFCrxJ2y4fG2TsBfiTE
gU/UhsFbRuKEZmj87oUs87Fgd/2ctz576kgn4z6SfXGcIgJzyAtoes39Iz7fu3ExRwy+QMycIDnN
DTMybfg91ePDRv7uEcw6/1Fiw7EhImQ1quXV6FeIVNuiEohWo4IPUeZDAS0T8j0Pj+HEZJTTEjza
U3VPJf4tSm8PYin3m1RQmJ7kxiR9ccO8wiZ36zRGqe9FPBXLXIxCBNYUrkw0BqEa4kZd/DZPN/AH
Tmjjxq99rSFB6aMl2swiXZXTuZb8DEdpkAG8BwDaOTKCeQGlHOW4hrkQHgl3DgJMtKolBOknY9rq
KnX8vVLkH3Oxvh0wMHtLvWlPSHf8p9yVqBFdsrjDp2k6NEQ8CqJwVEhYeha+wVoRsJKAsFzUc0/a
VSXgaY0eolIi/ra405ilItdOnb5kBPsi5KKI7K/KKvqf5GRnvTLQc2nQFKtFjkzuUvXE/XLShdNB
yPa4IE5L/7jK6nIyS7rVUnK7ASfnsPk8TNeIPPEnRvbozkXR/2C5U8cZGEaWpLgeQx05faCQE8OX
LrmIezrXU7+p4LN+3GYNY5xDHsQqc8ileZV440m15b3OwMGmBaognmOB7dfWpRkJfswZBkAXoQuF
TeWE5/zKXu2UKFs5Ff9o6x6zWccg+hZPdRwqDot9WTeAz+NAcaoUo7vFDdciqKqNB/fWPWPHSNOG
hDlG3jRi9K+T/x7hyUQFkoigouVKe2dzkpYprWuAKg8aChvggcCZ694lkK5llJXC19J3+GLMuPLW
HpEZn0gDXrJLTDi0K0c+wQm8/fkWrgEIQ63nAF+276a4oQFJkPoQTs0c5uQF54c625MPw0Tu7M0S
1En2sCddSYPd4Ne4lQKSiEaFJp9WVw/enpxm+Ag6pjYNGWXHl1htZVnqx1zVjj9xUZuzu743a/s/
cJpywKNiy/S+lNJufPCzE2n0YC3sik1CSslSUQi4yfeNqxRA+iHXf3gxO2NkGYT/rA+bxov3b4d+
kfYVMs01GD9gk9K/mavN9w8L0ia2fTSGkJ9n1hS30yUdi3WIRpNxfbtFCdZe/2la/h7i8yS7OzEG
0/HfPoJ6s3R4iVSiRPFdjraBooPisgoSRCa+sadR0hsE7tE2Jn9mvhLg2bunPNL6O5Pp68kLcJYA
5909O8lUJ2JSuqKdJTdrOWhklSUNw9n+F+ytHaik/LvWINHQOLof53mskGcWESYlZuV3hPUVJN/W
E/YXtKRH8dgzTDkw9pP6yLiBILE40lIlFMZJuN2SLlCL8V6Xa+GULzsaa9o2R/A5PrZuEkxN0WXt
nmn8wshL32fgS4R2pbr4Y7HEDIJLj1GWAu+PJvN1D6Ad1DIDj9xtseZtOxg+eAKM81+KHL95OcTJ
lvYidNVjnbyc3U03hIEPeH6A38Pet6j1wHcUxWobCOaGfXpT+oWhGHSdJfw8atk+cDx3yVBiS55B
GlHYWoZ9YWjK79+dA5y47xMugsR+kVUVblhrgBGaM0bhC62/OzdbzXZuFq01WTBccbPmfikPXhpZ
Fys2paWtr14V/RVsxJbc4p/3Gf5ewz69kPcNWpsCb4bqDx+Ipm+9INnAWQa+YwreuParHc4e6qsW
Ql1tceraqEUkNlgKMfHmSsMV23mr4Bjd/MtuXBb+bT2cwSGU67WLLrjq2CAjUnbUBeVCkvVF/AC2
L8Cu5bmm69gcRkOOzLwWt+VP+0muIODoURewGjbfdf8qylj//rjw/i2jOKAMUrmaFMmZKK3K/yE3
ON8mH2kxeDATXJgiz2jzygJFErc9Bt4lK2ccouNlpDa6fWSBaZKoUNClM4V5oPZl01/33tRWpSNB
FZ6veHYTEITjIP+4IMl+dZ+N3CrbCmkkuSdSNqZXjsrw+Y0oXkfzRjjpHSlDMEKesUdGdzFeoGWl
jKg/f1t7pWJVHYAJlj+9N6L3cwTQ4JNmba5gSASgbQLdRY53h6sSPJ7AiuI95IL2j2iQ4K0AdLSb
88xw+mtG5xG+wKgQTXllHYj1+RvDeeNjYy8CsnB5e29AHsv7NGJda9TQSg8RPLz6jMjGVymI+lg4
T4vP1EiPmIkB9wZ3qFj5eQnp7r+NvsQYUZPbvZlfLcvOKxDjoBl8MbuJ0oPnVRyzKAxrPExdXsRO
uDB3RBIFXQmfGaURI3x22+pDjnI/GXqDT/Fu81D9wn+F7KzEt/lsy2LEa6dAmHmBmOVsaPcjZXRd
3rZGl8rYAj/jLaFXF4pC3KwJIOAaCM4+mlhazzp3bta3r+rpRyLEebvRoYRAVVhWaBNBrD+/pg8Z
6RZefUZM4uAD7wNMaKXCX/Yfk5gxnOr7nrEyCtO6UnYKRd6xMFfyp1GfIVKqpQ1nGZ7XLtNkrz6O
POPlKQlGAQv+PQ4IOVSoKi6csZww2oMLUtqKyTz8M3axh617vxZEeYQCpuCPnCo8/JRYteynb4c8
rQMJHujnyXIbtzFz+Yd/m26zRgdGoxRrswD9wkHJ7tDgQzrGeupOMdp0XD7GSbFpCNaxt50RWjfY
W2bjdpXaTy7l6IxqnSt7SNGLIoMB/6o57zXSlAZM5DIPMpv7CevxwjIsHhnT8jKbyFqC/XdTXun4
WGBkV3m96+g8MbBsrSPtSPPuJNkq4qN+e8MZds7HXbq7HIFoxR0YFFfgda3PAXZ6c67BfrIZZ4F+
rEnCMfYOJyZRrapU/tpZZegARji5UqWvSYdWB6+17onShag3uZOTgCt5+hAKg2Kr9LPsVPeSzEOE
50WKnjdvoE2l/RuuRuSO1Slhe9GmMsQhkAQHTn0PYoG+kn/8luP/uqXE028vS2YLOh4Hu0+qibq2
Bev62xbyXNhi0rBbUXFVXx20dSek6yT+IxZC1MaBe7U/Bgvw6qMQTpMKonNdOseHpuoPvSK0jpGv
uYy6/HNZpqUm2UGwC0a90zVHsKCA/ObYokdbIqesj4YBKKAR1WHK4NpYmljtX3nklTfNJnsc7ezo
AMD6lN9whgw/Xp4J+WUuVzJeIy+XmdeEl7m3sZ4IfrlGtFoUSWQN4LoEtseZgaGk4xH83G9fR2Cq
cffJjpI4KeesUuOt9ha/f3oDsvahRip4ymhXfpcgnn+7+htp2ppcpbFr1l1gEpUkt52gwjFJX7S3
5YBy1jKLVLsSVff6iWi2aC6UMf1NsEE6Me9dBUShYnhpM6xE51TBzoZ1GR0YhjIWcKPxYqVlVHZG
Z/QG8AMXFD7fSFys6uXq/CQFGmsR1z70/K8Z0MuLQOQjyi8qTjjEmAW0skgXMDZdSS2RJK9iZC/P
oIDy13yUsFOeopS+GTcXGCxm7+MOONP3d45faHF2UGgG3LxxkhDEKBXUQWRcynE+iPRW1N9ZDFqc
ajExmljTJAjjDKRn/On0DjZX2P7dmZGdELbLMuI0mhlUxpp1LEkbVUCycW2+ZaKunx85Dj4cTv7i
rnIheKd9hIv4+Qv8NkZjJOUahDKLeZt57E4im+vuODAxtU0xpb7oyGnUzmZPXkjwIZ4fBI2dJy6Q
/T9jaDUrtJPdkKni1PuAa9GFDATsUSmWTwVBqVLNQbs3UtybVM4WElVYwDB3OB55qi/9GWgYYx5Z
tF9I9x5r8908hdTQ9J5KNbbI3m/ZfUQPPoXh0a5j2sTrVXVwU3iC5h3So5TWVgbuT7rcaae5CEvY
8TFmdUQjYq0lcXNGKtSZ2ZsF5j9T61EnPl4XCRWv+kL7JV6PYOuVQg81/00bwZWErDmg7NH0oBnJ
ljzTWaQB7W+xKPhlhQc/AR/7ROpGvlxDPU9vgYwMpzmys0VYXzNdr5hZXgWwWaduOqh5rwh6tl+3
e2c4OJYUlM5gMdYDwgpLl8+tzZU7aFEJFI0QEM9iLwYombOwD5JUABkGu5otam5B6Yxi7v3tZ/qA
hJ5qqmPbY0txfS8hH98rvsZ4vHSiiSF/R0VzuoojeRg/DZwcYp1mDOLlFN81wn/OA2K+gjvhpR+M
MnqNVZoy+0LTvf52uMtsGB2QRj6EfXZzUsNdjEIJwVNJyCga0cLzDyzw6d3haINu9cSOAvIqAn3X
SqJ+LsKwOB6qBBqCG3J9bWh+bTmEFqVjohkCOoEqdCyUR/BOGlI2EYo3EmuSaNsA28BthBnzJRyb
dW+Anc1JlmfbPiHYOwzF2e4ROjz5emRVqgwX0Yu6XbS6Ds1Xm3dMjHCb0UAfQIprEDnl2Nbulxg5
UF+IB9/431vQOmtUnTwAJUi6P9uSEPSsDXmP8RfNM1P92Zg2GQd7hw5Yoo1Cd2P/65lsna6hd9i4
wi95i9WsufUCz/ZOdWk8bf1jBNDU/QH5mL0WJfkA6NYhaJLO1ubUCUanftNLGqzopeeAeQEHN2bB
f0umIdAcBJgpplfMcuT5jwvLecu2VaohsdyGV6TTYMY1v1roOFjzojYvU62BG3UdmJ43FTp0PzPM
LPEtgksGlzwmCUFadGfrFCCi4PazhWbkytQguPOl30G7lpV79NSles0Kp89BUVPMqJ7s9Q8NjwwK
XpDG5S83jVVrbMujZEkY0j2q9jCIHJdQXTfNmoLsjschDwaeWP89lF9fEC3DPphzHzo1yhYTtIpC
t9TghS11iZa/n+IbUBgZMBGwa25OvYJGZci7wgIUiTaPC/LranWcsdG5BgHu3YMztZlW5mdbd2GV
MfIKHuAPcayLQvwGoyYkxRrZHovhIYSRAZZS6CaEHVj5T5OuNepceOeyBq73n/MA5waiYGn8XgxV
Vjf6myDN9Ule6TVcU1UtepGNTy7JxoDnAdi26CC/CXeJUhn683rfnfYHmrBbs6vOe+S1V0ObRbmK
y80sJ+RSstQB4AvPAAhW54NL03LCQxVIQ4/qyMA/lGGtjMRJBejrBIoF4lBqPpTsBO2OYYDfn68Z
zQfvPP36caffxcMuP/loDUZTUfv1adUzIrow1ARoKn+L4XbaxUc02qLN7T9QfhMnaT0ESNSYGk4L
dKddHGxRkwehZybgSOzGL1eye2gS9g7Ew5bmfrqGZjSPYZ3pVlLp6LWisUyszLrQzznBpQ5XxI4R
s/X0UbAIMHKwo0cRDA2ORLOoKJ2kYyU/zMdfqqWlv6PglPw29ODqK4nr449OZJkeOtX9+5hhybvH
FbPnuieFRsJPg73F0HUPs9x8zh0PrdVOpVsoX1XkVft2k2ixCwIp8MbQ6qKlydNKyOWv/NIdQxgA
AwhetwIaJPY/rdNMDe6+jcWhjdMQsKMLED1BOvELRnPzpJbNBFuy85vjp6YLvrNEBqS149klAqsH
NNTyT+IcWWAy1GdsKwoCkxqpGlM1wmjRAjLlwH4pLdlpT06/ZpbZZAIn+PcEkINqvVZWBniYluqE
Qp6XbYt/fd/WJhZtt6Lp1eSWsplXBGRiJ5vjS7CW235zGjpYO+bSXMxdQeVuCytJ/2j6rnFOPcNU
3E4D73brpa0PYx0d0iEQvGnwVcnecnbQj21lYt+c5Od59tuXn5BmVWVR43nlQ11sFcgRs2zkX/9n
td7SgW6iNJ0jpnfnh1dbtoGn2s8vdIG2OKIFiSd5B9UUCJrmI3HcLm11fAkCCw2jjyNd5wbAg3TT
uHL9pEemNxH5kSB+/30QIW7mdz9ZRAOxdj2TZaN/X6pCQI6Jv2pTNOe/4NyI9m/9V0tVRstmQ1Zy
RJp3p3DJM0GhCxC4xXxSoEdRJKdWLNGxVUqBegBWTcFq5EesxNxbcSX7+jhZcEYrtoaSx9wPB0cJ
cMW7o3RW2XPuPGOd6i9xgvcOZbq50UYksMGuOlyXK7JYaKE0AmThP5dIsTMR8z/W+wZX4/i4dUVZ
I0MqPWCKokcGCR36VvQdrY3St4Wxj6Po2SOu7/WRlp00I2fxOFoY/O8A0JPjBPsqrg/WaCAjRQ1t
ijOWBf8B9tE+oAxLYvceQI1LeLN13TEeDyZOALYfUGYH8cWiEDkues95ALsTRXdGAFnYPjeyGJUK
1cG3czFpCmDzkYM+F8ZaBkNl3Z6n1/mQnlTdZTtapzIcwWVtCobEHWQt/nY9NpedXwdOfw60Qn4Y
OVX86Uht0DwdiVgQJTrpgQjNXcUur/jWBG2iaSPcw5sY/WSKln911NweMj5bukgyERelTw1xbkrW
sP8wFN4Z+IirNT9FwEvgsdaTTgE7vdL3LfcLWZ2XSG2RiZ5AAG/yD61OJTYIV4O7TrYp+Vb2cbMV
GBDNg5VICdAukxmKXA+HNe5ykjYnNMgyka+hXwL1amOqdK9xrO79CyIpOiuIWZF6q28bSLn2iYbK
ZZyfnlMAAkGPmOHe8/IamTlqqo/9X5jkOMtUw4C+qlLQcZbCiupPq7jB3jvLiqZutwLvGQSh9mK/
AWxOxP4Mu+GlWYzBezwZ1LY8dwmsqyUl99rheOfoK8wNK4rr+iwu1xgWM9yFfFIXus+Bm3ot8mAm
oFZCy4LkL6p6hvZkx03LS/X7hNCjj5GjskBvAnyWYJyrLzQCzq+4Kqq2edmzil+QcOpCsSNmDB7B
83U8YdX1EVCGjbukK2KkQnMgoeALiq81xoA8wr3B64e9CdrcoWbyBipJN7/6l0qf7uAncHC0gl0o
UzO4+3kl+BOS4oyE3RLQz2sI+3E8gy3nwRuN64dozDgDw0mTyP0Z2Drv6WxCgtiT4CGtIt/XWhTl
r2WAybEnAs6x9dFJbF+CPBAJuBlP6GsAKuqRXZoOMtipt/WznSwrG5paMd0IuwbHdGWM5M8D2iPn
BWAacGD0aVplrIgAXdVpcAfjo7iNNvuQq3mm61mvlgEGSDvC5sUFgC9JY+WyFR7KRVTvQF2dp1y7
CdOgNq0TgXQtc2eF1wOWGZLt5xK9/mX6/S2rB8ffUCwBZ7ydiJz1u/LNEIoL+U7f9B7t+eITmz1T
v3TfLEBAgWLSno03X1It5S9b/KsiGF0Ov/E0klNRVqJUllpIJvDACd19xLRk5NIuSlmWnp/Aojcf
yHashO4h+oEJX2dPfxe/Lzi5HYQap0fz8Mr8fAeR/u2PjQwjnJow5zg7H1aSJtS+wRBQVzvpBuyc
vxF9eOPpCk6MV1D/UCg83scbdYjjT0OQJmNuNnokICyRe2frYYNKRIlsjNBdZ4PN6VdEXWKxQACY
L3RWwI6n/QEDiB1d7verA+W/iaFeal2FS3lGFoaolpqOrWV1dzTosFQh9uMdkmC45FJzI19ACn8Y
yj5ypowlf6pncVkZN/TUra08TxcEk7zzefH/nqS7ESc6hTUuQZIx3qJ7HqAuGzR8h0mFI3ORJvf5
g22m2n1BTW+1ZLrKxbWS+d66W4t9z0IytG45ydKSMsn4yFA7hHwGSwY2wqh29ns0w6Yw+9POD4fc
JsdL+Kxv4/lRMyjKL6vFRTfM+E15uc1u5oqN9aRlowFmf5wT1QwBozmlagp0LRtcsjrAMyj9ZZ7Q
gRFsXTW6/AX7wwLZ7mN63LOCdmi20r/L2M6sxO/C2/fq8oOLxh8sxyc4Ypo8JT2hM4FACD1R8FFt
8D/uXD1zUYcfhqMqw5hP3FQuSQ+sw5gJEaOqdnLvl9u8qS51ksQiyqp6ieIy++/qMqXpi/zgfXz9
bkdknaMNcXQGjZCNup4CqwaQBDSdWqsnLxtBeoS/YcQGHkXycL8Azh+ZCHrt+gAVsa320WalGETt
wDciWuW3jFira8USmJi3l96VYhwzjhpXS8vZfmP0FzR+YNTDoMhsHTcNH9sGLJ+s36sw+vNv5ykz
wgGujBxvSi6MjQ/S9OMm+fl4z99L+xaWxlJ3GzUQEVy18qEtJHpQCFXAoCv61Cn2BKi1Mzbijtid
3k1aIH9OCLl++hQTyKBri2TzXgfCd/SIjOm3kiizhjStuzQqJDFFOn7xgujtZ5IRlhx8Tg8k2uex
OgVAD2GOHJOCBj6w7hcgrlcZln4WTmI76hsztpbjgjt0NS5t+MRRmUjHPfBOFDGVx470u55/nHSa
2IQK0vOtwmh9zjPdXQB+KC1/xivOP77nOy8wZM0+ptmZ8ESSKSNqHf4Z4PismrlvBaAklVZFRbW1
pyVlOJ+svKaBOteKO5qag173Z0Fp2d47VXN3QuYsqZUk7G9HQAtZ+fCTRdaLze3wiyRT9SE8EAlF
sAAec2ujP1Jq1i3KHqhOQ7dogrktTQ7NOu1jOojN8kYM+xnJoSRnhqNxVvTv07J28RZkfosm87YW
Kev1V/vbPyA3kxzm0uP2C7x5zk+JwaZdh61G7Il+TPLTM+T/a/LkK5A3dfiftMWDc3JjTC/OD6Z5
SHCKWhjOc6iePGT8QDdFimUKUFaxapIHWR4bufiCvKQ7meslqVWJ7wmAMavX9sE4cTNTfXgFADUw
W4MBIGvgg4camyBz/IIQ+1tD1BiYmRPX85WWMEy0dU8U1HmOtYkGbhpnEWGKfnVY9kHoVUyk/bf0
6X9A6bHN8QItYzjPuhyQ+7wQ5w7IR6H0ZKdJ+AQzw0kAOBbuR3W9jdICVL2npQieNTJkFp7i74Yq
wlEbNoGOPEqMLrZ5PCs5OS1Nmz8kTvWNziR9931A7TYQVnCj47cwQbGs4kEa4qhyepeH2nDWY2nY
AdQxXHT7bPqgHJsnbx3Gyt8KEd+29OnWVYF5tgS/oC+K9kUDbuqC7ebezpeQiMuUQdVImKIj+HmS
KOLSZ2sF6jmk8HkY3ZCPDJHZB37m9p3bA+fYwUY6EBF0MPCQNBrhhzxzV8F0Xatgz9iKfbxzOjzz
fvSo+ToBb2qevGdEBxCfEtgRGtl2vdO3SCigkbnmZRuNgISpir6ddJFzvAKPf42ADb1TDedO3hU/
T4hbHwHF/8IMRkXccaeYlcIYLnj214kd9/mrKewEtILsOZezdhhBLbr5cfjRZ9j/WGnic3JvWEys
qdGDtnHShXOH7L7EBZD9DkB5067e4xBtd5K6B1ry88HHlQ6MjT3Hv562vovfRaZbAoNXYHrpwE/X
h2TPh99+ldpmOhwupcQIUt0sqVYeF+Z1NESw4MmRjPKOvYiGhdemL35Sg69anV+e98n8FjjRVRw4
XtXcPjErZPPImy54BGLgImhkcdWJBNmcAKSCpsuL6lKwfFKKNdeOERIkCMrMAcox9c9KQUK703Ez
dvRmq6cSzMgp8RQap4S5A2ulqi9pheR/NsaYjuO1ViOVibLGre3zeuO7wXT7c4QbBxZEpCHKhlWq
M6jc68+kSrC09iGH+APy8pDmglq62lZrYJmvvp5uubG3D5Ql5b3rqfDxCpRLeQFgAdbSoQHR8g45
mcCgmCMxHwMDcKv8bx5xg3QVJaCN2sqSoTPI7J2r21e0AX4xqqCmKLSOlzQKyHyu8AjJq6AB9wfB
psXqmTE3uUek/QaSHiM+m9hudaQgZfEeT8PRMhaJezLqU0PeKrBDXF9vagVJGvQ3wP5Om2mC98Ck
t0hTS+BIZv5x4V8hX/KjEz4MY9a/H6vBm06jzkYM4g+bV6CBKnJmvFnlc3VQk24Str1b34afEqXH
+G9vw+Z8ohKyM5uqiIIBM7TX31YMkpT1b5Stgvs+DlQW0uX5QlTrw4dYwxsfn05opu4lFuDWPfrx
iHBV9JjIQmIl66y/Hc+Wp9Ot5WDdMNJHnYxHyHFw7KNsduEG260Y8eAHxVjLXqlOW9pj98Qdl8D7
8GbKmUIr3Zhlwdcgf4iTNph9rSzcxUa+ulNL1y8xXKFKXicJW+Uj973tGSahIJ9TnZe0NdtdPHk1
q+5p/20FCzyDn7Wl5yvauMeNiS6VuYK8SwyRnrEoJRKF8a41+sedXpTAqqRYLSntmzAsET6pIx3k
j9ZjqEuKZVvUJPnGWIHlTsDkiBkcTdWp9jHKtjDkmR5V3cj7n60pTMyx3Hy7YDWeu7IyFFzrxHHB
8HzOBEmbT6lfmkTCGnPU9sgIazNJ+XDnVksx4DeAHs4gdsfDo45wc/O+u/46L5snvrVgSbGy+7ad
EGbBKvfKpJAoTpK5CWoUxexoYPk1xSqJWdFqtn5U2qTIIrUruMkwRYEj+BegEht00NCjV2XqdXLu
78YN+BdAJN/PFcTgusY0aQiN78YIdGhm3v8PuGNmLYrQTM4OKEKFSkoL/aiX+C1nNTsDr5MpxzXu
LGxV86l96M4yWlvnR4tJg4paSyx8HYz+KmG1y8PV/471PqMWUikveWL8vvccyLj+l4iaYv9MsUFU
eQyJF+oVhSOFVluDKFl6Jra/UE2m6WK/gfJ0QJxB8LnzukBmPMKSvnMlMwd7SwDV+AhufY12VmBA
mCjMzY1zpCsdnG1puUnKXiM7jTQ/1gzh+okXUXMaOrE4rogEZh/fW1m9+oYzqP99vwyt9N2Ib5M6
yrFqnUpAv+9iXYaORbHlLc4PtP6aPKxEzOIiNFerJQmNzZCffBYZHNLPm3COeZlMUCY5PRtFFC07
feUOG72mQ1m/ml/XsgChU340gVLW0OQZTb8/gAYa93azwZLgvCAs98JpCiuQSNZCbVrz4TUL4026
H8F47cT2A3/Oo3wm1VBk4APNKVDhd/e40gHVefnWmslJdvMDknXVVwqQzKGfZmsgDHtTydu9sMgT
5b3DNct8gVTqiVR80mmu7jATSZaHSzyVtdRY7FEmnxwjRndO4z5LYnCcWBVB6uA7Q39NmxY/8XnU
x5KZ0Xkmp8QUIVOukV2WXbcM6qc/wJdvKPdQscCPGb6TNllh7u/YYQS+52BXiaTx8M+irfHMbO9Y
mTjQ/y1GwBH5aubDFjlvO5w/OuGEmVToQPUPXAwD6gF8ljcpfvwnY0jt9BC0QyacPzu8WydqykBw
f1e9MKTAPSatUf8tCrPjNoamKYxylejc9tHpz2YZOweSR6krHZSBqFwkAghFwZFDcN5BM0O/QB2+
h0JRZqoMsaPpmsHEeHD/4NGnHRgu0A8+bMgm+TCMeCX/UOM9XtjhCvC5j5PHBppTPg6OKMeqDjVl
11QPTp208ceAaaBM5ib5F37n2GHugyWE3cs72PxPyDQEwT50KPKTtaJQqaFanaAeexANsHyO8t8R
QrF7i7a/AYXAdGvdHBku6RAKVMAeI9bl4uMHB3oUjMWQZP1x5RPuFNsVTsstnjjpWONOtxXZxMfz
n+FqTS8yYtpWuUq4iukHt65/n95rGIuuv++F1BQMSvlJQTSAEcLVk84ZY201wwQ0bRBnS4uX1PW8
18Uh3Zm0aAgc+8AZtL+cZJLUWZmCm7NYb38LpkPYuRnoV4ApPJej8rcrHMB+1UIeEoDT2KFL1296
xU5rOL+l7CGuev9Ci/soENIwH/hjbEyp+c3jsJRZeygWPeuatkWnIwFNEtCQH9qSHwekD8gr0/rQ
96qg26xu3Z46P2docXnWY+D8M8eNlCqZPMJk4GHH2p2ysM03CV/AxoMfyzLvKBC43fcKl6wfk7Ro
RsNTf0H2bU24uOjPSImJp6XZzNV4Akl4H9SvKSSzXbmpb627/HsIhaTBWJtOKIHI1z2X8IT6NYZC
+9orS7rCMS5CK6sc+4UVqhBBcFynESc/8wg+5nW0jfsig2oqmYX2KVgiOakvpkV2fxLUIkQg809X
PvogmvzsJ+MHZkfNsdf2AwgbMIgSPFGVSRJKBZk71iZ76rsTrz4O6lQkHOn5XIdGiiFYhQpi/kRq
Pmt7tploxegpRMW4LhT5rqzDzpSjESXv8B37lX1v7X/7/NZgCxK/plwV+cy+lD9vx9XRS2bSjuIy
IwHcVVlZ2dGkckThLOh8FQf6Pp27BYS/8FTdM63Gwes5GPyBWhgsaHcRm3VBixOpHDxic7CwG7Ok
sDe04iIutdVHjcd5AY/FXun8aNQz+GKk9JZ2JapcJvBUihMgcRJ0uEWYN+KalRt5ruMIBY7NzdvI
Cei8n/fxbMYqHc0JSPSwLDxBzOcqL/TyHAnCa3VyyRWzUpaQ0dvIltJaOIQ4EhS/4p8ZW0UvYF49
IQlJfOe8EAjFBZAi5rZRsK8mFJCkLWnk0TDnLnlcp68PiIIMMfJIYn07/vtdFcmP7iqiWddvDDSh
OWA6Mrof3EmSvYf5lAgCGhKQJqk/TLWONWOXZViErkcHzBRrnJ1Tq311FiQZSJeW1crID44bG3m4
81JI0yzGG7UPWP6wvPu/Py+mAJdKAxC/F9usuL2+znwk2YV64N1+MLNyCpc7syt70hqyY+1JPGWy
WpOFLJW27ttm9ZjqXnO9UYuEX5hf2cKddOJ8sCJKKCHmjvWhcXe++1aj5GbsFdpA1/+05qvZAIO2
yYVmgcueBBst/CIh7OTTVIe89T9OY3GKVh1vwlzilz9b/t1V17beD445ahuUZY2q3KKGiD9H1Lzi
CngCRF/SDD5gvMtU0wDM/pWOmvdoha29cBeHSGJ9cEOqQR7Y27SYN6z9PO5IIE7xuHF1gytsqpXK
LcCBnDmkzzKYdh2XIvE6bG54/5fKkjvrHTCp0lKlFXckA34OMaXUJVBcG9EpNphMfau2AuH6AeZW
maRJnyp2EhhGoa4ToKyaOVhNrwW4aviP9a7r5BehacVl55EsJzRuvlMSWeuiB9wSRcYH0bvHohIQ
34vUWkSpdLH4LSYWT4zyh48qmu1KgWs6nuCizshLcsmjt7a7TS/tev6UhXsD5c/psz3vfeucX/2g
cBdI6FUVxrKbXu/p4XadZa+oND78lWuDmcr64U41P0uLWhjMrFLqKan982WJeIVs8wsU5Uartvmq
S2cbWwgeX+bFYdZKSHsdU9TlOGy7ERqwf+Uga/zBGWMhxTLuU2HsAtweAjGJVmM2v+pkFbN5tKk3
RFdEcUkh2s/rvyNEZvQ8uG55is2BpXFaWjMpfI3OMYMm4alldMAxPpJYjUo1Fk4OedopE3SggImc
mQiwBjtZdx2tdyMrH7Gm9lZJXpUEXhN2d8BdDX2ATq04x/SmlRl00dVl8fMFsu1LTeYDD0GUugyi
P+IyYEPlvOf+MHg4gKKprdOauTKj2Ck35eIhrTLqdl94uCOMYsTOLq+7LEspMkMiYnvGrtC/8jCA
WfpnKsKOqEF3brxgv8i0yIiClOjmFiHq+/BObVsjfWzQRJdV+Y5cM/Jep4NYzFizhILIMEmoxush
FJ2GS6ywB/dlD+z3QqRQHqQboVB7OhAPTfAkAzKRDBQHPULmK2sk6bjbce0x/b6+5p6rBdkKhxf9
bQ9ksuqzw2xeDT07kiccAAQ9k6XXmi8g6Xrw64YykJMzYmZlRoqV9tU3taOFmnFw/JaHC0+ttrLt
DheWdekSRnnfJH0UsxYIc076ZCnwVsnYb3g+nrS8dKi2UCQuXISHaLLbgq7Jy611pDKj1Ew8cpP8
tT8WVlHSBRCohCDtJkTvCZa3fLWFD6HM7w+fplHucx+Q+vRJZFh58BFCb1U/ilHfzInZ2BYxkFqY
xcLcn8dD6WAqGiCcpLfaopVXCm5DXTFO6CErW8IV204fggj8OF4iyCf9eib57lVZp2L0iQLGHuOd
Nll0yG68PW707AVfOj0fjSTagI1VjWPthbKAph+4m/nfbo+1c6CZFcO0Zf8Hu2OWcYpSHNiQiKn/
12nvit1fsur5k/LSSNuqMBnRe8i20vXnlkQM1FhXCiDrTjclOgnArLjnbIDkzkmq7QBC9lR1E9qh
O0LtL1ZgKVtVgA7c4CjOLmh13HTUW30Gc4Szxz6tYrCXjsfVCdrSiMRtfd/Sm0BY92k8Z5/HJnBQ
k1G6VlmavX5B4v/F6+5t4szOSAymuPbIX17PXgduAvCaijUpWVTQ0EkjG04ACpBb+YEEGsByzAc8
CA30LdZhUSyI7xSjaTTamYgk0Dg2Vx8CydmE4/ZJl8xopxQJ4Nio4LEuDx+6iz++rW0YpkgMYBvX
wbNmN2zp5fEQ+8/oqqdEE8Tyln6lUKD/QVryW3t3YHpAlmUMonRz2D5f9AqCZDEy0Dpx3XspvJfa
JKYHaD5tzkwzlWxOVZNfHklcUzrIils3A1SHwgdeJvOu3ec8L+S0HgYdfjVKcFAHvni9VuBIbUYv
89l/7IWB44oF0RyuRCauisqKcAwSHg8j1hQ7M/ev7dR39MwIB9q1yKe+MrKwMy3c6vcI8toUMQfl
AH3Q5MqAOcwVYWQCB05ZnR2Ut6IvpCwjtwzkiGsq1WqqL/jGoh36C2nt1dLhid7g8G/rS7yKTCuz
rpXkNofNzwC1g6nx6xPWdOiVW/V7kY8Cv3kQ2s5HaehAVWSHJGR3PqV2Q/pxnzhkI6J3EHsHDm8O
3YCKwa90Mg237KVB60VvI1TqLqG3vl4uLks3tQAMp2bsRmXXZbs4wkNox5NFpvaTGzIsT2XYtmdq
JFr7s78f/jzTt311HqNpZ/C82xgRKmo/oZKkZBqipH7RQd5Sbe+zoHZLoVi1qSdMWNln0zcI9SwN
UaqNCr6Bu0aEPm+q1B0b+QLsdX2xY/mpVs3YE0C0WDZKVAYAfnIrMjPj8gGYjbMY8zhWVwzOPn6E
Jp5rIAlZ8EPhMRRZNOXYdr1IxSKhzrknNauprhUxh+nDJ+Oneui0gI/6+sC7feCf92RSnPZoeFjN
MQy4npSxaWKYwTPaXH+PQnGdLppGhEKab6bUvnjYrXVvfOCiUk0HMlMPNRLZFFbreRF6cF4woPwI
QlYJzcsFOTBvJ0reDH7zSopHzXjEijvpY8XBHtoofhpWtOAsEVz/dToeY36MwR8OfHSOFrA8qGhI
h5OIko8gyDxE0Ws8bOgaYI5Mb8OBbeRuRgvWkGTh9C4Oa6i7mfKcMVyspiBa77wIpdaLu3g6iWG3
asB4a5A3lBTqgfGM8Ot57phPvVsTTm2pEYDvv5LU+jBMMf0H2uhbD96c5Ss9LROIlDulhPoVxKD5
zpxQWntdyzmh+Q/79nFJ43lpyyTWkOWrXkUDcLGhKX2YKWtDSIB5MYgRMsbftLvjWIvcoRMwdWfL
AxhEqtuAvql6OAMPbibW+oDh+Azz0ODPF2G6QivWdH0C+i0kCX/ncp6fhtYVYlCbhhdReoqTsg8W
4dfESyV6u9nrWT/btbVlGw0pDZmUQrZHMLUDw1Mf7pWuV4Gr+4LRaPwTor5v/0hMOP22c9Mbzegk
hYycO8goEMg5krDRr7C0Pm9Nx5eHddcPAoSDxDlErWlPKGVuTWlL6e8gB11nmr8E9IwHYUO70Mzg
L7EnoI+q1uqoBjdbs/06nUuVq7w9pfKEzTPFcZ2CwBBMmeP/9+I7tr46wYqq8j7yEVrjSG867iZ3
e/qL7NZFnpCLkDUUX5aC0WIqxC2e+0sGwsBTVmomX2At4zL6DFQ9+7+vswT/w1bJC8v5ADupIDM2
W/ZtN974C+NXfg2MlhYyenRabVPna6qwRvYuiflZHt/FuEjuvCs1pi3AzqrWqwdAOLOOGs7LGZj1
qIp/x6g6uB7O1uEdhEcdS5RUlE8M78YCOQySmppXT7UTPjmn4/MM2AVRI0WVrnlkQNF1bCEQ6qBO
q1IuOQoqvjgpmDGzTu3b6hwqxTy+J/aJPcMilIRIfATn8BtP0gp8/8lq9gQia10SqOBSd3UtXU2e
JFVFrEb5id0z3fSlsZUg4cVgpmxzK5ueMYRx3cWqR1LPfgHSwgY563eBAO8fV8aOKgJrvDKuAE8S
42hJxGlATNHhU7vbEYvnIR0st3zR8V1VGL4rf7qbKxZpiJsgrvsbhCI694PAjW+COHTfQbSemlvq
77I0FtUCMa0IDm19nd9NLdJkncvlxpQV7ourkWZOFtGLDZv5CQFgiYScrTdjfinxtd2JHCGCY5Lu
cUMYQlm/kBlcxlXgfkhdB88gTRCJCCGcsObvaJDeuA7v71AD62PvoWxnvThY7hP4YEMZOZ0zv+oK
vc2Lobb/EakJvOky7zWMu79RtUwokkvU6LE4UVZGz6uZK2AKouI6NQFD+mbBSpYCvxdCSo/ZbBQJ
l7HbT3H90WuXuo3tIQjB3NsyAKIq3/Nf3a6QqYe6uEeuRwQPJg9+RDOoGOGIGqMWydGUIzFS8Gld
Iz/xtRWTU5CyLVEQLDuieHW0NrMqQoFZCueDHM89a8KAAv7b+Yx5S7ulLafiM8Vtxw/BuroUFHdi
yLsnfqQx++32NFAgARnJpwJUvHCIh6dFnlMOEVslM7f0ks10Key95oeyvefgZoT7zdjYOIxWUYkB
SPbRYFILfJPrlo1p/s7qdgYssB/+K/2HLGPSmEDv4xm/tQidIPZ0Rf3wggGpyKHnX0lvi2sopHaG
UAuWHC6/svrangZYGz9g5v8zfOGHQZBcqRoAhPbzlFczN3+5JvSC3dvhkgzjzeVMtjVL7HPvg/Yx
UC67uxVuBjpWF1rmzAyqIxvrushkGe4fAMLHTDtrgo3tikd2f8nYMqIEf4xauSBT1SbgqocW8PYa
UeXnlHEmvhuhw20F2fjFUudFCAXnE0ZXzpnidzCg64l4IxZrP5lHra4h++S3X+qErrZmf93KAve/
mQjez193dJD0ww2M5CWWofnvb5d0VXtN5Fu8UHaekksTxnJ1d9WmWB5QotMQLVHg+pPua1TtURM5
TRnrst3wgLk+ETpAyDC5uswaTI+j/4kxYm22CfDyKBf/s75A8RTSny0zmOR+XDs0wQy8MokfQVK5
RCVLKK10/sD6AS4VkqSH0LUkdyCvncO6NE7VfS29OZHsYyFAqtqV7zJfiLi6LGCMmsTGe/XcTuav
N8DdiH2GV+uDbeakXv3wKSLQRUzB02UN2bI6NFJ/GXy0U+Rh/JfD1TMzeXafAOg8cEvUKQPzZ0XC
435nbLJHloK1ZulJsCKywq3vpCjp6v7CpHkCGNvP2K3Wr3AAwh9ibxJJ0n9DRJjvt/75OLHMc1uG
4SVrqeYC/WWil/3oGFrJC68IGn8DSrm5c91pHYmELdKibtzMVy8VS9EnTb41xLuCDioMbR1qBcVh
tBM1FcGQCk4fKZmFVVXgxtWD/0OcS5ufOVmPknUKObZzqt37WuVkUbrKikstJzy5OmVwvthK2G8m
Qrz5Ndx32R0LgRKgd/tKqZKx7zrIwj447klq2QjMhEc+cXlsXf4g8grEhu/DfxhAyLaKk5lQi1Jn
2FmkjdjV1fmmmiXWVDGV4PrOvVuOvO9JDiN88DQ18MoocXDA1eP54x73jpwwPZeCtNSN4TVUQo95
SI2b+M82D27MKs5TOW/wCSyx25OQ5V2aMTULMcrOZpyMIm0nfJKBsiDHmak+iG1NfYqlnmvuY+ZS
Kq9XDeToHVYennnr7sQ8C8xeLUhR7bLke0CgCzP3fLDkR4XF+Yhi2f5Es8DLZUAKlMe1XBqKszC6
vhWlpO3PsfPVATdLChcmNr+wVMnK98mq7OHdtgl1wM1ROqbiwkQKgFqjcrtOAmEZEwyLadHxmtfm
Luzi/chiYLtndA0qXJWP6Guj1WFL8+4IoCuU7g5rSxvBTkw5V/kLaf1lOgWYZEjQe5ViHGvBjPh8
USnzWnNHWCTdpZvnjO0WLhvaGeQpLjO0s2dQ1ybslKZ5vvoamVOjnjIHtLTC2UcXEls83rMSauzQ
JGTwdi8j5rY8qDwU3pX1UJodgD/mdlthL7j3fO4olis8sDdz1wCnha+Lm0HncQKhvDOgg/KWRlGm
FLJ21CChZxTSMz2ceI3eM/O7eUhgLbPeHIpXgQjT8/3NmEkQ34IG04tbASp/mj4N+WIxKHjOtK03
eq+IHDXC1S6naqBSh+NgeQmq3TH/8TugtR13G6734rajKKJhFVuSIAwv+AOMhADA1DbvKwCzhQBD
6em4jZTiECE9uW5WhO1O+/b5jhr0ijO5ZoCPyW0k2tf31QxR++WSPbtiLsxiqxSUlQMz9Bl1614x
TEwWvMo/qjW5kk28CHV+2gKQTtX4NwVjkjOf4snTKdG6NCtJuDMnzn2dSYHRhaV/R+Aer7VlAb41
f6qtLslfqnsiVsRO0LsoP4NT4xLYPsWZox3ipGhs+wme9q7VhT7QM41Gn4ifKA8WJJ99HNBiiLJm
IVkg40dB2S+/gctP1xrEntWwpLNKbQRH4xnKsX9Y8PPXOS7j285QZkHdxS1JTDX3rgiTyG58SkZq
3bgmNP5+AsXzo5MMa4lHFw1UI/14OmsMJY74MpV3qIDR6UWAukWdj77w8FSPRPwWYmt0VwqbaUho
tO/h/fkM3yajxbLCeQ6agY0YJMS3UvJaiHGN4eeha0nbrmlYoh9mpUV4m74615dt7wErDwdRpjVJ
7uSs2zKPX5ARs7+ni0D2y2BC8BdyhYvsCdx9XvFUgFowBVNJgHOYXMH8rBt67ZAbmYiNpDV7V2b7
L0IJPAHpKDmO8qpXk+ILd8ZuD9A9VlAriWriqFDGmJfzapjnXVqnqV5jLWNNYZdg+jgQf4sUpHPD
po7BsgzEdqspQ5RM+WZgFMblw6EDNE8FEVjiaqpybg6eh8LWf2oNXkAjDR8EHQZIeopiXZ6y3lhQ
Ok51hmvGlGJC2p8DHtPi8y5THNxZGT53EDha60kfs9DCtNpbJqXV595wFznDyZLsiiA5X1/LXBsy
oemVTVJX3w/UefpnbAKD6irXZviZKRlaozPKnz4C6Z0TxqNu7nVxFmWUXgWHvLanpCVzXvM4pvbi
4NqzLNR/LkQ11pd64WhkzW5JNL4NpNsZs3iHMa3AwD7AdkJiijLuviSer1fQehW1AMIab03buwVW
iCjCiqjH4ADt9bqJ+y2zWoo6NdpQ1irtRntPtCxl6WQKhS35/5gsm4XNdZLPyF6y3v3Dnoe9BYsv
6vz+6+EvCXZJWRMH+aE/ReodKbrPxV0ljhGHCimaOAA5UQ7KomQMrAkU9z94ELpBSMUWCxXXRLoQ
smVVYVVPTEvaHn7uorv6JW9Ko5wuprkhrXzpBehsPc15reIazBQTLy5hMfQlBOSuoQEtjosuEhyK
raJAPFq2V8RLMzkmnXCSkhmZxsYOGIS+jdK+27r1QSoegB3He/HCrgIy4MwlBuf0nlyp5uGHJrte
7N+gkqAHifLL08zE4X5OTQXguUf+8y1tgbmAQEErFX3O4Rjg2NVnoredy8h2RTM85K8ilOMpZJT2
XQUvIH6AIDC1IRVw7cvuAgR6/uyYfZTjdqXveb/sPguHr6P5uhqdjn7mygsPKUYBsUAaQcbJkH5u
x3GmgR91eZbIBX9Otpf8kOYB9dUCCg/nfzUSOtM5sMKirxfKFkpaN5R5nRt/wHA8mfHOzs3KmHjS
Wf5rsowibv1XRhU7wJYXg00VTOq2IMxbTgb3cWmxq97miXVfA1SEXnlQroQdPy2yJRGHU/dRG773
kuRy4rOg8X/YwboCI/Kvedx2YM97Q8Y+A8HmHJ7ItF6SoeacbtCZoP/7Ku3hrmSKXy4wL31ZV/EE
U+8S0PJb8wZHSh5Uilis4ZHBRVOHJaOGOV0oHpmzWWBaQH7z9hpz4ONxsCP+4YJRRPHnirD3CRq1
RBIxS0F8bUtvLH00UIMpt22r9WhN725LAb2IroaqJdbg12Dk+Y5khtGwP+ALTUvAh4Z0EehNwgro
dlpiM7bTmlX0PBEuszHlhsR4fckidL4PdSzKb0BucZQCJxlEylNIPrJzrVHc9NNQypQEvI1ABar6
St5ZG9UDDLDuBplfthGnR+SNH5/CWLeOuibEZdHQ/G5KWjhdN9or4sclYAw8SPhEgp/SO7CN+orp
WcINafgYqXmLtMHVkXURQJhUeDbiWEWU1VPjvVybvNgxVGThKfq6YoTdD09lU0KTKh3RMiI/Jnga
URD+jDsmn9JV8TKlQqFygbCqSyyqNtHofwaYoNVwtUTWxp/S+UgLHi1GgneFuKTGzYefbBR3ZFuv
UQhRs1TcbaDilk4zaUej3fSQRtLA9D9ZeauWEk3QirM3M3ENBvCyY9IufXe3fKw6Or5lpVs8/tT5
tsqeWtBPCG8bp/NGzH1DiGCfkEZ85kTB9P27Wnx++8pLKpvOeZcZHoWfucXcCyieHQY/ZGrbmX7p
gPeqgmth3qpvKWaNMTk02wIQx88Ea2INvvVc0mB63aIxCik6emeHiAZbNzzW5LPWCTXef8uIa9/4
qKcLLbDW4kMHlYggmXSJYpSGLMKdnzw84gtn86CdwjEelUtOXmIbqMt2zHPBibpWGBqWWxluG7IV
P+hanb2M8HOg0lfMnq4/HlxZn+kpA7JHAOLgShQw4XtyErDEcU930m4Gvi1b/YV14Y0tIRLxhq1n
/NhIqs+UXGjGXCEXy8xcSWekfWcAWuSSskDrGtdU3+LMw88VGNCK9ndG66zjPeDMEDKDQtQtUvNV
pjYVN5bEIaodKKdAPDdxLHPDoozUrmr1u6qNrTpiHAEa/M+dQ7IiTP9I6iKub0+M7mveRYBxKNKw
9zr2khbpEL8N1TwHE+f+0lJd20gsRgN173JXrAMIcX04pKwPe5LQ1F7pSWSRZ4XO4Mq8WFZTcrbj
wbZGQn6MExd6SyvPqlh7Y8NfmYTzcUl5Nv7Hac8BMKGS5/2UDkwae4rMh6TUty406noIcGgsoJdq
JS3lrKYItxH0RoPSwWd5hDS9fHJwPQ4L5JU2ZBpsEmmNsyX2HIOD46+jI4dWgWvt4PDABy+l9mEh
Ze40/T/9T48vPctbJDMA0fvHIq70niGUXwpGxNFD1kp8fmREm3U2hiQzSJms8MlOBsaYC3G4ZpXx
omvouD23Njsq7llv/3s+G1++moUj9ZPvKuNxTw8djodrnJ9yLHxRQ+9EKVkrtz5VwqPiPFl5Omgb
Nk0s6DetIRQatPzuhptAGsyvwlbRi2kxonkklRySVU3A4tR1Eb6pzHpPtt0dlMM7IEv1Xy4gOc42
UlAp6gVe8vg/ATLYuju1STqNXgodaXG66mhmu4i8mzfI6bt939ePviMpBx/Pa5koNfv+GYKt3tuS
JChkQip4Whg3WkR/4dGpLpzb4LZVzRptIZOnZuFTEi6i3HNO5mRPVLayAjqQf76AkVc/KRpusExJ
+PwCnMzQ2HDku5qawQAN45ffDP2SOD1nShevXmOAFF1XsrMu4RgGNjaFgEAEhOfCwkA7u8jC3PVS
YPaYQO9eK+dn7Z1WnwkmtETEPwbvkQfmTnubzYg9/ZE9wOuHNfUD6c1cMjEerRkBZo+cJ6vx9yUf
LhE20wQzl08oAjUl33ZC5N/K5zxA2DPaz7rdkCoUMTTduvHcw70ZOOkxJxIfehDCofo9/XTcxIUx
uSqzK6eb2LEFjntv6MELZwnXehRuTc1ZQuo86IlISh0HelgYwk9NGQcc6P9EqS4lysOa9CqHwk/k
iMSYwSgjtNWShXzfk0pNhniHjlddQ5cLGCIbC4FPeBS31Da27X3YPb9ERHAQwl4eUzJe/UO8BbNA
/vnzgIJBlAn0pUyFyB86GUkKGPu6r5RJPtwHS9hXK14CSUd48BZmYpO8l5nG3VKbsIfMbTBdLRnx
4avVS/KwqKj6hu23FX2TQWinnA493BzrX9q3TppkzNmniLgolgqU5VZ29W+xb3+OqiOSw4H/0/hw
JGI00OE0W6LToBNjSF+p2ZSzun+2bHiqCUMuRDpn5nbzrFsVzB4TA3v+RQvVUW5A0AD+Vk7u0ksu
2yoxx6yDOeNdMCbq4lQgh0wbQC7JHLwvQGYXznfHfeI9KTORMrdV0sMIcjhy5jm6bDqEuZ5aIpHg
FwPpWZWGYBo2iSefkrpkLVSgTgGgz1lbBmaBXbCW/v2CYMyC7pA4fEDeanMqy6geeZnXXxyOJ5F9
5vpql0eZb1KLs+FeS6bjs7yKupYjl9ugfboAlLw36P1lSAxPygehlqoUGkk5v84FJn4sG6YdkAm5
z7oS2OVyF5+RSvagwZOBn/BWFYXWT1MAQ0Vqqgtnfs13UXFcD02O+a1Su4b9Lf3l5tuUO6ltcQc0
dKy8eXXFy9te8vKmbXpb6kSdhx1S2EQukCuCq+zR5jBsgePj2MuVvNCDXLLW6vncyM9Xj+mSMjCL
cpArBi9uFmlhIZsFC3hKBp1N+7ImEg2TvQH9PfHQwn3sEtM8bxiSqUJ9lkl7cIalaca2wZ3NNqRJ
b2E2xtICK85W44Jh/FCXhJQ+16dOALNA3XCPplIicgzicwOBRPkM3KLCRt+QldZCxGfTdDnbuQen
rpPeSYn4NhAGEr/V9L6Rk059cFfHMU27TtVqblGrBJhAZ5SRLgQK7VCYyAEKpZijxJ6+q5Vrc9hP
I+NsRbfE8tmvYjqTQ5EgNfLMSu5QblforipIP1UGNw833RqKhMpxWGyZck+MfJvzwIF6xfEbJfqf
U2FcddSZxO7oVFGbmnpTnTQMNId8pnXVxmOVbfvXn4LSs33j5hrDk4q/XA+iW5nPJNN8KXYMurND
9+dqWmF7+YhKLyocQuWEOsHOzxvYJgwYt8PvYdx97p2kw+PanhJAOuB4u8aPcRirfOzbkrL+PUhN
2l9FjIhWt6Tm4jLgpCauQX+W/U+vbB1vXlgcs+Dj+zG7waEwGnn8IMGspQSrK49UUkjuUR212ess
Ca1MUCkK0MiXeWbTeFCjpR82BRDsxgfeYjVfy/Ff6xc7/lP0ceubGigGIJ2n8H/mzVV6O/PABu7i
7bccEDkg4UbcxiT0MK2dBbQwSGLNGyP5hdEl71YTpFRU4D1e4FkflIHWnmFkIEkRgbYb5S+K/Y3Q
DhliL+M3OW1vfd/cNnIKsh5bcAy8OJ+BazGJtZH1GHcIKx+T8VOnKn9Xg+cGJQGE6NW/h94i6Iv5
H+y7hOyzjxXPojN47Wl5rc7Yjgc665SRBezt9d2Si4CECxAVMJ3O/yHm5qTwMNusEUSOWTaMnQGF
GZfySvjr5OiAYf1/gRjPbjVxWW4sPilMAMdiwIS5A4G/x3+ipi3dYHEpMABweY44ualq9WDZl+y2
poC+rjfmbOZZJfs8P7rlkBnavylysJbc1AN+9B4ABISYvOWydZXBTnZfQzDTue03vbxwdx5+Hzm3
mZdm4Rl3NLlnv55s3qDkGPo45wSojmaTp2bsTiUzpGk9GisldvA5p1HeWlpFP8SflFF8zp2W/Li6
Xuiu+xJydWsip+pePPk1DImIwt+IB67m6Gyz3RfO2vSX+KNdoLtvH6drF0CRvcn9o8gfT6346CzC
lcHiGdDpkA2s/VpKQ1K2Ss8dBe77d0Ka3Eu1GLynJtonLCy6QQJVK+R1OxtXEuLEuWtpSsmKxRLW
8ZOJvPvKdr8dGdMDgDLLDP0e/G2/NaxTfn2OcihXLtyH/DBbntrTfyufvk0nQ95SqiHThXcbHRpB
iOstegRqqqFRoozFgxeQcpkHlbzfNZ1EdB7DBpa3+GxLxUwGKj4zjy53kq+ExT2b3/cwLguDc3ji
xxykqoPseH7hZKOrZtQZg/36gw3h3Yuig29gGPDf2Gs+xT+71jiXQHDxUT+YRDTScoUQTAx6XCMN
vlmH5+ioF6AxcYBoHJ1eZ2s6+F+aYVaQz226ioc70lhwRcUy+m3V3WUyJoV5I3KpzpairfGs9VRv
UqVTpdiNO3Vk+XXzTC0unW/rXtbqQMSRVpjmIX0BTYW/UVJnRTWVhKqYi1sg6DyZrGr39pq81IfA
ljwMLp1z+K3ClCXaXW6Hfn2nDazvxBh67nYflwSWY2BxSfhcMXqRzpUQKib+UOAiEQ/iTeVhkQQb
OkFfUoofK1BtekMApuUBtGoSBQklaZnuhpNgVgRbAOANm2EU2mac3efp9n/ZSOqV37+9TMvNLMmw
XEplA4VBBk7sRpb92ivOboyclqnQob0ORyaGGuqiuZb6Z1JbXfJd5eCMY6B13wdM3HbavFLYDw6N
uQ0pQY7QJ+t5/WjvcilN4+StIm7oMGzt++fp72haBlUSXC75Ko3Hsl5jzWOLO/W0gR9+yhHKE59a
tjSzBto6wnXfmz4CaeVJTphmYShETAu5BX/kj2aSyhQHwbkf9UmJJLlroN58aMJhH4UBDcYq2VP/
DG2kpB4dEkyyXKYGiQA17FubB4SPj8RiSgjXs2SlenNP+vtHKQyHyMc0IHo4sDgHYQSyDQekSYIB
lmlbvk6dxeDU5V+Q1bJBac+xbnaAx3vwRYTltnAe4ieMGcheKMqxjARPys9y/uH+LjHw21uSmyBz
QASwdRbKDsGQRs8SqAEEPBJtGM6tyS8qS3Uh1s1LU492oXem09K9ze5dMjqCJQfqxeUThEjdUmGc
K8p4GhG2XnvV+cIFEC3Fp7Mq+Hl313MM9Vq8J+IR7j+1p4QIrWh/0mS/gvX3JwHGhtaKKE8rNXAN
4fVKvYk3TAVeZAZ/av6EpSCSkWKQuOQ5alPl7uGT+37aPD4JTMEhiNbxGyFBGyISaH650rxpiZIG
LRC0mrUG6Q4I+tnIMGOqGhtjKVE0u3Udn7s+l421clbUadv00INwcN7gYnU3sR3UZqKLfb9wjSuk
+nJClzPn8Z24Y9OkYxiikXAdslv0Z1pSSHPK/17b53hNitVQmEz/ZWPOr2/uWM9bTrleLvKKrws6
7txO1qshOSOTKwR8vRpwa7WpjTjxiBH+SwkOTkkPodmPKNhLnJi788Y6AYV/dKPgv/cMS/GJwm8W
yUXViuGf2RE0JFivEMn5ZCCc5iv3wUVcMdJnwRM2ZtNzhpBm+Vf09/AVaZ0smoMv9SGnLL+GWppr
jKLh3nTU1b2Vdf3tIomhFcbR4dfT6CT7Yu4ADE8R/l8Pjyl2xE4myaqnyXzPWs1k/X3LobAoqj6C
yfDUq952xzIA2VYm4iZZsiqJaue8M9e5+X0Xa1zp6MNt+PEvACq11tKvhV0ILYNk6l+CoPzl96+P
FXaK8LAwzLZtS3piHCAdt0Zqbcs4rcDLCYIfHKt/nFC0s9gdPq4NdWHUsJrGXGaALqtMr9owKd6z
1ndRhE9By/REmSM+ul9wb3kZTDnmwaVWNuOcnT53aPsKK7x+K/c5mdd7XYXd6Ij66Y9LJLtkRY7W
Tkj/oCUjKgYCiGLXirXwxOEMeR3MVYiWdMea/ISdS6pCn7wSpszxp7HLCnTCtFXNwnToUdKnvwB9
ManQtG/GsPhRwgWBhsoD1OYdWMeVagCEK9iiFVyTHfeaIL6RiNiy8uXxQkqp85flgTyxDD0UKlPn
/3QkYwaoIReBd/baa6FCoKegIFz4UGwIffD/VuU+8M2y09PF/yhJu5d/6Ltz6qSfziv7zfnd9klP
9jtpOdYGktabdkRDbu7NBX10W5U4EKohiWyUE2vbRfJ1pP89RmepjowBeqdUGJpRFeEEJNkwvt9p
hhDdmdTdFEGPIMbqYOVUP8UpYSwPDOyld/cLOT9ZIoIaoCW05Et7ZeJc7AMYcNCj8/211IfRGd3N
vzbXm7nf+dUZvuFWRNP0BLwu+mTwoUMTWPxvea/znzbGlq8eKNIIBASAcIzflLEBr5uWWsXSYi2D
SRb9nj/C1avIHVc7Ge0um8+I3wG5N0eaIgiiDJuqk2++j7AZy8kp5A8GpCEj+01HAaVdof1gSLG/
fbOwU1NmIuAmWZKp+FrzI7ChCuOId9T0b/JwrTrYrJ8WzoVGc+FMuq7ddCg2Ray0jTRQCaxE67dd
i+zb5UNWFobWIPs4f71PuUHWBJo7iaxBNxrpuq9Mp1/uR53MQa5lKdVC4E5d7ssqnIdxnB2/x+LY
yENBjdCSA4dTeECeifnsvFGgijfBUokZwafoJ4RGtrd0FC7KcQlnKSnqJHy0YtPJ5piul0OKHZ54
WGCCLuKy5R89yborrtBer+Vx3lo18wRkounBizZGIyBTW636lpZ3yvv56U1Uodis9hQXuIgcJPX4
J7XrqCoUQ9B4Rdv3OSFWc9a0BJV/qJpZws8RvTBn67jzkaWrwdDKdxQpnVGtvKAiJRY03oe/JQZJ
rJmNmEx41f6i7Q57h1zGKHYjw/dPWtnODC3/JBY9acGNdlPF2ri1HdW7Temv8+WLzdDW9a54b+XV
BoQsz8USvIRFXxwY0QH29SUjxXI3hHeL+0FjDD0YJT16cBdePS11HK1kfeveiC8e41GUCVeGgA/i
57LD22qhZ9MjQElcriFmAGGDk10qhzLvRPIHs97EGozgO0goIwlTF4ck9hq4MiAnKc2ep4mqepoR
7LiSKhmIiTTky5zoqeh1+Gv0fAY0NNhSRCOIHyXXvWy58jke7+GfDYgEBChLBYxBnVcGQqwNiX5l
wmB6oJDwWYs+F1QCGGLIifYyGp+6Le28aycPpjYlYw4k+UVRqDQ7jrJjOesl3gxMWS8+bXcO1sn1
nM9H1P9NpYyGaTUc1SAelIPHyFEpjUWkbj5JpKm9y61c6WO42GO57h/pEyL/alPP0sVSb9fP39Ko
dx/l9TzBTWdPG9w8XqXQCsOEzkS273uR3KfUpt6U7ozY/shUBWixqSOQNaEcvl+AgGv1qid9JHiy
qvVI5FeW3ucTa1BWAtlJcLaFdfW1/Dqc8X9j0E3V5LkzLAdSGvIv4f8hRB7Bn4OkFLXDS+8pBGyU
VELmy1J6aU7exX8MhkVqjtuBmhPi7E1ARfF4B5EnEaJwu+Ew+qYdK/jhYXBWX/S/jJ3JqzQS20F4
r8F0v6wqWg179qQJUejzvkHAPu8m+D6xgaZJ29Wsx8f2spR9uLc9jYwwAC02HlPtlBnD6JOkrrHg
a30HtBISE/NVPtUfC0KwLGgGSCDeG6fiRjahPEAbIzzHvHfXG4SYa0o+bxgx7BqPLRaIWKCPnZgd
KWgyRq4uCLW/jPJzoKakiBlJdsugom1uKRLGjBb7x5q+VKSHUctRPZwJnjXmg2QzM3PTHejYfCvy
d8C9ikXFCaEW5cdUVPQAwv5lb9Kh8CEK6GbwSaDeeYg+XiwCrEiGfLa0yqnJqn6QYIxbTyz8nxJo
TJjJ4731rs0LWbKuKpxPCC9CEjXbDrWhLWZquS8ua72O0PxvOE19i71tCP/6s5PHYPvUxTZFhbBy
Ztu4DXl2mqFowel+5ltBHvZCFMG90uE36sQPAP8evuhkhfKJkcRx9ryLUU4kGzj9AHaQZLKLEo2L
qReNRaMSk2IB+m25d118Woi6gmD5dywgEXAEP0btmnrXSXK18MQqxKv2+SGRigswFVlE+risvzEt
CCPsOgQOQYq+hDrIsxan82pxAwjQDJ2sROIpet+O6vHuKuYeZei2xXnOB3eNfpzZQip9zOGoLP2k
G5aqyriH7RRcpHni8COAbnVbrum2imVtQKdTBJHzuAwKdEQGapiZ1jcpsCh7rw9GUTsUdPtsYL89
QYZvgTXrlu2+Ozo3FHues1siQXK6ckr65qirEcsr+p898QYhg93PQ1LDKqfaWQHLTexA+ZpgGSxJ
a/6i9HPYjB7Xl51vWCYcRZPfKBgwhHZ5g1UGoiGCjy3dATuILMHvKk3mZC85Oh+N8LoYJWgCZy7B
QBrTHJqW7z11dB8lnA+fhMfVsHXwSCtq8TZ8iXLZSAqLoex+/Cxis+COhKkpvyBc/WhmpZIftoS9
cFbulChLAit8W5ZVyYnFYTVgCy6LWwx8KE9R+vN4yMqO2Xaky0whdzNXcJ6Swg6z5oGYEoyjmZOi
jwHeqPPf9ucqkMX62xlAiZLBq0lM9gBNRXsFPG+5xCf4jmAiF+byIXw6dRzG7S+0sHJ3ygvNwrPq
e5LJnX/Hg6lRWTwdCf7lgmwTPbI0a48Y9ExKy0UsZ91t7fju5uqVUoFsf84TXiZgP1GP32oAqCwS
OY1z1KGwQwomm52KcG1NVuQ04E7dDMPHxid9yQ8Hj8MTqwOEJa7y0hfMtc2SpdDLi3mAnxPLtcUO
WEiWe8pRBYlqm8dhZXZol9sX3XIcbnvjOjkeyoQc/9EEGNHM03szTwGBNWhyTwwFEmDI/bcTAmFt
a9ium9HfjlAkhq+bHcpRyAsWzhNG9NU1lGMnVLdJzEEqnE1JVf9/z979FLJSIgKzqeXK0SimLmYg
U7TNccjBdVUpaO2CdpE55BGs/DXBqu0d6QqHhuqVbDwxuXWZWbHRgRKebPkaZuXfzUJZpTm00vk9
Q8s9SMu7TobDxAeDPEfxHUNEpZJYzc9Qa2Oyn1NeM11AHx2Efd3ccee258bi7uY9P2J5gXxtFWDL
UKQLcq6KlA61/LjL2OIKQid72TYzg+B7zCPSS52g8vwm5XwhgLOzh2hE/+gOZT8zTAnjFWgCDUhO
+elhWfwkg0AP+NqS6Jtc8CM/v7b5WqkSXDCDZLVVFUuqldrh6NE6jt7+OtIvmSlhsgXKG9Juapcd
lP/t/Toeiaw4tRMk4Jg//GVWheGiyAK5KkfWqhrrtqKWgSiFNTsHliNN6e21BRggLOqUIZbN5gX3
uy5oXUOMe+ZdTUBeoQ4NHFuQ2OTUO5/bRvnIwBiNWvC52+ZIGpiFDsdkQIIgyE9f6cyD2e3sr4XR
H7xuq8k1Jl2jh28NZdne0uFdwhwASSDZ5VGIDkM+XyKSWSyFiA5nLTTd64x5Tv4JfXcFwYFXe3Lq
uzaw0UmepzlJrgIkG2noDdmEZaCWo6jZ1sdK+CT+u4UYdvoANiofyhLuEV+C2Fau95+7FSGD21QS
OGjJvKLrhQa3XjiM61G3zogCGOX9mLhp2cDs4sg+6otAExOQCu6AuZmrZnn72ceWN/tQcL6/umb+
D7/umNGrBgUCwx5XpNOzAU5rrV6zoS4aaXIe29Tbv6tnZW81WsaZ7ldiqd+xko7XVuifd9dCbW6c
4lwpO0WOOAGZTdRmZ7i+YqA8F3lG2jkuMj4uk9AFqO4FnvHW/MJGM/CkBKgdH8ZzWYCSHYNTUNxb
Tm2RvqTpdXsHuLxvyZmT/t/3fTaO1QiCedD7rQgKnp4wV5F0BWE2BcF1YO2oXlbfyDDvVRdqt+f1
ov5J0vsJpClS05U9RFEEyBOQ9YbJvNwG8O89QJxKHKlNQN/omgqYxXXNMW8tRQ9X4CovXAClQxwj
v2Rmc5lTep93ey6SmKSD4KCCvT71W5mSRXsOwCtm7eijfAUkR2heQl1P+ZFaDhOpQ20JBuUgqHBv
87L+z4bOGWF0oLeTNE3R8ytWfWKNsao1tToBLpW8tYacWh3el8+/Xa0YnunLkkdYMksSfk/WXF2Z
rJfjJe2ytYJ2TLjV4ZGSmJ9vN1TAkuEs/kRDsph7do8XHfZoDCaviF+l6al3xH6LNnnvQDTHiIcr
yGnlw2vrVxSp9NUJZ5SANGqU4CgVZtpW5HoOQ6LNVZvaGGS+XU/Tl2rH5a6DmBbWYUZ/tYNdqVh0
UJ29AOwYmrvr1nIXfga+nLrJ9ixfGSBhxscR8yiQlE6bbXh0uC9WS0DGSzh614kw12FVKRqudCoy
PTWbv7STJzFlse8ix1MSQrUzUaNOCJA2GVPEGAY/bSgOtPoulNczsVkeAB1+ntsm919gBp2c4r0s
16ZQtSiUEnngaPnddBBSX8O5NaSSVwJUlPXF8YhTvSYwvtXvTqpANLr9mBdXBpSebZFGrpprCp1A
XHdyz8vvZuPnQ0SVFeLVbiUR924BW3I+TxhQ1KHe8NUCcx4vOttZFGqgYGbrHwotJYxyWqqmzRuK
GDl+fTSKRb0DPQCnVyRSd3SuM/QYf2zijU2prAme+V4MYD53W+e1Bun4mi086yDvhc6783Gu4Igp
eo0S9nSycoSVgvene/FLIPS+xvtw1eG/kqbr0myrhSupzjxxB1LwI5rXEO9I99dDpeXrZ0jWx5H3
93i5Qwnx0/FImP5TFwJ1Q9x/TY9GHIDT5JDfVzqmNLPBOroeLFyGv4JOzEXmQbWOxSsFH/ZPA9mL
4WPEQOzYZf9Ud1UXDY5uJ/JIpHAe2Uc7x8sXScloyJKqigqfXSO9m95zv808UIS5vj4VqMQQLd7s
kfKZCYubdBiXE4z53an3A3KtsF7hMk45v2pOhD34QBGvBd41gfjbNJPA7atrRh9WdvT/PUujSv+W
r9+N2JXLTTjtLHGjHrLbcg5ZkZOIdqoDOsFqG4Lz3LVwdsW87BbSWyGvaVM+z562B+3Qhb+imggN
nlyvgb2D7Y+Q4h1PiEVZLsdhHL2BFloeMVPmxEeb4oUQ9vvLKSwV6YMgNSiZgK/hwOBKdVs678ET
YemwOTk/7J2PfBNTHNpof3yITTat28QJ3MCGWR++N15RH6IqRaAAnxjp8cxdCjdLHZEJU/F7ohBy
ACYew9c1bvWrOnG9CRgJndG0VuX2hyLRN6cSXEZP4A5VkpFASakC62z50PFjxso3ZPjRbrwAR/yZ
6htNyX8IYuo+QjTZN1IoVdu4vA1gulL4jz8BM+Vb0ebS9buQpLSxvmAdMdSKB1oXE5Jxim2yQnMJ
TkrjROOOTP2Ki4pEkxLtJkKaG/DIxGVoa5VavUG2NEx2/6GxsxpMW57lyZFPEge711RnhPNWVuVb
Wb038+bJqU2/nMZ9fyTcC3i7wGcWkRibYw/vyzN8MLIw8+na577lvkZsTbTd89L6g3ZVrR052bMv
wiPKzbbFnZPnDSwnHfRzqv5Jt+CE7ZeC0sn6OVKAsuD5QV8/ifm7z6pL5StlSxbBSRoe0xGH4Blt
zqR4h/VFXMSPSK+hqDcZdLqqVwsQvpnylA9NNJsNOgZpl/RDmjLigzP3qbuk4mhqMNbG+ZlfK42e
4lSv0TCDtcYnha8LO9PHQ6r0GkO2VMEk9txTZHwTFe4MCN/EceKUME1VBWlCOWQ3vHy8BzYkdXwc
aM4yAFCEEFU00b/qaBysSAKluqu19UBPMlyWHmb8qEhiGMCF2g2q+w8sLj/aS7tp0obKANMyEGE1
6fKp0k9rp6j68+yFYMRKkpYzMcCV31fnHInJKNvkK0YbBRFQLPdLYOseY6taaiIhrKTp4uh/yY/C
g2dROZCDEqu6XUxbr8SDAA9bDqyhPoDET2Qkfz9BM5gTDEEdnplEvMAwFO/brC0ufhT8YtdlYwr8
aTHEr+2WUE5DtIO8CB/40MdpKSckEg/fBcJDzYJkEgSJ0+WnSCQ87fsRB/8QlPE2xFvuN43GpXvj
sFYhXjZmVECmtGjeN3C9S/7vRKEV9sV/9aKOsySty2M7Tt6uE1WT/NQNfQJFDWl4t5tHqoevSmb+
moDgWIkH6kmNVrI9a9AoDa4p9eojPROEeDZf1iKB0ZMhPuXbWIbFfRh/N6w879QlkaErxLXaIPBI
W/vwmsthRucGmrtE74VtKaXR+R9XfW5xGVM9R80iWktAWrMMhLhzyEvEqM4RJk/iFiQrK0QPDcUr
PKdHfnaAOMCGkxyr+SWzv2Kyo1lRO2u/74SxgKLWFDhfvSTzUO+L3w7+c+5+3iNyixWhHTk0WbjR
l951yhQni3IU2qr+lwzxzRFG+4cMGqashNSrjdVL5jmudp4JM2gQY4lR3wRsSRq0Eex1nhUQoO/e
6g+Z3VLxWArVuqzsSV7HDeRPFlD7KAWYtEF/rttuOdbvHcLYreTc5l49MYzICXAoC5uce2LJavNR
zum8Flc5k+Q/UcFs9weCPFwnBCx+a/HZTJ6adnRhKo3ziQTveAGq8Bx8m2XyjUngyBAw3K9/JZ70
BabAAWdpjM3F+KpdwB5UM+czEC0toi0/dZH7RXNzVpr0ql5W20dTy7ImUxUfv6ATI8AVsydtc62E
X2WpaIVtYoOkcV51xja2SNIVp3NC/AuUpi2ALqnT/LFJr4Uw5p/Fqzbj0LD5xINCmek9qbZmivWH
OwNMyXq0ARN0/qxVKEhnFmuXzZ+KCiCqmw7B+RoiNl3fq5WAaE4qFoBgOfpDPTC8QNcvAccuXAmQ
Od7EnT2TFds+vQuk/sx+Jy4NF3DoTjqBt27q+rS3FvnwA+6LCdB7aWxeqR5xpiWhuy7YECt4prPC
Ogxhtm6zYCE/L8QP7GXEmVNI5tCVQgEraIg4DDiQ+CAnPVKWKZEN4+BuSkhNvpK+nARV1pxWpMot
ldzF6H5f3uXIQSDSQECwEQdJs21jd+rRvDGQmCdM930iXvJkypsuijRMQlJqBUjS4LgkgqqiQDXV
P00X6crpwXYf8Zx2CrHMXshth4y0rOYV85wQ+9zz78qAqtKsSCvBeUNnYuQIadhBAlicZBvnQM11
SmDaz4anPP596vhhnho4LG7pBltnUhkCCwAOEl7NVJJnSTX8U1vihYH4E31e7MZccLprtAVCzzaR
J/QQ/DkjwScBqmLCIPJcgThMSDortbw2VEKra2tJpKgmRYGgQ7fwKmZQnEqTykaO+Ti6SOl1XIKi
NLP7ybpUQbAvScJe7Dp2m/oX1UyUNfTuGh8P2YqGesDWouH/y7AQLoHkRMVX12pBzC5cCp2zK0sf
KgUGzWBYrkjFL8zbSaDKLLYJCr10MOUYp0fxixzVQgeJ+J94Y3hlmuIYcTKkW+IdmRXnactTphFV
imEwePp9c2RLyeRqyIqhMIytBLxArmfxp6drDZgAlMGVcxvGKMiM/DZT0rdfi6bfm9VbascWX21J
+Y3IdJUjkJw+vJcg2vrO3yySs9PdDU9peJfjbn8fG2ixaehlO+/WovZZO85DcguDPZLR5g4SbL+a
xm8sTPwvWPGO40H/4eEdAvZe4Ib7NZAUkuVqpOEGzbSY55JfWte/mP74Uu+Msc/z2+Z5f2rElvod
l2tDQZp98rOimjKwab5yC/Fb1EnITAGVfv2LSls6TOBCMuays/hnSQYBawDDPFmEJuuGtFt6+/Eu
IPI3X3sg2aSw+8LAvHPDFLX84HOZJsjGuRnL0FGZTax3VFLZ8HO4ZBeVAuVLkJf7sGs2lnCYgVfk
kHm5gWtfb35u1MRKBsOZvSky/pZ4uasn4yQKihBOfHqaYqxGN/3rK6VcxmCMyyYg/N9/a49zj+Og
jG8t+rrsp5FXbnihYvYrI8DvqmTYvezgW2sxL76Aq6cazqbFAP1U5ppsdtPLEhjInLdTLfwHvXtu
nu7ahPpwXdppJoOpYyIOBS1GltWAdNWu0kOBoAuXTtjpyLObAInucS7L2VQzemDx89zQeF4WFIZ4
LAGbXqdXnhJGq5xvb+igq45WYG7L8qgZNRYkK0c/0Yw/HbPDZ72gHfD7gI4uUNe7CsQ3MYBjfAB1
hVzGy6rVUlFqcXHhBTJ0K6rw52QEhl+CxqNh49pg4mXMBVuZ2uAyoIJ6vPxiEqiicGGD2UHAPtkk
VFLqVZgN4gwlNXdODCUFRiAzPOwF8/VOgZy35GhlHYzS/tmtmXIafL1AQyrJDAN4ypH9WbREMGXi
e5iHXVRM9p6kJmcXabkwNqKGfkGwGRcMhJCmq92uBxfUjZS0nsnIWTXOruSLElFmECyQRCyydPzJ
8zbdu5DWHVLZ5OtoGKkN6ZZ9kF+Y5yjvnx5e9vJUihFJeBp9pqxAbQ4CbrHGo1kalhaaczzO6xx9
DrJqb4jIVDKDosZdrVKEcOhYksyV/yUzRxs13udJrqteXTxUx5VgVn7D94XHtO/fvEhtuffp4Anq
H0KKVjDRe9x0/DGCVm6x2NyN3ejZzumSxpQ6gigfIZpXETsglO1RpRBlqy2GnQK8O5QjOLE5x52W
A+C0hK0PiAwhs//f6xV9GZZzDUyEqZBIWjCoMM6Lnt7rDcT9dYxA0DCct01N/ctx9JnUdn1Yx429
vYItbk9Ec/zEy15G6Pbpu0GoFSYE+eHtm+B2Pmxho7G0mtHvLfbaTKrxRnDJr+CDDolxTYjXv6B5
mzA46NVQV75DnYAE9zYk8XOpoowEeaUESNM+2BCGkKwCovknvqVfNJBwCVyZpGFMp82jmiF/ZKeK
8Q7kVNL2Rerj9vvoaSZQMG5f/rV0NI7/31F0H7XBWchvfAsSkUAvy445vYNfxRKO0JmcsH2UojFd
g1GrBxfxAK+9hGHvS9SHubhXGZ+dsF4s6GBfHvteeGipbkwYslZTTD5eJA9waa5WghOwZh9LTI/4
hOilJ/RJt4wysM/aC1xkh8ErU8C92oBhbC9q5MD1JY/lXJ1B4uC471D/4LWe5w5g69QVqnDVh0bq
4DCSsfgpKjSiDA/cHLqm2U2PEVQGLxex5irCq+Yc3hON0YWgaTTGLzPVrpBeI8DeXNVJ5VoG0jY+
fQVJWvyVIfIFDcsnZwHRyAi+WrhbX3PewXfyDFu44hR2y18fuL68lTg3re5N+dKoXevWglqYP5z1
qd7us7Z0tqMiCJ9k4So6TwOSYxXxPKMqJie48VGl0WN1UFT+BYyar4eJJevPYJbgH8iO/wVs3BBO
1NU2QoSuEW+mvTVBOfynccG5vhjJi/JnvQ9UZ3eOZMPV89wI2DFtG+SDIETI7wyqZMGYWaxHk7Sp
Ln+ns6o6l8D6fYV9Rwofz04qO9d7I8UtM7ijTvQa7aK29FHiTQ/y8XHFmvdHNSZuchiv9S04OC7Z
W0jCjxJonDxZQM9fkn083dv0IZFrcINzf2LCkFcQLAMZ18pHvuAbE1ssWTgoN7Nl3ij/9/M6CSvi
a9jN/sy1mChnH207BscdU8EKnM/djwXmcgFDd/NeoxhV8eo90aElTumBDMIhTrnbhpAxEYXVBJUR
DfUlVhlZQYeTLYskyFzqFyGuLM4eAb1Gd+i/8IVh7xai3tNim3/a2EwaawdDTsLJqVCSdf2wBT2i
uydkg/0y6Hi8ScZfiufja+p0KNUDZ/rDh9yasvkUi630al5jQQrfWK31HCB7/XjqQPTnPFP/BXkj
qjeSM2kxv0/mD0Gvw6wdIJ0ollmOGtntfV6npFe+pD8NFGXp+mtFCVwltqswrV/lP8PDUWjkhop+
3iEtrygbQicTy7621SpNmfW+gIGmpegEWYHZDpiruuFuFV6GopC3qyfw2wkkCMRrUeQw1BVhiYN8
j1VJg6NpaQx6QtXyKxycHrnU5BgS+YAYuuouLgU2dBnzIEb3YvnhBOHPeJCZh9q0rxgvcjeNP3EU
PYf6YUB6XkUna9pBOZUtQj9lVcSc4ctOeRAL43+D2oVpdh9YlywzoXlFSJ9RhFZlSBNhPdFSBcDt
ySDjLIu/BTL6Y4Tq17ylD4M2/PqBd67pNrNJb29ZmvVRPfTTjbzJ3oCnONkxh41V2mgAG9Jx9mLy
fdEh7s4Eaq2b9AV54CBaQiO6151LVBhLHvyCInVMeyZh7fnd9gPbOzMs3YoyPcZArhfl+nKn2ksU
0R8CRM0TG0fA0R8PoSM7jtwb4vti0033IHMfnto8L2qsKYKQi/4iHgg4cPiIlh+t0oKgACgFdj5S
4xvo2rzGHHo5zVvanTba5mUWnjN7M6MCLzp1yDfbCwBvaIDRXbArCUmw0ZTutroMxd6buTQuqnZI
OedQwAFl/YA91oCMeK3El6MDaZoWtfsdwIZkDABW/FWHLNkvrrBntIuJ52yuLJTd7GWXKqQjReA2
EPABXHA1bIT8k0gAX+kbJNIqC9XA1ZVslGKAi+vjcDr/475w3SXBUxVcvxfjGP8ZEEa8jKz8oVx5
uQP0Ca2uir9qOAmQcsTj1B81y6Qu8A4NAAylsb+zzdHUI2Mkj3je9uMA6iSx2gY6VHRspz1TRDuN
exNnYum+hIydaoezjrmJ42fQovs4vqwuyDRx5bF/sBZHxlxH/OG52rLjOeFuLkAW/tDZKu+b4wHG
xG6CcshQFNBGp5WYpCSW59DT9v6MRp9qjocgIuj6q1uF/+2QvmDUOAF7QlyH2q1SBD12OIfs+AyH
lZWU8i8DQXVLOL3e6TMBB8s4WINhjQ/rOg3m6wuhU3lYsGajjpc3n41tEzOxozfrV04rjKCiDhdm
my3v7ztFLiKxGz4Af/wNfCEZDkwUS0IV8L6Amm9hzva9A7ei4xxUDvjUIk+hDlmyCbIw3hKH+sNJ
7pE404rLumdQg8DFZu5yx39YMTdCLKbROG13WSLE/BnfM8fRqpB17UG4vEbblC2I47BdO64SpQ8d
j0zLisqNLmSw0RI6Q1KLqfhQZKhwKvQjuwPRX7uIpjhK9OQVbRgzYE4knEWQP+onG4B5LX3cRrMm
GeegYnIo764ca0Ph2kSIHBuWCNpJ0flHyn6A3plvY0lM1G6v2jhAHDIGl6PhicrOHmiu9Ae+pHaA
a1yeFRAk75y3lBxfqCMIDUfG0u0Ua0SqOcTkWhTU2nX59Jb5hyuzomrT7ASGYtHriIr8X6klaR6t
6l7siexVPHtzugSmJ7KuQrFrIS0PvBLDL3vZ113zE8hAgdR67YHDwvitVUAjEBGiBDlDsXTYcvQL
0ZoTBZqev8GrWUmpz+loEYU3zzKQtG3h7Ef0xUhIHGh9rOTslBf48mlhEu/CZhqm2HZ2W19a/b9J
a3nf36IHTsJQgUVykPT8mGJUKFywUufsJo0i9iX9QkjPZwxs7+Fk7dp4PjrGNzcq3c0XbC20lUyH
k17Xnz82b5yAJ6WNXibkR5W6lbbUN00qMDMmPEGCh3dKr7mPBRDYqohJIf3XRBJPpCa7Q0g9aDAd
h3dmJ5zj9VUckuc9jeQVlaB2FVOh9Qf/i2jyAZHXYA/5JpNZRtoklBcY2H3osiqyYs4I0hgdUV06
8TNatmwgFKeVpaqgwlLErnmzIT4djpsvbN6mAchiw6AZpHeGvxh/O1WxgV37cK51xgYVqnRVCRIL
F/ym0UACoiBh1uJd3XBUQBurBJLwfsIq+0Vm9jLJiuyZfH1KInPsYrLJuZZTEV5ogjo422oJPJZa
0GESSqHYeu50Er7CPzL7cBWZLsTagq3iItOZKFaQCq8ms3FOIaPq8n5oZAVUbnvtN6Tr4DSzgZNL
QuI6yWsEiSx4SKzx3+0kxqJ5Zc+UMeKA9y3tAye4ETwqHk4nxSJdh0LixkffgtCI3+DUtJ8v8WNq
/WQg3/KO8y68nD9O44KosB12F4/wdorPjMzK9orCZ/xOi5EnLtE2ntZau+2zq+v5SN7RUMRiB2sL
hthGceg4Ah9faY0X0IYeTRqN/Z6An9C4f6bEX7n97a7nE2R8/tQlc2H6CntTTyEw1JWPPwm91Pvd
+0V3aT536fmN/fibodONtTMPuS9KrOgW1YMdqyQff//BvNIroun93vHykWYVIWogBHPmt50z4Bf1
GeFwmTkhSN9eDmnMePYgEheJdirLpr+OjCb6yqzSD+u2VoH2euQGvKlHONbQYotv5ZMpgcJ6p6u5
1SE5sRG0Ay5sDotXEbXH5dEPDw8BTDepanQpV+SIWl5y0LEm7E6srDoANuG6tiDpbvZdj2hx8Kba
zSQAS3FUwBHKqk4UY/aeUGZXDXfkNRMuxBIeqW1tPsmHYwe9v9CJ3jlXaTzmDCGk0pHBS2MoiRUo
28Q6IDUZZ+k8Lw1tqvn6GWke1NLLT9W93rgvJV6OrFR6bCyJ2jbNDCkuvjt8cagMScJgTYbFtE4y
aDQjWFLS1tRUtvVG0wU7ZH0nHQc5SqXOS1VZsCnJE68b+ghy6hKT7vVR5T0jdMfqSJ74P7hIL7UH
u1jrp6IO8ZKOr8Wu9l7iz804wO0zL3K/72hkOyARvQT5o4B4l/R8txuFAKQ03iWnoK9guj9JQJc8
wxQtD4ZRjhzQTbQ9WG3CVTCk1NYlLolfSW6AdSgQBrYcgaX6fol2h/p2/UncL7dkcbrTQLvFvdKZ
cxs3mOlcDfJedI5frx89HGjwhxQM1a+o41vzwAba0gZ2vHb7TVvVePXAMa92LIRP+4pvbaEQGAjI
Oiym2DFMtYbeu82FXHmtdlF8mfJH7s7PiXQmyUai70GdI+W17pwKHM+UrQYN6ldLQG5srOa5YU4S
E4bDu7YTZ3KYSP5Thz6UbCWmun/XlJGMddfEnWnOuaXNQT0Vw3l68ioP3NNFK3AjPlLRQYBQLyUW
j/6TF0yBTfrWih9g6o/CB/34+bArA9uhiy7mZsv9FVqbfS/xwPHkFr8aC8HhYZLjYV9Rlfu5VoOV
+9JhhsGYEZ9HkSwCu3cQPHUlI9etlITIYdSm09EgCVzMmcupuDZ31WunL9hv+4W44aQ6PABRb3Lb
oQuauYyMEEwsGyPVf/bTbmPQdc/bEDkeytGlyO0W0EbXWOHM02wxJe4a2D9L/yoAgGPFZ3KXniqY
tDgxu6rchpPxG1dJDeDjx4x/DeQuxbpByON8vsRHwZpUsaE73Nu2y+naXfklWrvVkmNXVW86j4yn
NuMCpN82/lnTJjUl0Tc1HT/OwWtyQBcplbkR9EoXgRsG4XW72Lgrud75Vrak+yWZfnxg1ZuntfqH
0u781ND471oR3oJkihaBDdXCG3An8+8BFIR9QcFyL5fdx6hYr6wDt3oCjBpI3JJorN8b6exxXM80
ZZO/84zG7HqHAAFzMqXZSyQhjNHbx9h/opNAdMSITnrgNcQF++k+l4TWAjL2Og86giFYNpPPJU5P
izY/5rNHkNySWWiSjgU4SEBRiHVs/cQIy2SkDvQmCdATtofhbctUw0lqH1l+FrXrHp24z993BzR5
SrDgTbjKBJOj6gtOkVKEQ+FBZnByce+9WcwdLMgbqYMpURAra0F/VXKN87w9mhNX+Y+V5oMXQhHQ
lWlTfEozDmc3OIs2UYJuEc5ui9ZgQDETz0uhb1SUi53PqfZj7cfDQet7mUw17900lIfNB/zvvZ5A
El+0PV0p6Wxj4SREWiKhoz/T0VXzxPDPVRn1m+ThoSvu5oT5BVF7MKa2/5T5YnQbo7JFFk7JAXer
VhbK7wn5D/5OJ9ZkXrIgkPHeHNak4Rei6f9KzhgLEDnEhonRpWyXyKf+BjlojjIRzemOsSZHvAh1
1iHcomTM1/LW39a6vY5S1+83MxHdfycF4AD7/LVsNSqax7Ir1qwllL9k08JFz5Bpk2u3Gqh2lx5i
vpx3U7Ef3wt8aYQ8FuGbrCXYviFZNk0ehSvY7wteFuXPM7j9wXW/39A/UOXU6A+taLF944gemvjA
KeWFmdsK9RZsw4qmhyKKSALPMxsIVEp71/aUHAIhVxcdBmgPpMlrtauPXAH4JizdVcQXiNMg3WXA
C/jUusV1JaZUzNcKA6Kp651nUYl8fmZvJVvJYNXLkxxvkMNiKic9XyCgQb9xODMihsyltfb7aaN7
xhdHtdevbT3NohqZeOXUH/dAXncQoIS2+F4uCu6JCAv2WxIVtDgLQuVKgjBy2O9HUW/mfwgYjvoD
+2tLTJlrFBsaHLVeCC/X4V/QREULqLLLAG1aWnWhr/vRGkQ9+7YxK/JYdPqMjnrf6BT0Mw0YU/gQ
QRPYddaHvuLiQMDwlu9li9VK2dteoY4AyrHdV0Wim4MszrWlHzLalBo1IZm5jQCExd4IMZxo+kPh
YTDZAM/FeOIcvxdK+xdvU2pHxw1AFFeoWWUOyGRHS3SVD5qhlFHfa/bmUukv0twyWuNqOk2YKW6d
r5tObYvvsFCQ5Jorno0v+7K2NECoZWJKAgQJFcdA5g/+7zzv7ZSpnsaxrmfpI+T12hpza6qselEu
5C1DURle6yZV16/JThpoCbx+daNPTDra5BLPyhhr9OvWnwGrpLWs5SG6nmrF1P5qxI0GccazD/BG
2hnA3OwPhNsNoZDZUOluJt1TyxrqJRt9KFvDtssNN8Qbe+E+EDtjgqiJwQvnJLwnd7Fayk9XOj14
IAI9uvN1YrIiOTHys/bbsn4XC0anUgCx17fdLxPtr/Xdr9ykxVihB8Koe9Ey5YhbFa1X6kNQ2Ibp
wiAEj5togq9Pf5MsIr0oOqTlE9KG/rv9FAKs952hfKf2l4LcFhHnurFMY9Zvn8QIGIlqy6kqMBqv
nSECXe35JEy+apSoiWkTMMDWerjza1zOFjgVdwHtQ/P3yL4klnoPNzZLyz7DsxKSOPsDmCUSYR4s
AW3ER5LeFJJchT66n2+3uN7dR32E/80yK+OP0WRFeTp4VaDK+iRX5UnJZLWTw4VEue6OzFsYwa+d
g6l986zOFE5MYd3oTufNr+MsOnqfhbSjk51RHftSv8Y/jBv1j4cgujkMRZhETnF9lU+OjdkVRT15
kCPxYVZC9y8gdekRVgtHhbY699I9oyvOD62UGY8sTV8/x5GDtkvg232myV/EONKtOwag+y9q3QO5
oMFVowy1i38VSt3fOyf/zp9jZCe4BaydV7RMwqFNTSDcvfuzhqjGmwW4eQfD+m1B5IxwXDg9l80Z
Riw0v2Z0yxOY6RNxsMxRoYj5UI6IUdun2pqFYq5Z+VlUR+L4z9AO7T4Nq3g4PWZOgBuKotcJ2HSn
uzN7LwVEPKHS59vuqO9ZLc2gqRVN4CINlXA0g81Y3DcNi4s8TUOK6+XTXaNbOTf1qog8O3AhcNOQ
Nh46SUqtrj/VGEdhw8bts9r0ttoQeRkHDkJW8Zs92lTegG1hEz4yrWqdFEZtcloPi6wqu7Xp/N1O
T0BgM5EBXFe19g79gYVfd+88C3aCk9teoq02DtirmLyObnjAayyX7Gk811msJWDqS5tVpzCIlTzP
MyXzXaOnnde/q9m0Aenbyhyh/oaCVlh1L1vO8yFxAP8mvYY6QJDjgX+YgromDLhjbOeKc/tE0UQB
idb1lBElcz7kyIIBzzryAW4mjjYLGF3NGnGjdYJCFsmR+vDx9v/tuZbCc8ZUd8VBFjDJgQVOpzGJ
OTQYOxYkYHNFL6te+8098QEzbB9COY26W8F48Qt5EiWGb12F/WwWae7hCRisRYP2fPUSL4qzb3IV
Lck2FDf0koleFrDgdisgrc+3fdQ/EbLwMl5vksmCTaPb+6Jn1bXUvFQJmNf4iirXWmK67Z5Qpx55
dLTN/viEH6aQjWRsCMaZBgBXce0PLudy7Nm+b/0sw1W3w1PChA5Vs04DDgoM2QxQXImP8p6mETaf
LhVsAkXKljGV5WycoqaeUDFBPzyp6tdpkd4c2su58id68+73ldGodRTIuMZIGPG0j/B+JRmy+p37
8OCqRRinqk4awbK+6A4+2PcvlmdhkJgdzzAmNlpA0dyXAuYbao+gD7bVv56Ehn8srixkfqcuP5Mu
qnbVN87yUyVQ3yuohZYRKeNaeLbEKAE9AWo7P6HMx1Dsmle5IN3kdF99ag5KHE9wgthxqOKZfrU8
/gliHpMe4avRosl+Rvu/WWI3pcfYNCl1JlxtNRyLoEu6oS6AvtpkQMrfONaqqgC3mfOU7ipYC16b
fMAsOt5h86I/NFems6I+4NWgkgCP5igTLV6K4UjB8AbHYiT5QIa908Bf8RD+YiBNuO9j3W37Lngi
9kBTtlUNiZ42N0erjhth+BUUd2Z0mYalUNQfzGOcOPnwsPmV5PUYfIZEbNjiZqRJdJh4MSZoHsrH
VJ2rklOy1I8szEKNGvInacc9w4ADKSb+ErrmjzWr8a3vPhkLqFEjavDkbl8nLgRY32Nd43xS3PFf
TxojpK3R0FUeDKbXOFJx5x1dX3AH+Badxg9/5wkS0QLIvbRW9hI2FdleSeUTIrnnr5yNx5wayEP0
6wBh9AnLcJKeb4OYO1KN/nacdsmaJDFFmVnqRj+renjObjYlpyj8zay4LCvn5kzwqiQTAmcX+iav
8EJI3gsGfQp8ewRKFu++s/oygr5DiyNwo/QIVcDiaRcemu/VP3tM+e/szEKSGThEd+9pLy8hzQvI
HztN9NNQ9Ev9YRtzOXoLbMCuCh0xRv2kcQ8ZS4NHGDDJ+Zo5n8zC1YbnHcrG4gE66seSksE7YWyd
oEhQ6Kec49JH04VnEmV+w5Ibn9Ded4q9DAEp7xFIbKLKQ9n7hNftA0TEBPhXaM/LJTTILoMZDLPs
6JN7YC20MIrZ9/k/TlI8f8klnTJKi2mrlBztwwZ1lUlk01dU0z1i0rlWh6jJT29kIrZAkCj/7FnY
uIf6E45r75ho0mX3ZQPuTIP05h0j41XFZBuxOOOI1PgxQ4mSWeXJ5Xn+zg/gwDQoJGIicSjAqgDX
XsAs/4BqcMploxugyFiDEA/bIfkCk+IymDoEuS2D3GAgY6PXhPVOP8uDLao2F75lwmHU6l+tGLA2
2k/MVRGqdPAAwvOkYf3wlbPbXC/OPRb+mX9DyERZ3KwBAIXImBaRilHVHza9mgmA7rc1zHkaIhkq
1PTTQB5+IzlOfDAVN8/ccwhzKb+2HuMuIFl7aqkwE6G4CNRZH+JpvLFRtZKD2J0hi3BRBtWJkr6z
CCRlbq/BYmnoiqQPZ9T0mYcLznaCNNbdiKsJclGf/c1FtKknAdYnFA+NISNfhWocdoElFDz1NCri
3VD5qF60DQRVcVaQHrgIp8/Z6bIuPjqp3L8iIkTHega7FIO8g/WWoiNFH9mxOlWG/thx9lmCxYOO
gO9GOyzfmThzGlp8lcwFo/CTDxTQZ/+L93aqqXhh2/2BMiHNsZ3uKjYYFA77/kzHZV+qiVbz9M6g
x+MSu6Wc5g3z3N+qUEYQ2CiMZlGb46qSXqnY+JQsnpbI+WjnTyDH4THOZ7k/Kak7KaAVRaGAoRBI
hr9+a+IjZ28zpZmLkpYu5m3Gyt5n1DOvi4bscGUJCWjZ884QV3Eu1Oon305dLO/QVMtuqu5xSQKj
vSrQN1s7tHPlCvw4VUlTEpdjTLj844mEkBetxwjaCtjKINTwqOxk3fIholZiG6xxAMLU/s96n330
94fIdLKm9ICSfe3+znwECkvJlOe7byKH6b1pk9Ky1mUwDwh6PIlMcT169+edW4sVDXck+/k26dL/
MDyFvfKulwMEDoumR5L0VSa0LGYqM0L/QSuzSe9ceWkokCTGyzqNBFI9EuXsIBWdwQLttIH/WHdx
C+Dw5p07NsBih8+GOJ6bJZgOkyeQvMSnVXgx3d5QYT5XmhxvUExEV0sAwSvhSLI2AMcrC/k4VKlD
QLE9Pc88Thrkn6hT5xEfOxIxiHGVHfTqrETdMDrHc0BkhUx6rJwK5dXKPMJp1B1Nldx1lRcuFm7j
rg8ZSv9UPNmXIebk4Gz+NVu45RI1jAbsH/gybHo6pM2RslxjJ4EFfbD+nn0TF35MOiKu4heJcQYY
ipvWf8h1VqaCmaersTlPraxqBF/y1+/6dIVE41M7wKP18Zaf76FIayT377oR7GQNXjC38rA4P6Wt
gLLat3aVZmbtH0lsWLxOacjTj6qY+9b/48MgWIgEjHFQoc9l5NgiIEdwh8ufA6lRgfX73nozA0ZE
RxRMygkuI4kBKLV4f6yLNQcAlWzsfEIuHIrI5oBqPt74PnfTEXmyPjkf7f47DE/CHRFxbk7pP/Pj
XMX+Z8YPcNw3mupSLwTyyrF3dxznWT1mpl9X+QhXAfHGKPuw9y/+zMtjLPCpWEmY2j9KwjENu3TN
CQgy0FlF4UdE0E6oYTSy4nf2jI3CpywbUj8fNFykKCnxnn/xYHdIDzJMu6xFd8143J1f7y0ceO1C
Lk/p9j2v5meDtodRmhkiONDLrO/8m9Y71IPSeMo1Bwub5seUKWlQ4Rqah5Dm55j3/5d2VTZ2zzMi
hFHtH/5+nzmufCItitOHIG28/v6m3MKj9hpCvQCiQUCoDzzTREW+XUxS+PUJ3ECAl90FgCU5Vk7s
JK0En2XKBwNT8x8mFs5XRsiMH6JUEHQ+b5FhWfQ149n8fAUaNvhIN3mP8wdelDmEt2u/Jd5dxkBm
OT4uLQx5rBySbHarS7mqOB/ygK6K+XIIDPEgFslYEwydpzRNrDf5DXKj3fBptVogUL5mFdDrX01x
RhR9/wtM4pGHYDgaJcKKOkhnjMqSH5dE4acA+TZVNSis5K+etobdqwYApboKdty/bkWhhemV++QX
5p7Hy6BqVE1X4GMg/682FnR/YqcsxJEYKr937K4HIo+glliLNZhLS9MTeQci0h592YzHppR51Qb/
5zbSDSsKQrfizrUxD9IAX1WhEMDUXoqhzzQcCgEfae+rjbcJkwWt0Kc2qqsqgaUzJlC4sU0eU5lx
NY4EVI0jyomjOIBYIrxKWMjWYrqaAtF6GQPFJNTW9xD/6/EW4sWijTHVw0pK7FjTMIP3wKnP53BO
A/iBbhpjVRagny62YmX8/caL18t1g08bcEjMaUgiJ9jrVA+YYQHkf5svDBfYNSTNoUUm4NERotyb
5MswujFH2C8/TDQNebT9HECL3tOpMQHonYrhs0XocIDSAvSIIsLemHhzs7glqJPFcgWcy0AduJFu
SYgBbHbXJ62djtvN2C78Fz4NgkyZ2HmcSkDTUgo11yvh1bImgCWUX/ZKQG+BcfnhIhElUkoO3AX4
dNz5HKlMtQEr4PJnEk1ofFX9l3bGcanHTe+W3FFl658s8d5+nsjeioWMMM1h31HjB/AgVHYA0dGz
eU1ezS67+Xv89W897NZLPRRGas4m7FVGwmmRBBjo1v6XtxTd8JOkVrVp8s8BRek/8X07bEBg+dta
DVglKCeWR7isGeERiTmutrbm6LTnzY7+yd8hbi0nxgfyW8Crf99wzxUE2VljCSL3XrR2fKFug5ZP
tqrWfq0Q/QriuSn1hnueddNDXqSrqlxtY8qW3F+ko5OlwkvkExGq2t349jrmACKdj8FjQND+1JK+
cjRnniWZO/DM570Pc+4hiYiQeaXPaH9nryhQARBFsX0jyRTC98t0DOCYY4Hq56EF0/lrxNKCe+le
+YOXrDrKyrRFNBFHYtoyVwl7sWt6VeE4drGfQe6La244iVZPeE5i/RPwXZbySbxbsB4GPEDRd8J5
8z5zbIqj8mPJAnTO03JMgWxApXd9CxfKsMCBch0OGYOQcHKdNf/rB1V91IMeDyODJu1pw9u1dJ+X
n9li2g85WF4RbOiJRIJssjp/FekIFQqStZAx+3PKbjIwBJH8dwseLzAmvx/txwEjpLHuxZH3LzR3
xtIeV3u9XkaKscCaQtayd1VYNucOBE2U90nONlnTGukIzdhEaIdHZqKDvkQ8upnhwj6pCSQIgLUP
c9D1fpwYxWgkaqgHdu8vsQy6epuGII9W0YWvOhZe0sX5Qr+y2gwFE1dCHvkO3MbDuaPwBucZEdVQ
9SRf+Ra2LAqu0R2sDu73CB7gmdCjwEXAHARVVqW1UpL4wxTkKo5bL6EeReX2agMCNV6jSlcNuUqH
uORtzK8iuvYn7ZzK9JUKtJOrsxq6QaZ31h1L8En6YxSrx1f4wOb1+eejXYDnEMLM4VEBUs6UYGNV
hJbsRIzekOV4969GrLLI2ZW2YKANcapFfc5HjixmOUSVjajBWRLGO9myWWx4kFzkoxxhxhi+oS/n
jlD6KuJpTy1Kt/QgY4V3wXHYikvJnvrcNrhmAcSR75ZgTdLXafYAMY/2uIgpeCzQpU2N+QMZqPph
oIsSr93BwnRB6ydfObCfk2A6ngaEV6Bqy0296kCGw2kfR1QPXHf7D1A+X1siz9768JT9WWgrYeuq
7su0YnJCXDwJLnuMPJCGoHJqFgcTyYWZoekF7QQjM/SfzgmQWI6hwVTa8hDHxSToBku00J+THloj
eYI2NdbdNCAuTItYC8JR9JM/d/ojzqFfXoqKhaxNMgKjoxkGAZ9RBjDjhQL5G9wM8VBooXx9UynO
r9khnx0dk5IjrjCDcO/Bw7aTzelVXI2phRWx4nWO5VEYXKSRAFEqyF+KV53OGxikr8GAxlr/Hy4J
Q7oHJFiCe+tyUimLuJD4Lrv3EcH/K4VGPZKxBsnIxI2Lxmi+6P0+u21PqLHXNrrbaM8D6cjhU+B6
hENZ8+aL+7divhHGgIDKQbOpn2t3v+OC1fD4tfS0udLeRsoz9BBHws9OjV6WBfUaeYPAtawqxnIa
BNLh6yA/NGRdGd9bEWMpbpNH2WQyZj/ENfXqcjyWWVMF/x754qZylrcQ+VBN0NDare0ywjL8ItM5
r/X4FV/OtuIZE+8dBxA9HYzRNwnX9Tzz5+XcplQRg3zSXmwSSBGaZXtzJJyM7To1tCOqz0u9acqg
Sy45Irs/XrnLDHYdh+BOGsii+dnc4DtRF7gxP/DNy0xKTop5EaZJCow6R8VQ0TF7OxdLaXX12dhJ
HNHt+RR/0CmZ69NqddGKPhvu4BbLYUB6QlGnd4xCgYS9YSvsZb8RM43R1lm+7D0FmeFNgwlW4vZ2
NxZcd+czG8D8RiK1uX4/Sr99lR4Apu/ZDdG0cZO6viL2DVbkCp+Dzd3t0Hu2MVWcGmjHpV9hhtpC
MyVk6448vA870QoMXpcOJC7rbFHFwq6CoRE/aFbtaCs9Tv/F0w2GdrD2o+qdPkH25hjY7IPAqbh4
hipsqX8MaVwkgGzbCaWhUvKS5/tY8TU5sH7yLv2wzLWsE9O9QLaZ3Nn7oYSU4lw/NUPSdBr7Ah7A
M+f2Unwa0NBcd4IaV2QNvKP8IdteU7/im7zOrLodZka+BGzytP+y7IQxHk+zVN0pu2rP9zx+pV1n
HjKInfUmBhZPc+/th+f08uRIg1mrDfvLEFM+XiNT+kaX2a4LDGk+jHX2TNqR9EYCpNcvGplwoCSE
2yHqCrNR5enG5Im2SH40NlOzGFNolYs9LuCHtcGqFRsgkypf2KmoOYjjB8m1yAaeXU0m+buhXbhB
lzs6SsZ+zeqBSZiwpijmQw46P3QWCDTLZxBe3wQ+zWFxVyx070akjoR7cjXyjq7xC0QOcN375ygH
isMiiAg3GgoLmg+mUiSSNAUgq9yUAVS73mZXerHE5Fu1HfHO+RTyylveXZ390TdhNoAUINtmgM5E
7A819a57Rcp8AMAEqJNy5CcJ/uWrwHztz4SVqYUZAuTTl8QJmioOyfWbmB+P/Z+kG6gwp7Hqe5CD
GjTXYVOIJksjo94MrzIXWO3eY0qt4Z0ZLWSozWow2ux35hGBkYb49FxmyfM+7WUJs8gsdEgFbUt7
QvId8npwxXG2j751ZCN0P46inC1H73lw61xVpUAZWsfGIB3p0JymR99M67MR1s079G+gDoSzH1nI
zbWNgv3fJ8khp3gqngY8IEZd9mdGRhpWf4Qnt78AVBSAFePmCp6/dsQb1AG/c1zqHG3umC4fMYXU
bszdfQjSlrnKtADZnlJtGSOuBRlrTe7u023hmLHhomYXMKpzMSA41WaX0hrNAe0bmoE8PB95uhYQ
9tFL9Kv3UhenP/7vwvra+Qf+LojD5fKvAggfIBGs75Y7+m4AprV/a80SlGMORDCBzr+lv47PeojG
232hZKdvJlTF8gaon47LrgEAIs65RZki2WiK31/ItE7zmiFpwXvUP+tsULOFjv4BUmVviRILm3Ws
n7tVp53DKT+muno7nTaW0YxFo4lTHMx4AzMbJrnv3VburXwy9B8+i5esVVQhMH0/dYqCAUJenaTU
wzxkmhCIgMTop6O4WFZZcvkBe2W7Rb1/UOBxlJztYC7smAEIhomctWIDpeG8gMkTWwWLVEPabcir
jWuzDOSSbR40LcIGHPrwNASq7nva2lgL2AQUoDtC6+2jMC2tG1tFt3Un3u3BNj0DN+hL8B2kKeDJ
htmTF7rGx4UUCBSUGf9MfAxtEHFLj3HQ69sSfLhvQKwNFaTRGZ7SPfbkAqyHZ9kFqeJKa4p+G1B2
HBxd7D0P8JgyUUBa5alkXXvgZLqcyE4A3/IN081Xxd3IcuTazASjyNBPCzmZuGrB9Je56gm5N6W4
vfLPwufrbVzeJDE3ovhqC/AUuUq7Pl491qX6anoQpCNeiEpvXSOvWxn0jQUL70n428LGWDZPMa1n
XxCC7NLHFWlKq+dFTs5OppD8c1PHF2NZpm7QenK6WGO7ceoqNgaZZVu7pgvvAP1qcGynLWmj7o6t
Dy0ZNYI+r+RmzscLm6fNhWoTti6aGxEr40cBMRHkHmtdFEPNOrfETfTGn7xQ13cBzKM1jeZa8p+v
G1w/46eWkwycj4+VBGByBHSTpdgI9dppm5F/nD3k4za7WjZvAyIxQGCBfpjU1IkmgXnz5aZ8F+GS
/WrC9D53T1qHh4wkjlVgGMCAb54Rkmz4HT0893p3Xygw4dV9ek0d8uW5pUy4bHSIqLlE74JpWULv
M2mNcW47FWWCyQLUCgHHzY0GbM9I95Tiqo/3Xt/Uf5+dSEuEhUkzTKtngFWriwXb8zYUI9HMS8oI
FpQkzG9jT6F7xoi6cPEcH7UvnIvFN27712N5Wya3Kuqgyl9EsyaijHMHxzLDV7uxWLbWyyIyViug
r8sDLnmYqbezqOs9TTKtrSyYQMj2UWBdD4UyeI4oCFRF5/RWKBRuzsKf1Ipb9oQz3/MiZkEkzkos
fKhUn1NeQmm5XNevV3tGRPvI7IkJ8m5WBsdNo27jDwsJ4Q+GQL97+OnlOmu/8Ht0r7yYcXp3ajRh
GN8JPmXOrOqKqie4R3T3EV3NlMVoO6+l0mCu2jACtEAAgoqu5Veq3ru5SGUETsL5frAA3hcnvbgk
d92XoWhdjDH7CGAF5SZfNSvMwUKQV3+mkQrjntkZau7hq0r01CxwbVDpHY772BqTSI1mhjhryuii
Iq84AkCRg8lfjDoJICeRTshpHgxATNvZ5gBr7KvnV3bL/uBO1oZfNhDVdn/D7HTJm9F7JlHqbIMt
4LBN1+8BC43UQbBlnpaAlhemT2YCPsvxCGk4XyqyGHQKU6lkigR18GPLxOojxmkqchmAT3SALgBR
iLFDXFOYoXY9VIzluWL6TVNcE/DXrOARjGT+o1NgtqtOnHeOgvtWvD5pbRSxfZqGVIQxl+gQ5gUl
vkuq7bRm3x1mEx8I+VMnqhJDbSx1DKW/E0umuT6sAfPind5Q4g7yUD3ZXRN1qHjP97vnZpoZdAeA
9Xv22xe/ZC4Zl71IBI2ZkA8uWuHLe9Q5j0wkPxB8FM5luyfHxOnqJN6oLC/1IaKRpSOflOsN1gPD
w2cKktXbqcN+bw9PfL+cJ68XMsdgvviX+FZIWaovSDNTNXjYEU6cUEud4gpdN+VdaUtqHOPtXDtr
F1jgONKv5eD5CWG36gjPf5GM3rVLtDAh4Yq/CFW9jjdaEWLGTo6iBrD9OnbupixGXrxmglvycDSQ
gK8e1FN7d8IPwwtp1jJMJcjit9OPlAKWVUyANq3wgEEZmtD3V3isLOfyTMBCEvkMesLRp84Nw84l
/HoMoHACDl1cx3uN8pCXRmjJjHeJWph5dF6+yf4vFb3rURc4IVcuIi3UzhZ2fGnn2Jsx1UlhqmEL
ZOyhLBegJpNvrkubCK8VB5qzK22qA9LTiBapdIYZBJk2Hl748dEFIZELOailNCF426KdiGWu5wif
+GW7+I/eor/AWTUxXx53zYtsqCB9Lu9war6hf0yUh65WiTthgPUkWVnU6IMqXTNPoRh0QiBOG/Eq
sgXKU/wBcs6B7/k/XAcmDlliCjXj3Fv6SjfQm1z5kkmuqCSpHFN244mI+aNrYkuZKfKR40PpdnRc
eqYwb+vYu7Al3nAXhUMpgUzfcgs3ptDhSDaJrbzqJBL1gHca26s+9wU65WpteaT9SkKho7sd5PSe
TnsoLTH/lK+weEiOfqmojBp4zVMSBSC6uGQrfd+pKHB65B9AQRjqTcY13soahVeK5XaKPfKrMWps
WGg8/j4kavvGIN61k1IsN+2lX56v+m9wbZ54CVNl0SFY1B5usewYpSv5t4fzCrQ6jq3cMh+cqmOk
BYa1d/39O7nbDPSgLz/dz7LhgLFU0sNt4W6uKJSOCIKgqhon/EWnxuTA4zcq/cVVNqHcWXH8/znt
iEbe00+W9NWwwHz69I1CAhbEmne5VU4JN0cKl3fR0uX5TGqE58mbr5l7dLEmZ250oOWC08vK7f8j
96HYmoVYfvkZpliz6xwnHAnrXKhwlR7sYsI/XHzW0AJjMsUfmjU8T0ZLQ7ZNeKn4BNrkgC5bvjoS
0L3TeGNg+P0rnE7NpVgA4BCON7zKG/5xca/mniUEw7raX8/OzbM8Gd2hxTh94xPNQn6ui0srMISf
z5ExseeADo1qObDpjhnWQRNhzjWLBquZjNUS+HI6YF0rBIcAo+X2xArG1Fchgd/f/psBO3CMQrfT
GB/rr24XsASzKqqMiAr+6eYoLInzSNb0FWCgX+8WftTQHp0IkPkgllP2skFP/KOrZ/XyOv1J7J9k
eu66fmcHKwe1njwdPKaqmruT5Yb8CL9dY0zm07q11iBaFvQAyMKMpqiSFAOHJL+DboFq4Xj31vXg
dl09Kreeo8CZPcF/oXYmePz23/4hUfgzyQfhpH8jpV7uNvGiphv2FNX3hHbaIco/6ddr7vo/5Yhg
ceKh/hoM83cvtGOooyOBz0ffq5Eyegtx16v1dvGQbN1cT0TL1NatAt8YrvPs+Rte3Cm9lrAEg3N+
b5JGUB4VbP1peRHoxaIxdItAXL1YAbSftJB6h+k9EQfiech8w8mG2mS+AmuYbUl+erJ+8LX24wum
QsHI7lgec2AU1D+UI5YLv7E9cwYYzIahwuBO7Cocvzq/Lwj9Yxn8wW+m83/QA/f1tKhRuv9XwFa3
cNlRFtw2AUE0HF4FpMjpueHzJCCbK1/6l3ffN3fB3zM9f4ueRZl0sz/kvzoq4AIhpeJ9fAhkKuHY
02SqWj8vzlnryu3fnuO/gXJwRobmoGtQ6BuEDgS9aQzsG5ag307PfMwPLoAA1lkEvmMXncAonB+m
18ApzIoZJKZpbHdy0v46iQk8woAoQdSPB/SZaTCpmJOTLwjl/gIuvvMmGyxbvu+qNBlYGr38r1fN
DeslA1r/ekg9cq3mEPI/nmtf1g+ygCAlX5S4+E1KOv9Lip/6847kRkztmz9TliQw3y7tJ8Mw9Rg5
oF5gGBhXV4+Sy+ve6qZmVwtGee2BGt3O9uDwKOnZXS87vErPqMaB3TMKyUoB5Dd4bYZ7M8Cq1Lro
awl4ppeTZ27O0wWMynhuX9NXUNODbkFH5MIpaoUXhk0FMnKdjAVXGDaaeaiwJLNyVt9oGd3Ljiaa
rf0F15tzOF4OsQSdFrViRzdMlG+XjUeVFIErbqxA+zta6Kc0spA4DOPoPhuDqLG2qUCfrRhALQue
lOcNM0LiPmJNggt2xN7CU3poy1hmV4ZWLN6UfevYoSVVoi6GjHl/IpEs3tmd72YXkiIO4PtwesA5
1m1UiHm6xj1iQavQhcnD/Vk4LqE2hm+Hl14kdPgMFxDjfie0BI4ylH0Q6XrtkkirQDmvESKEqu0Y
NtrJc9GWsDG1KR7nAeseD8ukuJHK9DC9nkGk7dxoqjq5Sme0pGxW8MPDejVkb5d6Z9ym7dphxDbZ
tAcQ19tagK+FhUMW/a03W148p+8AUT6dvpwUAaJp2RefKgbn8mFw2jDWRHnbKaNVPG1QN91xuIHb
eDpr4G9wpudXPlYf6MgF3oSHgz1GHOhJf2lG7ylZiCsEcr1t1sgG1wjNKCzy5Y436aOlqrYjh7sp
Fr2f6bc+LJ7F5a8T0w5BH5sUEiEQ8/VeyDy9DaCW6rw99cunnWw2a+K2D9Z+kuco34IrwBquTihw
eZBDLzgaP2DK0WRTt5nT2G13zYDaxA31KcQZewFmPJ1DAH7q+jJsYAW6rDLYlLM1YpA54wYvfhIh
5cmoQNqm/KjRuUo1ReVPjBeJJ3sGFjE3i9zA16UjCxAtdnoXomLQXqBeqzQXGyhw2MYa8yqu/QMr
bzBF3ENeJ+crqlPUgcv+kdFzooHpUuTZcHtWwe9kFPDC+DNqStNXc0WGTfRl1m3E/tY+jkWT7bUw
aDJ3oLWBi+LunNC1kwRbCBCFrcf524EbeBApaFh0jXoa/3b1QfU+DvnGlRCEcKHGnsz325gl/UBk
Om+VU90o/vyMJSUd71ERFwOGaTf/C9VF86R7VKegKOIKMRpwkb9hDI/8nPCZ+2bJavVbBt196WEX
IS933dRtYuUdUAnPY9IVlzhDANsQF05PxctnBSCJ0hkGSLQAehYVUG3+bWhmB5SK8z9T3TaHwjbX
TDVlzHeJjr01YE7toJ9Ex5KpXSkqVC5BGThwaXrG4ZZellUIFssOGNecV/YMEiXTe5WEET7f1T0C
NRZaNY7hEpQmEFmhvO6+qQwlbZ5txZD+uMph48vZeJu+/6xY7ypM55WEBM9J7HCR6gBh43StxhkY
1UnthWcSjphXpoBtUJ4JVkWN05pQsUR56oy+///z/5XkSLETd64dq3Xgx3QDGc0lhO8VZ1UtKDHo
jX8GWA9X+XdowdFlR5InO1HLkjQ92wR25XMBX+8MLt7WDx0OFUq9lZ+8UjlCCJh29vY3dvZs0cAs
XP/qsdogVauanj8HknrYoyJ1EqhOc10DAJzV0jXcPTlfTRAOwOIoAkHf17NHRUPaKoSUVJf6nt1Y
VHbY7KOPFCPnRNUNXftdAqxkew/Yff6jSmMy/y9i8pt0VN8pkcn9SpA74cKXgyGeUy4FuE5LWT+b
RtOxQC9SoTzGfVpjwEn4z+E7QfH0VqBym4JUcPp/aIg9LGCdln40xvM8B3JaKUfXs+5dCu6hBIGJ
feyPjqDeispgfyldHeZXBV5zp6/qoBHnyGiw7AHEDS65ueQRSqdqOUfekVQiQFDMxWkUJpwPNKHW
mt7AtY/XCFiy1ejBkzFm5sSkYR4rjjmJrWTG9O1pjCqsjyhsUWsq7+ZFaT7swwpAU+f9MIVI/Whx
HKb4C0IxM4PNQBs/uo4Gwx1gZ8jetdTYwPcXpt1a/e0RaZB4ADkKGJHPHy5CXC1Mt1gcaElQhDUq
zrWRSRVggt5DXSJ4ab++ku4EJdFlsOOco/dFxeIF9k41tYRoeWCI5bXwnxqXDYxF1/VLT3quxeBQ
dZbDdq7LuaL/vxUDG8iDX/KIw3Z6Z6YDYkIfCjDQTFFiZP7NDFPMS0HiGRYXKjmdDIAhMcCX83SH
QSh9cSpGKbG8gs/GXiDiQZBqVE1k1DSNDAluDDxvn2Bh52aC6KGs4CcqzMda3/TIzB+zeRM0v3bN
6+i8EWlKNWZ22bLJiDfkB/8eIU6C6oDYCIf/eCMwu3VM8xGrV8SQkbCa9/B98ISQvHm60hLDhAkj
ZMkzh2uqz44sMvElZQDkOfTELbcq8ifw6mcVDRaOtH7/nvROCNpGBsOfLnyz2hm8TFM0FQGNgNTd
PDqvKkieWSMqrU+3hwHtP7AHKirAe3kurkk6EuJHkH+exjYfOfP9SBOvj10wbiBW/zDb6bpIYq4e
mN3rxWvoXgZ8khc+mrbjdIUZcYS9wYv932hp4HxIlA6z6gqQNExu3OIjx6KkHFJPyc3SbvsCFdFR
joJx+VbgHQx/FP3Y9Xi2EV/tX4e6qWlsvg6wD1SWVhm1CKlI0+nJtVagjzZHBp0Nf84DAOJzoMT8
7PoTbo43zurRMDu+wqqD/9YDbgiE2jRKc5v0xMnbGrldvfDUN+VREj2gGwF8iJZKWej5pguHDID8
d1YPcCULfurW79y8ZrXqFO/Ibh9C09caJmXiJHASEc95d/AgLPev3X00GpVBdpkvg7L3cXqdmyKX
qrDgqJWwwomgULfbcukybXKXyMOZ8d6dOs1UrrgSR5vrPEjkh3jqIlf8jWuj9z/7QslSa0GKZNV+
HxEwPz5JkJxBGW7ikulVj9t3DJ7qLLKfM9Fmo5CGI9pzZgF0Jgn7dCbAsTksiUB6JKSKekjZ/UfL
gB0PSli7Ie8x3k+j0VZ7PxT2yd45O+uuTBVprD+JLeU9HbjdsOUFa9B4ujtOLpqK9JpXe9Py9hVQ
vrQScxgWNTN21nj0iz6ROkjDcfj/XM4i/r7f4bRkAJaAJ+ApqY1d0XG6JS7+GFrWszBg1x44F52W
UDimQR3XIRB4TRdphUSsW8Dj4Mzli7U9kH0PhjYr3sumyPWkws9fSrMifHhqh2aecwBk5FgA2SED
2VWG8bKFnpbKj0bDIz0hCataFoBTQ9pSjtfMMBva6VF4SpngnrfwVtFqBqiNDfi+G+1q+0LEtMny
k3kcYhXCOEAVeRxtk45n5xjgpD1Cc2F/V/Iief1GQ1jOeIreRnMs5lsW0cxUC0ohXKTbpkuL7O6K
CPvnFDj68lcVTySRAC6xsxsX/oJnzNYuGi5SHWvtxriy03wFI6jBE1OIAqjODU0+SYHbD5Wt8ID/
xCmSBZc7xjv2iIWb+qR5TqTzfod3igyDJTMvnBaxYodt4msiuzxaMk26NHAkH1te2EpKsfEwBcVC
oMpSCmBfo04yuARMhtSUhQlkrG5lT/JDIFLUIhJYX+baMIQacB0/ixzHCw9s+qfmwD/8IC3GshDM
TSeMmTR9ip7yXjDefe9w0RhMUuWtLNq+bAHD1HiKYuBiZmG3t1CK6qWeRgNR2oX6YEsRUDq+RnqZ
MP4flj+0JA6ohv6/Q8Pbcpk1EUw/vF52CXFCKDPSnfe+/CL/D312SJoQy+WduEZwgm2WyYKVmP/U
epCgVs6Od8FEOUEXXs2OCLsRklHoi4dP4sdidXpwO3jdzlRmQS8hH0SopokP0Mc3wxjHxwgKQrqp
pEnPB27BfouKzaLSaDbNPpMIzcET01Eg5U7gUB6Rdho3a6fNg4F7bf0UvnWVB32DuyYp/eUf2QYs
Vjv6oXAOqrFfAw9UzaTl555TRCBC9CS9EWZWefxf2LM4gvo35/lwXW5Z1rhTlO7dOAwHTErWsWWh
tgu2kQTtwecVYNfp4WK37sP+SUL3pKQBYjrQ7FqzdteqtWgxkgs4uvI9vVmYK+tIUj1I/vdwHbvn
kPxtJAlcC2pSUb0rwSVNVH7usw1ArEZu/JiZ5I01yFCYeHZc+dYTVWPXjPBywij5M7UCY4Cz4Ifw
FRgpxaRzvp/JTJsv6iPpvvg+JG9fRjNzb/Oi8VPB8FEdatDBNhii4mdCSkP7iYc9vG7BzixCCbRL
ghTscxrhNoGnRc9gbndZd3Qw2koHH4ZrB5OY304agOqEYKevjfhDnjBLMbEYSOF35AaaruGivrjF
aJnOaEpEXyHWbuP807+lhGmw2zKW1PT2meyX0Bv9JfK6IFM48YOS8JivahgeBjPEVDv9lKzURfH+
53eE9wDAcujvPwdkFMgXaDfjWtkuibRbDn3uKW9uOUNcf2hID7Uq6hZ3bqYeQCg9EVEkFTWOZLnp
Xpy5NSD6/sNjAfqnhK1fU1hIt1Zn9kpkWqz5aY302A1FoF1qh6yJgDkfByNEhJD+eFX+C7MD2cwP
wyr9spLV2jVeNIeyAKYdufmy7LsQ58h94aUJCy1k5KEC0ZRwBQhSDtlk65fEcHnZGPt6MhmB0ko2
mgtsjKmc6czEAmZA0JMbKkg21thhpMz82gH8brtI7ibZpDL15aY9Kcatt3zz0SWQre7ShSb8gOe7
4hEnLd83IkcBXBjX7BGs+28wvKC9l3aJDtDDJeai3ADwYclCBf/aeA9CuIrE2CJN7ljYBDG93sWR
fnO0hOkLexTPPhPQF2My7yq0vWw6oIK6/Mg1/aw/S/ejsqNmKUETsCqaFteXxgLQE3p2Z3PUbFiy
EudAqBXai8eH2sXaKk4oRWmOB544808woVKu7lM1wu2+aSsE4L1j5O0hoInPlklQp5Reg9AczUd+
HGYqduiGYCMxmZdJ1NF/i5xm3tuMCohV6HbEihqr4leavK6ohFL4cJL0k7CKsFDgEZ4w5GXpAcV2
Q8impjDf/HA8jtVCViLIUR48xXcISFX5gVZgS6Mai7mqtGpYMo4G4cn1Tj+9Eq6qE02EqZ6TSCxQ
pdjKpsLX3Qq+5NeCZsASp+rV4bN6qfmK5PnIolJ2C9e0FFi9hgdn+gMqVa/Xmw9VKrc5ttu1pnNt
IMOV0bVpLiQceAucYGmYaswxYXTnCeI3LMxWtxWeX22R/4W/4jLCF5sHEYbSHxSu3Y7drsdCR08S
OYwZ7oyJyTSUkYQuM7h16UpCWQoEGZrqr52i7FBefTHQV15WpMF6ccjSSjQaXUqK8rVpVo5WAoCD
arBcoBkBT6iYUnQhd7VaqeBtceZ1wwFQX2kWrk5NayWz4MBGGNBLCcVDRdNHYSDyEZ1yG0joPxvf
ttMHjJ9Sp6zjC4l90U9AFjMe9ZyA05VxL239X+HEcTyY9DGiGzecrM+srw1bPNPhjw7M8RwiqIqr
tzOaAE/zUrH2+42vmlWTfBj9DbphDnkqtsa5u587Tks1Z+NMQIF4ODC0qWoxF75yG7hTDsN9JB+9
WGDgOgCnIOfffDEo7Ca/sV8JMeo8NXDlsnIYWXDNeisIqV8P+57hu+yiYTKR1CHIzXmHorVpNzNl
fpI3HA7FYl/a6KtjqlWz/R9jGjq+9js8aFfX9AfYCeP6ZVMgYDyCqyu2Vwo7D/w12KRZYoC4wpN9
Uam/pL+Y3j/TM0Qo3933FCyfmNNdnLg795uESKPCa/W0+5isNzQ7Nu+z15OVAju8Lqi5p3nu70Go
stPyrR69tMxA/TSnnWXNDqudlWqoNi/4JOjKkFYhbTNNDYdKTVcemq2dWD/KZBk0mvlBqNFhrmUF
TNg3HrRxUbmXRufQiVGcfSS4Xg8gRXfatI3UomlMzsmy/TJ7ObQzSlY8J7MigbKgYMolT/gIZvvM
6e1GzlYR6i6r+OKXTsu67U51zyJAzBAQQvpTDK9EPXnXSsJ7XNcWXJ+9Vo99ifND5Zz6V4Henpa9
cAIyAqrkAJSStH8hEUK0wdHlGvqzBPoFD2S+GKvmBpfv4RROXe9e7kecn3zeiOh6vMlXaxqVliVV
nJt3eEA7PokZS+VnRgEjOqJ7JtkhXKzDlaCnFdLMF2ms2VXBjAhjSK54j1c3EZpr9HVG/VP5lyfV
9Hkm2Ce9X7i0oAY8BzMT6ZeIquptRr+jeQkm82pB2Efgh7w7rxlmm5PNqOb2+M9N0cODL9GC6ofr
QKhusXASkX6yD9uT9U3719UeGm4AWSKTNKDMfokc/IEtrpPfV02mLwky/Mxv8SAg1KgUsAqe8XqT
DlmUpYlHmDqIbdvvG1wwaztAsvK9jfE6UhoP5rkke0KnlRt/fT6G1jSnEwW22DdlErEv7A3Hchk8
jOkfybfPzOjCw09mkkAZAyPfzaDb2XAdG22CuoEd+fV+3T2asX2aCKvQn99GMi/EMPr386zr8aOI
ooMwwzNAG001PZOLMf8oqpet6PdjqCTE5qbtKaT91P9H0VmWEDHEzcaiiMFSxJAwaNT8AwlsMCb6
2SY6WGev2qs3B3SjtosuyHTVpspJwi/DGzmoyBrfc4nTo38wwIXoUO7tERTVVc1Atxn+5xtSI0dm
5k8oZazHBRa2GE+lobHrtCccFgJnWdTJOA6446XwnKm200MfNUyVzql5lh5cSngQHa5BLxPUfIms
R/TKg3IEjREzZA7g/U9JWpCz43+YA3L8YKwzW8ULrFHznWkCnM9b4wZ3R8F3Jckwgl0Hu9/E7qBH
gp7yGgyOv5clPM9lHGw2DznXtwaRlUw1pa9TGQhB7b6BQ3sNwRN1KRwgCoHgJ3Q8mqA8OZIERJ86
Pq1bqmeOZ73q4hLoYAIA17eyywXmWzo4tTa7fownVnp6k8sIEkXWhBe3QS4aMi2iC4GfKPvD811d
MAdJP0ojrKaQVUu/V8/jksyfpU4aFn76PENrthsl6MWCJbP25unDBhjwzLVW/vBEhvgWPO+Vqykc
TOJROdWraaTxksTNyUpYogFiAzWn5BhaeLV/bRxI1NCovepaw6eM5iRoKcuszXYIo5ORv+59h+B4
JWmzp0R+ImQsvuDV2Y+ANFyMjAMoiUe6GCjIjX4YOCiTYCPbUs7Tvakdkac0I1bROo3aPnjs8tsd
NXwwkY9OkWKl81DLrz6lcGOv5HXDvKwED+5Rn1tQED0oHt1DdFV3jL9vNc7Ce1bvItRUmTi3JIW1
lZM7OyuUJF+Ju+THNgxEzzfEcBboVgsSVLcDQpeuuLfLkV77ltrdcWwyo1jK9298e0ymhbY2AD92
vbPXqkvEtj2ydyEPnWLGrupJuqwY4NkQHU07FrRyu4ULQ69Gmg/pPXube0OukyCDUpeSlgit/j24
FBqo7evfe/XJ4RKoQm0RO5xoyfdhzsFFdr19lqhbtJSVvx89kS/NVkO2wEelmTM7TMiK91K990wx
Khf6myIpRwW8oxNIhgP+D6lUkATSgQGl9WaBKuwfXQ9Ld0Ivw1NAMcEEUJE4SDCTFUeKZqm25yiZ
OXA6bLm2BxGtuK3b/CiRCR1GQbWhpEEk5fw9WHPpM2egLk77ZnrXA6LzaDOnc4wJ4X3Q2JD1wdvG
ThuUVyulkOZdtW7eVB5VLh9Vk3xXCCVuNEn3YLsSLAVZXMmfgahaj4vFpr5OALaGlpoHQMi+a0Ns
K5yl1uFk3+rHoME14Ppf9lcQSZ5Gxv8zRna1iLosmjTRVHIWHDBkawX2i8qkCFl95g2ThdNj8zVj
IsFh+4Rxj4yu+4KgY9b9cifcl3k01nXi3BZL7EB3K74b2WBf9sGcTBfDB1J326rkvTPqYW6yQx4v
MQK9avmrlRhxK7HDvDvzwE9Zzdj41pi7+4LLzLinKIdWb2guAk0XezliKzAUKmSRvM60rGdlr2wT
btkuHNczmridp3xO5VnQdRT2lqNhGHT4F7yqZcmIAxqnn2oh2L9IP7Ua1VKDKeA7lnOUiznez+R5
hZz6JkAMapW7F1dF/w6vipONhJmphOR0aPEUAORg21oLv8vA9ffe9GqfWIuSKFt/BOJNSAp8FKEI
le9gS6MCNC3Z46I3K7roltAR3x8NAeN2fCVd80b+ZDYsp4A9xW+zS+NPkpiUB0w3OGMXbErBDX2S
GtpaJaOkpB+AMyhFPOKjqx0lNrSilWE1uA1BvFSiqRwXmCz5HmZohA6jgUzE5oiO+Buut0GqKHf8
EcXQoxh2xl3iul6WkrDX9kU84tUfelVi6End6wWrh2ZaKS9LosECMsqnk6wF6yBvezyk5hSETSvT
Z8WdmZjkRB452bEsocfEz1xG1jmy9zYB9QZatW2th9CxNoGcFAYLO/nCjHV3CKyjXLE1KKpXHtR5
nBt98vwmCMhpNvfcbZMwR+5+2xBk9+PQxj5VBOPS+pOOaEiQnsEEmiyYwBwPnPfUnI9/SnhL0A/8
xN6emBdrkIUIyyf83EPOf08ho6ZzuHHtz+EC7NuyN9aipjebgGGsyPVqCGQ0h1ODJZPD6uhsyNYE
RQHSFi1PMMlODEKFyoMwPKUeAwUX4Zhv1L3nDJskpqNyuI4+JkInfxIsEgSBdB/jg6EAN6Ic/5ME
knQVbnlEhjHQeclt0F+7jWmiqHGZ4R98isuS2CVqBWcgcJEG+VjvFVEnauJXU91s149GOqzAvmbw
w7g0re3DBRCsjBp3wVDY8vhX8+mbU/6hRXOm+ZeQ20l36hXWrUEy+hZ9HND1JHb0WuA3xUcaZgB/
RNTy18AzQ3WOnWoyjJ+6zP/Q2rvy+snUS3h2BSIydXS26qhFUMQlGRdy6OFSY/swDTCSxVKcC+vT
VzeInasAg5HAABSIvhjRBwT+Ra15jtxA9YprIWbEQ76RqFOLZZYKgJsynGLjKb+MTcuJkAyKoxw3
mzyMPJvuXfMjGPfxiNQVUuXrQcnwrGTZXe9c6q2ctkibxM2z4xeX3H48nUeutV8zz1KxEpY8mRqP
hr9dDtG2V5AkumYcIZ6Zsa2aeopKdhFXGzeAhBaVxpCeLHQfb+MaNP/M1X+UmpwyfGRMHT2Eqvtz
CBrtKSR6dgSZoddh74rmBdXbAIdLWfQJf5LCxvSBT5zxH7gAs4BpxgRCfWe7IHPlrOyzWaQ6we7y
e5Xypn9+DiDht4joMD/bpBwO2RPP0TlUE9WddGjNut1pvRAp5GYPPdum4yucyFfhGrIM2evfYxth
LkQrQ1CHC5xAUCmm6CzeQ8tENgHp/InHhv8GkYABBQc+EvRWdQh7pLYt9tRVy8TjSnCl/uI2EqTV
8r6Vn3AcFQpwjV9k21ivrBraDhLZ8nQww86YL/wK1jQL1k/eRtuEyC1wRfnWdvUkyoLvlkTUM2Rq
MQNoW6BimXgT2vKsDJcJTd+lMouByvbkXul2Nt9HpmxUvC5TyxU9v0UBb70PX9FhiCvGVLiM7BdH
JlM+YFPSqS8J0k+KqDSkR9TeGNHyeOtpX40U5gMf4uoY55GhuLMKFCPP6lbb1RRgk6uhHWk7gu78
ELDbUoMc3FC4zqWsZqGgfo+w3wMm90qDwpjyAATWRg/HBtPM2olAwKl41BbSQKUMbapLTqp0z50E
CS4hm7f/nK9l1LI2la2SQ/UCs4YcjmuQKcKDtd+2tSW2czRHMaBR+75Td2MVrlRWQnv9yBF1FFBu
mzKj2KdmPzPks/AVr5v1e7gQjEYETYfcvZZNy04Jh++6kH92re+NeyyPepG/3BnoZmW6sUATyHpO
gn5cWPqgQXwDqDoyOhry8Spy+k6ZnP4qpRoGyEYDHvc4mgZyfw8KZN2xVwsySjVErFTwb0Bf1Kvq
czpMRNkWn23xcyDJ2bNz/2jXr6R1WXOr/Qzxl+VRc1n95WWagxjkAAKLQRu93xUkl8ybbP67hB4W
UfjyT85l4dVoCNBivR6KtlPqwgJorBOHtfwJIoJWExmznP1+AKgZbaKvN4ihiWon9p2UA5Rz0ClX
xFqxTPeAfrfZKbYm4++2nYW+d66A5PbfRhj+nVe8u+SnvIZX+hKtsiQ7GS/Io7B2E8tE+gG/fxUR
AK1R7OjdLSskaXGtcEta3D4ZyVeshkezU8Fl+lBoXIOd8+Dk/j33X0ajhJKwVE4YCDW6hppcLL1a
ta8RrW8fyuNVsa6gSN0EfVFwu5NiT0/CwtcR55jnEGRiclheDu3s4WIoG35HTQX6tk5xmy61wS6c
fE+DXR1Es9jCejmULoCCybkLkFbbifuQHJmMeiniztbaniu2DrRHDZoOTZE4uQTIWkCK/0AGEiVN
mzl/vhuJhKwieCSopWbuUR5mk40LiluwS6N46aBpa6LkdwrzAQyC8rJNNqI8rl7bRFFs3NZSZDVP
IXPznSMVJqSmsWYSrzeR+Sguh8gjb/caO2RZv4pBZ06dxjZqgDvzZQqwjSfqPHRWg0K8DE0oqT/M
wROl/h0crbQ+C3XUeps+NBjFAVb3/Pye01lE1nTfFKQN9k7jS8IcMjcP1zDWP5QqB5xjkaKqeyYQ
fWwOctMY3NH8y634M4v6tNi6d6c/gYU0IFvngImtJ9D3pGzeNWbvr2+XWQ+u95D/0gLuHUDB1uHC
XWzgdLOeR131LPPyopfBwPjdzdTw/aIRQPC/8GCZPLy126e8pGolxXP6J9w0PLa0kqo7VtwyuX6b
8CqGH6e9EVfHiLBQ5mEqaDJMCL25lLeoDgZeP4Fl4grVstiEYiyaly92s2DZvuTFmHeDpcTdA+m4
0EUMZsC8kj63O1PuW6jo4JYgardhVHwvVTKh87H8FFD+AHzMTuTcNeJw9tnsNMhvc0M+hSOi1wqK
H628ipgzfT1/JoZjI8lDJ1W5pT5lvYYMeJygvN0A4cct084uZEsVJi/OTHvsUDamSOLGe84nivOH
cHQMhkoOYZqKMRCqtzLWbPX3zB5FZWV3fh934h/yc0n0mtVaObAkFzYbwjvtS9ApiRlRSgLC+cBG
PgZFCCA1wZtLor8glsE/qM3WcyW1uj192grV6PK6Dk3LPWLlBkMqzpJuD2hkD2E0gDHbWxgQiH7M
x9LUCD81eP1QRYSysIpcwOJgW0ppHWilCDNVszLhJYCLoVY7Vb+R16xCYgg0NaaZ6sZo6fM7sj1o
2BrMh+0kiTAjYHVFZX2Y0rKn6V2IB1W8bpX/tlRisJJSp25BYIsBpjA7TG47f2t8rYrXqj8rpqNP
z1rSBtluPohztnmtpJ4hOmEfQbXeIPLPFxzWmTVZDMZDTDKP9fnPYLSA7p94FSLJHz3ksgDwLUKw
ICI+BpAXVRnwL+U22V2LXeczaQejHm0e7WPVPHNPvVA/sHbFGjuLtj+JcUeWHl0H/xasceKE6jbX
sYYA5ymHqimt8kHA0DM+B6A8nE52WBB1NKuxrOMuaOJkdi8Cqrbne0GaId9Dw5NtNf15HqjkOkum
u9jBfCbohk9vt8BSEqDnYfy55SfzpSRvJi15qBkUdiyOFKC9o6jnwLSkgxIS4AYJ6wec0SJ+5M9O
Fhm5pb51YdLH4CacJlJ1Uhrt/9vtCExPdcxFQpFsEbyUq+IT99x0wjFAJG+/4qCAZYx+9ZF5pAxG
7S5agEZT++FZJTbD6s4L3k5NR7n/lSXfuqo1qi73mzfNiAIHDmarKbT8ThfuuI4EupcwyKPDV9Hu
S4k+d1vdgB+c+xEW1lhQrTCAVaoL6CuZ53/UnmJgkesRXseTxYH9WjG1ayNOOIPHLSkTh5Kpp5RD
IVM4dnhU83+oNWfuLROeW9gZuTp0gUBI7Cf4+iW+AhX6JEo+DFQj8wJz/CkjlKKOvBe6sSTAUCzi
gUBz6cTsffaJcLzrUObRv2DQQAi2ikEJbjnavtRBVmfDtXCDSt98amg6fh38+JPeEsw1e2l6MSWr
oigiNdqQB9D3EtJgocfmH+g2EZRKHTo1UPxzmpKtpwm0s6aEo1I0Zhla1uWABY+HRW60yaUDuo0+
hlg/8tfZnDd5F2bnII6pBFWgbUu7hBQdPFS2bCNM7SlC4LgvuIkLcg/oCVfyr/guaLYSicWES9KF
l5FpH97ZmJO/ZNTrBmZ4McLKwiY23y68Z5WvzOJKsfTzkY52I06Me4w0PkbbfmEd4MjCITQmNwnR
2ZV8jzhMtYByzwweoAIxU/GBVlSiJHZxHUJO0ZQPYwucmtRivhz2sMybhGPLO66fVZzL7kjZkPjE
Nw9Dy5Pz31ifIK4Kr4YAomMFhnVfE1ne1FkG5DuT60RL8vhhngF1Tt3e6HKUrqP/Ev00VKQFmo3v
Fxkquo2ugadAOAdtZUXZSV4M3/fBQxQHqohMx4ZGxjXID6dSkVPNHXle6bxp1CpI/dP7kQuwDtVX
t0RPan310sBSAhUscndrs/PBy9WtMla5MSBTxwQdQwdvOo3i9J3ctObbPZqzqXTnGTmTfFDCdjYn
Igh5TPIXs9pkjGw2FxFF7XrCweduEUqtXYZZ2FT637oqdc0p88jrVvw0enUEq515Sg57NzR67XBr
kaeMAoMo24SWuoGAT4H3igp+rXLIM4Nygc+CQOyOa2avd8zVlOiWgYtLEMnBoMKns5zvNb65l94u
3KRVM+ngN/PFIAE0Wsb1tf4tYTX4L0V/TyvkeQgygs2zFx8skZwE+eiCx/AK3z9RlGV92L0gQtcd
yFBqnUDQ/H92Z7WtR+UTG0TGmAZWw/N8YNXtyVvgYXQGiURpMy6gL3SKlAO6ib/xe1202zdmTwQw
dNBL5mhMwHp0le8hvYgvZHaQrC3AuPvR6OcmvoSmPDwTxch5pHqveE+dbybyM4Jn9jtMJqBCcPBJ
3CFppUIbdo07k4ECJykR9itY3vVGIzKaiZuQUDWLTHNScvDmHfbzVRLjX6BlAr73QY+TAGIvJ3PS
Rvxu0j7iX3QGP4b0LVFiKKEqfPuyQ4syW9SDW6N5FVLw2ow0FlgYypc09qL+Ho7Nbcq9i/qGpDvE
mVXqwtZZcfLiUcX1IyLLhAi5wWPg0/OlHQshVo9HN1w/KUK3BzVqkJqNl/a0n5w1BbsMhb3nPsd0
8GYa31eg19Kb40xEvRo1AgYa79GQ6unbhiQQ0yaB5+85vVe0rqtBkO/HmugdaryMXEHbZ7wMCUyb
1sh3lTYi5DZ9ODISrP+FHFTH+BZLpaamiu3s4prpaw6q69Fe9agxFhJ3iYK3OdMhdlmmIOUhZ0Nj
etccb51sS/jp+/DBvZ2PtELUhRTHHiO53J0hY9lzGHG4kVxEu5sQ/ZIDnlZl0oU3pZfOvssJW+SF
YyXVGsGmjjWKBVsNCNYGF3nwsGtNOOd386UKqmMMxGBWw8oOLl/1nNvReSLKDCSU3S8n7nS47/hf
TGpP9KIxoS8cLK/lRRv6PKGhl2mgTZAGpky0sJZweu3ZQVWtPvREisaKlfuX0bGuvNa8bxIMpsAj
1m1sMq3GzOrbhyiYODgd96BrbnrUJsqQI0ljeMmLDtxQeu0kYZ8KKZF3f/9M/mCRobVxWixOsa26
MCsIz7T5iMOuU1FsC0Q+earZN66ZcK6YgB0lBnKjqXuEAZjgwbXjCOMN2b49lUW+yNRke5FQEhrr
Rc4jMWKybHIjEEczM7ROK5L6gVfGpBs8Y9cM3KHIHXsSEh+b+yu9fokSJvtqW7NUk2qzw7C2uqoV
3npXdQfRvCw/GZJ7sbEu4H5J79BLQ1gR0GeQonbm8TcLgp0216KUBPKY0xCydiW2fblFjdXmlyNx
uC5/EZKBBwzn1mG+VJlJu3tJgZ3Befb8g3+B9cUIkCggFSQHy49CRQsPlA0vV7GjcumoLt/VV2Zn
iyvrEILrgEDj47C3JALQoy2Likx2dH21nS0NpOGy37FlvouELorLGm4vkGdYZrJYyzq8Vxh+nTk3
L/OoykIPxslapuHpiHggs4DUPLfFA+cR3aWNKsn1LtZcengiFlc4FkKuycpsU2rkfKKd6xGmV3yw
TXaMmU8nMJf4pa10rdeNw7jfgshSWkmZOuXW6YEvMjsYm6Eelrgl/H0TDNxJto/FP4SrcILgP/Iz
Eh6H3FYVOT0LIz6gRhJSelNs5Uxg5xNJ7FyA6rpiIxe3r6MLNjbMr9bLoqhIGBKn+JlCV9gIrMQ6
hPZUvXEfK2GUWflsn9tfZ19IqDmg13vQkko6OpItc+Hqoq8x/r/6H3Q+20g5hPs4j7dXJHU0QRp6
Cka3uKb3v/S9l86OChLAfQ2c8mPY+9Hh1D456rZF2Bqo8GKV2QIPi+J4QQbpqdDTv0aJzgnBj4xG
oFLzOVVLVOY7mnYTuHF4ONZM/8XbE9BXqJVFV4fqL+ibVG32xlylXbb8hX3SaCgtqvrylC+mienf
LPz/oPm7e7IZVNy9v8i320mFv4Xru0m9YCb4eQjPuZ8Bi2ab+HJLfP2Nx8ra4l+K1w2xsSG3/Qb6
OPOX3fhULzSnyCIm0VQGDDFHsAG9lUUlAL0NgpPASUacysXHEej0n5MEPPvB+g+CGQoFFFR3cybJ
JTtAqLtmuCC8ZBqyt8FXAodG7QgxlZDMWuVR9I5A0W8CYG7IIAWSBFReNk+WxqWKg5RJRZytipe3
3Cj6qZEh5b9M6oTU2yR2lYKNumNz4xu6SALCkqAWFMTOSqpN8fCZFMN5c8b6/r8u/s4An8zVOVB3
RogFmtMP6N6O233gJtG3mr8AHKd2HvrAmVENpsKlSIYEErjhEi57VnDxCqtUfyffGNyIoXc9M+Fw
izEjrzeKI2dFxkk9JJP/23yvwpRLXZjmchSIfww/3I1KhdX71xkJZM1InSa8JUeqwFrsGlua0Hsr
5zVg9Vl73JzNv3U5novfgFxVNo44APfW+LS7syjFn82kpI+msnRCY2CNaERpZ65MsApz02J+KSou
9H35ClPBuYb8DU1TvGNk83xwP5RdKMpCJuLu6COuIAy2y5eZA3MZ78m+lpg1DSb0JbQiWKkNzjpC
0RKSrBL1YB/1iNOTyg54Xvq360j27JQbyreEQmcndHPHgPos4WNX+eJm8hMyHMsAlB81a0qh7cti
trKqcspuRT+bR9ZQOZ+scIn77P1/Rvn7eJQSeJ/nNM+ktN94ERZIWAatj5NO+lKyQOV06do56Du2
O5z8AK7zwBH/YyzogxUCxe4AdILFIWyEwxEfP/EpXaqcaLbM8sIMNrDK+kbO09VRFtiLLsXoVDTR
WOIK6FYB3nd4cDp9odA5LI+lg2TvifK1BYDga4ttTIVSHUqIwgUQuFfZorOLUS2Zz31utiuz1T50
mzb05dlXZyGM7ifipxEBhNwbde43bjDQ0l3JkjxVGleZADbuxYO7CrazjPh7BUQKjJcdp7/P4oHT
Y0V5+qSL22TfMw4MBtsYiNTe2Dq2psVP86koNQfRs/STtD/CxaHOhXfxoCV0YRdvD3utcn7XYpLY
gorlzCxNoCIjPB7WlqoOUOoDYADSRxxP84qBrrH1VDCa/Fn68LoAaxTpGMP7qk+coZmhBT/ubnpC
Yh6w/2EXcWTP1Os/xLN8Xm6iC7kI0Jwxq72OxxcrxN+1HypR6GuTv9EeeBgjknb1cS+Laep9NW1A
tD4Pfoocd47jJPTod7lht4RBDWtasVtB56Ca8XrYNvU0Z1Rrzc8mW7FdTBHaH19jAvLc2bLiS+BW
AuNA8TJrzdlrJ5xWaisj42qGjiWv15m96kcYrpTgjm2RW80WMfCSjGeso4Zdb0PVuwpWy548pjc9
9dZLqj1OaHrT0bjjeJxlyoJmSamNwM2g+XgIlksVZ2t0b+pckPoM6xTq0I/zjRBExYdkUYKepmkg
uKvzkWynqETKIy+zVTmSJ0C7qeaM6Hvkg5wBPza+MyGfm+xNXRQAIsvI/49uKZCNre5jnZ0JWVHC
s+cYApmtUbrWLeLYUXdZvCkkfJVQ9R/o7wNEfAXloq8HQxR5rRJ26fhe5sPVvhIVy05feq2zPY0/
J+nG1H36qVPtg6Jsu7Ivo25Rzt0Vmi1GudDfcXxuyxIgOVdbtEzzvynQHdBusDedWTBvxd6yrKg6
Zb5gBox5pojHRMmcBM55gW2adHEfQFhYq3m3e5k/I2kTUS3VI+oXq1xYAjatbJAzgM2JYBjyAa+t
gx/fnXv9Jmwl6d/8yCPpp/LifX5xI19fFiKl9lzz3KBdif2YCOjkquDLsKD2wqNTHnjemEVCKYK5
pN+w7dzgMUn3256bFWADToeMbd3avnbs0SvIZP1irGz6C7wmPolj6Toj5CerGjShGQWmP5dnQkDu
Nk5OnlkHrgH3yLeQYU5E2a7fE7/umtF6wSbXF5wXzcKx1iDT6sPpHJ1pFikBxoaE+t5fpQcRxWG2
ZV/qGqfTghdTf+w4HzR6DKivbqn7j+hFcGVUTxzathaEdzlNAgK104nh/qutZVlDix7JdyjMOkBW
FCj5t+R4YpNtcFKGIaaV/KYVGJPzAFKl80MLgP7bXjqIMbGvOydqNawTBVEfHL48I+GxAlgQgAEy
NtuiEMDtCAr9kFcGd7GDr7cH65MRjCyDLpeVjIHtoeCkQbRiICDpXdrkhdqR4NF96l/Iumx2ALIS
pqAgltRbW+psD8JSiNoXgV9ZLc5C5FEBx+Fbb+3WEUWDT14xZ/lswvxMoPDi48aHrgMW5JK/1OLZ
/vgcYdDY88tRhDPOv9ClTFN/X1dzvc3ItzmxVz07yMX6ReWdSWTY/ufZk64dDQ4vExF48gJFR77j
q1JwOFgmkTD4aoWDrtdsVkpRtomQXQpxe+7DTimR3Zo4BLr70MTMSIm59Sd5VZXz2nyBsQ3U2wto
nyN2td5TkCxqSrbzUn5tRncJGB09D3Ms6WN+NlVNR9zFIJf392iJaAMDLPvDDVnwrM+1w0zLyV/e
ISz1r3k3wFaeI7iofQOKeUfjsvB+nyLuFtYY8jE0CKOMzANkMdhgjQV8Et812dilL59g1JA7lmpZ
7jEq368/jpeOZszZyUf0xB1EswjlGp7i4pJlmkWt06LcDvNlD3UAj8XDKBU+oi2PBQ7WG3ErkjEm
jM6LE5//W+DRA6vSbqU+6Lm0IFT9bGp0RZ8MrI72+EnG5mkwBIn/BacbbtOARLqe1b9aB0hpHO8y
7nVc0nUb7N8fHLLDQwcO6iODOx+/jLZDGMh/IQvGjtBJ4dXbH23vbFDCi6I4Fo2oXxGB1ihGSzd+
ojSKuliuiYem0B+jcARhuE0eQ712wiUsnPyknmh6UmSI40Ac4E+O7AZ9auZliVPeypVSup0B+Abf
yJJjJ7Sxi9Kyl7F4Ix+Ah1KrLwuYewJQgNCbhkoQEtL9ic0WW9roUrr6DMSfJG95H6tkJFLVhZQp
k7YactGvoGnmPOPEYKd8d179gPqItza+NQt7DAZw5nT8JlO/mm5sR2TVG9Jb7yp2w1+eX5gopH5j
qE30p1NFy3059FxXoqvtvnv6yIxCmNrI9BK0QQMrkWFNyhVNRqFcoJ08Mey+4ekVNtSbKfqLXK3F
PTSQEb7C9RS6nduZbJ2jDOl+CSrmMStNKCpjwWU/heHYdagCHBSN207ycQ4bQRKbB/ur15fbU0ao
AqoprF1DSdRaL4dYReJFIwjwUSiWksWh7ogc6T/UGoUG7bt3X83oGGlp/L5X+WWxe72ujPFDrWOQ
5EzPaSVrgkdQbmKVrU5zTbN+idKp6HvaYTlmLQhkq59Fbb11+qpqItVSrqd+bl0dzjfvBalybevJ
WDtEhmWbBWWVH8qeUC4PZbeYluv+OQc6E4LTySU7ERwlTyzXlxFzT5LZfrfqVeTwMs6g+zC/4ltU
z0YkiMHut1CRWANSmlXcICyQQ9ZWJREO0x4VU9quzeMr8ycBYD7jTHb4Xs4+n1+8einXyn08qSld
huSdI4n0RNFT+35QawqsACiTCtISSHd1dy/RhV//oKQMhEjiFjuGFACYLox9XYMUZQVSepNdGmnQ
FqoCIXIwadvzd9sCD7up2s68boq44asPturqjpn4nE7xyZmy81c/Z6jvdULZLkG+6GLIO69q5yyL
07EzY7YP9iQKvw7LGcr6nCdI8dPAQahoIFNHF9t4zaLo4fbRmQvOBs8k3m+IcotogC1MFUkijcuJ
6VNNxWHBkC/JBseWN+NHIBTaPwYkE7koDl50jjTSSnsep8RsgFGMorgXI3BG1pzJ6s5+0prfJybI
kDViifK073L6a0EMsNsVcyobQMA68RkAmHyyv4raWB+M4IRgwOPLvILcRLWyPRNNLlWf6vFCCPBJ
mxkJZ1uCKXj7AtVrJhG+COrTlYTUNCQRkIKdS/ylv2HJZyHCvxNhsFwv0V/5T40BaWtYsb6UIqcL
4XLLstm2DnIoqmj7ltXSf6R7T+w+6n92lM8MU9nA60oZvRa90+NuU3GdiHZxtAjMOEHHNN0IHGmr
gNZ/E4hJ6BOi/4nl2DkHQSBV2YnBP+750lLPY42+drQznBDghxkMyT984tzHqgmYcCdnkg0WSRBO
Bt9jDRHPUV9OGR72+rBv7eeZHjdYW8cBV2qkLRpuJksVyDiTmhyfeSDp5Bp//IuLQefVljUQ5QrY
BMsMo2crgjT3iHkJD/1PxxYgkaWZ3Y8zR2k4HY/FvluV5uGIW4xjuQHGe+FJ7M901sRtwzxmq/zo
Plo2U+GxVETdQ/GACXOUPp+6Jl77S6IZwBNmzognCFhqbEMkMD8mfZycLk/tKiVRhq+nJl+k3RDY
IRLTsvhF/SPHqWSnBBnTaVks8JKGjcLAkU+jggv78TF6MpV8GiJmCpy9nw+UeG5neufRtF2U5cNH
ES8W3bBG6IDwIw8xjrUsNyRuabUuMoJ1fsrKh4zf0eKNKfJOsjgDC99rYBmpGdfEFVUGatrz495C
Rkh0Rl9Umd/9I5FC2fE5TbvqM3xuaEyEJROVAlzx3tYp8LnhmJQWPproahXJ3zRPs3VcsksZCitt
pkEY81+8ib/WYaVvjKWfK+zd/piQfi+rVWtGPvZluOqgLriTNX6caAlt+785TMXXGx0bUgeDMm1s
zYsPJVTsTOUJzWlEOlst+M+rKUGZnmVxFWUtPPcieJkfN3GGbIdnOMMnsYTg9kgFHlCtISkFYV/G
w8qC7G3cyrOkca2sGB2rxqoISEjkHsd6jLrHG0gnkAMuJ2jyD16iPpV5OqwSk13aFquklL4yU67w
T+b0w3Ec8P6iuHYVJ5araJOUGzqjLjK+CrwbXBrxxD6WGJHpI8Sr18+BywxJk5akhNOpkHlG48zu
4xtcUk/oo2Nmyb4SXctR8YmFZ88KNSIQ0zC3asviJTdlHuRMIlo60G91nnGsYM+97tf4/dB6SIa2
LFSPN7gWPCysQw6GuX8jMi1dsdkOqtOjHJu28Y+L3XijXKDedDQQPuTNNleBXLRnzUbJxe6hPmul
Prcqvbj69Kbt9sXm+D1mpinr9WrbIEhHtX8+XHyT1rLfXsFupSafvXhaWQI2p4RJoT/WnXYMGfLR
abeQwZfIRHm8T31cXYd/oJjUx7JGlnd7ccchuwOAXehba/FHxNuWOOlrVn6NUBcCipwBe1blEDtF
kQ+/W3go0ydTyhwGX7rmXrwhEQqMh8oTrtnBIFSqaZejt7didG6MdfAySqlRnm4fDVrpThcYUVQ7
Tf3HvVts3l/bRuADlUGopGxALd/NTH2e3998EhlLY5ykDes3HKHWG4VtCu7BtQ4k0VUltXluGmkX
p3nlHV+aAsdrRSWiVOfladpeRJdkV3FNeshJGQAbd3y2+DmCAU8Q1nJABtkL8ld1NOwgjCa1yc8I
7zUr5lAklXu5n9VVsUpYSjfI6EWxtqxLxxWTRDSa3UWS7qYbaZx8nO+/K16OiRrSIu0pHwf728rO
rvKtSQgbbq3KV+//RgnvWIrHfFGPtELK4V7Obo5M25ynconM/fjnbI02TTC1kg13RUYTEosdQ8Ok
z3TU1F2tVRKGUsbEY9pHkbukUHA7q/TQbHjasYsG9Hu63AOUz8FdLjr7FXbetZ1kWWeoxLMeILE1
Qnk9bMNAwakfx5yhPiu9dkduLF1TVyUDipH1fdf3fJ0eYTqm+CM4tum9Ex3Gk4JgMEQ8Gyn3Cl1a
2PR/M89J0umgQPjQtNNKQLK8tlKVYLLb4RZbU3c02utI9IHTBYwVvQVnuUJr6dqGdKVNznLL6svu
fsFz9IfUrwk2SA6+S3kXacMtctL5l5PLeHIwCOoxBJuqnJki7CkvFSFOYWsfXTEIlVFyt0lz44Z1
CvxsuL4hWH8ZIqSZTSOxknwnIpaQH3IKo707ZlZPhGHNmpf6bPJVVjV51ZmbtQ75PoNHtFeOFMqa
1TU3fx0A3++8KDm34n1jRrTPImR/Tvb1/GyB6cu9w1zWtPz0B4NrNW8ZM+F+jtw4wDOaDjuhc79p
Fv9c5ZVolqRYfXVAz4lXi0iO3r+taxff0gEEQyQYJF1bNF40FIf8NZCOrXg31VBoPm4LCswgXs4I
SMFP6+5eGbYqI9OW9RayOhG6BePXXTtnO9jduAMd+fDZv+B3RYy2XBUddUJKyhjtGRZi7/4YOXsU
H28walirT1KCWjP5CUaNMGJ7ZtawwbBzxF7VoHSY3jH1VkgnQ3iX63AJubsPuGF36zY+FKYK/6/h
xbFGm7ew59tVTdN7tV9SOtLNHtDuo4XsovPPawvKu4mgS4L+YLIT9pUN35Rd+W2hiTAgtfPsn8ab
KMgox1mp4EAjAJXmEBatmuy89V4wQ9OU3ZfxsXtXAT8rGb+RX9I7t17CGsDYx5oTjs2l0sZB2Jbb
TnW+TfYfBihcHVbBToCF1MnQARkwi/60XCUNDZJn8/JbzFXjzY2S1rfKU5TfF45+4GGijKa5fNp1
36b6QHGxTURvzc/Waq8OyPezPG+dQrz0XMDkOBRSjzkadU8VjiMzZGqe2zafr2Vuf2ITws5CseY8
FA2RFsUFvdKNj8JHMKaAn+hBCNorHVk9w6qXIbtZWm7ldGp6KJA5WJChXT0dyOAx/AaSf0fis0EI
xzmVUa6JWb1ejgpr4rulEMVIokbKPX1E0OO5MSLsZbZLqH/H2nZSrdqlTi09Fqmk04iTjDbaXz8U
cOpqln88TgH+VzN+euKedPXYDUAe5xQIqw9ZrE7CVhvA2q8PqzL1goGfiyP/T3Xth75mSZ0NXbBl
ynKwvqkMMAT9BuyhCnBxcbMxBtK+sZOipGLuY8kf0JZIoLyK+ryddkgtIyj//6/SEcIKAo8cuiTv
sksY63lSDc0XvHK8tb7HJNVOPeKW4/kLySyU48sXUn+iO0Vh2jv5zA60fqwZL/IIvRLa7y6mbjGg
ZlzYo/eTiJ6AkgtSwTB/cEl33nbCQtm6DJ76iJhHAQNdfOnpKs+RzFXCYsqzzVXcSvU089G6nzeb
C46jX2o8GV3+RA9VTrjN+hggEMYVcwigxkKvJ7MmQFohERJIBQP2utYUPM1epWpAEudmR+Aps1Mv
OIWUCuR5mnMU1WtJaOiTRl8d6CbUY2Nl+w327dUgi+VU4zCK1HfvpE+F/cU1UpmiLoSkZs/dZzFI
v0HBuisBE65G/nHas1zLDAYCwnnrunj53gX4p0CHWDoAuavw2i1fNTWF3azUHTPbhXIORZFPlVPQ
1O7Da12t+1tGcB1kk40QJVse6d/xPQWk7w5ODQGOMC8mBJMK+WfMl3DXOmlPhlw5QApGoGrv2PEL
kAN8to09flAvaW0lZpsXpezl33L+K9pqQf1nRA3uTu7COJHD+o4AEuiMPXSLScjdZVXS6QZwHFTO
xuNagolW8m3N0CsEPAI0vYLNPQ4z0h2mMA+ZMSTUqJkmOAzy4qUkWneNAEG6uMHK9ur/1VAZ9bLg
lwcwmdr+TmJSkX7hYDdrETonr+Ldk/3/ba24afC8pfiVqJW+HCdku9opbrGrZbVKG1O6nTCB0EGy
CPx0tfsYzaqlJ1MSpNNYUiqpK2l2tPyO3it7KD5fc8nRM893IFuihz3BeZ5mr/MlZbnIeeer7qME
FllQnJC1jy+O77vgYvJz2TnsuhhDSbByvcuRC19RNopVnFWIu0tfF9cdRM0cq8j4iS/4i84R49kD
20UMLIXP22nYxUivJrftcNwmrNhC3Pp8WGTkBhHA9DBAc6R6Hqz1jBuwPUP5yHmnP4ITTO6mz4IN
LDIrTQSoeXKZKvA8uaFFcP3L1ZuOnwa8/64RU5eq2EQLDP4VnC+Mg/20BMPi9X3f7cApoJs2jOiw
U4JynMYbHiA/kuEbuarT8kHnVH4HA1mrT89UyZUZWz2wR30Xx6Ix3HVvse0pAYm1jVUZDlGvcNDQ
5JPdolP96hwvDQilPb9jebbw2s5gENF7qn5jAVMFstO3Z2qtmzWa1OCZXsm42tWllbvE3XSpGhur
iE+nxXH5mwQTvBwyl3P1QQI8mTG91Wc/NMAvTGB6fjYK2gRo8VRSsM8TKRtwXpZay9RFM6aOqCAU
7lnAPm65MOyWf6w6kkkdTr2oMrAxDHbrpW5pBFL2iiZXCANmUDozOKUAZYn9PdCvEM43/984ATMJ
HsucHK4enh0RiuTXsoXkPqI7QnsX9TXro2zRJhQKu7uxs/IBu5+pFQFbHtKfyKtZky64slALK1YP
SwSmmOok4COJtNu5PhBkbD8tiskOr781nH2YZ57z1hLV0BqPGqwKGVqQdK/Fcshuq7HsX809DBOM
SMY5vLUehHryb24oWCEUwVcisi6TTPA6Tb4ag7ZAr21LyPiACzb9b4ZN1epedJTPu30E/42sZgdD
4bVaH61hXvin8ul2BOLY/CVLqDh1qY35d8TxWUoJ/CDT+uOxAHeuOEV1qn74Y1AqeXEgPlMFVPUT
7QFrEs9f15YAiTslBCh+pgj5TA5Wvc6aR6P88qHumd5HvOWs3LN+EGocaDrlb78D1MBJg2EEtm1y
mNfkmds7NHiMS/av3atGv3nikoHHCWAGRkLWGOPmVPzpQeWqw15kQTXLXYSsiBYjKBa9XjtJqdPQ
Q3nLX7N/+GwL7lcURN6Mlwz6OB12MRJSeqFAlaRR/OFXOxhCAn1+YOiEhS6SecWANwFSlt0coRJu
hTINbWy1Cc100+2c2PcNSXvCkU0bCMYp33K2fINosTkylOSEPelrz5jNXVDUlxVWP3mTAO4hvH+s
sELQwDzf8U3xAqQ9vzldxO06OcRvVnyN16EfBmq37cnA7Pz0FVP1l0ZVQpcGEF5EeV5GbzS/M1Aw
vTNncrv7xeoeMr00w3OOWyzpOe0iB66i9MPkK8AdHqjV65mmNJ2jSd/Z6VKbzpAfNWRJL/a/mml7
H8/C98CTXqqfq8YNPvux4A18TJPK16OxW88OP7vorISibZ3izMHkjWRs7bpWG3vnAUehQ9+5sLpz
H1Xl1ZoOV/PR1Z98gPHr9GmKHKmK+FqB7AMoBN2pDEe32pPjlDYFAFBM+1oVcbZ1nMU/3kA7egf2
Nm2GGV+rvBT9wMJL0OVvHOhKv4YyeVrctZ+6Lf1m/E64IQz1iaRZ9dJ3K9Zs/ILRQOjk8MNu3x8a
d8LMvPse7kdOkLdGu4yRlUengl1EkeI4I8nfPScRoxuWG38d8KoxIT+Pz9Fo+LBLDwt4+5QgxI1s
5HWlIEmL8tIwTcbKwdzqQlmTqXtMuN73Zr21SLV8yE4m38KlVIZdYOW4boIeXyszlaElBt13PAcx
h5G4oUO50WZrGyrt9qDugVW7+WhAK8KJGQACeOR/Yzg39pEhd18NviD9NLrvsSA0ZA11IlHusuS0
eY+Vp1jpaw/FFb7qfVuG6s8X8SMvhqyecL08Bih5yCbCjRJFfA7t94WzwEhBA4wJleZgovHsrXsN
6j5ufJ5M7VMQCLh1+3l7kZ21BufbhpqzCu64S1foBU/GCL3VeD1/W+lmH1PdBRTUbHkZ/eQZzcPo
Z+cbNQ2MzO6gXf3NCOl41jFisbIvLh5smizXOAL4mwy1IFLkiKwYcaSctx6EhsOJ61OSnn4bXy74
0z7S9XWeo8jA85F3DvdbItGQt2JcSDSYwa2pPelWyFI/tu74MV1avn/kbq2XVFHjxaDaN7sTSCWw
wUBlT8Z3pIWTp31PwmLWzskNLk5ojSumIPhCK7cdiz8pBALgWlGOt2gYuCw9m650cZwT7LVPruHZ
jTXR/LJyhPMQNeJLhaqpDd/RGrCEYe9bORYCAmXjzwwuwmVhApxgbtmUXbjtMl/Y6MWmJTm4jq9e
vn8RYZRDrKZwB7tJJhXUaqnZhmUwosM4wBMKyQb3mC86KnU8r6r/51KBcjFfFb/yoN3Ddlf/10CS
ZLP0GJ66mEsLtF1PrmumX37HkEm3rL87uhKZCKXJ9b3zX78w3NlDfh1Cx3JUkKu/gKx86hEGV/6b
8lI5c0ZLmn9vOBg0hciElWDkKb2sfe/bBz4DQ3xHy+48grZJMB66XkXiOOp5LtTY/1lSyugu1RUb
GVE/J/Ic/dqK42KmWVnCQ5NA1UxuqfDbnnpyfCNUzlG4dAUgRgtF0NFkAjnsmBKGDji8uOOwLZ92
vX9jGraDHhT/H9+xaBaG3m60CAAroPDA0Q+hIprQS6yv806tHR3VzgCqOftx3O5VeNX5rOcWQO4Z
LDroyDNwuMwyFHYfkMUG5ddXItssWcZzwKyF0I6xvy38ZWsRbNIcErTRtnt/5cY4YIL/1Kf5+LBo
PIDXZ/Sw2YqptKCEUFxI5nQ8G9dyn6S2cQMyPGXYw4Xbtg7kXchniIANore+azBP3gW4QrXk2ACK
alr4oMMOEx+U7rNWjuGcD2QbbKZlKCOoVHNpnsw+v1KVB+6t+HkIKsZhheVzZu0eTpeBWVbBFC3m
Gia8LaXjLSMrBBcv/dJV6y1JpncPCtEawIMvndgbRiIYbjpafMp+M2nG9oNW1xLTJ3p7l1HlE76R
+cMp0ZbCrk5PyuMcla7xHFgmY6mxLqEqVYK82YcL7DUtYjmZFwKCLevMn4fpMwad3TRs+97mixyz
uBCqXYbu6i03ouUTgUdLzZmdI6RcU/bsi08pfpglUjDGr3X6zwmvdm48zEA35/lgFUfFl0rwA4qm
JhuaZGzynHjbQnBXsGCP0R+08bJ5OuTWzGz0fUrptApVO8bE979E4BQqtPJ02cf8NLzAsXdbDgsz
dTGLNitjI2hnZpXyZBfgIQndT2A326464zxTNJHW6DyJ7o06YOfsbx7Ni7QPpcSLRcMk0wjhH98+
oawYeqS2G8eD+pStqNJDRfXvVJBYvsDyeo6C03cZ4bYPFFnviNo0SNQRpmnBixiq9va/SGc0MVvK
lf5bN4RZ/29IF0l43qGq5hDmDNSjoUZ4sQv3BcM3CbJbo3xMsSj5LmLSLBpu0fqnKhwRAmGcmlTp
8EJzGPI/6WamYPZvPs2YSpmJrIqlWjufn2uchYUQHbo6GmQpCF7FdB1vd6tU616XMsmrMJK+aLSA
Rv6CHdVVkqG9gDVh1luutDHxmZo67P6SY6dn8erdFe51IV69WBMEiLwhGMSZcwXZDiqFpqFWy9bi
NM/0fqzbLi7a6AzJ0L6geAdlqsUCHkUEM12TuYuLyyfKldiRGDVtEM9p3whzTYDIhlzIZJTrlIM4
JRVtqql7YhoKWkNqDz5t0gvSearifQqVr3QSqo6MW7YpsSLL/YfwY/er3/IB10izZCIryjDwnGXp
b5K4gn8cnBLhrT78TGqyqblSvy9fOnw8y6zUeiYFGwU4EWZ+ELeIB7qDPNDI6qcr/Yh+fphHi4j5
8X9wdPnpjBMmRk06nRLZQ5tAIQ1YmE9H5Pkekj1pM//zUK/u6whzk1al2XOfeXXU949Z0mu6qjJy
uay9C/43x6gBsNlY1tnQL/DV43Js353WhdZ/vdjd3XYka88OWrtwbQYFdGQqGEyi7b8g6D7JoS28
KLtkj5WwrDSA/ghtUcSnWKcMXOP4ZUe9/knY8RP7ceUE5vVnArStnYMBqdl4c1hc2Chis4El8Xwm
1DeKPV4zKs0hsTt/t0xDkgJEtasDN/zaYQE91+wqGjHBp3AKXGlxK1QzDQi+q+v05iNn2DYbeWuD
QVimX01tyoVL9jPQcWB5h9xdYkwW3pMMIsbxGr0J25CLpnzUmUxPiXMesAeoqBR3mgC4Tnf6AYnr
8RzZGVqi9ju+TkL+8nAXCHLL4JeZ2E+gQyIVXbzbOxBW9Zx/p/HtSfTYKJ4AJAT371ENxUAtgOUz
OUSLmokdzEajDqjfWkf4ShquqHbrLX3p2lGrxtyo/rUUDaQDt4Amm526fkpWb7y/qFqwHyFHkT30
DWN8vETnniAFP4OFSejGHMRitfHYusiJWPB+uKT+tGWfiw4REZJyGG8SbRbjUd5B3sDdMsxZO7Aq
Dx2umEWAoBVrSMTL5TlEX7OzyOnk8yb3jLTdC1CeAO5UR6u02iuDyN/ZM8pFJeTwesjl8u1oAvGk
JfWSRvTfEVZJWoWnkcNf9+L3dw7DhGLa3EnkQ3SO8gS64fNvxmiwG85Q6f4nsJPAfmlsoDTCgk93
AEdHYr6ZCFbk9ecmTF+PDu3I+V7uCKoqijdxMKW3fnwFIb190W+aoDqnH8XFfk5St7AhIvi6NEKh
Gc+sFHzJBv3213/KxWcGaTY+8yv7X9ZW2Myq3IUtEFR1HDW3BHoMT4q6dTkJOXAuu0haVjYnDsDR
wA5kx/Eq9dabpCzj6l1QtRpMpTjpIe3KnO1GUHxjzxCvS2Ntmqv0/kdWqIUCbKb7ZmAJohYamwgI
Nhm0etLgA42x9B+7NuuwHUDEUbPEhuVRj1lPUIdiy12tdN2Jx3eopndmrlFmHoYj/rcAODvNwuUM
1fjNDOd8byuBTM77wik1s3GUYDBVqsrN93r8uxtrTgHhUUHj+s7rfCmy/5jBv4sJbJGLdL/+Nump
lIz7gi13XNSqui7Ced9brfdwEp4C1EMzOllu2reldrSzQJ24scMhxzRXUSfHlZ0qS6xUR9+mqQHr
mQR3NND48wjoWDxw9bbJq/SfPvHKaPUZBaI6T/OiXopFemYOoB62PcP2c0TjNz75Gbvt7W/JUoQv
OfrmRLbqlQIT2xDzpoU2kIRgM+fjuLTWHoEyvvHY0+ZY3HzA/bwQExW66tu53QO66pUhGUtZL135
TIbJoH0SQC+3J3SxOAKsIEQ2Q+caYg7Bn0L9zJfMWuOMWbtC5eCggbmsfTBRfiiuF7Eg2M6zUgWf
U4LYcJvwaipd3gnQ6iCmrpst6Beqwilz7gOSjEz5KdwUGOTmsz65MpQizIo8nfpOLt8LqIHBge70
IX0kFKF29h2+d7oJ3yKpsqvOWuigVX24z+V6rkL9J9ebv6LgerSIcbHRnLBx2VmRdeJsRoCXi6L8
iGeTWwiid5aXh8vu2DskUZeTF+8vuMDs49XoT9kXTabzY3YRGgig6YHmO76ZEZCmpk6oyNSlhzuf
gV/E2PVg6aqeH8IedKAhJF+Ykv6e4hZSzfFzgGYHaTkaQ3x/S2exfGs7DdI1IFRB5x5UFFJwkrr7
mwmycilmuG4TBWH5QZnu1GLvSlFPVddJDFLLbnzU1eKW+f7inaSHKECIW+9mtGWo6+5s4iBzIfqD
DLS2E5pwfM8U6MhXFcGRLp/sQF9KH2jZR+gr6qWNvDX0J1wRDpK1yr1+Y6pKfCGdgf61vQOKjixT
HioCAlz0X67q/s0pAtSVOZKLYwV58hMsSOjLY67DZwkceGcfaDffLNi4jsoAs8rfZv3APLpUhtzS
dZYjSxrDim80mcLCUEgm6mbWT2bNSc8opTxUbtg8mWiORwHMRSPhlCp0zW8IpyvcAm4u/PLq+Yly
x1UHc9/c92UQh9X/IO/zHQH8IaBfLE3fdxLCvC1CCzatQJFQa/fPT5VIThs9LlvO0F9SuRQ7MVQJ
E/yOUowZC3N8Vuh1ET4o7Jly03Uh0Tn4z4StzIdhik9V9zikaLtgPGyjvgNAJ1XL/uSBm/9tdU4i
S7idtd5sKaHw4RJyuGOaKQyaIkfhcg/4gj/3Z8/1qO+ur6hSNml3kseYQbcgPN/tQ8wUQgb0beFj
6hAOX2myJRzoy/pdDZgCFaCuRXeV2oMGio3pR3JHM0JZn2wQDrnYl2wtYdprtJ5uYT3NJok340Xy
+T3EkO+GiDaxH4v4/X0SDhXwFHetzDRKBkyqn5wIwuwhE7paJUpWG2MH0VlYVIcHsS0eZY3HFrfM
w/ciimglmR26I8ZvcIZmo8X95UsobTJtCwZRrFEH5Rflh4/5OjOP9pwlPVwcrWXhcdEFC85gVxHB
ZddHtjRQRXnet+GPjWuEBDIRuXeQZl2arAxeQFACkDia4Q5pQiEMuZVE45P9cLEy8LOtWABEaRP8
SorhwvzrYJJdRlATgXBpOQ3leuAwJumpd7F4mNWni14HeiQFrkAyerlsqtDo8W4pGAMTdmZ28A0K
rhSPfg9X6WHvhhOWvDLFfgdTAWOEwvIRU6ednC4jNiMs9zcWyVlW08d4eWssJuchW3Dv7UlDvxGk
DSWSSr3CzAZG4lkKoYpEm+LwrDLdGYJm1kcupk0OC3RsH7nzIrsBIOSA7pUb5j1XiD1gdgMd52ZP
3pNN3vE/w+p/llkvx8EDIov4Ncp/qcpyIYVpx12Lvu2U2eaysSjZvqIIrDw8V7c2MhGraM4imLnn
pBJMTbfDMkuAUNvhYQ431bCunl25lFFTRfkR8lhxKqexQ6NZMyJOwsEHn6yz7ENdEoAn41TECS0U
hi2Q/imjFqc1mTR4dMCGpZEonYEm2ILRZ+ifSrVJyZ8LTt6OW4cWNq1qN8KMT81vmkb1nCVl8fyO
S6brshTVlufG4rjPGy5y8q7V4fGE7Nwe5PFSmA5aQhtJt8cCEtc187XpUiYrJKIIRPfb3H02yX0f
P5mDU7OF83Ryh9wzCiJtG1dSgk7v/MhBj0hP48AqjMnmCAmOjtS5+kzh3FMOO1JI+BsPkhjDzSFw
TSvgK8JsZQcHiuDje1UlFdGrKs5c+BdF+a2iW6ihRyIfCovB4qZPYLI+FmnH3cPxWA66+ui8RgZ8
Pt0RrrOz9Wbb0Mb5pb9RkoKL0r/+icPH4MToLD30SmZvszaYxhIPrG98t9EOz0NXQGa9Nd2fmK2y
VOSapZN6bYSODWESApDl9rg4OiGer/+gO8oDIqGrwbrEvUFtlh87EFSzZ0AdAWrWR18pNrzFUGKn
I9iQvXOAho6XrI3NLj+0d2rtJnbwPIy9I4L/gf0bk7hTq7zqDl2If0g+O1xAyk0WKN+Ihc4KwRpg
o4rj620V+iRn/LlqTjAC/4Miz9lGz1G23VO/z+nhh9++5HvjxtD1VVUYNnnVtUjFYXpkD+r83//3
o3AW8E3lyLsAOSQbI4BwWjuK32boJs8ZPN/IORvmPgiQNuFQ30e+G13K9iHaiPH0xIVINH3Fp4mU
wwJoD+oFgOME8j5BpHpDp2Yzn8Td32g/yp12fA/Lj5JajGeJZMWbKXiEpxPqnoI6lt3emYJx8bF2
mDA031yn73bXSjA2tam8mu+XjWfYWpDA0GKABKxCzfI7phMoCc2BF6FR5EFuAK3tzAmd+RkG37QU
j0PSWtNF0lKUj0SbIRf8lGX1knzDQPc40db4Vf0ehk7bveFTha5PjkO97Hm4CnF89x8F6grrevDj
CTubyKNdV/D6pmPXjLZbS34OfxyglC0418BLAHemH0pJEHXGI282r7SrfoBNLH5fT4gZGsFjWLjL
bQOe7Vz3ox1g1P3PnD/Y7NgDErZr0x09KaLofeb2awxAeWd3oEyzM+XvAt83np4bScBZjPFd9VBt
OoczCg2l5HTydFAZtmQcp6fGcMoHCD3ru3bkuQm/0ylN5zuDah7SwRZ9MxiZ54X+S0Uqhq/M2hkn
kB7uAiKDRPvPEddpt8jRikO4NdMqxTesbRZpKUAgzmRS3SYWQ93HyqzceGorSZcZWSbkubbaRBT6
iPsIGPRRhtZ3bSQkpEveQVqKQy7SUDmvEiyFiUVfP4TqF+1ue36w23aMyHOnK71m5C4tVk6oolcJ
HMhtD6RaqJL6M0BP9PmcnTiutRiCYItkOp0sdy449RbJxSDpFygf8leChXL4JL1JNnCWm/VXROK/
ulc9ICrY2biTrXiJRqzPpG91BafMF6LL8ZdAHEZRavjnmNPdYiiCP9/UGvLr83Mkuj1sqTvSiMYu
rMWZQ44ADrIuQYavkTJP9PWg0zjFzLUpLkA/qzTBORRd/jmFbfF1fENEGFnCDzvfajocyYdD05Bq
hSxsjVorF6t2fB+EK686aHYRFFjIK+sU2EuL/uHQWx0bpNJt2wZjYrixtj37P6LPVqPpfIPyrBvH
+4jEKozKaq/zo3fl7wZyo6xfczW3bLBGW0xykavQTlTwoG4Q9g/hksSWxntMUtkbYEZ20AASmIt9
6n+lCgKfktg68jER2vtaDEefs1f9oN9Q9bQ/WtLT6Z5IhQ10c5uAf5l+TAhAEdmd8ffEQzy72+Oy
LBtgrxq/HFpLzQ0AiVBeJZ9TrdZvepnHEbt2FgwVJmlodgXz9e38mQo50EdvbIKFVCQwqXm0jM8Y
iWVw3e962QmpaimSVP7H/LTMDIDeutZVgfBgE0lzgvXJE7GvS/kyjgHpsMPqa6wGiVuS4adquWyJ
72WE+3l/IR1YPo1wVxJqCvn2gyYdOiwrj3fyKhLpUAykxaTPGcMG4SiHo6yTAJ3gHikJYA7/hUd0
3AQk878ApNu2HfxiQZHc1jzYh8ZTVwiJexcgxM3vz0H8EcJqjxnECV7igzIApJbtq15nbsWYfz2/
JAmkHtoqrdzF8AcT0hUXXGjUbQc07ZvDIbZkf0z/BNCEDXB/2pXOw1zc1POrEzXOifM2Bk1PyziK
39/rnV9x4uR89oHcqDBNpUJzAF5gcch5I3ZdPNUMW/aCdglnys4FCd8c50q1kCwJM+DaOsaxYUmR
p3gsW7A7EiMWfmo2Gaqg9eOQDCgg75j+nQ+solADtOBrLMCL+i57SvQbyfSxbxw2Me1i2WjEvTw6
TK3ng5+yZMM7m3vM7sOqwgY/l83rj7pbG+QM6dQly7TjdHCZBYWgRYQNgD2YcSrE3M04EvtdkQe0
iEw/5NX9Iwy4cbmwvId2ROPbLBjIUt6a1/Nsr4ukWrw4x6f49dtnEx1rIxLsg+VwF8uW54mBv+sM
QevXwP8iuwXRPNc+vJtkt4HDAWs8BIf4jefujC7hQ1HR2WHTbFuGG+kJETa3B8NAQ4nG4klNdctP
Xv78jitdUZhzj2Wl0KKOidWccwBLmb5qPNdYmVyl8KLKOJQP70DJQruMklweDjxVLuzHPeFOaYQQ
h6lQjeHzCD5cxX9yUAOpBCzgOmI+udHuIqiVA1s+bThafTmoDymXazsiPtGVwpMoN6Fwk1+d9dwb
6hfEr/g6cKwwqvH2Vpj+88GCxks4XuXo0FaxAml+BfOtJBiLQvQ4C1hbsUsNAMBlBwwEl4dQU2TS
etk0BQ0YmLYflabq7RgqIuAGQ5gsfwMxZzW+jUO1dqNYmybqOWBCTjvATcpv0MkaALGH1f35VZCO
YGfnJhJPs1Z2DGv8u/kHyUFPYGktkZW5xR9fKDWJnJOnjJY/5rYrcj7cjRCQke4BH58MIqEkytZk
ZhrjB3WEWqdwIWcgKfpaZLr21bys9kmquw3YZOV61ukKYeWdcGRIuVtXNUt2Qn9khwIi6M2va4aA
6aSFfsIg2LZZr/eBJ0OqCMC2YBWWP/z2QpoIHBnxcgSMq/Gxkd4wCu1p+rKxW9H3K8f9+YAE5oS+
VLGdhTB8Bxo0rEP/sgIuX5cF3umXAJFQz02kzuZljr5Qc0EI2mHDoBTfRiym9qImqH+55E02kFVU
PxG9KkzAvDuJnGx2l4QbNAoKbg/JnfIY8QubYEIzGMGw7FyEAOLRLWd4AKkDQN/EvXy8VHiNiTkV
NfCy8IEjTYbsNrWJqNHfS6p/JR9zFP53inRmyHZotRksatwiyzwy2/9+8h/OfJru+3Hxn5gg1Oa1
dYaJWxe51ox/jDYXBHsGpUCkAB1usS+cWfXEmd9P43X6sbasLskd4LOB4fHlPl9wmcBIBn9ZsMCR
mWPZ4wnU67WhJtif0UTNFdcXpKEJGeOEx3OTJtrIhx49H+2YjVFFka/P5t8VtiWmLKwHomN1hPTQ
doahFll5Xg4uD6RlmpEE8l4SXmY+fhRLOltCRpPkkFpNiQLfmFd8H4xh8p+1z5x1iux3T1bfe7Be
sxypc5WSuzcJehcD0g1hrq1adgJlDmhD+5QOHvu/Ga5Own7WRjZ+2Sh516A3/a8C3ku2LmUdkT9X
LYPMy8xE4MrCBkeUDYouQVtcurDnLdq++HRsyXU4WmoVNPN+NQjn7HpaECEeSfRlBs/bOJSi7taU
hWZzTK8PgKgIDG27oXU/oM1YPO7uCXnC3jRbPE6Qo6UJmK2EPV9P8I9Lg0x9mlZkTgbFdTQE3FNp
o4x9+voU7YP3OiIj6WXJHrAUzktvQ2MQH30OGoZPxy/HA24on3OBqYe0ngAPVDoy4pe3sg/wHPFN
MrfmRLxlJlOMh6MkSYsXHLx607+kchd6M8/hxcLll2bTml4AnmFX7itUAJPu91PrA80fJNY2R1pi
zDPW4XFZLqp567UvujtJx/66tGUqf/LWvQPvQOTGObKsOf+qKtxhsXYBy4qGvOENpMtUw7lZ0pNA
trG0lBta7h4zF5lNzjykSuln4p3/mLOLRY9ax/dDm4EmfTSEkS90cZIfyHzzetcju+teK1NCJ3Au
xV/gkoCzh+RnuTNKBjoBnRElR8A6pqmIDJzOmwCNmWVNjb853KzB6mL4amwwmjW4UkuSddxfE7qN
siyw3wlGVzx++9AF7mCxevoJOiLe/NmrAVjqx/hLHNfm7VXfwafaA2oUZld7mljil4ojg7WrRf6S
1mOqPc6ThohPQwx10L+p02dta+ThG+CQezCtj1n+vE7ATtPK5KuBunia0CeDQlBuFvky1aGg9Iqq
Ix2MOqi0jDz18QOtY49ZKA+FX43zAX3mkKN3MGiIfflAGgRvj2CPRmni0mpJjlqJAI3vy+neSb1f
9BTy/ZLUECQXTPCnmASm036JI85EP33HbSfTm/WuQ2EEO58AT/+ugFblKGNjyTf0vUD+X/F/cXOH
fIFCbjU1jr9V8f2KgYXVo2zXr8mRa7mvly3g7k+A0vLBeBnEZSn/0aQiIn6A8BtFMazpr2nGCTy7
N5VuH/6eEsAQwHzoN69GbO7Vfr/64mxIfzr4jCNvmIM2lJUVDxfn0nIga9ITEFbDvB+sYsdhdPKO
S0MehEvJ7ogA9+T/IedSJmbWq9rEpmdonLgyygFkQVvRDJoF74REHkt4hAxaLVAX+pT7+uHR/MAn
CALBrNHb+K/q1SFU6krwQgu6mqC/wqDBw5W/2nw7a3pbZziThA5hVxvT+3C6371OIWSrci42P1Md
DrEFPyfF50EEUq+7mBnuzD658hPp1oboAtkNrqb06HWcgwRkLqGcO4jebbp0earzujzIWeRxmzbs
izs6AYMAmiN3e6CRpnFNqrPV/cTzVjq0vKHeGgvlrFrlxJxPLbj48IIerwMO75b503q6FTpwAx6c
vJtoKqagQLiAMpVYO/lY9KoHbeKR0YaV3KYxQmmRDBZSv2nVo/yaoJhU0p8I7XG5h7hZ54dwDofB
aiICmn1+dpQJR4mRSK41wOcZVeptNr9j/TphLi+cPaKqeLMRG018LB0MPWHYCFrUe6oYs36vOrdD
7y65q/Td7LWp3JZvUasXoKKcKG5sFcvk5A0X65pX2p814iuovlr7rDZ8WCbYUi5IVXQhyERkVZFq
jrTyBpZjcIZlToy3nWDEj4r30V2OOX49b1K6mjIGl8lpQUMCQrmZVwmBUcAWZ6l8b+6oXH7TSJtJ
XcmEAlvAlEdNWF7Zd5/Y3rhXUscpCCMCiDWJYK9dZz/5fpDZ0fGLSPGVaFdosYo8bVt0R2Lo3UVq
LI1oqkMKV1NNqn/6LG8mJsRxL7vOuygvQJ7hiCjfwudSMvXUprz0kjWUZsgE+S1H0GVT2OPtIu0e
0epOA1jZe/EDcTHRk79AjWFPiI7xTolXrTw1pm5Ux5bk2RwDqy5XdvOyBSxHoZECPgZBXerkfcPy
PXHCrxDAQMB/ZTPLhHfTkPlyLjH7a0H3MVvV0MKsho5IaPr6gPsPCuOwIbI6qLLxqdSKdZ8iHmiv
56W2c1ILpHVWoS04U0ZrjDs8UeyKhEb+YvjDlpBDUnAfVS31/QY436IgbXccT1ZLV0bCe0/X0eSu
YBmPYn5TOlBBdMx8a+AkGj3e1+V+qEi0dLCZyKO7kxi2vs5h1+bjBlRFn4jCovRAdrUktTzz8E5J
OOFHBShNdi56caOAzYUfCtbc3xbw35DpBtgCh4VGk2tY5cT5Arjj2/hU/aMZuLTVPa3airkQ5y1r
mqwnEhKkmI/15JS9wMdr5yS0dujOg6EmzLSWqeKXxE/SovSY4dUkt1TQg1mkXQE4CCtPUBlokGvf
eYEfOCYersSFTO+GcZ5luS24+mGkIli2tg/qN9yD0w/yv/cwJHKGi6v8sRuvslqjfetlp8D28zeV
Rta08DcgezeZ+39N9STnmd+bzFmv0YjvtaQWUbe8jEbWExsrercbytqhSCif3BM28s0hJPs5MVHz
RTZGjM1LPI0IYZ5l5mYej2KvTi7Dur6k305e4iQoXwHAjK5paJvqIMT2paUsZ72pICNGXxJ+FhVD
TIII1qcG62RRTG8Vo/IBj6uPJ5sQsSo2vx+A2vgDiOZniqBjxNFjaFjTJBS1ru0BRtttChkUe7U8
R82TCYxM5csF04K8pUL+7yyIjBTvDh4jU9BfCNJO3OkOUngyCPr8L852g7R0pQd5njjao6P5qkXA
kX/pgue2xA5DioU9zXybTK8G4Ip2DDOAhvZZyvYek/a8mysyaazOUEBY3OIMLCFl9/QSz+bhJul2
tkZdJ8oT4VEPwQZF8WBOCN1F5oNs5Aik8GYHIZZOW9t8wD9keTbxfebpOu3Mcav5X4QPzIzaKJ9b
ORGJrkZKyodYD+gKpvaYa37tqQL/oeSZSToDtjM4nY4lcVKL54VbAVpQo5R/hDJY9Qdu6yHkw3gx
f7hjogZJAmZWTl+6LWhWUxb2/nCMkn73V15bvduuxVV/n/66nhiE4LREQnmvcfdi/Cju84N4TxzQ
Dvf52isOa8QFRKVPuxSPAIlEWLZ0gxQKGw04QqbL6FQMzHyWZZ5lEtuPdgpF2WrNh5bsHsZ3Xx/r
6ftCw2TnWtJ4y8d+sR+0s1G2G/1EjR6SyDpl3WB7nZ3UmiFcy4zcrsBdYo4p1uPf+H+tIvBbtVzR
VsRXL7vUaNqgVRgPJFTTciVPlWJ4obcOUHyD3nVfrHg3ETflwPrUEY7YyawmU6C8hJQIgg3XN8JY
KhMfZ41Y0hVN839BwQ+rc1HDv2sB7kJqTKIr3ahWDlTylAclyIoi54B7/8WSLUXqIGI6IWHpn8yV
fRaeeN3yO9F5dIkGInGnzkzz7rNT/XDdV5EdwNzQdhhdl7cyM87ycMfx4phtPMIr2KKgYQht2rr1
FCibPepe8pHvIvFCGwp7OXcqXLYggImOGBg6yBIrHe0iGA7mZqTiFf4OU29Q8SBcfoPoe4rgqGMX
RVXdDg8DDkic+IUTDDEHBybtnWG4WrZRxYBTlgaIAcjTmnbDZxy6ooxCX8r6pe4BaRSt8WZ18zsi
B2Vy8FO3+TX+RgRTj31ekJEQ99CU5bZcvJTIUeIx24yfLBtw0fWnZWpg+iUeqXfN3DlNxZO3qOwF
U4W7aV9HGW0ZBWKKzy/RO1f4qSaLLaNzhRAnoLXLxjtc514elPmRe9f/8FqvpbwZ2FwK+T+k2cjn
LXZzRgCWEh6lCy86TtFGwSJUknIFR7J56aYSbp/12iwanajNE49uMSe8jEObeEtX+/7/KV/Atuov
7vdMrKuVj+9HeFNOGiwV0M5zdWy6ibbAwNJIcXds+uq9qxjcEkMrclAhaRm1dwNAf//GfwplWbva
/0x1pnmtvSHsx3d5FAzCexrPMijHxarPTKlW+PXNvcC91Fo2g5DaBOuCQY8fk4Pup4wbO7uhaVbL
hB9wjLgENU3adosP1YaZYiHn7329xMLEMdCAfqH3Qhq6y9AblCyhs88PvAmxF19ix3dJGxDJ9rDV
wv/2lR6M2npLri7s2rCUk196J5LcvzgAv+bwyljnUCQucLuEK3IkVZeWGwKq+GtIswD+irYNISLt
WhlPE9gw6hYiXoIwxmEszdYYhHb2q5nb5J0N5N5SCDPhn+YHvggHA9J7gvbeqgsH9/5DWbWgCPA7
SGyNGzLyWK07L2B7ak01CjBzm4LgfgpA63ZvXZHr1Fj+RhhCjQSTy6Lz0JZblOGN+VBPDIPk2q6H
kLiCDmvIz9y2kReSgDYIzyvtneH9Ldd3vRobpvcgi5w40+Vx05GxCKPGyZ9shXEiz1ZoP3D3/ht8
b/z5kwwitf5eRCtyyzAtIFEhSfGmX02jMl7QNS+x6bZgW2sB7CCdBAfwY+yjntx7xp0aXFIMU2S0
F0fiW0x9dvbW3u3R4QHaoMbaVfo/b4qlir0/AL0D1FD6HjXYn2eF+UN1NgV5rSdkZu26P+/D5RWp
bv2bWVeznHTwAbwIgIc1ENdow2Yg1bdpcPlS4nEnPBhKzdq8Qv3nJ+rZfUnJbpIk0aA/7V5x0I2H
gnZ+aUzIFWEalVBBOrghBx935hOjgmr2S4g1YGFZIpSyqqB0vSfOt/PBGhbK0SBmDgJUrCEYWi8R
l2aKa0B0XdKZ8jc4EE3U7qsMs4GwWaHGP4V8n0OyPNbtSkC8YuHfjzm52oZD+qqwnW8K2Zf87aXf
M4YkwBfCYrVA1bNi34d9ZcwSmtS7kDQC1rp+0/ACp8MbKf2AiVu5SZBZIluAEeN0LrdhV6ogK2LW
bIXEVYTyD4bH0rw1trk0Rq+mxtJ7nw3EDJpUMmonUsfVq5eXgm2HHDyGt4ingdgqO4uTG2rk6vOT
ZXGV5Qm1hFNt8WawUyZ/aEcaxHKs04UOktMIJP6LAocT/i4Yq2turaz5wOca3ziYYDk5Pphv/fi/
uTLez0k4jofGqQsETjrqfM3zbU6PHGAJdHHgBlDadHMlb3Jo4igEhNvpsLlonDvawl8DOYbrX9q1
ZcZrBSx7nJ31IWs0uacqGxKlGfpue8sb0zAD6GbUQJqWmDviVAQvojbo9Rj59xBMN4y3KEdNxSv+
84zELb+0zvubr+Sg0D0yoNW9IXmL3PAG4Cgw8HU4Fy1WTeKZIh9EuXhaqBLhKldtcgJfS/qfmdcc
DEiFe505bn9742+kDJE6qyi3zF+AziSjJ1iklWgXfzKO1oOLID6cvhOzW0DxCQTa21JHEckDn1+P
of6BST3jrex3/WGKIkWkbF/FwMOViWX2VN1Y3KTyGGSBt1qQ69D4IMv+7lEEJJBH0bYv1qA10Esa
rC8q/bSskswDaa2UbTq78IQnnVyrbXrgj8dLOXvf74HY96kPsVTmxwSSU2Yz+cCOWk2NIARtqI2O
NVHfSYRNvjCB5jNAo68Vciw0HVFoS5tjd1u8wyBpGd/tKLBZCic1IRV9e3r+wtPDB7sGqnpoqv/e
JfHnLGBb9doIFMHbDp2LspPfvIzrmnV0374ZQJ51x6SycJw05PcGf2tlQtoAN/ssq/JXyJ/iVNKu
HCzdZsw0X/mz0TVvVk/CLD8WY0Db/Gh44gHMnD0EAlzYziJH2Xk8wsv/b16DgllkUlhvPxwKHDae
KDbqqXSA9cuM1vuEYWd20R3hp0Rnr1IsjwxwISA3YcJI6yRxVx0MPD+FG7rCRkdVgacF6Dewy0SF
wnZplVefJ4FNhm3dXjlQz5Kay5Ed5JYquc5EZRn7uPEyiRStSsDSW0IjuBOolrlxwthm9uvxZw2r
o5WZylfgrcScV1klEbslThANohmRGp2rBlcflrCHKeIGVUqCBwEXYM1ngeEGfjkZkEBt4TuWNOAQ
8fKExfBckILU28t0vgGO1PHzETaU3n8zbkC7hxXXRZsKTCmGSaPkPJAv6xb2oj9Dc8GjrIjP+66O
nl85LHJV1Wlqz/HsLmQWL848guWMKaMLZ8ChjvmFePxiSGxhT8SmJd26gifqfEikle0CYjGZNE3j
AZgen4EIzHizWdFXoWva05bGmdPxrVklNBIXuuBaq91k5EwzhrrVocelNGsR6/x4ycfefQi6kwA4
ZXy4CH2rjB/zaLU9pXRvhhQzkqSTzDZN6nC5Qs5t4uot7EY/N3IwqJ18xgKG+Msipi6jnCNCUnLR
vxQrAk5rAlJzKp0sWqmttZCCG/0V5h16zFY9xoLmop9UNnhs0GQDQ4hG6D7ZDcG3tMNvyQCzNQ5f
2+3MOsGLYuuNaCUN3VccX/OwZ1u6qk1WuIVnb/gQppkD+lum6KN/8LKCCa8Wq4OZ3SpTnuAgJHrf
lkTQqJiVvBfY+Z2fW1dY5D/A44PAoE34iFpuynGoQ7TlHXRWsn7noVlGDfPPwIwzX9kywqxsVpIt
HocF6maRjpYo1nlF4yNEDGEF8vpnGmpzygvVNSrnIfi+6jB0HR6PS39ivl6Oh5dkqchfdBzVCMpJ
XJAQjf6n15G4Q9cVair8DVn1iaCcUj/dP4P29CrCGFf8XxT4dtJ+8wg1HkRtSDl6C5kDjzyzIIN1
/DLddyYqTw70jTnN4B3pUPTGm1/9TXsO0wB5xUgWiSJMnD255K8fVfBMzuOPNfNhFx3unyRg/w78
DkxldzZINvrqgvaiyQdr5nUI2z2KsuoVZeslYZ+XOC20Iq44754s/Nsys8hVq3+WHKexCvMU6Ei8
3GKX9gWNb5Vwp4oB8Gl0mMf/UnlF0ffd/V8YTG5UFqGwlgyS0VD69NOxpLH4VlUjTLTC60mYpZNj
RXrTKyL2Jj/TgN9/1IoK1OE1lyIXTWkJoaCRNhwo8eY39LPy2OXxAK1yvWTioOQF4+fw6GNmb+8W
QIDYOvkYFYrMkrfFnNPmrx5B0BAIfsjht6YgD547HYZwlGX+tgTtn9wN4Ari6K1/3uXYMsXmhCx/
BIQjh/wALitiAvL+EuagwiqoJCPJGNUag4IHG3KvUO4MAucIHN6QOkNoLPfPbVk1cHUBqSifvtw2
MQfbiTmU4T2f17+Lzdykm8Wtn8HPksiRBGLKlXcB6sT136D7Y6l9y1Y93PWZ1NRu7AVbqWSk5+jI
HXQJJI7x/qnej+ODmkvxaA+g7IUU5ox7QBpO+yvbMp0n3ANDNLwKsVIbxGsA2i52C1gzRyhfCZem
SijyjPMqw031tgHsfFixiDBe7HYN/31RtwlokI43aUYrg0Cfc6u5sUB77u0dImG3p8gkEopkhcyZ
1Sg4LSQRFJ8xj6AlTEvFj8svJwt6nkEMCR3ISnsbpuhQpxwv+QY1YT7g6FAgFhnv5bxAOxJyAiaw
btX7jKYqeS8QrgzQF6xrJj4W4AyMqMtNRUc3pHCqkgS0nMzKg5AahREWhcsG+2Fm1hgghi13dqAC
X0Kci7NxRnwm2lkwgt9trtKxyvemMwUqsLDs15HQlqAlCrAhzaPnCFpGGGEmC9LHmXZy7aPLAzdz
EGbaGl7ZINng4iZA5mCQFZ62FZxQyzA3BCit68abKPWKl3FrV6eYw5BqmNW1PV4FqOrF7ZaPMfyz
+XnoIxVapjBNM5z9sSAcr51uNM0lHpx5oWOxduXQB8MK+D+f4hri+Q1zYAAAa+4OQ7DSwzZKsbbH
921EIqMEEW0kbSlKsj/zvCGNiWv3tdFpvYbG5HzUvx3FxzeC23YaZHlljONFyCfrIqBRbZ0Olz07
KuQwKqtekOKOCypqsI+7H/u/pRa2RHOPxYD7Ni3rAMvjPogEVF767/gF1PToIsSN69UU29R+XWGd
niTZSzafcRPeVxotNb/1bZfeSkf0cCy6RbENRxxDyhr/9VGieAssmrDXWWYmh2ciBYDQIxYW3h7T
mF+eFmuAVYg+x+gYif1TTmxaq+P6oCFLhhWiUpHBsYl9hCQy2Kf3BfP/ckJvoQ+ahver7AlMR4my
zS87/knvlZATfrJxVL9xVc6KDMzISFEdnrsxICxUPzSYf/JmTOzpxegthF2ocOi+vUNz7r8Bb8g+
gHPpEhjRm26BP/8KyFwVgT5vXna5XxXui9m6PA/pkGhb1dfaAL+PxaEgB891Q5NnAwEd+6dqlz4w
5mVCUKqJVKbd2uGKrQfP9+8q7F19OKTCokSqtSIo0UTUrVDguCpzlPTDMCiQvo8Yusgi+2z12C0L
YEsFDlfugFglTvBF1blHsytv57OBCTjFMaC0fMcf1puaBzIM4o8hegvHAgvTreWE5/FAWrr+5NSG
femhT0iftJJc8ck9xH0FYsBdjLCNNeu4k32I+RJSf5dj0gSTf40kXPGpVALKuRnmbzyFthCDGGqi
UFLak+oy5mKKleT/NL4720Kmw5HbLJ3rGnKJ7+c5ZvqIqjxCqKZm2bnGe17oEawr/K5KW8ejSk2b
BKpiDyYYENndz6xguxCCDCFGVaVQVfnh2Z2cOqxfwr71LRDOIxA8vxVVVHVDDo+eOvxV3MnNWEbj
uhusNjKgx/WkcOUyQuK6V6YCFcEgrYaPNAdx0ClCrBnAdOcP869qFHllu28wSrweaN22JuMpCfCO
ULCODaXsdIfgBDwDFTw8s2s3fTkFfbl3dRA4HbED7o7TqyGetwlTmT8JiLnWw2TO8iioXJqupHSh
VxNPV7lymajSqnO9//g3Jy7yz5doQ1M1qtJkdrWILvp4zfWt/1aN59cv1htpUT6/zDGrTaJwEbFB
J5Zk6N1+pJqqa9Mt/hBYVC1s3SdCr/oXdtDv8dgubGQk8FDg/jCspAp0/cOrNEkqMtM5V0Yhisec
/3xvdFBqW6FxibS7ovvrXmXfY0ICm4QaZWntxd6N9z+Gfh3q84GGROWl5jxCaVMjEaUTxE6MiF+Q
f3Af0zlfwmKgpQYvk02F1Nrg6uWdZAg0hmD5OCe1PyXndlFl4ObwaB26iTFfcMzvKtq4fSEHUD7I
2ipL7WCl6V+lYDFGh5kBQUs91SLjo9Qi8zJkjAKB5zUa3/3aAc3Yn+duXFd9M+VTYXN+YgKb8JHL
q2aF0n/5JdK9T5idJh7x/XVPQbKQcRPyZqZIDN5O53fYRvv537nQ0/pX/7/MZQUw3AsaHvU15s3K
Qb4Q861lDdQ/aXvZ5gfM2GoBKYaBVqwviXt2aMRKRLFSfL7WD8PiMkSv3FGG9mYiISGAxeQk1Dww
08cFOXRVNKCCX8mlTrhDyrgbdAQV/ZIiPeBq5ZCzAN0DSIQdXz9skubcq+55PID9Db01diD+eQyG
N0sJv77S3ix299UJFSsUiAvFDptEJ5mpK77+27V1hfuZJunoYztwujserKvmbdha4f+kqKJjtRHz
qq7GMvMyl7ZkW3GGg/wOOgCGlZp2bhS8wtjRAZEIX+zvYIUNhJT8svsZYYPs0HiTBaN6eok7GnjD
lP9kQndKqhz9MIxIq2KnEvdWsjvTF3Dl6gUHGTh7LZhU2X/7QHQvf97vjbEHVxtNw9iwIQQCsKut
FQNvVA6LqXHbaD5VyhJ43wzdxrIRB/EkgCf3MiiCmgpLfXGze8NcKPejR3R1x1kdmWYiXRttcUHb
4JOiffNeqMT/qWNh3Sc0Y1WJoHw3K1vEl5KavtrLIakZbwTf9E1wqieUw0JRzDbhTaeBGqrLf+mL
37cm8A6zNXoIhJJpChuVbuqZZwDw5+s+/mvi3pDQU5eo5TWw4GOayIYIBDqPN80yCriXTdgoz9X2
S2iJm80Xx/ks8T/S/iK9vCCmQ56rU54886YaOMnemLQkvr8yHPe2F0Qdm2No+rAkbyqtLlldbyfh
l/965G+kXu36cl5yOc/ZNm97yiJ1+Wg83o1QPdNLVGQVW9bKlLG7lhZ58mxJfXo4Ru1O5qSs1/rf
tcIux7b0ckL1qG5076kvMIUQBk1NU8d/iqt+0SeTkVHQtXOYfOltEPwFRH6dwUUpav3VjR9sMarj
k9nH6biAVBjinhLQXLDldsctv2QYE24cwuCuoOEYbzBfDFLlvX1LSjNmro0o7jId4+yjO4sniuzF
fQIFMsBMtFjrTK/Zm2LsNzHVWce0S5OuALNQt69c7vfPXeJCHcABnpsK+sL7gE8g8wiM3viAwkcO
zGyNVgDTxO4vFhsOFxtw8MdYcg9lcMEs5uvWiZdmxiGdDIo2IN3AV4r/r7MjTzYIJPQT6NeJ34uz
eIHur6x8S2ehqrL9/tsniagc4BM3VyPDXGjQ0da1ynDoxDlBe32IxoaW/W5Y377uGjLzAhPmEZ53
btfGL+h9xgjOY4vEBN2v3WWqvmZtgLMhGCVWooyhDLaaPD7r+KptEQoEMsly3kNF4YsIbFhZgref
Ww501e9gqn6otXtQPnSGkpI22hlofHR9DYpTHwfj40m1IemkM/RqFYe0gO9dSrGzyIr4xZbu6Ehg
5C9lXtIxSZrh3dxi5xlEdQlxw/63ZoIhl02VkQlT3KVz/LssEz69M1OrU+jDE8HRSXrQbBj0u3Lj
OXV6Wc4Ific63lM2L3jNS01ltA8sE9kYW8aOizKHHzB/2Wgb3YpKq2JatCeKwDxfBp2Fk/YJTBEX
KYIOXMUV7rvBVjA5N/n29HTr82OsRc0tSwUxgFFf45Cy2RODO+NtB+29jLjTzCPmHipKkCYOYa2u
TyhpR8dJ4yPDTWil3MhlTEWf2xQplwtFPPGe+WX6PZszJFtZOMFUxZz9XtxRQOKdc5gKNjnO8yzE
lIPX9e5sFUl+q21ItMGT3JW3ueQAMJiXz+tl89ZhhSacLiCkhV16ZzLmkPXVEuprx+Wz7mcdAtz+
j16VWDSjqOoebCaqOE3LWBfrmLg2LoX5g8GcMfbVZXaQmaTSyQ8s6E/UjkfYafr9G1x2TfV0l/9W
OLu4WkFc00a/MfeJ/d4X4Pt/P5P1hkLAI83LkDtRyDv9jnp967ngTqtUigV4FYcv53hnsRgzcjvX
IPfm/cdruN6pkjMxK6yESHQAQxbh9RTzSWVzkAbv0ttz6eGDiXES8X4oAt4nXEHEGy0OKTcmKcxH
s9JOjhSwJtPByCq1Yhpm/UY9ilUOmRTdM7ifhDgAwKikwHc4SUhfv+h3U9V0KJ3VcS5ldVfcXAq2
r2b/MLANwGvsVRRWBexfqbT9SG1kHp7UPx915JvYx4RFlS4SGlMZ4BBuuMYJy/yA1rvAUgc6AEob
yrAWGiVEZP6oAhdutBaaC0z95BrDObb2ySDHYR4m3zZqNRAOZiIG7ztLq9JOhkGUxqcFgZDEVdU7
4K0jfL0JVJi0cCrnx1wDU+1Qo8Ja250guxnpjx3n0PSw4Z67R1rm4bmNnDxgamH1VmDPOrF6vQF2
10fXinYhNhyNkEne3mJ/OYJiHUQdxEl6+KOV2qH/Hxr1E/c3fXTzUCXC75hA/XDZIBu6HTJSol99
Epqcyn0LNyAQzhegaj9w6PrLn0OA0RmeD/ZQeDEhZ/inn6PGkIpvyvUYpkNQ6ZAF4LC+hLms8jMD
ELslIqHBUaDZgu/p1oG40iuxnv4fJpWw2ekFpTE7cZMDnzx8PsxRWt4ZMzwVqvMyRgJDW/lG7OAp
3+LKQQ8QVlhuIcC9gs/Cx3cTsbhei/nuFnS9qyIFEop1fCxyHjsdo0jVWjF85wGZI/yYBiQjp7y+
q5tvxvpuoT0YWnA49AKFpW3UPn5LPD1FN0dEwOB0DK46KkDMY4uIUgPhzE0zZ2rrGvR2Ho01wbkJ
LMBO1T6fHnm7nsq4aZYgdqZ81GUKcSoC8Y35D75KzioSfi0qOOvvWXe42OE1Pm1Y1jV9VnV6m6CD
MbCgmzbbP15gLz4q0gnHjEupOGhDSi/OfnOVysUUUlsyg34/R2I7MXEMZsYCO/9MZ0/1/HNNL9B/
AsZrm2Uqya5EYpP2Nlk3UJOKt5De3q17qT7fKy70sdy/WgK/aw79Plfg76pDygK5UTblyYOaDgEu
0d92Lkz8TiDe+OD39zrqF9tepTn/F4eIpYAz5nJKcT28tjHcsiXj/XqfhLcLlG+CSczv7dEbpVP3
5KEhuubXMX2ylz1xfAgT7bzBtr/HmAidPELO1ILJDlznxEDB0jVBN1+q3TzIQ8H6FlAcR+2dEgYw
O52RtWz/M+PaXV0/T32pBXxFvFFHV/nBY+vVD7Z70WXO9y5l+naP5syC9XQPw+66Owt8s2UnuXQz
/IiP8Zjrxb5vZvPHDJ29IJ1rsqKsaHxQ343N1EIlPvis6pbCT462VsSjZQ9Ykn1IHeg5y9t0JR78
CA4DzrStxW06hKCcETQaBHS1DRijkx/hrkKwig6KO1vkSf5Cp95lEdlXCbIm8kceHQ09v1vactzU
O6nbzHKiTf5GCFUvTWsXO0igbneBYjBNoCnDl0dhCPcWlawsC5I/qlPkxRQV1mBp3df43fcCbU9d
14IwuRgyUkZ681zjt1UcxoiXhfIUeh5+RFRjOarnCzmT0/RNn0oOcL8GCnyZfHdVgQ4gWbJW/jNu
gYyd/T5h6SAgEbufg/bSqFZKsPmx/vm2LxcNe3QWNNGZFYXcD5pIktlaSaXWn/8NZpHROm9lbMiF
YbpIOwwiMoG4ngsRJb2KU8IdvIpHm+IiNio9K/hSL4zmpZYRi+tKP0tLET1DuaoGAljjrps6f2yd
p3LtPW3LaTT0o3KrGuFpybedG052J0a+Z2h7Cw7HI0YDpBsrIVLdxeHuicdAQf2aXkhdgRUoVluC
uWXlOLL2+ld+r2FPYhTcA9Jr2h22kpIPQ1ILIGk2aPCP7YyaamGUUveg3yuXibux/Otxxfk5muWJ
nGyiMorSATi2EQvyS2KFNdWgpUekgAt49LR5pqY4PNWYZNCXEn/FBnWDsCdpYRUpCQ95eHJlGfPM
P4HrNRSZTNzzRqJ+dh+D6tVtXGvRiB/Ckzd0kxPimYW3E153O0mEVzmeWusMhe95AhPAlfp/Teti
LIh5fWlDK8/iF+eKGCsxFRxKrrhfrN9jTx5g0IPFok6jMOl+FvUa4RLB/CUkz5G7Fqb6AQVZNekX
JidDgarNm4EWc7mDmHJuJCgk2bkYERZn5cvNCs/COczEO8a1HHZo0kpLpIlChmkIj3J+wTBgK4zi
mvVxp8yYuRsJ4Ory9bKEkf/Ti4h1IBv0qAarRc50EnfBF2g5NVYBWayM4cHChoDtE5Omyb9B7hdR
bHMItQDRENfRZjMilgbZNnIQclxe3dSlz5Kzz3cI8dQzJ8GJs7+YHPfzd+DiV5i3z3LuSY4hWeMC
FfDeTPrDj1GxHN2y7ByfsXrzWPR1j6j5f1H5OyIeHlc9Erd9DvEot8knX4anEqUROYUnJITTKhxg
nSuGQYGBYaMhllXVkjSGkU2T9IRQTIpKUyA+2h5NNIpxhrJLM1FDN4mQGV64UsfYj+s7ozEaxP52
KQWdaiiSf6MEwrgs+VTtG2CtqC6L1smTR0c+b9C8OvRWAXDy1RXsQMepQi+aNQWOaX8Oy/1OVdfv
HESeOBhseAY9RVEtv43if2EVrEMFuvCui8HE45isBmsgJdcQg8EuL9Dd0NarMJqPSQdCscQ5srng
QbmQGp2tOK1SxLSlW0fVtMaGxjoKMyVDT4gQNT8jMFuJjHsMByR6zjG8ikK158Klh8fxbHOklOVT
mVVPuwdKyof55pShAN3gYIk0NUScbCuoeqrAOitVZD0QV2jJh6YxoXyunHyf+55AVNFgPI0iH/Ja
bTVgtH+1w0vmpQXNqwjfaFNZ4cu/0PDpIk+Dpjr0g0XxILgb5wzH4GM8pGR8NnODeHD50rR9+pxJ
3mR9gwX0VLfGXqo6GZkPJUCULKa0QxSKjrN8CZHdL6neGbhk3uzS00OtaBCrN8g8ti0K9g29Hv6S
i1dgHD1ImLGQCGoiKxY2l4Gmdwi8gv3ob8ss3HVdLuHzNbl95IkpdNoILucQcuISoZG8o6161vvb
DPvrR9U277cef25joVlDTEJGaV1AUR54aCV61j5cs8ljAyMdI8gv6EmgkTTQ/oFvMxa2StmACP1K
jdjDzqmXeUwBfNRX8vQO0IOWxBqAB0eRIydBlCEiTj4Mb0rwzX49hLljSNJIAM4uA1omJo93Gfwl
Kmw0qIx8PycyluoLtaUCXzwNBz9aWhBHEIOaGDua4WymvLbHTqrmUlZtxDS7tK+M+JDGYbBV8Ng8
O6lG/DoBxgt2QjT55QpNgnY9RTHpLpRo2VDFtyWL5liG0qoycLsREkO6grI2NPRMQPAuTPQinXTF
aB5pMBYVcT/I4AnQ3Las9z+MQJ4GnMHOZXFHg1bylixt47hku9hShcuq/VLPYMWyvOUghzD8AfUf
KIMBe4j+8tCifFw+0bIVzjBS8jc/2ugxWad5ZQlFNDvB2iYUzIlEu8Q6Ve5/L0yELZIaUo3isG3j
AtB0wxOkcttJ0wCowDg5aVIYxsTRvh+hbCyJYnGAXUpW5QARY5KO8Hn3WebgEWeaCWf0EdbxYWU3
A6XCoDJzYKqGc6UuqT4jHEPLTaJ09GqchTMaBt5PFm/p6pI/MLFQzTIk2dZJlJ7EQZvTrBmBG+TE
oR9mwuWpUCTC7g0hbbp8brCpipQfHW0WPKcvwec7Zl0GlY8Nl0YODzmxNG5uW56AVSLkrmd9tO+k
014nxZ9Vc0FY25wsTSNNhiEF+qPHZEuRg6WW9dVr0Nrd5f6hqfIq3T7Cjt/ORc/Ffo/FZP1pT8Sd
npxfxGC8MchxmidS2OWpAwhs4gwSfPTvFjSSizvz6lwffBVSWDEWR1fo/Ys6K01UdeXbw2qqtufd
xT9tlcInB31NfwosA01845vuIGAUiibzgHZ8OkU16jIqIt51hBxCoAx4sqfyrT5ZLFUk0YGqtjIu
WzWuUY7yoHpxYYtHKZRx4ktYchpTs9Tm0uWgojYIvBc4WxJHop4lxZ+By7EbJiPnv3QyIyvj0JUv
7SI0Y8n1u0FfEc6fT9GpROw3jau+E8TP9uodtnpyv7/39KV5y8nh0OVk0a+6sBqRD0mGClT3Vs0P
Dp1BzHqxJOpiB2xwbQRZlA7vUI5pZKmnwEjfcwHtRS4TzZP/kCo8u1OUv8LrDqkKqa/wsrjCdNyz
bXT21BfVqaSbRvSjvBPRHcNqiU7hn+IHWFrZTuU/lNgyWAD3JmIwKh7m6cFCTBJGWdSR12dTFqk7
tcaPjANVgtDqo0DOFB7UuaCk/OuGI1eb0+JVP8+UloJePWSMlE6eLSXBUoPA2eqUpcvDhsmTSikQ
jA1H0vmcOAxcUVq5zKb5gQnf5DGf399To4bkgWa0Y8F1Wv06BbPGeQYn11yr/znsav0DXf1ht/9x
ryD3FCrj885PGZ8RiqcmqrxUlCqcnxda/8alvZm1SxxHXkmT0mAYmwMFcDzuRuyvyXOiqMd9iS+z
EZo51CVqaaOWXJcnOgRrJhEtabS2zv+roKiFPwR7xynT8S1cffNdtK7HII7el0VSAxMEEyS3OIQU
+uGdn0xyCXqhsfGtS5PerK9nqDHMHY65I0dE7iTV1wk1hbBmlZBhwEmNqDTUqf5ux5XzLwu4o9Mk
UBTxcTW75Yj2NsZOdNKOI7N6TDiWIk9Rr+LIFUODsDeJgqCHhGXGFbDQXYmMvQsHmdITLzhVtXUJ
3MOe4LyYa62N9vnZm+TRS6rGBFcd20FageXVrMSXJc84aOrE71qat7g0yNsDiQiseZGT5CwSRtBS
mEor7G5FSxj33qFE4vhzHSoe2g/IImR8/njxT6bVngknkJ8oAdi25Rt/k7rtr0DhjO6kWOZwB33q
XaWdUeyPV3OvV3eU1SN6mR7PGITxuKBNQXTnSprvh/FIm4bMHBH4O+MT4sm8I50ubq/NDLYfvnKd
HVqbqbV+dtvcsDIdj74OIIa624XiVGxqdJIg3lnpp/MRZJeUrgILmCz+BKwRjLNfBVBDJIsOQHzX
sRFvbukUJq2f4m2ohu/jEA67spLtBCcFAATzB7dyOgGiVid1N1u6EwRQEp0vrZkFxnhuXrUgGfX6
I+Os9uafz8Qvc4ddIU/NjgElpTf44duKOdM6MdqHqAdCQgIYY5cO28BHT+apWPz+56CBs9zVi4FM
AjqkxjLK9mh2qFtu6qkCT0gelfrHSPfnHrzId1t3Xp6GZCsHsSKflDOcG/sPOskVoCqp+4AayTOw
i1Mnb2F04DHSB+j8fYZVwkWvRV4zKuTGsSxnfgm+69vDfkoZQfZFvISPglKGAwESDDCbLsTTb9wB
PjsAtRVfQPk/f5YCwBGganLf//P7gYzmwWBThXh02WGNyR9Xy4vDO4WMN0J9s01j+GRI/5ZIsv7k
Lme7V+x2LufzWcHxz78igBKV2Zxss1rV7bHAf2SkBZHU9ea5BDGM3ki7lu+CqmsGGcuA991w/3Jd
Kx/Vvi2cjUwHLWErGkaink63yHAiF7Wq+x7ENrO8MpNhKjVVbpEbY9S1/vDzENZ3tp9XgCH38KfV
cXPKCfKmZLEc11T1BRIEnE9knCYb2FjVcrUmrq/OqQhVnzzlsX23sTqbffAbvrSl62HObifb6x8y
jz48RwfbKZ7aod2uMU6J7dNdqqOQUXUm+k4POs6KiAnfCm7tHfzHKMXTIDAaTvUKcCM8ZHpdkwCZ
EcgrDCabMAiRBfyWGuJ4s6q2M9dR0WAvwF6gasrPoyYcZ7av6DpzsHnRmQLJzf7nH2802hhSuFta
P9K/ePwqeamI8yeVLNJGlVZWRBIB23t0Y4mb8k8Qc0a6EJ7BFnhBukxaToZDmfMxsehTVFwnNA6n
68K/VALO55Pfw2Cv9VTL/Afz8S6bvJdAA+LMCusLfH6IJovKzqXw+0/8lyd29xXau++EZWF0Rf24
2ao+HVn40IvAwCkpm3eUOtQIk0mXCpDazMMHSLW0Ptwnn9sNJSvdEzZfIUxkRVxQzNDgDvHo5teJ
bh80pMtVttlSuQq19KdKsb9R8o3mePCvuPa1gzWbBvwoXYV70umhjTtCiacEVOxluThHKQW/tw/s
MdGWqZDMHtdlYDmLv+lyvZnsk12HLASoFMdSIDx1scJ5BUgRmr7IwcPC9B4tPUmtSwSP6x7YnGG1
d8tv9td6kN6kJ6sBpiUZL4TPaIIRnzZXKi9ojJ6ZmuC7afcjkbYEGZk8lnzYHAXy/8curkiiuTfG
pgUdi2wZOIgSL408z4LYhXbEaNsGbTpMczsqWbRxl5k4IBaWQ4GhF3OjCXLvj7D65J05xGUoAdQd
yYIRdzlZi5SHifhRC+xWQ0IpPl3fmp2UHprkMNtRH22KyrkVd6fpY48pH8xcoZ7VrpzIlP02rgpv
eEJJMeuI3FjsGC0G3KDeSgV30uXiRYFhS3ItXyw3VzWVRzrNdIcakV/AGjYlpHQy2yDEAZlxUcyJ
17MNgoBas4HeIRmsdzL/ZTQNiILodY7hzlBlnfeWIFzTd9QRCn6+cPX33VNFlGFwFRkiIHSJ+968
8rAVqy5EB8qfm18/PwJLgmNbIXhQL7ZYQRHvW7+mmUssW+AGBjIZoNEp9kHbXRplNYUSnyHPvBnX
adu9/FOJMsOGAAHlybsMDzUDQckV+lWiiLzjf8WftAeNKA0dt3b2XhilerVh+b2EPCXAFLJnmVJL
+O6pB2nXSeuIWsp5N6pem/NDs66Gs+IavcUe8N76XVW40HaWEut2Nd9EcGU1e3Fc887p/f65s1A+
g+h/ZNgjLDfam6gZBf3kp/c/RdlGXM1wA8NwjGWkDXUhCexAhae3Cs+M9g1cBqpUG66icnLx+aTo
Qb2HtzuVm570yE+98Z6vXCvc20vFebuj40QYWpF2fZF0jEa8wYDRM45oN8/z0CUX0TAyL0/Kqbmv
ccI5jdaYvxrFI44DHcqcdERqmQRnYcJYFWqhDf6VdyGcxo8l3NBqN97VM8BoyPBCsBzHdCri8L24
cmaLwEjMv7HDc6erEMGWlV5sHbJm6RDFMAanljnxizuZRvs3DNoF4mp0wqiJTGGxxWbbVWTU6Db7
gkRStk/jRXgPRfnK1Hp3gSj5AXvwaN00gMX2PJdBZT5KSHNhToggZ1lIOHQXgb5SKsZk2PoIncLS
yBBIThuu0ljeoXPtrTsxAyXbW2PY1Cn65MTcYLJkMm2ugkrQV2atbSAc/Jf3dspRmi+Sp1Yu9PTa
QSdZFFVRjccE6YOb/mSwXzXi7ZOFjLBAsMGgpPSNlJm8bD8KTbKbgaJMWstI1px2Yv15qO1glz5b
PF9OQ3EYtV28ace1jIj/A16grGsE2EpTwW7QDbHIVUPxgAzz56bSfpioqISoqpT9FPzjy1oq+yII
3qN4OKEYqK7Fo3gUHRXoZQASL+keMQjNBW65d0csy/E4Jz0UfzuHH3Vk9Q05adguHLoUWMAAYw84
N010KWUmzGvLSKnTmjgooz28HXzGy3dhwsE1RFS8qD65ugxB/lz25Yw2A3V5K+NXmv6p4/VYZrW6
lI1OpO1ezhQSixPYysrUCyV/eenk+GnhRPhT+DsbMhsGpV5EhjZBymC6lz1bMzihoNOkEHLWNkYg
tJFzF6M795yk9ap2TXDKxc5SgWIA5lnP34HP6UVUnJs/W+V1ZqYsIUGBhwrBaWqhwkg/Mrh/qCy9
m9kPN607Ifu8mQNFgFVJOG8Gp3aMo0j3RFJJyZDsr6g+PPSmV6/Nv+UqUeqRvd5vOwJF9eDQWZzX
9ZjTn+kGJcgrwphuGd+IXeVET6Y+58KWRUh17lRRqG+y/ajOnDzLrdbXjmGSMhNXC9mfvO9DTSDo
7LPYtaLSCuBlFP+DCLRJ15FkRuJ43pH4qPeCydR8pPuU32vp8oUX0WUszv7wVD/k0Nk0YWADxDnc
3gZFeMLZITpkLGwPfRUv0uOemvFJrnkygymuv9qqDycu5drZbf5oIUFEXEK/rRZ7dzjLH+4LLIG2
zdbcSX1yo7Qsd4yPMfGIKZINCT10BIefTrz7jvz6jrFdiFIiKUzwGNyoEHwprTNUkI/2rDlLdKmO
l5d2k9s2uKJfC0S7zsYaPXY2IOPvv+rRWbBtkr4WBE9xn9ElnaAQrPqfpZsZmyim6WiY9utNh0Eq
O8RFLrLUAZumTrajBUGRynWe5Kke+yvz5NYUG1PAfw6cQHO8slOn9eoSzFquMQd8S343C6fqK9tk
Z/f4IprNczKT80Fe9FdH8ffipcUVwnFFICDVRAJt37MDRfbS4XkzQlmivw5bveIt5UrQn4XWS+Fk
ne4pW1QzNBM1aJ6NyWj7n6xKfMCbGfc0Om9bG15wf7ivklZ5aQ+EYs3KbOiLc4WLUkvZCE6Dd46b
t/G8p/81mm3k7F6vjdICahaDjXD/i0eprFKltrccA+PdkebBDHGACENETeEs2cx5uzNJ+T9FKBJb
Gr39FzZGYxspI0vRZf1QIeJPZewBIKjg834jqJBP4o1cLdKAltN6vivgl7pcb8NRGSvUTeaWovdV
jL2MfglPnA9oSlWJIQmwLSOcE5+l8VdZHjsFIe8ppnDz6Ppy/ep2R8mHfxPofKnXe3q4kfEsNfm1
YHaFxr9vABK6SMvVfX4GES4gAL7t6fXLRO0T8nOXazGqDctGj/aGLorbI4aKG3XCmBqnv2HLRXjM
xsWhBTNOeVkUO50WABKLe8ahaPnN+sU6MTSRwL4q8V1YCym+gDFj0IU8v+kt81QQ9LHFiS9UM00p
ErR5Zjzqjlnqt6kFakOXWubDkKY/KT6a5uNWkO7PWYPWbBYcAHk+Q/La2v9V+39E4y4p0ZuhmdgD
Q5VxaSddYgrOvsZ5OYUu6vHG5UXtuI/i+2LbOS2cYEYc9fyCEqTGvSaubCIB7GKLqcHLx0bMaR9u
mA++moIm6ZLKJyoydSQf3zyAc/pZA/MbFIZQrcnc7u01iDkLcgSOf3P0lKXSXsKi7lRANQCRv8Oo
VUid1LhHvLkTmA0ZXxNXN3pB7c5LRRpcUuV2+eKCUX0DXdFTIYdJcLrAsGxpiXLVPCYF7pCUQHf1
5CgAigauo/q2q42cKCU4xtK8L9SUdBZAkURfxlDX+uSvN+gXI0l1/W6CWNZ7i66kMuLxJnWaFyOU
0qQnNh9RiHg4caxmXt1UL/grwgbU9Neya44vBEzCGHu7q5QfGhoPcOYGNySaDujKrqLXZT07n10e
VzcfkpumQZMRDYsgd//rbiKrVJO6Z74Qev57HmCuZUdUUgoslTxCPEjj22ZNjwE65y4HQFIlfe3G
vpaD8vBvu1Cb6tW2T7sjz+k6mneHZblOenxeTTLC7hSNXiLgOpHh6Tr5OsVk+0qeiZsBGVCoqqly
6eDCY3kImAvvWB4EEI2k0HgiYnLiOn3w5UmVO97WlZ5gwzEYepZVDAKA9+oiBvyTUzsS1zLIUHMl
KGB+86u5Q536w99AQv0HMmE72XBccPuWbV8eRqNGkxdca2gabHSLqgOxaVV06JhWd/R0zVRnNzcZ
jHJjWsiuHkSXMx4w5C3qaMgGxcX5YNE9A2fyAbVuzKECzbC74dojcKgAnN98UkdO/DxfdPh63q/w
XSlxpGAd2vgNvyc5SV8BF+LLQifNG4jiO1feC0dI2jjQMQxlfFLQECk2KyXRXRRwmZ4hL4K+gouH
eBzqPcjfY3wiX5qS+hI5WGmTy6eKecnKlFLBRbmLm4ARzI2lF60TaAkz536xURLhMYReqOncvXwT
x3iwnYCwU3DhvohoZqlwNKdSnEEpWZkmDR6FppFRGhEnYqjOQAxzuHDu1fEdxIl2R8CN6b3dHL0b
0u6XxpiG33+ZFkIbCUbPmFm5Oe3cDlkJ1izNJW7BLjdQYLoWz6+9s48oiO24hbAEZSM56zC+hCKQ
hwYGD5w87LhohZAatawyr4pyTD5hrLDHwJi0/lrH12ySPsdKEPhKWjHry8b2txMX/a5eHBrqYBJg
wIikkpHryGfjYqaewq6bG11TwkpTzcXXRDXWbLNHZmU3pK6jX+RsqQf+qvsjV5ol9pIro4ry+mX+
FZGjowOuutvQHIzN0JKU2DYGVau0G4VTsTAJYPXkWc/1O8DkyuMUMWFOoCxSvp3j5L4IVtPgiA0v
8oTD19msCHlBMml6sATsgyKMK4YdT2p7CZoiJdSC02Rt8jEd+GpiQJzB4A0agXuVK96nYVl2CwrG
o4LnhS/CxO/flmv7quGoPP+46/FNzLd/4yS4rMCMQNiYNOwJxzDXKpWdXR7gSKURmkVRBXPmFmTA
A7I7IMA8OWjT0xR6EhJMLUiQAsGoIAWNzb59ZficXuD4J4IARuOWJiAMEQW5frxRE3G2zcDVFPmn
kA7UXEzwI17mcif+y4g52koBWpnQWpNNAw+7BFfsZxnBLUjAI5Nfsyf1xOXCXzF74UYWUTZLT9eO
xxma0XuIQx1Ak2tkRNLXz/Gq8BipLPnkpus9ZToJKQhv0RozQDarWH0d/XEqkMvwkZtfrezSi545
GmeWqUOIkNWvQRLyi91ez4MZ/M6Uhbdb2BWHB9arc3DfB/5HrQyzX6KH2q5Bd2BkIFgJMJojXbXL
PcWa1K75ul8Y/I4TmODcnl0dDYCa1teR8bFr3kxEsF6AEDZvXY/W4AObJwudtvS5ZR9q3ObZNV+0
31AL+rVYmOycoKY8g2DOSNXLQ32zbxCnvU5MKfoPyCkhQg+zcFX1SZ3PxRhVOYTKpgL6wJeqYQ04
8ss1eJChoEdFdRQStt0RgciNMuROWX/4krUPA8W67aHLJNgayQnNwJfbDcY0Sjc0eQGDajZbRkM7
U3Rpf3xdXIxsjuRwZgdsMnxgqOKBt60nTogt1wKOqZvMVEa0++nFJ6Ec/8tvHdbGghxgvU03NmUG
w9HYpcJsSBZMmA/XdgKKg/vWCxNKi6RpF0tL8Cud66GQqsuS+onBeiutIPRi6IIremeHKD6Ya2Za
vrMJjSjmbUkZPmXuCBLH0PfnYNTbJPvsW2jC0z1eS2tYLmCBK3EO3ZeQIDKSO3ePzJ+J56a0+1sm
TeLr4dV/72HeSIqa81Pp4dj1Ok/t5XhXUQ8z+OQQZ6m7aGR9gvvTkZNwfYuvaDWL3V1aJ2KJCr1O
W6yRKv1s3uDItCH2Ovt665aG4oTiyKGv9VidObu1VGGq1kEz9gI3lSX2vzD/DT7WUfKLLb1GXET8
pU7Vov1eO+N/BsAYQeuGkcaX8vwF5VdtyINpzUiuDxULOfYzjXfY9wPxdKXQnfANsQQlI+9RKYqn
GyMXJhgmNS2MvNyBFdDLMEjFKLi54uHSDEzK3Cwh5Z9Cn8PNFo4Mum0HRsLfZ2A8TAt9JEuqsWW2
YJAcCx8IUQzqllPt+QI7xCbVBLzhXzXYnq8sD8te35UWRmiMpsMJhBWZMm9i+OUdTQvUlcMFNhbR
olWuAYHKFZ/sNflWU3U2CSTl5GIwu07w0T7rVXuHiSgxkc5+SjWHr1y+co1z+kNOkg09uS1C+OVd
rwgLsRE8wF/Uu1JeCfMSKkA9oZNX++ShNjWeM0OxlMMeto7T6MRc/aYAuZbNweiB4M77pjgZYQ+u
hj0ggZyR62Skvu7iTDqR85xCbhwT0r5/yddnkVKOArb3xevbwYGMYEJYYcu7feV/70ejqLp4LCyh
i9h5yPPMVjH84aNmnNL9d/h76CGTlrlQc9zknUp6kUCqPsEUTZ+GpfIyFiBt6RvBvgaI1YaG7PhZ
xiGvEH5SKRFM6thueWXcFAR1/4XK1GAYub/L5PX7mOMnRWn5T1dQtx4yexq+NmrTz1Qpkrdsajd0
Jfraf71gzVgBDtfjBBkHaroX0ySzBrnCjmtIkJVlrBtBcpqG7gKJVkPAkshqDJJgV7bhsd3LrF+e
mTeA2Z/2VMhLf98rEG+GdjouchXRB89VDnqWpCA10AmET/pg8aA1xoTWnYHATgmk3bLR7CE/YOQp
yYfKIHQDlZkAgirpSw93VJs25BRItFhoinBv0ViO3n8BVx4N77JP8ndi3mfkEwChjWAkwWwzruGg
jdMsxBvzZrrkPpT/5uw4gBpBCunPcV7EqGyYCVJu3Erq+Vu3vEy73Sb93rlSHZ0N4k87S4Eutitl
ORCemSdCgwCxGeJcbLonRj768RPv5K7+QftS28Bo1Woogv9D7j9hPoO/AkgbvcsREMAZK6rpL+mb
RWfo/NrVoun+SAa3mnUXltMY5moC2HVSLXE5fzxO+bFHv4HI7fRTJcFQr8drQsIPcvPTCuCYipZd
m56pvWj992toMnxbhA2X4KTwpg1KjZSFv/V5tmNfb/mWljVgNl4sdNNZWwC4OvaHqf/yadpmZsgF
UWEuFJ8IlxOydMW74FiQiytgIC6yS+pHQjKY1mDB2/dk53COn9GKBbxfQ0/BbQJ3EwNu6mqb/Cko
s7wL3tFqetGsDGafKaHR3RMZCTM2y+Zzxn8Hf/TiI3SkptmqeI5Af041Rqi7z5fA3w8YHgQqf/l0
w/zXOzyd6GM/bAgKrA2nVA6l7Og+Q+f0F6u7zsRxxGSEf8MAgjYwDOG8K4a04kzFw9EkDKqty4MN
yjOK2covaW39eNWc92vPPMUI9nhl10YTNd84lu8aAYHYr3eI0mRvUZFWA1OP7XJStXn0MTEXGbwZ
tL1OMpQbXx1bVGqihAkkcaTsXq6YnhbqH5ykrR9nTjC+L4xhp6w60ZATqoS6iKkLIALC3UujWv9v
5BI+JTsktuFBfBdJEG3qsqkoijkPyJ/T+rsERd8qC/6GmhPKN+mi3nDaPJ9CUCQFWIcXXhjGrma/
Vcs47p/8Ne2HME/1omMM/xzW0IzeIDv3wKGWyPxwuNf3zCZKWV6U5qPV42BK8J/iwf25GrshT8EB
BZEHM2H3lnkG1HCFbmkMF+ToHyIJ1N8s9gIe8diPuaBaAly9wJWJkn5qCT3VYvdGVr0QbaSPIKZr
ingDPFKNZGSsD+LGSRTjS2X/bG8vxXtk2W++aBPFoU3OioRQMTR4MHbNWKL4MJvpgRdk+nh3PKQT
JSTcBOMJ6+OIk9w2xjv75eKTpgut9g8iV5LJ0r6klT/YhICAODrUW8xFoIAx+HoFlf+Us48uHkji
0Qjrdu8PsCCTCiNIix1W7Idcf4vcFdWOLk7e7raJh2R2kHqrrTe+7fqUYmCzyqQB0nvvmCWS1NEL
pH0VgHpmHpCUsd8BxeCtOCNsJk2Fh+IsgD1fRaV6tITfnZ//Dk5VKn7T5k3AGcilTJubwWvk8jIU
NWYHw0AlAvuaEfI8FtCqJmeeKHrhwTZaTecwLdvKs107eXYNgo5oaX6Nij67wpx8bCflJ0B5q1Js
qJ8xtWAjoF73EmizmIKEdij/+y97qmE1SMZwsHxhJZ5VGBCP5N6M/8VIkgXx004Bp4aWOiZy+Pjp
9mHFF/1ezzQuyLCXFQBxZiaKyHPziystChtxTgyv7NHrsGxaTaePGs03vFv7h0187cpxbJpFVzhi
+Pmg2pI+DwiP0uMsTcu+q5dQEqPm6cHh9i2TelpTWNLwtXuPDAEcJIsLecxL8o/dMr1Xp7tcFnqK
mSUaUk6LiGJyMWNH8+LH2t3wvCMg3XVoU5sJTzxlMg1Gj3sQOU4N7ZI2j17pSLBzWeQDiAQHEQRQ
jwyzmxoQ9Nm7ZBqJJ8dQLkhoiwWvj9GFKwf6YNUZ1AleNOBpHnjZcKBZKaE67ucKF+jHUZRAGdSI
8pknqhMDybhCLgy8m49YBgMcNkd8MH6UG51wj7hi3i9gw5rbNHMoGcHnGaYuVLpxZHMAx5UStEXp
kskHRFAKBfikLpPwWGxdjPa7bdDxytAqmz2/d7nW9mx6aECv0YFBD5xNALIfliAfGeso8r+ZzwBX
rvpO4HE7qutzJFViE8/VrTwzCUa4/0eXV1pS4qleLw26KB/Mf1AXUq0bQpnZID4jmjS7CM0pGOR0
pw9JPEoNrmCdBSF+01RezqCExuoPZzhEPKrUauOkbo3xiFbIJ9dYDhGgFsbh6bC11d/YjRiI7kgT
Dg5MAgLTPvwUMugvaYCU5SfW2Am3uEPZ1ZPCudsQ1H6iEQOrdf3jmfFyFEftq1g+cZJ8DbifDJtu
y1QnKT7ljQL303/IpXxlXJ3JJLGtjGZCMxaSX97FQ9Op4J/NBqnOwM0aN3wLWtN1vlFeRL0rBWOx
oM+/r3vWj6dF5nU7o+jVQkwDZ+8MLq5bNj1St9r4qR4CNtvM5GFZdBX0B8wAAsbqBA8shBxhM0dL
fKOzHUqLOGkbumL8hSPhd4istu0k/nBFTsozcqOoeSQGHpc+mroCSsUad4RMC4jzYVbFjnta4gfE
/C470e5Rt63HO30u//nSnk2MhoDv8iPbthfZogcSleV44qbyb0sMhkrevk4cupqoQ+EkCY26wEPy
x62oHrX0YjPWNFbH6Zw10+Y0y11DQ5fU+oCF/nm2YvOXusKXPfOns6fbrjWcWCtNEfcwiFwaWbyH
8EBD9+ISUaO5S3fC/ZBAOv8CF8I7RJpInH7VjxSERjBogcUkS+TF8EkmRygNiGXV09+WeIFBU9PZ
82Vv6Jg8AhHOWVszBQddprgRx5Qng59Uvv4UV0gMy2kGOrfPbozgivVXoml4gQ+ILYWwATJRhwKp
SSVL96x3yWbAp7enXNA79v0tzPyL+aaBg0mQHzuEhJG1zoOMlAZ0g0j+fYLHEYrrOyjrICkhLkHJ
3mkNz7R2v7CIZ9KUbXlmUcALRF/uKtFz/CMOKTSMVKOkjkpHc43fJcxqowKIqPeDcje0DvOowN1K
Po3t6BVG+UCPKDZk8B5SYyc3Rogb6TzLtWg1H3mu/+wk2gtWEDT3DicG8U2BMjmtY8HlytHWqB3p
xxCsUEOD+kzHP12tHof4l2patIfJItEwPOT1GWsP4Ro84RL/AX8IJra75rcYDHhMpzg2uZoYFnwH
WYgbCiZ7ybXswmwHGb41Bn8pkaT6bRubiqsvllIAsc92+hHfV5uMUyCcZ2a+9ierfMoNcpvGKks3
+GeQ/7EUWeryUtA0wbJSXKhAAyl3KFhgI5S2hJ41qQP8hXl9KzGicr66eSn6wvwMl56fSLVq1U0o
EcT28lySCThYgOpV28LTMjDfto0w82632nRoK1WVtxfFtca19vDTUd6JA8befWVo2JpP/zFwvCkj
C1tJsiEgUEuznz93O1p1K13yo6sBiokmkKVioV9sNgzIkj3UGM6VWWBmPpoQrdg+L3XB2WduFnEw
9MFxxJC9wZ50mjSGSxWJGrCe1nfR2hKT7WJp46hBJNdcB5f3E+mla+f5MRM8EOv+j2BCe2e3bPCr
h5ity28uH7oBZIKxB9L8ddmb/7q7BP5wj2NjdyLiDdY26LIzpSf6Z8YEvBEJIl+PoD2gtgTkLZ5u
vpqS4l5+tlDQYw2fvIQH00zfiqPxGO6Y1UKSC67qe4TI99GaovgGYYgk2sQE/ReRP+J2o4RPqqny
lAfG63PaFZXaJWrFJnwXSrBU5hNGBI8zTD4zvX+IZUAEWfTDSz2YKsmzu3r7Igm+kc8oKxGFqDNU
CGz5UaAK8l9HJB3OGkJAV8z9fenU7ah1r7r+rUTJ0Xruf6M36U8kRzR+HR+vWK8K4oh/wJ+gzzUd
+95RtYANSXtUF1HzUwTEVw7Sze59u5wVIKUOG4HJQjHfgtQWY4Xqu6q0DgVxxgkRnIRzU2Sro43d
A98ixMG90dz1/qDlKntWa9CZjSKBFcZjj8hRh+5faXllUbO1b6+0YnmxAOCJov/IPOgRkmJyRmXR
WnMUSPeWFVEYbNF3+4CJ8wPwUSa1CnGGERABs1hZ71hvD3Qn0inni7Mo0AI6QmWLOCk7QLSq1wvw
r8H7PG1/Qod96uEYvipHGeKINP6Zpo81N0k344+N1HD4bwK9M27elahw7K58/J5tAEIvm2gxgrGR
gT0x6MoUl6C7eJXpt2us0QYrYdD8rPprGvPZYNLa7LPkQf88p+GYfVyS4qKGnLRXj/pEf/6T1Axx
yY7wGpkMf+sSt1qssByiEVmDIbXefyRnOu0ypw/U2NYn+tFEjsTz6VNtBuxETDmWxqBfbITDqqTm
SqNwZb3MftnY39uU1ynKybCQKUhtw1ziF2uhdo1iiRIv7eiF6njMa7lr26ym86PRdUOesBq71rMe
+5y7bufJrkYgANrvouXoRVXPAyKPL7N2ZB8DDx/vcVkSHFN7qbh/JCSTcwaUreSFSg4XasHCGay0
Vzd3O7qUP9WilqR7folZ3BeE/hpjB7KRWxjubSb5/1i93lkUlhT6Fcku01Bcq9rV5vHvUx62zGMT
k2ZSWc1J4xj4anUBso6/FCXvL4smQRg4VQYZRqVU55D37b6EYTJUWSLSj4AfCzU26AY6KE86g/80
XjKfp3qejvgqENIqrGBHA/OL1pQSIQgOSt5dXIiWMyUkaUOnJQRNAgXBNETrcX+DGy8YXq4+hfdk
dqWUk/E8/6+p+Y9CGGZMkqx0h7F7vBPvnS8FE3tp9iOvf+HRNkQ2for31O/iRM8sTDTrvVW83DhE
Ji05RK8ZaGW2KVWQm7q1xUs4EQ8bP75FK9gYMAb7+uxQ7g3pPsEtEd+SXYvQ9jNxhKaWZfiJ6zSV
gfsrV7OvC5+7Dgr8M2Z910oRp2bQoB+IpPiPcvbZwf1xHiEuK+dTR6I6zv7FB99z+fUvDn2Oi+W+
8fs3O17p6GqhtF4PR81t9D3XImm3bmr0/VbeXpSAyyRC2c/1gyy/dM7QQ0V2VwRD9/llxlRPt5f7
/9MtLUPOMrkcRZTOixV4tauiPvI/SYbnPOPYC7LYIeMYmQWp+wqg97JeoqvWENLITDiKFsBUdXWN
hAYnft1ohYg0TBqSfI21e6acrc2/MlnDE4PjZTCTisXey6AVtAsvYfmflChABDSfvtf6sWZb18la
wjGk00o9r1r9mzI+ed4nt2a/ANPnGaXI8JlKOO63mU2HL9RtEsV1vsMRWPOfg8avCraMVn3rMKyZ
YHozhTgZEUovrdFlL/wmkwczB6LIweLJodUS6OQmX+So7Bj8ao6vkY3PYkPieW4Sr59Ka9+SApPk
6CerdjEVM76GMG8suu6rBLol/Gkt4bFKe9odIckKFfx3SEQDqfZrEiQIqzxDwfNUFtd5cpTlUbot
Cb3JW6drOtVKeVHUcTs2/RGRDRcFwfqa0PLKZIsZ1377lt/OnMBLKyvO6YBRx6XGeUIO78+4Y5kX
maqZhBs68oYxQQkxmayKtBhV9DYxrF6u7xyjSdNqngulYtP7C77QFe22QWfsRVocDO7faTF18Wjr
xfROlAFmjxufbgbGr/8LgdvZGFmGGe/r6zhWezCe51a/fna5Di1pLOjZG1EKQdekeACd19N5tTbj
Nnsh2dhYMV8f1f+rNeIgq0Gxdo4NT3ibnzbBJarBlAjU5yNvUEe0MbO2q7sJF6PRL6+pWLXaaUjI
EdA0p/g/VyUE47B9I+rEEUkMb3iM6ES55J/eb/GCvlMxzVZlSuyZSib65k7QjI1noxKxXFB/zrER
FRgZ+5tbeEiNys9fppUp/r27C51BfgyVqgoYwKjigwmQBN/Ipz63aiPjjpUeD7Jg0YN4PAFt1P62
1j6+Af+VXyU77YW47TrYGjod2VnJLeqqARAgxNMjieYvqVov7G5ncha2ty01E503QOI22bV5nq/1
p1Gpqc8yyurXj6glaCm+7d5x4NSvW+LASdUT5JzZt/sAnq1ZaCZmdFI1CEc/JJx4NKy2LIVOakEH
uy4g9OGLx0jY2BjJ5ghNcWXbzbzHMS1dXUx6kM0D0zTw3EtbEhWj9SAdrZYkDjw3yFaIx/tZKLMJ
f8XBdzWXyyK8N9hICEZLVeipxGlLcy3JVmA30ERTpPhZLoBW5IlXitHo9BjTyiWnIm6471B/4dau
WLBRgPQgWnW2647lw8GS/b6d7CHo0m7uFhYOmTmChQtebpB3EMJ6u6aXYzY9n/dBRV8xnPwBlrgf
1iWUU2KtkJkc0PkixeDqgNlixSq0s45nJiQfSERt2+dWqagIpzsTeh/g7zisxLIV8j5fVwzH/ioA
4i63+wc9B/faFKc28BCMJ6FbU3Dn4oq6Eyo9OOkWMgnb16iHgyOYgnjrr7hkoK+ygvEqrCFj81A8
/l58t5Wy5rONQ2fHDCXjzL+pE8lMwnykYzyp5IvslH+4X++PV0kUIeAE9Cp7cJm01MhAtI8Ei6bt
sjgoqQFWAz/zHYpl65cZZImbteWQ6w4M97OkRjcdzyoSod7vnMf5RQIaHWHO4RQJlefD++G/ZwKl
zLplOdWgaJKvj+loHOMuqQ+0pjLk9kAGD7JONa75GZZt82w2hIVDJPy3Mu8YPBdD1WRQt7lELjNN
cPR+WM3JxerUPnF5M3eYSN9LXcqEzCTnz0ngHobVAZVe89gH4TzQ8qU6DQ7CcgoLaB9fqKDYyv3Z
Fu4PBYfdOZajitPXbEqufRz7aLhP29lAei/DNGWhA3NopShI/EhHYvK79at0N3SxZOa76WMRwXbU
PsEv1itoXU7PACopWCXDfA+lp6orhwhGXzsg6zElOc1qvvKzRvVfcEPh4dCRiEX5zi3jB2yBMfi5
QWXCUGAZ+auggCwVtry354CL0yytmyr1xxf3Lch2Y5fya6+AmS5IB9oa55k8ez4r0JB6aHTcwLj3
7hF9nxiZMceZNHKmjUe81avZOaaBuN9tkSi/uGkMRBPXHGK4dTU9Sb7LzOdUjxTn6dh6NtNg7dNB
X4Ivrxr5jGM3ryUlHm4k7u83/XHbf0Dd2s6F3aodrrILfIix67AC8d5XbsI59BXUFx0TvSowVDLf
ARc8bGkisZG9b0UOQSx4mR5jkFSWNs/NIchZ4ipOhxfoukh6AW+gUJoP8ZNalM18eXzEp4LAMcK4
eaRxuFLZgfv4EpdtMKPzNCQhzn6WenNTXrhc0rywngawDjm6Dy1ZzhfMk4sHYZgoT7B4Mz+qySL0
zzyQ81H5xYMQea9rSYs6qsRnYzf6lwYgzREDh0WP2LFHuEt5JH2wFnGrFxUCQeI8ul1ryOHxCxjX
LX15brdLSZPf0B9bjtrreqMIt/p6USmJTW21+RR0QLPFZ2pgPqm0mty+xi+Hc25A06yNNC87j10k
iSL0+Hsca/B4JxquFU7Pqded/FIPesEkjUMgXG6CYoutxHPD4WcL/WpX9lSD/9qI5lIiipIiq+LH
vpwudPcM6Flz+QiHd+oBANPBPCbC5HX8DIRZm/KlufY5dnUcpOO3+A8aFB8FccQNDxuzPzbE5FLI
Djzg+6VvdrsK3AA4G9l3obdalruwWgZcAr58kScvJ9Y+eIoWJgx15crx9jgclKjE3kUqcXAb02t5
tS2QOhmfzGVcIT2wGKI3psIftLy3Ko3yMZpimuuXNfk1BW/1QGPtSbfGvlXGmLl42IQjjV0srfUH
yiqMS26nqmtHkwChJHjnyO3xJ2nWSuhU6L+bmbBt/ltDYTBYHzrmVggp0OiJCbT7RmjNPaLUfSls
vOJ7qg6z8e8PBRvvjo+XUkrcNFfhTEuE5xiT86km7KMxfICnqk5vCi6v95KBCEBHSHgWkiF6TXBG
f6klTb29nQ8t1zpvXY5XydMLgLRomkpsMOMzGBRHS2dMRGV2wbfQj2icTavqNW5bSoZC6K9mFxOn
OsQ+xqvVDUpXfj9jvyG8CwHIuht6NyGkkeeGFGpPYm91RBaKmW7/V8xNuEaUI/00DuuuMw24kfpl
76eS3ISL6KUqqOqj8k5QLH3Y1YBnTnd8EPgd8RXCwinG5E+7ArEHtJvuiLSyAk5STNE+s6V39ye0
uFpmVTKZOBqFmMvR9E1GW9PR41gjLHfD6yconA2Zzm1ivSsIyKuEYRYEMScuX/AZVvtfREdv2azB
iQEyQ7FTRpk06uzVQD+IpKGw9GRhQLzRdPX2+XokI/9EeXnQl2Y5+r7Kac++l+F3VVkLahdcwoF/
czLH1QCoelxbG7MmMjYUnox6NbKan7223+4WH/3gJAAx8EZovCZPY5J48alnjm41hBiY6ffg0omv
vGz0uh3IhCtknjXt7ohvmoevKA4WDReijHefSVSim1zKkplYAkxK7jzVg/yr3KW1PqkSI4cDlBKk
4Ub27paSJ+rjub71XaJN6cqsehn+3vimmoHzQiJs+e6B3+oQcH1eE6tyjGuv93rt+3fviNOw4Wud
kRyZAwg7Aj+HQAgbkt1vSQSUj5Y9/CirMXEwBWB5vM2oqX6Zo+t2pOT58hfx+t5fTYigB8pgoKZV
SX+CaVo66BtYUhQPKwXkoTvXJCX4ovlrVZ7ffEw+U2ZRv26h5qXe/pm8gHmbaHfUMTS0YdnH9xyF
KXB3Yw/E11huAHeU0k0SfKb1q9XdCTnWymibBR7rQtG89K+lHJwGMEAhmMgGP/LvXFrn0DAVC+sz
VbTTg0egpPIPxEQ1zUO6lClOdkom/MA3u1Bh5ys3IdfLCxz9g80N0fmEYS/tp3znz1PE1HBT7sPZ
xaOARaP4uEiBU5JkLIQDKsiuvz9jNg2AeTb3nYeG483aJmIIhGoEDDJ2vVHk6mBo3NSre4OCj4f7
hy27WMNZY31uP5MDEsYs6lzwefWiSdcaFQSEcc2s5+zJqZO5rOVs2Gb1fMAhix0BEMTQydb8gKrf
+tBrbEthGZNhKplED5IskvRntEdDWFir70hKLrZ8LdLzByLNHMIIbUmG7I4Vpy2ZyZHYoY5FMHO1
ACQAu+79UOBGw89fM5x87cSmknZPAIkGe9z97TXQB6NbmWwqFrDty638p+mNM9DC+/6MT8oaZMlV
MUxCWeVDijF40FNgwBQVXneHQFb52GVILSrHnhvv3J/XQDJNjWf2vQdXx8fGrbK/0GFFr60O9wsG
t4lwjEzrhyO/2CC6jBush2LpwKsQ7wD7zssStjL7l9Aj45PLTm9e9V3VRJbSQcInYnFNGRsjiqhj
RT0FuujnzpeGRHndWJZPZM7YOGS8bnB2FTahDvlsGtqPf9KOz0Iwyr0N03HDUtQ1Y6kqSSEaM2hn
7R+/CCe2P0Ed36ftxfVf6um+tx2NTZpvhwm0fBCEJSa13Mik6NR9AZxuulCWE38j0ktfn2ZRGHcH
h8glNjuFoBpdpMQwFDgI9QrCiobcVKAOPNuelYL7JLflrf7AxwB/RmTlxAEw6VGEOTpwQA1KeUTf
jKh86yCwRpv5b1C+k7w4qPMuMAlZHa5jMryZEGoILzLzJzkwMDXhGTrbqIaqgHuhR7J8beeo7tRr
3zeW9HcJJPbh71zlEh7KbBqQ7lNIpycQKI7UQRLeMqzdSM08SZXew9FKfcz6s13e6xZhSv3ScMdk
Eb8EqHzYVVrdZEx9lhU+XSpE14KDE9EdjWxkN7Fdhyia20m7wtd22gcmnhPbLx54XdOaDQDE+f3h
ejBFl78zl7mUxl4ggLPooQbxrfRU8tLgNc/d4gCgYQSkq5PM+rX/+lYz0Ix49CUdL9jqfa5CSymw
KaQI+V5ppfkXi5F6cFxqlY2/On2qs1m1nGzuhU/QcHOk5qaCzWWm6+NstZEDGcTBTrabqZBoBKXz
HRDzFNK1WsLTb40OLVuSPjj20W5WAS54rRlzlXAktVhkjh/sLJPlW+bsWdmRm+hpPqOYbpRASBle
kYfTpfsBaShz6yIoABaZ8QTTx3LOtpdrTkuAU9IDC9emLMZp14VtN+aoO1EPSbnWpKNZR87MqI8P
92WlkN8xzAdzNDKJl7aaq0nCSkwt5nlKF28wBThH/P4JI8sAmO7sWd5vZhPdr3HTYx5EQ5EfLWYO
Fgs7k06Ju2YJNOwrqc8CISQ9vkPGe3BQgjkvwdF2ped4n0kpZx6YWdS3nSkKDMKDk4/lxm5DQ9Wj
f62UAm603CiLU5CnMp7RgrEHa06d4b3Z3HlvE1NUT9lGnz89eihbsWKU0/mhHuhA3eRaflZhCbMH
6x6Q0BlPQhvunof4cXM+Lbp+ou6RsFfjJCpk58UKcJalqRCobpcMZOdwefuhBfBw3e1eHA0WsH15
ShwyQ4kFx3Vm7SOyxQ7xgnj1T+ZAFt9brQii4m7CT93gqGe18hWN/FrRa97r+8DilIPTtVvxS7Sb
oGlVxq80GZ1s8838ynuwYwLEX2HzJ0pcOyEuywdwJ5G5GojyozoMoIor8UX6Rmh+L2OIgtbahoeB
imuFUCgiIAzhkigACmYgIMwKIdH/3TK/83hBrgNIOFWLPXEJRPLQjp7x3fL7fCC69j4scFvhLhT0
G27ZKT5vwt0eBN9AMgXu/rXGCSvLzbV5BCYhRIrstZ0F7k5944vUpIwC5UPsRQ+3w13hBsTK5PJ4
V22ClI///A5rBT3l7w61dIHhqWYYuxP51tgywdQcaCR3kQGK6ayOGuhjSKgtcS/TzNRbNqwQ6k60
x4Nq6TyKvZbHVlLBL49TimFHS9VlUAjpcm73e9PagHgIrS4o4ScEsZC45sgaIgQJPdUii4YNGwzh
FiBlXuIuMTrR/YYHFrftV52cgTR8xzxzTjzt8VSmTJamfAN4R0TKPRl+zfIBgqzQxGZASlpYg5m2
Yb6SJpmXexiCDWY+mGGjycTLP3xD+3xFEOyQKb+NNybhazxPk1lLuGMgS1zwOfCuBllu8iJkCH31
wF17VyLXRGtDA+fFT8lvvrVOIB7UnkIoMhwHAhyheEFO+ik2ODM0oF2IVN3xhnvgJOd/s3cfnyby
Msq6kvIFh8ESqM5JfWCEVtUlH5vdW3901qIS4niEPqrhGLexJMn95yrSeekvAkKs1+GLGAZQyzm0
aPqyNng3TYZZjYQe0NICxW4ZYv2PJCzdAU7Xb90PfiOr0Gerrme0jt4fMb0u5oCg5ZStRccQ+GFD
AxUxVbn5ttoBOFe2OFLgqu63uVDBqZ1vy9yB0FQvU6WyAaVYkQixb3lDV9YXL+Ms/BvI9Nk7vmiS
kEvDFYCJsJosKDyiD6h2DNW1NMa20+g0J7pZ3+7n4KtLJG2hN2viwTb1PQEabDShJ7MAUMjkgNp9
Mk/raGqLj3bbsiCwEHHqowmWpP0C8P12XYTLQxBduhft+26d3eF3tuqbyE18orvXq8CB9931J3NK
0M+AKOEGujIMJE3+gSqSffLrOACWauopNEG05nWuLc4F20nY3xsaxDNFknWFiyhhoQdixL06dR3q
3AfVpLwpI5HTtCIAizC0qVj4/jBb9wLwL3pbqmkTSH0ME2J9pIQpbVWo5/vnaVjUVm1rdZQVDkgP
gcxs9kOcqkX9K6miKJh8F4rxamcQDC5XiYSH1GM6MQGQ6+Cl+vSfe5/eTBY/LqcKASEDmKs/md8c
eW+dDUGPyUvtLWnFw07r0QVAr07N2Blx5h+2nnG2T6frsx7LiEcuT51OzAzcI8qzCEsbz4gMh0hD
8RGhR0V6p3cqU1BzCadYuD0iasaCl9p0uqfe7rHlHMnShMGZnqaEypmai0XrGS8RERUDKy59GNd7
LF4h9OSG+6cmEFJjf/VBfFCCQ0CuuvbWTCu24UOyZTZMCGNuLPiFkwuQhJtan1iVOacWfONPxogs
eenJSwuw2Lq11QSYg2j1NWvtL/gvO4i2oZXyo4j4lXkAlpYygnDVe3hBnldjp00ZNFMJV1/pHxiB
WPskCGAU9dyL37GpiG+HMy0ttAt7hD4vdwzAmwHskGOtiUp9pJ51fu57Sq6BCNaQlpEyvUC+j180
p4NZlYxRglfu30S8UQiRyebMTwmsbIEL7pBFOxFkOxIS6mQjeMMu4vc5SMzJyc4PjMVdHvmvCM3P
MSuHhQCtOnTKsP4kFbMduLgKWeORXI/RvIhCMLI9NE0zf2+2OmZuNEYPdTL3W4mxQrnwbgSZ/Cd7
LwDOj3hJ94n+jp67dCx0KpqmHfejS9J2Cpvw+gdyiel67T9pKBX3nZzkU2b5YTWzBwh5KqFmzFss
QTKm+fKZTr83jPgHcumUiz+aizhevHDVGYPQaydZ+UPhBTI+oyRsd0vlrN0J2hyUUd7rWIQ+wy6F
uSZB7vNSbN06DWzd7zUNZFiDY2xDtzpKi8FDMJ24Lfdqzgw4VpZ9pFOlGx1ZBB97W3jDm7uUcJXK
RMnB0f4CiV2YWpkfgLTXIsor/A25TlY9dSNsd/W9AmRwoK9Q7LXKSOYxgaBx8PUmEdBWW13XBL5B
gGkXC0TjtxYoSbbigU9kzrF8ROTTW6fePkp0Ykxwl2/rFMysTDhP293XamGXVQxVijqqyOO656rf
kmTZtydB7RwgWqu6JcfUC9nrO1Whq9dfNn3Hoe5nizi7QWGMRLU+Prwzc9EYMjzQmxae9jf2//mB
kCnTwJRTSE0F6lcYvplxd3FA3jnTPX5lDVa/UdRHG0Sck+J0XBkbVwxpiuXQ30dR9xI3T+73apko
cHQ4j3wKBAmlqicgr8nww9r+Cl12EttIikdQ3QRR+IchgQc8ZX6rh1Pk53pKC6TAI87doqhFFzq5
uj0zkz4au0PuR/rcvcRK5LC/QeYTncqs96U/OOaO6w43NEquZK81b/MPUksCgzIdt/1btT6biaqr
HrMKavsuJO0cCnLuaXPntds4rYPKjQfr9Uto4UuD+0HxplCOgqxQChBvjjMZWgxgJnkE5HfvbF/P
BBfZlhH0NJQ9/eDvsKpTq5RFttlzopu6MpUvrnwYHvIe7OJmE76nDtdUPyhlR/zxiqqYN/YXj1/y
YDssX/yfFdwip7h07USWJ1vL36Kzkjhvt75+1oNoZe8xXZgX6i71JlD3CPQZLuWeD1iOkrQGfii7
I4q2py9/nvROqPRe5prXAFV47Nk5txXTjDsSRn+RsF9E6M5QTvz8SHNgyO0TnRUgy2xhk7t9cksK
MN4ajvJ46f7lNHJXKsoEjv2eQEPp+4zXwUXCgT6AD2vqsbzYS1qA9UwMH4zJ6kdulDid2NU5c2FW
+QjCwoCJAfKugqw0rTLHCg57hsZNpvI10BRL5vjishesk50jFnKSdW1q94bDhv/Vdz6SxsTkN4Sf
Kg6lpNeDsSEW0hsNWzU/LUkHru9dv3IEpfoWJ2Q46gQJM2gokTeyFR7XSEggd5JNtu1zK8/Vik8y
kiuXxN09Kpab6/54tLYIZtVl0dENq4W2O8uyLXGYIG6MZ2zhO0wZ7596LmbsgsGdzi8g55Rl0N+i
TlePo3yNpaEIRIkQpUOLmNs6pzaXSWNI8+Q3uT/9jRCihCcXko1tgYFo2lYbUgW+pRLoGGLfMwb0
ohgOTFZp8Bh/cAMWb1CPWZvyAmY91k3/5eyNw0PN3/eKJsi+NZZDChRXd4kc4YRtRkPTnuzTV29l
CvlfkoP4Rf2EZ+8+cH7iadsnEcKdClk/M0Kl6HkywwXqPjPsJbkuuN5VQ6vm2OVzk6Tt6kDwNQfm
r591F3sO0tfOYZDjSA3/W8oa67NCL5WXOqcHPZKNhSBcmX/4lzsxu1Uva14NKXrrpBog4E6Xj8hV
0zCuJxXOg4J7b1Rg626F/98/rioPNB38KS3PFFC/tmpCw1WOtbjstTXXjPQ76MLjPmrlGmlPkzeD
wi+Ig2lISOlpoPYDb0uZ4qySnr2qXDBCjFh5hjlPeQWZncJfyaYhfaIFFd8pXo4lWufKBd5CwUO5
jg2lhhi1Osz80pYVOOBsodb+WEAav4UsjLEOR8HGYvixPFoBfwjvCeZj2DGcWEW/sR/CHspHTaUQ
p4UclApz+QOlaWqFUXG/n+/lPucBVI90vY4qoIaRitKADf+T4LMgoTLUkrFWPGLrE1XjyE42IADf
FFOw0wblFMYkkbsRb4Snr53FOYJoV5hcV8rKpWFOqiKf2KMHmSsyr8u2BYAi53Qep8eu7JzGyPnA
OKu6l/0aUL0OetWDjMk5065U/4MfW0yKyRrXFXFuoC76YMFb880rQvmoTtG2x81vaBLxTDd1JWFY
v1s7rqlJlVtOYwmN+m4QVmET31PZqp5YGWx4NSOLE7g8CGH6oP4RJ42FWYWC1kLPPeQHGZZP/4kW
7Iw756u8i7Io9YQYUkp7rsHFW4KZ50lZ1IAEdaEB8eJxEqivb5ZbZNib3qKHJJitYU4mzcLgSLoR
4JZppmnf5Nyk7Qv7V1NmldwkROArnslTNJ+/1RXP6mNWJr0Gc6gjaltN7HYLUAlvHbkIkeWViO4y
8ndV/0JBKGiNkuQqYBRVq3/m3FxwzFq79gj54EmsLaV7XoD1nhVRAypt3GVTvroTmdnoPXXG7yVe
Mn3uMICmHfG7ZteT7gcesYlHY9W+/ZUI9h3bz6E/+rsfj63GEgJru2tBed6roihu6BlSgT/8FnSi
K+AXTiBP0lB6F+JgDVvjMAkIoVoY6OjFgtba+fTkhY9Vpk6kExTU/lGK8GsOJH0VCJH7DoZSrJWv
dcoUtgoCQwT/5qhdUNv1Q/hSbq5AQyHm1HhhuLGNLCXXlSV0wlQO+xoEOGuto7x1apCbhy3n79k1
d0sIYDugfUa+tzQLtfJ5N11J0LRjFULwuU1bZbWprC7CIQEyH4muIFbXklbz2R6nbBDUb/E0di0i
wUUbccBa23lJDQ4QEVPpKQD0g2zQE56ktjBQDd3WUtZQ11+jRs9hE/1vWbc9ypZZcA747GqOQIdZ
sm+XKnkykXUQ+tT1wILfQRLkp6cUaFSfnctBcvAZkN54KY2AkqPGAZJJBQaG3YQU3d9AAcHuhcrA
bf+4PLMK/+CI8MZJl08qn4ek770vveUkrVOCa9F1vDuVHS++U6CFTvNxmkdp16UPJ3BLlc5sEgWl
EDyNqNPvxCqXEC7qwwFh/9Uwi4DcbAG73kacwi0xy9p/MhvJHXANkKabE4DkZ2zjTYncaQq74wU0
mH1dSl46gCdRI/0/vseAVEYs25Dvnsx2K97G7PqPMpdr5zMIYdDBN5kgRYQQ8GmcOeDTBUyZHPvi
GiWnx3EEPZv+KCNo700uRZExgKhGPlZRL3gOcKlC4+dYjadP5lygWdYX2lu0lhQZD0ey7jnMItov
RikbnJQyfc06dK8iGKckL7tApC9WfmWfJjD3eyHL9qXvaWs/tpzQVnLxKmc2WkXTvXOpRh0cUq4+
qgERNauibHgxjeRvKt4lgTO6tx6VjLSC7d3oaJqSs7e9TcDuzwQG2cYzYsINklqRLP7HiKq2klWB
44XSySM/jI98C29ERzoQg1PCX3ZLzZb7u5ZLbVaH74eGZxFpStxeCJyK8RhCWG8xIpLNpt7BIyXp
fnVqgUYJKpyDkC6l/EiZbHI3I1YiIMLo21ad2uK2CiKnEiwANn8ljDb6S0vk+CW8GmcgGIdYtrwy
5UKXxDXLZWDkGtDVTWUGhgKIqdMwezQVpJPYuSgkxhMeFeEdf0nrr/naIU5XkNyWk18DBoI5QB9g
AIUjK50GAigrwBknPPwg42PEbx8e9Zk2Tf9BwEM2RjR23cZgOTbPnu5BcrooNxwhm1onrftMqN6r
PeV4UDcLVzptUzW3AjfhntFSKKpQOm/iIpvG+QsAOg5Tu4rlnJIH/OJb33XKbsGQGsdNW78l2vbp
9YCGb2EEEtx3i0Vv5qNoUgwDPMgq2g/iGF5ozEBU8b1I1CuLJLvSWeeb1VuO4TknKSTRK3sJgDQV
IO+Y3GXkj87858OKp+VOSzLdm1eLY4c6cOoRavegz0R0p2pVG1np8dfJ8+Y6ox84W183GW0ZwzoK
FD/1Gw9QFxnk9kTlv7m7jB89t+AMH7HRihqbQmQmP7jDE7IaJZu9Iq4skh+h0JyMK3YNos8igSHH
Of3ZqACPCh8NzuYXnHG4D191JNdgVhsWsJTujQgjIe3sezZCflM5m6wogkdsjv+tdFTttr2jm5OU
2E7GRWThOljXKUnnkMwmMKzYgLw9A4mpniotQFZtspelu8glYgjAlzuylgGSw8+ty2f46J5bc9sU
6zAAsa3//YQaQFNIhspPA2woCNVMFwB/Y79Y3ZSbUq0AjaCQjczfWnYmE5PulvC3LlY4MfRmNMt5
eWyDplux++XukPRvfnheQHLv4oCYqBQ636Nw6PxMZzLsF7vQM37mv2MWTl9Vb62zmt8x6tfW1qel
wJrQx4/MHbdOh6/p8cA5C0bMSSoLz42oPOQ0t7WGKjSnB4qUq+e2a+/VUOqjUG79TTSEIqMML++8
kNn1QcRTcF/BaRNW7LtdN1J0vXb2yr8+Cga/FBZ2K4J9te440jsWzsvIQfGTXumCjpfyqyXdWVzR
D+3U6WoiChcyBk3YZ72/RdgyA6X95Fo9SBelEMRwsA6b8qPSw0gJppUSClUs8nHkS53P1QH+mRYI
c+HfF6X8p0nVTXRJCvv1RCGehhu8AJNUFFfWogSiYxEHXFMaBBmSdT26BzZ9FTn2bK3b6KnuKL1O
N4EkfeKyB8QJbQmUL+O1jJW05mPC62X+WiM1n1mTcfeKiaPWItEFaPIkR3iRcdsZnsgvKQCEtwfv
wvOHfHZt9JlikfTUM3i1B3qkX5T9QEGBIvS5cbLtmbdm6q2pIbG+ZbleV7yUQNfoB9Zt7b9lEwJE
+75T9XQH+HUsQT+nCFUVGQcbGuFoOW6x6C0poF6oKphU8IuJlFqX794F27Szazqf5n8OkHVNFF7N
oy54NGG7fIXXfKMHdks1VHmrpiV0KqyOGnj953OhfVqlh30IWJHToiX7aup3I9DZMzk7xADyCd0c
/xFjZS6MgoNqiyvsAQ8KLaro0lj/OaSEtFsjH4gb/zqfH/GbgNCOeKZ3CGb5R5sLr2Cpxr8K+Uw5
ZRnhlz9HU1TnjxLKRLITD+89+X3sdlik2bqAx/LynAyQwKUVemEs/02803S5reWl4q055+wi4NXY
rcgdDISZsodg1xY6BOcUNc+wDKB/ENTEp5Gz4vGBpOTAhWoQoLRXUcDV6L4zs1P0rU3zmFN2gLxC
iaJaVsT3wwtyaD4expaW7AHp+fClj8XPc1/7K6kZmDEFz/pYG7fzpD+R8DgDwv4PLGcOylLsVoiN
8tuZWAikjBXnoFKjJkrOUvxMjq/OtnCHJt5XAEByTxql76hE3eS4USQwAVC/QfkIjaXVv0PkS3aL
vGA9Lamhx8kN+1XzvVXdcBggXOtVfQApS/ImGL0+ycBHpixxlXcry8RM9UzbIn7/piUXkhZZhpUb
GQhovktpZZ8ABI7TqNqzwxFAcc76Y+8ZkoU2XGKW5w+bLQmfJVDbWDNgSk/pdnn2L4uTOX8ZwPOo
ib3m8C16COHN1TcQLU5O/q+5Gv6hI1QJXMN6G5NFM3snkPP6qmdbGIpDEF8s+o/LPoRoAg6Rc+4r
CA2X7Z9Bwk0q6s/MK0Vkp7t8E87DBFNQKzWRAaltwtv3OOz4Jgw8SizHzv6Qg1dR6jwC/vIYkcbQ
uI5jc2Y6e0R8pWjO6MABIWjfv6l90XWpEcnr2B4g+dzFhcMTXxElkD7izqwsh/+3HsJf2GhnCdcK
VPIgfYtLWIH69nbYL9nVcmLTHgMo3ygkhL7qES4dY6ON61f94m+h7wv9cORbAt2VDMRRZjMMo/Kk
G1hIhPXIMu4QzhAtjQPHD1RnH+de7EF+CYiUNM/XDv9cYJ9+DyyLX6EIdFlgTXhldWKNKnH4aaS5
+gkjYfuwhs7jZAnxuH+275Krhd3XuzkBVLgVoXlG4QlHQATUnoF/Y9CZCgY99vNkG4PzFcPJ5uR8
EBL1jQFsuRxve/PBe6but9YIPFuSnHYgLMH0MaO9OJmHrzCQofic4MKcBJTaJcAkNd7hL/vpa7DB
gefsCGu2HTr28X/vDx6EK/v4V2PA6VYCys/vEBvYfLWgPZCjs1SLbtb8jYZWzVvRgrS5LTPtFYJW
v6wdkjkdQpWWCX6J3cR9l9wBpbgc4cBzVBZGK7ZNVKEjtspNNHmjkWbuafscm8PXuzORY4QIhsnR
MvAvhbd9260x1vJEiEK4DLCE0SFdcaUAvAri+29OyOrLq59gJ4BnRgLcJv4+MtKGEH/NgtO+wijs
sh7rSQUyd5/NOfJvDcO3t9bcr0hqSkUA/LbCFbSL7H6updaHATGncxynRWpCxgTRHNrky4Bb+7ir
lma3UM/P4Y+9qU0jNjOeD5WtvORQX4NEqynpt6KmH9RFKyAIp0BuUfPHfR3jvvstCcAaPEw/VT5q
/g86Vt5OGz/iryWHJxubU2GC9PTq4/3t5qkPBcTnlp1tMvp0m9NNMOncNUn8Vce0gjJ1oq+A6cz3
4OJ4McxFfeI9+J7iCLRlA37bYGrFUihfNtBGG3bC3Ju8Hx8yP6iHeeOTrJ7hr+kAcd/SexAt9Smk
b166VB28yE+go5hLdTpmk5cdp38jbO1EBd+mqNC7UBacJ46j1Ba0VqYBKA6tNU5OE1n7SNeWTDKc
I8YAjWgSdOirASDz+wR+Sp/tZiBU1ltiWf18ad/PmwZmT6k2Zocb/fhjIo9OZuPC6PqmM4d/tGLV
70RD6GUEYIMOTEjBFBP/mi+Bai3PqXmEYqTiL8wFbPdMmI/Nm7kwK1TNeW7QJ14O16L9MY75wzKN
VvkyPNLQMTlvkvN+PAWuw9CLX+qwBvBwp3zL8MfAQd7D39H298y/ym5YB3Tng3z1anfeYik1W0kH
fVzxHB0d5KDYY3vbiiEWYUuVt0p9LMa89CUeIxTUvkAWXUH59RAKMNlu+1PZWGjWJmFMwPNHVF/X
hVSrfteK4ZGhPpimj54tPcrd98CSWmZkxM7VAdndUTqDYVxnr8DMxHEH1D0bfON8jTrMahVD2N4J
N1hT+vM3gwgq5UzvFuLL/1x4plzdEKaZlAPUXocYA39VX0Bx+CLXwuBbOweTvfLGZUWNV5SnMQhb
zfh9Y/UTEX3BaUUeWU245jAK0ys43koey7lWFC87bfNFd/r09h3jDDCFNl2nFHwlqwvyrQ1mSuyo
e5bdcokAXvyGzUMb2bu9IRJI03kisssSMEpU/EkqHpXGAHzbMW/QPAA0D2Te3UgQkUGUm+jhWrMR
slPR4peQxVO91nzBgUfhcTy/1UBlErM0TqgBpxNPvdxOFIYvQ1hUuwOPyWMN3Xz69C2BDqyukYTQ
6jhmfSCJwdzSe21QL8+4XJMVeb2FYUs3VHt7PHxTxSWDmFMjtHMwfJfU0I2svvQHapApbb/SL1fW
NaW8suCNHGz8ZpsOnG26Txx/NiYGArTS1WUAjQv6BQr/kqx4yDKlLnmnRdlUuKR7rG0RsOXH1l0Q
6XORU33TtA/Fq3MmKPEBooWR77knJjcJENMupsKEFfKuk99ez2lGi2JbGxR7gf81dWO1rGnmxjBK
B37QG7W2V9bQa2O3D44B/ohIIMd3pqaUVO+Cj1x/k5qaCABEeZb0FJiZz4m+UrrGi12nhTf0RJe+
jinWmk77gXv1RVZCibAl2A9fGT8clgFvlXrBdH71LyVT+3OCOjaobmPiXAGpSaYBLApoZlUUl9i4
2cM9SerfcSpnLugvBLT3E1qWeI00SXUzTnaDKIoz8+7VPdu7m2nL1c5s9hCKTdhUH8YBNAJkxNpr
kvlz0G3xNB2RGYAmxzn2b/ji0VWyxdrMpN2KZH4DHAGrZLcGLgNikkJ68gofyqg9g9VBp8t1dpKT
7+lfTyUzx9NZhL/hseJzC9TkHb2iydcyVI1TuN8MRLnYiVEWaObmGk9POciXwL2O1448/Znhqm9V
mmFd0DBhU2S/E/mbIG2VsHTkOy3UyVt8s9DUpBi0PagNnbD+2eWFZ1+7qBf+0ZZKnZJHlR+xErDw
zL1gVIaGHwBys7HkdDM/y8jwVcsxyPSs4CUegyfJ6QydKrzFySM0im8IaEHQgXLI6jZU8MS1xryi
K2C6icGypgFeL7601D/vN/IAAsM4NHjcux78lFS+h5wLngoDiqI+Wngy4nRziNs+obg3dA8TbfbP
IdV1PFRyzK9zxA8ACrQMj+CgPE4Vt18GEZbunHd5Q0NZeETpi/G4f/IaWBHxI6q2qao80sgfrqUR
lk+PRZdzj3LHKUwLjQGoJCVD1cy+9cy3GJ0bYL9jQiOC0aN9rMdmiQdWTPz4Nc9HKMmgrdNJfdzl
IRStmZjx/vviYFAaXUHnA+otTiOUKyDxXkD1kaYjnjCRZvx3G/Qu4Ml79xErpbFixN0pql8XjhaI
wkO2WjQ7yvJLmFLwb3TLYjwZgIpujLaQGz+IgBpquJcRqyvWrBzBt+rNaOn7Fe19nL8gedobf8mi
mDh/Oe3CWQyrwBLYJjHyyS4Im4xceN4jWx7Gti5jFNhz/Ff7PrKYCoVNl1/urrmsAVtjftZHB4iw
9INM6pDRdoUSoYeG2MDodXTVz+PB6o/DhpVAbU/0qR4FSAgUYOZa308+un1SEMmbMa3eFJe0Xzxc
VBWGnscSMhijpTuD4Zzx1X7RodaUoExv3KywApKoAs6zZ1Vs4bLlGG3Bvm1zHsFGIOpBVGFwRG7h
O1Cqw99m6nUAxbTSVkdwBpQJ00mmDT2KcYHQtq517Q1f4qtGI6JndGETh19BejFHjO5Yp50c8kyk
pmaktCVEa0nmv8hSiKYwhyQH/LHMdWTNzTh1iehLYvsqmPfTUXTouE2N/Wpq7UOLE7/rS3Il4zDf
oedkQG6TmHK0hVqZM9TYJ4LuwnZ7JtHw1qEVIMLT2gb18+HGhbyy9CYGHwYP5JbWZer5Czqc+jKf
47WbLI8A1JDnY2a815BYjmADH+yZb+Mz/d7gruCsuqrapSkqtb7jZtVuwhRrRnKNrNhDk4vfEp+f
k++QU34Jk5IIVnYDJOk8nTXLfCLT8cnrnvBAvT9hX1hP5iH3zER23Xpsd8oLe6aFSc4DB/D2VpSk
Av56aWOILATfqC5UjXsH9lBkSEPDaQh/fDmqLImYq/wk/HCxMnmsrHIbUwkqFfDl7NPVFkvV0ncH
iT1xyIa2by2LUMuHOpwpqu3C8l9BfJE13SeRC0CRS5YO0OfZ2if/8tZxKqgJbPYar1bf42I9hLQR
j93fNE2t+KD12wT1EpTN7gKo4tsL8DGgAlVlecpop/GRqYLrjtddN8N7vF7oBjcO1RJoePY2q9wi
2ci9M+HeQmmI33/2+jx1esk+m6xd/d1XevwQxCCu3BWm0K1ZQAaVTDNusdPtEdlEm9ENvXfcNAca
BQF1Sliudhyz8IewOidlegUTrYniVwejR4X8+v4aRih00K64lxNICgEilu41shb6QJB46rAS1lRq
4x+5A34F2ELmMRPlfjv7qZkviykbc6RfVPTSGBRxGmFb5jahqxijjTB7VtGK2bXm1COf2S+P5r7e
EByegP/oG1nGYuM3OwlZ2+XpIslOxHTM6WNVuMuHCr5mKRFRhNEgVeyjsp652Hx0U69mbnFMxlDH
PiZ9zMIVKZyHENombYuNn6+ssH5atHx9jHC75N82lTM30f4cLRvRNITjm5Pdhk4aaplRGJYL2WKe
3UUTtWkR1OzU8eA01t9Ur93iIOwST/N2JzB0RoFopcUkWGGCYg5Cp0tq5YWam3XBkuSuSoxClN5A
f8Y6Mmdi7XMMF300g4vIeXsQPrriOjLII7cYsBfE0yjkt49T0PyLJ5Rv8zDfDT1dJfpqygitmniY
LkjJTG+AF92LjE2EIZX8iV5k7v/ONX7xFWrwdUEVN0UZfm9f8FWD3TW65LrWy5sLJAaZvsx5RIih
NonsGCpPKVYyisVEw3OWxnPaxeD4PUavORfroklttNGvbQz2QJEpcVPyDEtVQXRxSv9SZ0ISmnYR
SzD6EC+Em1lErTGBHSOxhw7bLeWuSawRxcISTGnWweuQswg7cLeTeoFRZ2TTwwilqVFSCbSqAgVv
dmWgA85YU9FJfGZW2t3VHmIy1ezCzsY1v4ti2Cw8WRpQGXZcnd5FmyY0t362cPBf+Pj5BqNCIP1E
I29CBLHwAcrvVl3xj5VQ1M+LuSklhAwufiL3boLxckCfYlfNseW560g5NZWwZm//+OekGFsYK284
ydgXVwBRuwD5BfOEmARAiwsaO17c4YUS9C2y9N/nDxyjpdXF3BhW1LXYD1ANZkllDzP5eM/3gWqQ
xbyj23tIRj63nDe3Igv7wlysAnLNL1e64O3fi2mx6oR3teKm++m7RMpMcFH4CnYY0HZp619pTspp
Olq17CYGZ9My8ilT47rndUTlf5Wf9pW5MNpoWD2MS1XI10UZaicrdZ/fDQMvXJ0pdh9lI5AjD+a2
ueF0gHp2+g2lvSc9jjHFicsABsuRYFVyp5Q6/DaEscD0J7YAc3x8s21aGPJJYH/e33POHggkIv3K
mrLTI8AkxaVdDlpSDCf8okTYc2ehQBW469qJw3a942hWtS+HTNfgyawVvZOwtwUQ3K4AC1Q6QqOv
BdJtRsU/jcZqT7kHIt/I7G8CA7T7leef7+cDvvUPn14YEPCm4ZNXqFofo+JNCI0oT8jzj7ycw35i
MwFNQD9m5cA3LjUcIaX1I64RXzf1fsh8Ar4vm/CEucOGonXfTU+tB2e5531Hc1vaG+RsAPuSfSHl
uLl6IQoXKmIFX6bAqn0GSrXbNmvcEhBtI0RnZG29qpPdP07Z6Z5cwCAm4TazfQj+B1585Fq2AtJb
T60qxl8je/JZWWBImXBmhZvkN8FGaea7x1QiJ0CKXr9MfZiu1nVdVJlIgL0SiXrE8qPyd7kzCigY
xzI0vvojSBNhYj645xUgrmxG2Z4eWE9i7gQwpWulAl7ySM8e1qaajjrgF4/Xyfrz3e34x4aOhDxh
UUTPVmq6gIWZs5DFsugw3iLgUz1XG2v6U7WQjI7L68dlffdvbh9L7CoIDRKjIsczkHozpeTXRprt
+Ki8WPID4BwwhrdIAexvJ3l+bzOc0Co96Gbc1A1lhuVUf92zOmnIbxBEVmfHNq1qG9oFH2uyz9l9
ley+W6bA4VIVMurWV/li3QIiS8u0IcgVINWfma1+mLIe5YejDWSuiomaZaC6qL1K3OXrkW+lb5XH
/izEfOdptVsf0+q0A+dqNdAeLbWaWhjBbJ3Yf12lO06lw8vPZRUGK4mhTjDzYVwHNsUGrE1MOXRw
N97ClRAvsYv50rfYj7X7HXpoS43UAF5+GM/elPkoqz6G/0BczOiGvkJQoGn1GIS9FU8uLu4T7+Wt
Jj+M8cp5WlFzdzKWaV6SIf+AcjOqBBDe2odD3r/uK1NICqa/qHs6VdN5pQF8nW7hJKRTA0Ve4wKy
j22As202wZvoUBVVzyyLHvGJZT+H2gkjf9SZqmo8KhqEnWd2IXBdpS8M0cxZJzijYgFW5YJoD1te
VV1wvpeBwCwGyNh/o5OQ9jkhrPptHN9BmuWRTGzIpziXF/cf2mUfob21UbGbV5t38mqs/0oMpxmD
XWPsY4/w6ogBqqqjzIqDICQWzZaBGtltc0G2mFzIKwFJBkT7PHZg7tUDS+wHIZIgCKop8cUa6QQb
F8ISqQp+1SqRCip/YqLdgIQWVmBRQFzutCvG8MWxLSS/xv+7Gain+J/xNmrxUG7GDRdN6k7CSd15
uPug/w6EGYup23C8GYhjcyG6niYpC/uzK2B3XhJzSmI5tWNOD7/SRIUf4e/h8aTev2cJP4CL3PAK
9SKGULeQbUTShcyrLqmPZ3URJcKtGo/h2QMroqGwXY/q6zc0w38K5wieODsflvIjVxMwkf1yQVw5
w8sL14h21TMEcJkiewRJ9wv1rDDyOH2mJOlI6ABLkdswWCEUEM3HUO/Tb+cHaZMUDMmQLQFyspmE
/3n4lOyB9WO5J/wNALj266ZxTLJo6slmDbcx/n1Eza7XzGGWGYEBWTVaJcEpFI9964gERaD88Gzv
YSOJzKpBWP6aNrg5YWCQGbPlygEOAFT4OyBKTsIuHvtfqXCclJuM73khIeYewnaHTWJm5WYF+HpA
dONa0nomTonu86YcfhuJ+EQHMDRwoVp+iWw5SsvEKNmDK2+UYHZg7+GHeo+a76tOyWOf0zpNJ+00
e+P5w+87DRlT2p60lL3EZ1ZSyz+/bhkopDm8oc3pZfWIgN/6pC9AXAstEJspOmVq14hQdhv6bX3i
/wKOsMeCkoYn3B6O37qHqr/1BnEl5hE10wN9oMEoucUonicF5xShkkHEG9tu5Cjshv+OgAuZgLS8
5bFBr2kWE6Ze56Ar0k0gIfj82x5kQSMNpnSxt1y9Ab6yJtatCXsJF8nXDtXCziSaqJX4lYR6N61e
rkCKsXAmrCkrk3qpHxvD8vMoNtVFUJoa/V3fd9Br/gLS/OibbbCuwoZoiyL5U5OVDUBS9to9YXR/
3oCDP+Qy5hJ5Kof/BMmNXtu5iIQY7ycHIUsr38ks6uUji6PuQgyso1ND1WyQeDocmNuHwi7oyKP5
uMv2S0va/S+8kPQY3TkUzBDSGNN8q0sP5lC5/Q6AOY/YLuu0KAF3vtvx0ZRJeqJ7txpO4y/aVDNL
qrigYn4sCwfsSKxPbWZkA3NPBlZxfew2HxYRHrZiUoF4r8S0B8KzMWd7RjZWaqkURVFJwSRSqxLj
4bONcnHElsI4zvrcu2/Rw+XMgSm0CDN85w+Fg/8bb+2FHnyHhJvEt7UXHHJOqsYnmrFOAPMX1CDq
yrtB/l2JDEwbJxsOoulLxE8xo9Ww930pimzi7hjnMOn9nv48X3RUKl8aGfE8bS0kCkWJtc7csXfa
l8kbgM+lO6q7UbUOH9fs21GC0ZbHBpXcpr8EExUzvOanU+Cst8GRZHbeM4BRxbYAejQ4Byf5dGxg
y6xAbhmgz1cRd49wvbVakQqq5dXV7cVXvPiidJHu8lBN/xKFGxV78bBl2T8U8AKRiSK8lAaVFHu+
86MG2RoPM2V7NIC6BNGx2OVOjgr1iCXFBdGSzc++N0lZ3Slea6qOf5ocEcPEya2OX6UOqcambYMJ
732uo1dBLVaij3yYu5D9YOJA0vrj5XoPBY2AkPjNh6FJ9tyhE7KkeJNu8g9uHL2reO+5H0Q4jy1i
gUpN9NqRzeoV8dhBRVHHxlTl7+erNV5uApgELMk/yKUAqOh384Brx1YqffQl8lmqHFggU508Tw23
ujw4BZCOx2adEcxqFnAJOWgvMRbNfIlJjgx785+m3AknlXKHGIq69gy8h3/7No1CdxHF4snlr8hD
1HMN+JN0yi6PfR6SSTAmutuHvOH2FywxfG9VakDQPdtZ4LD1g9Zn+84j3yu/OY0T2M/vWREfsAxO
4n5giBQmX9VSaOLL4ztdifxDW2OvGetdq4TWpE+Cha+dtCx3j6SALUPaMmpXz1yr7xtFyu7byL/S
YvJ4n9hxBdgbGrMS4llGSOi709RqVm5C9bwREffVFTF09G1Lkmmzz6xImReziNB5qk0Pofgl3bxo
WHy3Il3pOcVy/hDNedYkcGq6IvuvctIYPRwRfwlw6BlDE3zQ1aAo9kOawiXgSzmz0LkBoP5/Wfee
QyD31rykkFGQKL0cXpOclfJZFyVcvosBCdKuZJmtUxh7fr49GexY1ZtU7kHAvjzSdGWpubsWZahV
O4BOGFZK+sTz5DF0tBUzusRuw69zeZi2OpexE/J7NBNclggdhq7oTaN8v/PqpJIe+BliE0LNY8x7
WM2M5ypAuCkKir8WT8PaO9XhzzVo6Jutx6leoVlBsPLGd8Fi6S2y1Yfr8DRPnewcL46M2jCgTd69
Qb+UQAKOHLe+QPSUzPBglYqoL2k9MRdh2BXBJ6Zr+ybUb5MKE8uhf/eXAAFL6G5LlJfmw3BWlHWa
YhcwMa3mDuZH/mx8M4ecfxIz+WYA5RJJWbkh7uQsDOCgf6sD5TSTQ5WfQYtobSdI2v4w9p8TVOhu
cwgBmz1Pp2bf3GPvrHRNJ16phBbmTtWJAMDszBeCbutmxtJVUoDtbPVhx3+VNbW1d0mP+JjSWOoD
Gu5Hti4PQmCPcaYK+0gyfLRP3yAewJGdlFXf/mXOFgiDCK44Wcw19O3aKwVFYkxjBZogzgMlIs57
uFGtLL6U0HyCGgR5vVzL1+5YAcTK8oLQV6E1tDjIwqXFW9yURqMYXGMivH2LEUvmbumrL64bkqQC
Tdkyhr99kK4GLrHMc92MEloNgyS7dlPGo6GZnpTKGjTueyImj2OwC3BN6S0eE8eolq76Dhagk5xL
pBiZdeeYvthrtgef4YinYW6MAzO+4/FMr65XuOr82/cyLHJ80lImTp8TcAu6AMcQLJ68Q1XRGZjl
/MR0ZvkKEy37sglIZCuoJ8TSupdSqIxz9bDQPAEVtwQ108Bbky3poHIA7n66tPTpHXTOeqmYecJV
/eLbPTbDm5g2Ji/EogrXKsU3w4ytX5ToWqBk6j6Sg+9BpdZfe+AaMSzAdFMqpjcXiP8n/LzaTYf8
tgzqiqGim9zt94Hn7ORHkgIU1PCbS68fBRHbsQjh7ZNVIW1MvQ93350lbA9XSHPURAb0N/mGWr1n
0yFemXhn9WsYyWAcqAMqFw2EMLsch65KQ8xNFn82n7IrCuicFiqVycYfBUZClSQ+L914FXlnYqQy
dgoC1snsyP0tecbKobdH5FsNxelH+HqCxYFONsIs7m6bNnXItD11du7LHK0BsLURAOuzNpkf5O0o
lJ0j+q/pxfkNY2FwCHYNEpGtr/qbgrr8EJQKE+NMCUvLPZgLMBPEgZen+rhBsFelwwplZBPFhY2T
5Aw9H8txajwvDnOyOMwwo0+EGTywyMlNrQhG051mmBNFd4ryx7x9lpcd4dQbwF0YQO/MvdQofE+I
bqNjWdRs03jM5ZlTgR2YHA4ihvKHHZTLgveWjOYkYurYGPN8Ua4khtBK/K5s13F+Jy4fNMpL8Fex
XK+SLX6t06ZOJ9Qr08w/dvbKIbz5fkMR3okrMiU++ciFhf8jNv+TiDc66PbF3nKNxzBbymSyS3+/
PuP5uO6EPKtIKTJwUQmFZxC9284lpT26rquF492nLf5mzQAgq7CXSIFEdxuTA3NfvZrQhxgf2TeQ
7DZIBJ1OP7qOjU9exoArVAVWDt92735FdIr68HPsVYNlphRQpSC+Wjvqhm7wt9QypNE2MtTB6iAw
OsYAzJJksrQ/S2n1QWM1QJ3MO7pa6WkQbcg9Ke603NXnKBDtaeHUv0exYdg9Ir+Gt4nByU1kbjaF
7T2vvSRIdB7ph4zj9gUNC/F8AU82Xfh358vvcUN8Q5B5irV63ksc++0BM71xtChkkhWq7r6dCGIW
tPuV8q8c95UlLPIixzHxIAiLTlQnPZrHqSRUctXqR/tS4jhIYUp2ln2qyK49NjPg9gVHELuAJrR6
vp+ZCMw9zHKeXwklzBP8Pmbb4spZ4VEr5FAUrMd8r1WwaK40tijVOYiWRjMuOzM1gDU5qwDX+u7e
AVBIUz8G8iz1hLc03CcpYZ0XbRK8BWQA1xO7D1x7b2BXe/X87+3g4tHYPyujQLrXFeBVd4lboi4z
dDI60dtTZS6eZXHV8pluHO4HlePWou6FoQYpnJHf94kDmKNazLs23/WTqK7ANiOW5nOg9g3jX6vC
gaY3I1WRO8Toi5RoNdxDwFRnIrupfR24uG9zpgvaEJ4Wo7Z6uGf/ZH+AuonjkM1iw9jNTbbHjJRL
aHJhWTFhs62ZyjASEgwIo7iP1u+7M7LYcZcL5jxMeDGHSAnGnirUFkLVDZmSMuPqnxqv9t78ARO3
R0lqvDDsXcm5SFT4ODSaCneC2rJS7lAC9kc3lbg1BtwufosyviOZbCADYWstxpfk8D27xuNo/vqT
mPnNn7Big9qE643qp2VF+u0R+WbQxhAKK4g6lJv6wmLPjI/8VvQPNCWR+hyJ980NB/WAkZiOcWLn
1tuhQr/1w5SqdpYgKkITHY9wVnnQ2UBeATRJGojkd17/lQ1kcp6Bih4w8ar+Eml4xUvO5SAopilB
bQG9sf4ixKK1Q2PrZS7g0oixZZJH9Q1TW/q4qR1f4rryhR542B54Nnri2l0otlc3DoO0BTHN5O1G
VspT/Yd8xWpXEjkKMqs1k9e3mCsN5FxXuAKQuRaLT2TOGmR93+/oH3REJ39Lc71lV4sQwpuNRP17
e0xb2jn4YDrnRJco/9cvlrR9GAbLRlzMdHCWCPA5nK9mbi6T/WMPd86huvvdgZnBoC/vK21Lx8rU
dmAd/V12yk5xgRt8BFPUOtKJs4tjKFyaXEwnv+QVbCndYj/8JGuixBQO8q48COZdyPdKL9VbL6di
YKTdvZK9ySJEOaDhwtWdpu8dOJwmhCrVsTiNUKiG60M3XhWZMMWNV4zf7qe7uwfpp7qo0uW/Bfys
zPomIAd8aoli5xh0iu/fpe1IbYtevG1ntziKBgDix6HWzq3M430GoYHi2YGDs6qlHyzbC+CVZvqT
9aLOhfjwzBro/N723IMYUCkqrw0zpceht2mujaxzVkD5PtV8+a5gKxky/G+4JVJnPrSMADZEL/GQ
2ddCdlPc+vJ1iOjjrKjWBqoZdaAk3ycJgdQr1Ubm/Pf7sCZoqpSNt4fs5xyXTgYhg3m6qxCJZbd8
2hVFSTibo7yX0MqZzj8r/86O5ZR4wtXR83mr1+Yp7kuKeqBJW2i66hyo8yajNYMCkbBPeMdCKni0
mzOAg3x3yZSJyjia3AX1KBISjRYswTS3PxYCRDeEgSV6bueteZZwiWfO0aVR7bP418thZKi9kc3R
ujO+1fECG9Czg0yhRvXUQBb2nyU7Yh5mZqaaAO6gRteXOXI03pBjELeZaUUHuMcC2tcctx1LnuL3
SeBdIZWgEM9tzvqAKQ8QmJLvBXoNKOjso8TvknkTh2O0YtvAWeiyYhnwH9E0RBaiBg7Sdi2f8jBY
/B3yp3KAELS306IzdE7oRkbHjNZtlAUw54v4atMqUjUkDdXG5BlzYo0OZZjwRJ2tBrYiFCd1iK91
cMpP5Er5qraLRVmtCNZbYZcu/hbvD2ufD0YNfcwRj3Tx2ew7Q6qtjJwtBkJjhwPlHRgX7oYuxPeg
l6tlJE+WL1MBwxsQPHRmkuo2iDrQ7UrBXCU2eKrcpJiPWk1P5ZcCgjBvVTgUKeu3XC9Xh6NvG6aa
nsmNCYsMbcu8GpZyiZc+uzi6JEcahFNNyeBkyUNWPNuJZLmLMYHqAl7nFxxV3Um19bAWShGFCu9p
z4V36v1LAxCXWWFTT7r6jbBCV+Vwu7T8dNYuXchO4ACCIao5gYY7JfqE5G8GrtOiPPs0sXxC8SZp
kvP81ces2OaFaNt3w7K+qnZH74nhTkI7zMHL1LdMQqnfdpxq4bubTfVBqBAwNZEpSNhUXDeGTu8z
zNaVqmT2fTbSwdmf4s40wKQoNVb3wnR7uKQfOROVeibDVw+wCzAGXTeCVvXFzsStNiS1rx2EVjqz
dgHE5KSdIrfg6BG2IaAqAsseTLIXKdhPIg3RF2a9Is1Rl3w6S0hpslB96Nx+dJHo9QS7x9laWxeb
uGuxeH1gMyG8G+dBdlhEIg0152JwwtSzT2vl1/p0HtzUsjm2NuVx4XI76sVX+roI/b9D5vVRQMsv
k8kmDet6i4ZgNlrAtMIZVImfNoeV+Y5hwMXuJ05ar4hAWR5hA0upA6TbbPsjrP+850GFjqPxLzzL
cF8Pe60VAivR82XTzOCbYpSawUvEKqaPuQqcfXPtivtLNyEGW+lMlOMDEzQ/x95TsDsAxOTYCInx
jlDk3mQY/n76kgoNtbmy3/amvxiuFJl9ZtZ293w2tOtnJ2eyo0JoGSrFxEWoE5H7bF3NwSwFzIw0
FYq5X4+Zmv0xp6DUV+pXsh/+DCUpi0h5wlsCW/1UXaQmVgRXu5x83QzG80Ssv+ciqXENOapfzGFE
V3S/26jfLx7JOxjEYa7qQVuRyJF69bKDqdpCW3DMO+Jmvt2weBsarvfF7ZrFvXvWiTslt+h5apQ/
k/7LMh7EQp6wKGwYdW2WONb+4ICElDPulp87TbvtWQe0ef8E25ff2SQcafF2X4J0Q6hA/6L3c1kG
yXxkrYKA9w1m9APmXJP+Y2rI7xB8z5+Y103neJTd2XgDc4KAYNlpevHTImxNj7Myxko0r3YqCQIH
xqiaYF4l/sEWV/FXrtHIuayNQ1Xglgo4k4nyPvolPpAIhIl/0hp5Ey9zQmtNuCJXcLxWKXJ6w41C
mNXS6eoQnNu4biDw4z39quYVus/jBMYU55gGpaXDuOzYyClb8iAL8ZawkjHyqcGpYf0vv6hQg+7E
Zu/fKyITOrNbeS+d7mZrIEu3CBdLm0cWx3pYopFrHl/eb+LkY196whA+FidJDhKyRKCiDICjNaFM
ybzG+6UYQ/M/xBmWA0K2lsPdDlt1mAH2Vpu+s2jSBkSrV3WV58EnRL+VXlhuy4Wsqewo6cElgXFp
0+mCa8iFVMt47Ad88dyi98VLtMQPES78BIqGo1PoIPj2qwRuYf6n6BYIElcbYNIvstBF+h/pBiOr
F8zoOgOjLYqXmJidq1bx/nHCUM4X4wS4Qxj9/iTTcInyL3NbdWtmWCs7xnM/JRWIznTMhmL0b+17
13KbgRFtWSYs5nIBBNIem8P/IpVIY15PFmlaxoAKtcg0BK2bt1rbpzgHVH3gY34qd2d7GiaGp3pD
2ekcK/uLYKqVxPFTHvEHkYg154q65R4hxO1nqHrGrKBtug9LeSrmnJ0SU1cOea8gWb8Ymvx0rrSg
VUDnEBdFYc9Lf6Zrsf1ZOHVMrR6TVAbAJKFdO+1p6UNCEVtZcItz6n32kQ1U8C1tsrhVaejs7lxQ
zRLv02JvOkVDn1c8vzyya53PZBrTjM6BAd4O/7MnU4blBOiUyDJYyWnJ7h70Sg0RCXvOiAij7DnL
iiinP+tk/W2KuZIRInebw8Pb+hn0hLqs/lgEs0GwjPIdjBtcAe2Mx9bMo8SRP2yQjh7L2S/5G+xg
mhvx2G2bgFQJ5EK4GRD21M6GHeee8Qdj9BLjy3dD7elzS5269EreL811jLuqwhBzl8BdNV4DRwV+
NtdtALwqLyMH76Elh6zpdmCeikY1ldujDcG4nXxDBuEASRXVmdgH2+cqX4kKZGUlwcauKp7QBXoX
Bc48jwACHWvpSc0XqQbWb5wIgI0Q1GcO7F0uIldyZ63d0kMAiGYjfacyp5/0cSHKVC8MX+uzVyTq
RWR0isFLVhJSoVWibqt5pCGTXrU7rYk7g62khWlifvVBipIGu3tSPaEUfr5f1C0buxdRX5J1o6HM
9raFVF/RohhZDSwIIDKO4xbJT6dhRRp5hXdaWo1UcDYIwKbG/rMEgjeVxJfV+BxB0sNaNZ0YkFJS
IzzOPKAT3oUh3VJdOHO3+Jdr8fbEC7IE3XEgBBXM8m0y26WvdfCID40VWaetPzIpRtG8dRAxsjDe
fyn2scCYq3je2TJ+NMBIW9TfTvk9n2G1fSzhxYETsiMRTkLR0DltGAsiEsgZL0sl4YV2yrwuRuro
FP9PXLipVhkhsWmOFrWqBWYXYOF8qxsDo7HEfNzl3Ydonkh+EsOLtCsnnNKh83HtdUNEXCdW8GQ1
zRzg7SLQ+sZLyQrElLpu0uCoHTwmk/TTqEY4LgGSKs6zbQShWMCcqHW7H4EPkjaNn9Br1x9+7Qb5
qX87BjN1VQUVyTR9uAJq7DcRmnyx+FJjapKZE4BGmdumelX0xYxXFGoK8VgCt6gCN91Vhc0IJJ3m
W18s1Dj9uOzK6425W0/x2dU2EisrsUW4cel6u8CgydDSh9t3xIXxnucZ+hfMVR0AxwROF10R6p3f
Kbj63aB7XClevEG+sryxDbQFw9GwqrNgxsLwJjzlVH9sTqU0P5YQYve4HE4Fn66yRwZBfnPYkvf6
/vLtGDvaTNmD4T756SJQRW8+eGAFqAQ74NTW0YtHIGLPosXWjb07/+PqxvlHO2nCGCsfn/lDLo0C
zSD+a2ozVxUCCqyPinrGIOOfKsHW2cMQYLeeFHEDunSCJLy1IRWarZsLBEMK40y8Tjn4LIn0NTW2
GEW3vUUc/toLWgerxVAEgNsMid8eMYSDFQ2iE5RDkUJ1WerCSRFyIbyNs89PgyfrSaJtGwaMXz1J
p0iVAyMgwM+mP59KYTvOrYTIuU3wZWWZMT7+sXkDLjQAKTElts/7hZVOtNW7pj1/Lp79iJinUltU
toMjXAaLBeiXbZNh1m9eRXpyQ99heSHZTS+UUpeaFejy6xTlTYZ6olr7CVgYz/Lnt2BgDxaX3UJC
jyLldKy9HuGjkYp9tZWucUrfEElIV2uuLYqGV/fc0v3J89OSqXSysw5gsYkRKD5osegkJIjS8SXW
z0SpTDMn57oPyFEFTi+JSyHHEPk4sdZ3gfwNl5xUOAt3FfCDqUXMZb+2cRptR/OBzuRNUgxJendH
dOZTdXXK6bZBu4I1fF1XKyZqAgQStTI2qfv1I5y1iL6FbkG4f8oegJu3vkNtVpfiFrA3JoVi148u
DkJn/qGWdZHxBz2rRLWUupUuGTNRS8aAnqYfc2qLnVmzROw1E20sP48xAkPFBdw91dXsVG8y0Cxz
s77ZrYDW3Qb+F8GJYNw3lCZr8uB3PXz4l8HPgjPfrMyL48iazAzY2Qt0RhOe9MbWxz6UbOTCzKMa
ZvjmN0kXbDI6XWuQgPlOPGhNDKvAj/6CC3a/C3enOXNnPcbKBoAmd2l3AMxTPy0lU9QP0HYZJpcV
tEC8MMoJNwfNRV60Ne+oUreeg9K6T0J32kERbgm7W31EADoQHgQ2jm5Od8AFHgIbY34cMfg/5W26
OsV99gZxR/F7cPX6IjCJ4mSegNgTrOvkuZzETthU3OcT6nb0b6DxBTYyOMm6dVJpvGZatLH6blfX
nUJZ5HeoHGClpQjvQJDFkJ3VKweL+Hf/dCKQR5o1o+NrcHtDk+MHYN2BHeI/rLBJYHtxcGNOMYid
3Cf7xzCUncuS7tfU3SN2Lo6GmUIX7K7j7DRRH8j1ltqaqjVvc3AY1rwyoBmkdNwY3bpmlavXFgny
+S3y5jSdIZNsax/dSAGt940ksjJ+5AV6LhZw0AsLeCk9U71M6HJ8QVHyNh/+80R/qiRAaBN6j84f
6k8N/99BnhUS3NQk3eYTwIk8DBwk4XbK1xwnYWfirwGFM6JjeWJiJpKAHl/NLH++zuTkN0HS8eGi
F5S+LyHUbqR3TWi6V3SuCBYir3MzEMtN11Z/MBX3+5iBt85IK25htRHk4blRV8byIJnRv+saqhTs
aJ1hXv4LzakC6o4uGb2FEvXpNzTAprQ8AdCm3FkkkhcJyTmvFCbPW28jVR/Z4rIzUW+0LsdB7v6A
1uBB0wtPxZ+8SlyomWzWlWiakn53sigyGmTekl2AqXQzNzGN0pLbg1Zesz4cJcD1T/BeZyNsjCcM
VDPqfQswSQ0z0QVltFepTUnz13BBtVIOYlHkIIrE8ybqW8jHkXhVF7BxTmLSPv8fra+z8Mu3RteD
HSms2sJkq+lsBpcpRiHcHc1akvetZQE+rrTrRgHkJmEioLbak9ZkaXNUdu/6VMjk0OB9+Xa9zYod
7qFOJ9dqkkIgwKdOKGVAD/X4UgzRcoXSmX74pwGjF0ZJ72wiwVVyv8Mp2N6q6lUmImPLvPauoXDi
Xrx5zrm3/ll3wSYxd0Gfeog3Z9Wx1nBsZ/MGS+M//1vg5q4hxc+IZ3Uwxh0zOPRlnm/CxDdRhuv/
zPZuhXRNfu3YgWr15jJtaewedGBv5kiqA6/oWL+cTAa/wjzGrt2q2whSe9KlSaGmid8eqYamALEq
1UPnskkI29RO4fXeZ13FHhQgRuQEGXeOEs7U3MGe8ZxPqK7uV1uZh75TKRg8q+h5g3/BSCIdQ6p3
TzitnzNPeADxoxKN4WvttQbWMmm4toaHID9twSZ6tFJGvEMehRAwWhHD5QLmJebfJe/R7DnHRyZO
PqkOv1ZPgFYeF/u+hGGBeZOImx+nCVLZy+U+Z6LsSPpTFxnaFNglD3mUwTxCXaWN9/1efoU+6crT
F50bXm79DxYWBw3zmAdzzkK7tAuDaSVocx9j06d42yLS8TYlv5fhDb6SdlEq7DmSbFztZTQ5AzTX
MO2A+dE8ZMR3gzBQo58/vKUB5qyqIYbtY89QqAX128oZ5UFue1Kp2zmPKv5IOSFgKySFbjbGrQmG
Z3UIR6hSb1TYqlp94lbWpaYTnh68bwJ8xJsgoH8vqTzEznaVLMQzevEIO2pDkautnTjc+M37Fz0o
7ZtotwQOyALvoVAsk4c6ifNDpOn01GJj397Bk/Eq5otMEzeiKzc17uu8PKohQijJHlZcQ3v5yZhw
QxgacGuQ+u9LCKMy6lB6CeSC29fZrGKU1enq0+0AhCx/FS6d6bWEkmvGoD+k/OTnwTcC81Z29lo+
V3UG3t/+GS+ctzGQcKcs88il6CzQSuarLt/XPs/TH48JjxUihwznKN49kVdKrcghuquB97NI9A+L
jMjcwg3X4CJuJosFLM9wG6QkOlFWzyVrLDGsS5kmQHa2XpET4oc+SQOxrN7DeQlSf27MzwcI36Bl
vTUrLcF3WPV87Fy4b0J52lFKxFLisjyOLH3cwsc3aQjBmAmRXSlNG34OdkeI4N70iEjw+aAPE5XU
m+i4TrsBaWa9NPxrzFwB5T1Up36ADiS4ha+pv/X2dO3E7cmWt54Qw/76s47pkzvHeE4UjyOVfIZR
WUFi/NTfpzAhJNHHaaNsRRsmulgfzT8S3Zy4kyWAwRQ6rXntd02VtLAUSDu/BtShQ7KRC3pFOrH/
kGp1ct1dwMURE6LOnNLQ9sKzu/xV1oNNE+cZSIMrfJzSMWhxN+Fbor/pLowSsgnyjZqfPYJnNX4p
WWwRFE9aVN4DitVFJxNvMhD5kr19+/CJtLAhTHaS5TdZ8aHz5POZkTmgMF5pTthumwv1yiWwaNWi
YGAwg4oz+O4m5pE37S2e7P909mWs/WV7gbVJzN6pO7FthpXyHr+4qbPX6x4dZrVbenITHO8Sgisc
ExksTs28qPS5sM4kuuUUtvfqG7scOPgOYu/wTWkHhdywVdT3hX+rr0TNaWltOApmFR9H6cQ1xGFN
Sa6xBQSm7kVU9nqmJIgT8JvQuc7xz2yq69912gash/tq5U5z1lzNeQtOE3pecaxWLq0fSES9rTBo
D5JUdUdoO1j18fVmujRxea06s7ZyVaLxbedRWrDQHy6xybMKur9l2rf/xWnGRThA5yzLw8mJQdXc
2Gt4jfjyjUnlY76UOSMIsUNfifuZMcb0z3mzNtf+86PhFibCRUD+x+zP4FVeZlpjmBpgef0CC7ss
cK85ULdbLBUIvK+pkW9p2wUf2jWwiRCtQCjYH8GOoabIE/21Xzksxaynh5fs/cwX+OiUR/sPGR/Z
zv/hMyFYzts7qqw4m6N1ox2Fp8xUni4H0Rd+jr9G56CipHZ5a0xbsJacShPxHZB7gIALAWHS4+LT
yLxneJ7eoz/ErLt+wAlatameNKr9sC+IsP1Xy4sfaCc9EjEz18azPgfQMG6gqDpQJDb3bor2ckeh
NJAxL1ghj6JqUvjHiRVd1srAEHCQH2uyM6yDS0NddVBfZNLShF8T7TYmjt+ekzjhNYfm14xOEW4P
EUtO1wSya3giPLPCcwkORt6rJdYGW+2H5kLBQVaerA3lvdLegicveTLxcFSD/89MWM77fJ8fKNVH
N9ZvNubGpHkTxXiwIIjCbJ6cCOa52qlygF/4y8gEHPEgJi1cUBCpVSHjPGQEkBcZ7HY440QFuiRq
5cvEjuvzQ4/G71R/b6fPr87VLdXSgEIT0nb2ujVJe0AKo11Fg9SMZxQ/pIJAJL/lgBJkrbz02Btb
3K8Fz70ykwEH9y7gsvj9ENL7eNTGQaZ9quogP69eFLG7K7jOUfE6zOlfk90n7fZ3XxAY5AoL6RLl
52VHebvYHdRcBzmAJAhqMkG36w3VBDIjmRSA3dX7p9xoHFWkT5W7IbtW38Vgv6gdi6UyCl44LN3f
eKB7dPsEAtqFtpPcTTcDF9RIGJPytritfm1J+b8cmG3EL3Axj9nV2JWNDH3LYGHoqyEVz6wepqpS
WbyWJivy2dsLMVBv6wl4CTt6aGWeKvn/9/hx9hDTFd+LN0qzj5dSLYhuxwonQckmX/UTE1DiHTUB
LzSO412upZNauAxpMju6cjBGrWlRqeAUN+H6JOH0yxWZO//AGf3LvPzSaB3SZk6ONnUkKUW3Y995
jFt3sqtUBmkaVmV8kL6Jw7hin4kapnIfTOM/ZdAiDn17tRoRHK4tKupGm571vo0G/oW0VKnla47K
yS94EfiZGmEh2TRoPJ7NH0+z3WG4vxltmEP8wr/Rshr7ib7zdhXXXoO9hDdJRunaL1m6VKdLiDZw
xR3xrIOCpEF6F9NcQPOmPz73nV9azqiqbIp51ljaiTEgol4Gb3OaHDfT3lnPEAzbrjY7yCF0T0TX
vpSFVsMJT4T/eDG6eKCLKGp5erFO2XvmmiFMR92CN6UvpqrYknYrtSYdiMtZJAvAFk8BUowSZY5C
bI3bb9FABQTMkqNsdB/ydFWoKwT9WDuv7XH3K3upbjW0VzOaBV7DWUM4VnmbY9PLMcy4aBRL8dY6
u1Z4o0P8T0TQR69uAm4svarHBVMaMuSmXtf53NfnH5g365i6qZVt2dC++qvr9MgIxYaf5UXMYacT
5wnkmMUvi6pdBUCEogSnKVVbYWt4w3WtSmrbd4bUidCa336Wv4ljsSSisJzi/580Vl/wQ/ekLgmt
R0GzEg97/O68+abxleF6fvyAbUL0e5dNYxKrA8iFOiEdRxtPN84lTTBsUEg8boFkk41lRBOTr+mH
EZvt0dSwzsgTpw0k69jYZqTnnlRtz5hSALR61NoG1zQHNXWcokdXWvz5qeQilJWSSBuTs6wdhNdt
DMxZpdBdN0ETuqlXxKoPJQs/wvADbQJ/xmNi+8+NkiTHd+mRuPKxMrGP0yO6lgEWw1U7pCVhjN35
AE3XAVAhRb0seUCrPNHnfgEdw9Lk8X+Jf0rfVqw1EQAjGBlj4nsqtPDQ3Ivn3/QJwyEqtmtqmNdS
R5Y4H/ZRHnm+BrBzxRncgyIu4g24L68bwjPLaJ6NeHWRTbjVfiW8B0BixF+V0e2+CN0omh1wdc9x
x8ds/9fgm4U7JqGPoR+9rTdbU0LLnfmeGEyJCuuBNicj3Ud7zpNWvrP63qepdyFaqq3TI4iBJXFP
VQoiJZFrB7ODxAzKzZdCFRhOc20d7T/+ktpbC55mnd5Y6l95IubYq4ZoChV08CsdurcmKfnJwG/4
Rrjg9bUV1uVF01sucfD1pbL9b4fBqnUbfv1CxX0SK1R9+FLosyYgupsf0z+Z+YVHSpm9E0hQHEhD
NsztXRcNFpzQ2xaFm283Qh3h3IDdjH9mpMr4gsC1NQe8B82QVwC9LG5BaSK/eyOVdjV71+x89Y8L
lHzljuwGJ9e6F3LChDYrqDfuf+x0O3PJ1PgTLuplHHo0KOOyCR+d1wNs3Da8ymMitcX5jIeinTgV
IqPCVU6K9yKUXfgwu0zXZayqOnPWUvE1k9eiSaZQQDTKcHRhbkPBJMA7r5kovrUB9u7kmIgoMbOO
2pAX2m2ZFrBKPf853ShBi8Vfcsrp1tyQLrT7RsOjbJYYthi5M/iUrNlvSEfYp5Jp2wyTekP4qmFA
s48iiJfQ2uDRj27e/LRsEYknPXylypUAaaY0ogpRVaUE8/FdU5FUEa4sZK2rQEpkVmtwC0HrnYG5
ULuSPc+oPTEtga/+lgmGTxSmZYGr2ESxFv4LWULyjhrynldxqKg2nmrzcZGLFvsUPE6QCb0uLFxe
tWoRj3NDxB18/KsbTcDUh5EVx//cbr8/mZ7ORxT7l2TWMLuFfgkmabuSEXbcH8Rcjd3RQJcqzL4e
Ff8Y3Qqy20dcwIkiXMEizaePoSW2DfYBa1pWGCxpIpTZn0c3V7YTat6uldYi1aoYXVl8Hrzjf8FW
QASyFcBplDqDaWbiL94D4xhrwsBa33MUke/ctdxRNmO/Sq2viHR+25Q6XSe3TTcsa/r8M42Nq5kg
NKIxNFIKSZBimhI4rDKT8tjl/+0r+1OMvgh8TYEcg+dF6H+tMj4UDyiDScHu/MU/DFakRkyfZstS
JskxGyZM9GolwjX7CPljlHw4vXDbnCnQjpnSvhU3DbONncaraJFNadeNWWjZoWG736cHHhNUj7at
amS9L8sUKA7v1p6nF9Jfq68VOePy5hLTYaiEfiPX9UV7dwllnl4avN5j7JnCq1kCEMnRr8U6xQKU
6sUOI6tJuBKkhvIE/8eZuk6NCE/2s8G1ia4DJakLMJF5wNFoSNmIyZ5YWzPwjq3vIG80JpGb4/Mr
PUqE9uud9A39oQ2vQW/Z+nk+KCpSZRScJcliZBDIh1L58uYsRoN0eKrhT2j0DJyb4Npo4n5ZP6FV
QcX0MzPWut/CQBCh3G7831mJUtLz8V5cy4P8TCHd8xU8kT0/PtfpjN7J5IeMxYjCH60vA2csB6H7
DnBgbWy6EAj/IKQdb4WyFuk+tvsQsY0eebcHiNNRFK7RBNAPASZ38DVW4OTYK1VZCgvHkIWCiHdo
Nvy3UPuaP3fsdwjZirOgh5LA3zDBL88nAX3PMCZaUXVH9UKFrmac8Z4uT72hopujAkQ2DrLvCZ7a
1rbY2GhZ/9h8nMePyWcFx7pkEKz2bsx8Ui1fhXoUrttURjOk3EdiRdfxKfmakKrkGXR0oT/X2NNo
VfAcK2HfOvlgf5R/xrDYfIHv5W3KQKmNxOyFT+Nb7nkYs7usa2c8dMXxVp3rBqQJ5mIiCSRmmnPE
6XD2jHfOTCR9OeqR8hh4C80MMS+msQxh7beaaBjM8Zy5lB/eNnBbhHVQ2rg74Y+2Qhr5/MVLQ9D/
HeXSA+yVcOH6isXPzywuJ5gJBmXR+2R6E/eyaVyvAPRDX1hrBmNKBZwPwXBXiPr6dT31Dw04rhCL
nEgF70Zxi5sibDE0qiy9jav/FqRka+Q92pmUDH7ivAm+50NhQ7ZVDJwxC3QVRRkmmrR6kpu/DKJl
SZSc3DJyFFFOOmTd4zbtJ/9lv+d1VD0hc52vGyu1EyoYEPpJkzgFtpQ+OzQfnfBtmJanKOB3sCHB
QWA3EBAmZHmYgcQEbJupY1xcMvWJVC0QycAs3K1mJsnXHIgybQ0Ep1MaIFbrw78cazFuJeeGvZ4o
t5lkkwYIJjYCTewvGs1MAq0U0b20T2yOZUid8S5ok+G90NFA0I2smyJEGksyNAqVQ6IxRafikQWU
B3yGuwCkf40czHSJ0ew+tpuc/8Fa/C6if/xU9PSUQUBxSJwc47XXAAgKBm8REbs6J+6Fpdqi/sFR
pNfjTkDWEkdfX8qWqzievXA6Mgff+D4cfz2RsKFYPIsykhSJff+rG0xC+jtVkdRwRUZ5/sChiPVZ
n57K6yXt5vKZOLxaKtepKvTtNe40zHDdMfQcpbUP82UA/AjUbnPrFAU8jz5xb/ZZ7NV4AQ39i4aC
dtpuItpr4E4U13ilxhkdDENZGFg6DRbyoZslICiGOcFVv7gwUBA1et7qnWdb++A10X74hyUQmxJp
AIx2wyaYMOn3LJW5eSzgj1iPVA1qwvJ7hPyZMKD9SXwqQvRT97T1tfe/39VRG+WH0yS2r/LrzY2F
BCUQQ3xfYHEeGLUCE3lGAZQHaeI/WPLXtbU0I9MxHLzSBHt7lq/RrRmG3LaI4sKYJIDUVzySC3uO
P66vGr0P0zVOCrgJo6eTHOPgxKUYoq15dbPLxzO0rvYvCtfmWFf9fHCBiwTDNgrwOa6k1tANxsp9
CtGthDgiAspXjcjcmg4rhO6XQwAs0SLtTBIwQLSvsajfhZxl10MUAjhNN69WFquZsS1s31nGDAz2
aUSRgJDuX8idzToeoQD74bqvk966T6hQJMQ6/kJEiUmguJTKHNF9AzHsjKWXxA+/KewKvS3r3NyC
+Hsr3d78/xjMzAsVyJBWQCTOvgEQxmuzn6KuAJvR4Jqket4BqpJbLVxX3Mc00o3azy3WMEOJWHTx
AZJzYMc2h7/YTpc/XxoFdKoVYvmmDjjv770vhez3mfM3BPqppb51tiLMDpG7fdyIBQY9qs4RJFvj
1vbg18oyrxDbTiwoecpSoEYgrvmskjzH4mRp1UWsggTWsdaU//+VNNLe5lxTL/N9crgoIs3hdBXW
HQOyjnWm6IKNHttSuKOPBQMYgzA3wzsPP9R0YqzMCAuliONlisU9P3NPyvcOiUP5d/wAHC8FKpZm
CX+Z9nNaU03/yyO1Lb39BociVIEwC/lqfFbvqbSDQi5Gr8/b6DVfJCIx46ccH47r0+jp00huJYcu
GlXGM8Nk4iO6JAhqOV86a/H3QeVOIupUT2LaCD5Zw23rhAqAkg1EMyxadjQxhiyuWD3+jqLKtv2N
Oz9h1vXKhv1QpOB5v9juhikP96CI8cyRdt0o8ykSN5IP2pLqqIy3AqB7TCbRdUPYKuxHjWyV5o2l
BpppcnSf7kbklveFiRCI1lH+v1oG9ZR2O37J97QjkTp3Bln6qmdouDGOLfSCEjzSg4YE7nODcvAX
eNenqVC/sIc3YpxJcuLyTtyCNlUBf2o2MmBySAXMnf0a7hLiw7D8T2G7BZgKyuKCKKYfyOkMk/9S
H28SljfhHBDo2gsmG81kGYXD/JxUAH7ALKNQKy3DH2MpzSQXYUyFaMKi0S+P+PWJXAGaelg6tKcV
FJ7K8WG6e3r1qzdKafHuce+ivUuETp+DU1Wgiha/Nn8WCACpG/5RXDj63RCNKnc1vMbxQUGJiGcU
4FOubhuPwgkBNTFUHzT5gaiNdAkoexaa7IpEGJvtHvlhY1b+cDbKVf8biNC1Kq6jXESi+VW5cs1p
AZEIzT+a1hlCGM9iYaILyKa9eavsE8lrcxVv+6b0K3AxMGuB7KMxdzWfbL/uN8C3hvG4/DXwQEu+
bY0xbZiT4dCcPuX1DaUIl+lS3gl1a+y8JXz/OJVUExq9fIqFFT6wuzN84n+XFOkW80ULD//gGb9B
3r2f+5yCFYOnEmIBH38b81QnH8cu9a3U4wui6l3wpGGBfwVB9tBRpFh+A6g/5Ue+v5MDnBvp0hjo
qIonQNUqr0ALQmOq4Wvj+ObLJisv1bbHcy2wRtehRhBNmcq25qVY3Ev7Al0FvzmiwPXhJqxp/+0A
l4iKjx7as7AehEYL668KXUdlHVRXUZRuwnIcB7IElz96VqiJ0Phs1bQqJeIrEj35cA0PnrxsrKtS
/cm1b4wixy8qKom68Eew0FiG4C6zH5v1qXTdCO5ML5mkyZk5g6QXQkH2NDA4GevdsqTuLeL95fIA
Hb14pHV4Pncik0Z16ybT0Aqjuzaq7o0q48tE42panovC9evuwn2nkgbNJcZVZcEeqosznuYvXSgC
ufeNOvLbnyOaT8cfpCH3bm1Tlm84qEqD0JnWqYlNT0vy4a3XFPNuPFi8EMS+kljbDEzq19Ict107
y+oiqrZEMPjgjtDCSfsKT/Ypw8Ir1iWvQCsi6NZPm41ZMxK+n0/uWPxQfIxO4EJbc6K+8eVTvTsb
UXee5mF/x7uFR+QUwubOzx5CyVZbZPo2e+QFFL6Xjuyccy/j4ZTN3Q11r3w7ELjsjB/cDKfYkAdV
C0U1QTDTs7bTVNRj04aWFb4FagEz3WXGZpBdkfxgP1HrGLngfD9v9kv3/TlLwYEOLHtdGK+xQMWv
miegIr0SqZcH9222THnC+t3+ji7RrRm18MPjAsaDjNtfoPHG6lBLxnm0KiB15cJloqmyFoovlFWY
V7ghOTS9TH2Gy0esDZqBjLGCXLAyMW9y4jRqG4GqXdzfYrrP3dIWXHWX+8/7FiH7HvvZwzQ+sWmC
7bhbWLAYmJA3cYUqxVVHI4yJ4UKG9Wvec3G30hITLyZBRcxDhTnGyeKxRtTuSAiz7KK9vLT7qzed
rWLWFWBlDWH+I3HWlqJJNud98WiA7fw+m87ALtHaqdvMruP877s80707gXRHniXz2PWGXMz/Y9aK
vhgb+M9duLn1pRy/0PTEyKGbdhyHfFQhMcBjWRCcuYqs5Wc/PRFOj2Zc73ejrMZnvZpfI/RLOwyP
EKLN8sbmHUNXcQHepG+ZXAe1XLEn2DJEOkr6SLmh6xxxVHx06JrO1Rx6KwVNaBBqHNckG2WKWUH6
WFlDQNWll7w320XNZPc2PL6dLvSPUr0qe2fygLI7yBaWs3H2xFwoeKAKvmqjkFzXbgB5mSqJEj7j
e1Qh4AYCL4c/bB/H5gzHhU9i1wOaFNcVwFm82HgGK7R4B0IguSPPRiPFng4mrCkj0JcZF8+ZNc+9
ogYbrnNGj4diFxZolBEj5mb1eT8/C/C3d4R8Vi1tG8Ha51mmH00/LsrxzPiWpGKK3T8W4yKI0NfI
K0RcW4fuCg4p2cHuM8UkbpOxP80QBHhW5aFtpA5o+zQAeqVdwSWRv0Pl6iwxfEIEwMCZBMEQ3q1o
bFOz91i/EylyBHM0Rp69F760JyH7OEMrmUv/8ZOPRLpdA2+WInSVK0kGD3bG63Id9JMwBHCQYt98
PfWpE9wgmHgM/nENRV2SXxXykpsl4HfhsCpgy3LhWGqZ7ggNyCAnaNNBYZnJa2ZaoGPcH/RnrvoF
/ZG1PAmr2qrlWUGGXOqce3fk8CTY1pGAQ3wdXaGVeO5Zdu+M/DAkgQKyzU3mKWF+0ksk/9DGcjE+
tXOxe5nQlVielu7EOa59FIh8WrxtAb7pzotEE+bqLMVE4V0hOWc1RJ+Iq95TKhSJ7Ngs0mJLqsXu
/PbFo1N8oLhZ41t3QMNlIWKz2RcINVIq02TjJJn6dkaNrqeVRNWjcuL7ndY4OQ+FBCk+syd0vbNM
JdzHgsmCoO3Efgyh6eGxxznBuikL6hzibr2gU8dYm4mnXsYs7Dip1yCTu/N1weYL5PS8NgACY01Q
soSJM0fuUNw0fuZ17QFX5g3LWdiIWH6jFboA5qs1lj9dmNQc6fFO/yKNxSdsb9d5Gc5a4X6rxPoB
mU9KEnzNE/GnujJukOnbJESxTqttUMrunJWNRRcrkdjcTOJnZlTp7qhslCIESzePlpjHH6eH3h3z
EPNGQKBG0ISTv3LzbD8401xG0x/4qHAzAWViSELfgL4MM3srw7RIKJhDUN94YH0EUocZQ7ekcHQg
5uJWO+65Z9fNGbIX2m9SPT1f2qxCRe0gX2CAGpGmfr7J4lrBzGenAF1WnLkMWIHspflI5T4sQNkP
m/JEv0OgA6Tty+U5elBK/ciRDgsVtEaIT8Ld/sTAWAYXrnvBvyDJM/quiMyeCVtsN7J60MfAnMKA
BeokDkn87leM9DuuKJ4COxNnaOiGHuAUerLbigSZi4pgBBpVeznY0o1J7YUykPlIBD9iuPJsnlpI
DLrLgEkaqDkru6hc7QE/4VjgsufHnfzs0p7i8ITpWWHujoSTz/+RbuJREqeD52QRQbEy2PLDmrnK
WlSA5gjZnvIEHWAe8N7jDxI/73CHsNiqKPiFFP8YR9c8nCSayPw+ss8caYuFYVg7vhAAoY16W8wy
cT6f+s10YpdzNKNOoDWoNqasU/QUqqSPcdsvkACMOH8T58t6U38cF9CfdyjQlIX6neK1dlOVkuq5
xAaIyNwc87gh7pLYHQNO9WBBrJMebCMo2vEntRn6pmF1Pi2Y+8yRyDJ8q3mYpzVkWLP0epYq7tFj
7wVZ6/QggPOID7eQV6DNf9Bkl9jq5dieWL9d4NQ5i4U8qh7I25ACLIwVPzJP7/ViQDpedUz4bETk
EvZ5MF5KRUg6ei9B2F3iD5MswuYn/lCF4QdOlopjPlSxmutgQSlEZo7Z2ODgPhWt/glsZW7vNJzF
Xyu18T1/tHkOk1N3HJdyQ0i4iO6PcjpnRMSKhG50G2Bk3lIW3AC2OsEKIKQaVwlMpWSv9G1g8mQn
yzmFfhDYBItz7rPdOaTgi52jHLKTslVYv7Zksm43auHai6ZzQmc1Mg1bVOkS/k1hrEwCDrRuijtg
lULTbFvXodZqWq/jbdiTep25zai3bm/Q3aW5qTPdSeJRW3kEMX9Q4qsotX065TMmLlj378Ta00d/
oNmDK5Nof/kUjXF/4bHZrgXNhZL0D1sGwcIzBCp0svFeNUN+7TYBu0VGsVciAnAokAa2DAEUfw44
Q/HEksKxGqBY23/3yrV+sq18twSVaSaXNvmaAWDoIHUyWKLScyXeEvRa9xl92TqfkTq2f13nIf9R
lWRm0/QgdjsyEC/CQcwl3GAKgpHTyxk7Wo1ZiIxNfDL84GjRFVMBksU0dUEzon0ie+Fzrl+HQ8of
Dh2EewmWc2gJAUNQWwHkfuiLVGU3Ckg86u7vmtph+fe6xKaIU6nBAhaFPoxcHnOTrm1cN2U8fccM
gM+o57WXgUFccA9KLDmOfaCZ8YWxCNZwnO1tNobZX+zNpFLIzDlfAaGmBhk5BI2fKsxDPe9uOCxZ
BX43/iYKkxrsdgsPvpQIb2TVdPEg1p+WfgKTWQppIe7OuH/6bftpCYs6j13KAT3c9hB1LvN/SS1m
FMxKZ5G3IwVWkb9x/sP94eB9RAkWQRKwMWG5M+Domn5lpLZLfouJ4kJk+g1CkAK3Mf5WQmhKnl9G
sNUy+gfLg1vQrLiACCT6sV1GY8KWWL0khlarNFPkt+SH10e7dm7I+B4wcoxYarrI3HmQDnhb3/Wt
gqOwkWyRahw14SdOJH6JetVDuzQ2hRs8WYtdKbq5S+nrhygWIqY7YBAQvkC7EbSmxMJhRqv2XPFv
x57VcHMYAAETu8wAU/mpJGAVd+X48DjNLKruVHNbUC+LYd/P6UjcjXzjJzWZmKIJIa3Nl/PG9QOQ
vm9aQDUXzcJpyV4hgbohXcyocjmkmQscpuYzfzDP3cWs+ydgc5kl4tp4WwBHF6Nf+QoXX3j2rium
XDyT17UyzEv4sTd0i78CKelJf9p/AytHa6HmkPQmMv/oBnng40i+K+opAh8zowv8pHQl0hv2jL7v
yvpnNe0PeWndoSkyBhAxXfME0hLprdSlFym3HZNmnQklDYvIIwN8RoNaAAffi3so2A1/ksHBwbf2
IDykP15SVuX6B0qZ1brSPMR7T95SQAbKG0wYb28/kuh9/h1j9mbokmR8Q2vJ2klVq8U4dVxcJtQ5
gYYfXr2IY/zHk5ZeIzpJYvUfhaK/hYJxQl4CEhP3bxbh7X3TIte+cHC3kOrMTbDFEkhndMTxLNLo
a4IHD1jlUmppaYspdE9Z/7o1CtIFUaisVZsq/E8y9ZQRbIRoYiYWs+mKQLfGSC/tkHH+8I+UwU0+
9phGfqkyrlvIhNxHq7btQ1COiUds2wEbBfokVC16au6zTO3hf4c/S0+FldPMg81IaPs1yVaPxj93
/bCWSypG9PPawdvdJWaobyYscxxWSLKwGT3euXu6JU0XNmvY1SfSOqj50dlQdxu8yao09i2gthyW
lhgSsb5hq7qO9wy6BeNZMiJ0qXaIFAY4awRk132h1LDA6GjyMm0iYdxRRWWCqVA720feGD7ilXBs
baWn8YJEuIR06vO70+5RjFdc6Y3MrJWzhc9oexBM76Z1kLcpzmump/m71FB4oBToGkkzpaAyk2GO
zK/8QbnoGdUbDoiY7fPqmGiO6wWMMYLSUx+04iraFqdANLPuRA85rDcvEFvN4NhPHIF8JCsd0UrM
Njwc02/Icma9op+aS0W4L+MbhCCb8Gcb1U0IebS3FBsj4gOwuvsA5wH8VUAa3g5Oh5CR6Z1hGawb
KlSX5bTS1EIgehGA3mjyENZqm2w+luDp3NclMa1w5ggF93vBZSZSiZ1+mfU4MKn2n8kuNxNheS13
yqjpxGVYFZrhJ3oNIgU13w47SlrE7KQ4JD/hySlDU5k7IihTvtyPT7iI0OFT9Twg90PnqN3JX3rO
hzx8W1o3Bh3v3OhR8OEH4E8NM0uaQoBIPk5CdZh2Id5sI7w2D2CBtn7oavvSeB1K3o/df3fTtUh1
mrj207EokB8A62F2Py8Jayy0TYWWCQQMKf3Vtr5WxSrdgKWhK/wixmHkL/l2ONrsMKi5/Lj0sSE2
VPQYOYzPi6OrR5M1llvUIGfLJ8eIXurgd51wtksznVWuF3xFkT4rrs3xQYRwaZPk4E8f3hedAemy
T3BEVjLdBJFv9X4ZMkEtq8c1mEABXb5Oy96VQRuNqpOq4ME3sXGc6b1ta3PhpBkUamIMNU06cepB
7Po18ntmbIlGYk1pHhJ5YL1hkCVVkJ6nwMEJY1lzM4mlUY4s9FdHRPkE/98rTRuszZ8nUEUnQGVK
F/FX5i93QCBWfwylUgOtZkidFtFaYPHke7lPEq8CTVLGNxUVYGolPVRyeKzS5uhVMWRKS8OYEBb8
LXb+bPMAioFyFmUrkGeVqFMVAcdUvQ7YTOXc3pCMDLAH+YFDJs6PJ0KkEWOXhTqgsBpVdKtyWCdi
MDGU2wX5c9J+S+0krM/O/sBy6ogJYpahR0jWwBJfUyuwSm+k9OeuYe4TKuQdC3OuEZfzqtUo1LCY
jhtCZcCQX8WrdQZUqYYT+2H7cu3aUKELzjt3Oi/pN4+mIPD6f3ysJC+7cMVgwLpqZ9EhzG/Htwzk
NjCUWHglg5r9f/gHz/mCWBaZ0t4NRcXuTE0WdQ0pUTp2E72UDWNP3HJFzOu9aMm9dcT1yrUtxbx1
eJToXOrPwbH16/VO5RH4FRApnggeFHVlYLTv7W+ZQJmh8SVLtO1MOL0+Z6W0LNddBjN6UleJpmH1
doGSHz+GYFsMjfHffeoqOQ9A89jB0gAOYuzokQyDAXljeB8v3mAfRNes2Ox0uAjmmzN523IPuc3V
r8AJn7PjyqXI2se+lLHX7fvSbSmZf4SAph6lj2BJ64fFq+2tHJ24o48Miyzhog9HLqj4YvG8GbVo
2vgCdbps5AmuRwS5LPTQ2bn9jDTdTyqbatmUx8qRh9E7i52r6Z2iIbP+jqSePp06TRsIvRsB+K2R
pYVp6pr4yVWN3MFcMg9OU+KBMID/uJFzWc5P+SRX7clNRAZz46nuHQ2jIwqENlh6nrARfpxB2mpL
cj1rtPTWb/H2QtaBCeaz5+a838lgVSA9nHqJ8VWWLvY9CjuEstUAwGj4DPWNRkApL7sXZVR+xVtv
R9ggjEhxneal188A0QLcqJaJhC7zK4F5hpi0DfQex+EhFEaK2Zb87yBa+LXC/tAOLNNugG77nmjW
kx4YtQ6dIrDTlGIhshA9tosm0ss3wgMtSBdGt2pUm4wR0Q+Lqjnmmp+E9KiNHZbgattWeTp9cK/N
0UuES2Vw/SaOmKOL7kXVh8XkufRVwDK8jBJBG1gckdSHKn1zrhZAZLB9gybw5B4vHK5nWdC8kBHZ
ohPq2C0MMcrruROkno9HWbUvptMXsvAcy3OwEOdIEUwANeUcvn7ekoWd4RNDBsMZ6Y64ROiJ+MI0
OPWqFqnVsJHhIIv3zBJpLFlkOAtQfBmdTNDa3JHUwayHGXwBf9jc4I2M58+VBeqIGS6sRUwiPUYb
3/FsEPhZZnfPeyavum2/1SZp7QENKmkkWA98dQEgry5NTp0XZYMMUgJPuc8lsDYXFFXFAIreeY6U
BavL3IYibD6bhwXpBQh0BJislJ3KovtWsjxSEBeDOwIaQjtiAWtvl5RKw3zOfLuX+NVy3W8ihGXD
Ifc+ZVPJOHAfa6XyinA2/1IfJe6Ut6r5uGS9Ya0sZIMcvOisXDqCXussTxjzZNg6nMjMT4Wa5Kq2
XGgWYPpm1tTZBbl3QsZwlNrjAEnpc0BSf+iPRojvsWtD2bL7GedjrYLq58iawpypbHCpCa/SKm1s
1gQaKVYWdm+6E4d1oHfi+us2Uku0THfGfuW0ETT5/J/b3Nu+xVGAJ7vjtHtYrm1fzJGwQ/fqd/xm
g31oL8XIFY/IHffHnB6vBaH8mUSKey1h2iefYm1q8SAkDDx8KiT6GbfWFzGB3Ct//1bOpIW1C7pD
KyATiRfC2bD3GkWTN25r7TxcX6EuR7ofnBqCTKoItWQsek+GEb1DSk/oiV3KIil1rwU+KBYTmoGT
e2aafVb4ub8ZTZyBlAOrJGwwVkkm/m74323MGqyj+VlU6CZhohq/42JKtCeuZD2g4pJXaSYSGZiW
UV3VgFvq9RLHukO+Xw6yfL5w0pkuINxPO0Q/u9UUdI0Leux6yJF0UBBxVLEtD+TJulDcmpo6bEcX
QUCunAt+CbvWb4/8poDeMi6TGNMivGbJpMqtcVmulXKEIFltgGw48gUsMJYmMqSbl1Hv+xtFLUVg
b5Y1w+xwlkSfrIT/ePIdPHXQhDIjHIC2qYjFGG1qX2iTCYCwE+MJbEhBK2aAT102cTA5t2SCfn20
mkZGOBnkglFMwTwFXUXqHRV66+kJtLhxUTpxNrxr/RszcJ3uoxWSCho3SqtMaFTvU+MX4pqRznvk
arWxmdk9L2nDhW/UabRP9WpK0pd8Wf/Q0SjqiVifZG28/q8YxqCjHJsxpxPHiayJe2crLFOi6Pr6
ssJjKnEYigrb+yyOyXkp4T1DclfvAsSncVqxXI3mILO/qVccPpe78hIQAoo5Fd2Uh7o6dQrHhGxu
GcON8e3UGokpyWRQp9WOT+2pib1MbSwi2DzVqKbMJqXN9JutA+uwxjO0FBfNFW7pxI1mlD14riTe
G5bbHpBc6g6Xjpz8Lajj+1iPIx07AYtFqAmqttIkVIE/c4gh/wiCe9uafCjFMzJalwfNZV4DfH24
hNmMRZK7bMIKz/yptwmdDaNBvB5RY2mma2QQjwGLxtAWtvTQ15cNi25IxW01xmgRHGpL+4iUFU+8
Nk+A0ge6DH6FSYtFlKffD2dVk6Wj+xlI63TdoCriLWv+yrPJkchb0UeXw3Rfbn7X4IZcqxHYajK4
vSxspV+gsx22Y+gbb3qKQPAKvztDue6goPq02tBWcqutS6w3p7WCelvB+bqOlJmOO/sCH2B5ay0M
XGOwe5VyYbW9JCBGeQauwdu7m6lbRUOZrcOot+7n0fWuNWmaewb3A9IbFAdJWIBbMZfHbC74iV+E
FQKo9bv49KHRnp5PHaQAcJvwMH5SZspoAZ8qph6CVgQwE4XykWGxUBghu3HwrcZmrP/BIrTL4iOv
HdYWGuD2asf5EP0iYm2TnXIYcBfgLp+DVIGbLQxsPxdsUKQax5eW9Aksb2epZdvBd8xAVNmRexR8
98YVEalLW+4j0vLHgYZJi2d9py5v4M4LmGRIeEaEjYQKWhgKzlCAWWFPA40bGIWxDyP+00tR+iXZ
oV0Ovd3uBnlKy+q4m6CFGjAoY3t+tirG/js3j75QRx6o47mQDlxOu+41BRcXe9cmJncSxUoCVTTl
SVr3a0m5jOTbx6Llw/1QEgUkfP6HAdSqJ+tiWvEOBYEf8ITJEI4Ly9EyMyQ/glWL7qiSpC+j3L3L
CbzRuraMomn5sku5FZmyJGExXrVHEaR2A63Umbtc0Og9qWHOpVK0uNjIEszzx+m7MjUsyCMMUilU
tE91wd/mfVf5BNGJ/FOtkeIHzUzQ0qdXb8qrK4qzxUnZxHrekNL9g6bUishHWqTyubVzy1zAslb6
wHpqURpbY+jiKnnC9bvcqCyLuiateYZbNSN+bXcZZpfDxzqK91FWzkPM68ey1szDSW3akocc/wBE
5FHtU4gcoPCksz+zFDqJOOgYHHHsSyzAOptCqBaR9OJrD8FcgWEXjxHWmQzoMqP+K03W9oGNlNlw
glK0EZHyAAFvjxoxp+nlUtVNwrHPgz8c1MLDV0IvPFktLP0k/ph5SN6jch+MNByExoDvFLgwbosi
D4/mEp7MHiDM2KYxcIadpaFIGTiSXTsjYhvDH0+kRqdBAYt48tDH5btVncNwJwrrTyZouY0Dd78E
cwaFE87DntboeAGcDNDYCSWsjxJOFGPyR3+arVtINrmHBwG6VEQ2h3iLx4/ushhRyEFcfRdAPqC+
/i23eSxWoQ4ejv2M10IKc3aGijZnaqJnJkZu8RlFkLj5jk4oUBcs2O0T4YZjAbR2TOzEJn4BMV1T
DSZfPdAyHyHQkHf7xPd9M7C/s9iywOA6N0rLurrrHkbl1nAZNJv5G9iEJU1OfE1yNbZwge5G1C2O
9A5OEp4jOIH2S3lkmOrc6PJcYg/tHUw0cQ7HE0Lq9lQ/ra9DkumIUp++dIGk920ksRGqSEu0M1dJ
R+UUfzch9NO8poybzZHJYTOdOsj8urLuALsq1JXHyv72QJtMGvLtZfNTJN+U7GEUG3iK4sShoobY
CfO5S/Y40/nTBxlU+kz3QvjN+B44x2JMr8c0BqdJhmBOMA5mdKH2lY37bJYKqDxzj1/vxiChFReX
LO6u8VJvU4P+wFwOYaYx5pnFS7C77fkaAz4BdA/bd8dSoo/QQAIyY+4Gl07p7wed1LbmmYzpqeEQ
1MO8V6QpvEsxsu1NIoj6tHcy35nhnd5No9cUuUbBx0NliW9afWfM7/ePYs/rqMkc0HKV21ZaDapU
m/uLxnMQ0dmkudp52OwDG81hRMjz/pEU4nyVoDouIU6g7UqWd1CiN6wmsKpwYxECrwL2xz9qGr7J
Cc1upKilaTf3Dz2POtFeo/DjVWkFn6FNMvdtzLivWKS1eyzHzt0Ej1Mhy33iBBWJ+kMMP587E7wR
dkRwXR2w6IUFzz5ph5iu4t52OijYn+EnGnRPMD6e29VFFl3hJQUm9Pwla1gQW8Q1veUOOHEFy4lN
NzGhCBLZ3VNr1DssRipVeg7PKINsGFOJxoVsleHdQp2bn2RZvLeVRqrnDj6ufEKfBmrFRrYrTHoI
L0OZRS6tMXrghM6N/ew9nwY8SgtK1VEJw5zXSQCDHNEceW7XCDJ9Y28w6hIvbCHqZBcnQPPqsAmU
appoEJXywwCq9bOEyF/dnuKtFhM7B7n87HiU90385M6tjB30pZFfT1+9L7KezFBPj4xtDIKXN0Lp
LU58XvUXexwn4aoZRo1uRaUegDq90sJiijX/0cpZBiLImgBDp1OOVZ6lQF0ZG+gfJNwIiXzMhTMf
lRNl7s7msk50bGXCvjtTiOJBQ4k/8pZYyYykZDuTRMc/hLqXVvxcghJzGGsf4kc1qfIAhsbqO7e7
lmX6K+lYrtaVuO+n1NhSLzuLWvHTmd/I44P/u1GMo87PnnED6fV3QSaTebgvxPxT7qtq5SdG6OST
Y30mUL7bvIHhyEDQ23WTK0eia/AtjiHk6dMRKavttcLn+b2zlaNH1WxvL2KM/HaN+V0U6hoSzj0T
u27WPFJ9bzc2xDduZ2eev0c4ZxYCL/umU+Amd8cOAdvrF2L1vFcA+LGH8rDcPOYQfzEu/BvpMDex
zzzp1vq2ieTVX+0me5DhMkrmoE7KPJTktqNROsrnHaag5dLeuGNB9v1Wiw9kWc+OXrG30D/9ufd9
/T8G7xZdhTiaxA/n0dVIrS6aBbusNWPA0A3hgcpH+Y0GnUzgoL5qAAFNsD8+noml3SU9QrQXY/PD
ziwUhewrZTXdwerIP+huIdT+lQ46CD4H4lPSHfPg+jGXLySO80GutmIAmg6LW3+pLhhaAaevO/PN
vwF9JUW79cqJZa6PSTJdsEu7dorvMb3wgVYKiyqyOBiC8hb9uxKbJMDWIjzuqd+o9eWGV0NfafDB
KBJbYLehz9i6M2EXKw7fYeSvpgzyw9gJT8IPY1mc9msJl1Q5f4aDEV+vWFJvz8LVNJNxcBmJ8UGI
Ob8mCSGoICwnBEbO1xWNhz6/Hkt+qWPqxLe6t/X/mH73U+8yNxfakWfCMfGZXNJMaRBR6oOcFXyc
A8OSMKTQTrx30UGIk8/gd+sv0/+WQd2zSrrsr28aOWGhAcTuYTuR736O0l3If9lhlu3JHx8erp+t
cRCniPz3+I/HMeuC1pRDAyC7FRf3rpPxWV8vtcKlHAcj9HLCAJaaaAePQvei2i53pCFCuNnz/YbC
pFE0IvsMFYD82r/qAADLU+6NpTB3gBWuSJ7jCVV/uBJr2nRhqoXdYXD/rP/KcsYDWDfZnjMC0Wes
mOQ4qmT344BBAh5S0TSTTNNOuUHM1AXxhC1UWdGurHOnDCHmi2UXAHxug5Ug77+/zEl+/1dPjGrG
4SkYSSK9Qe2QdmVZ9hfwRd0nqIqD/kMYaClRcOJ9zc8enHgblQJSYo/IktJ3cueToT/KU6c2mAIp
mTwh2rdFIn3GSnsXyeub55UEmDnE3WxflInC/Uq6WJsGMAJzKjSujjcz4dGQgxwCbu4ZULCmLIKU
0EPVwnRqaFFObW4hiOaC3DsIt07tCbxn8sZIrGBoojlbC6RAgtfx0Dcv7OnV7MoICy4VjXyIYpnw
qbjsC8Max3jTN+/FjDaI2Ex5z1ps82xKvvyBRpNWQKjD8SAB2v0GaQ3nAzPCuhaYgmOGcbCI9z7y
fLLc/ahi5L+Vfln8jeVgYSPuIVuCIXHHQigs+gkvmudQ1Jq7lVhfBoxZJJBga3anAsSbyjuKUlu2
q/IhRV3cAspQrMXHhCvYH7zniPqc1vaoDppMt6wwRI0qeCJo+F9fqxDDW9/hcoWI3J1Nh1qakcJ9
cBQFe9ckTPltvJVhDDzGoTsDgMU4oiLfKW4x/kD8Vo5nh2DHX7CIZ3hJ98+OX/8VCYig5YeMDup2
RnAZ9n6ezuzg+CFh4NpWF+fIJm6vKtAlt/iw0kcQLxugPFQhpz3+Ke9Et6Ruxy1aqzadyFFYSSJe
emCVSwR8YhoqRodNxYF3VfjXqkFZ4FbQ/VQXt0PU5dpJlj69AXuVRVtzCf5ly62hiEoQnu0pZ4kF
8T2xzb5EQI0yXhLfbaM4JgrLr3afxdARmbWrgh/v+6c0NAVz6ca740oDJCUSFZIwigLBAkGsR8mm
1cILcPr6xycW1K3ucVJgbpz6YOB7YNvzo6yzWkFg9HfzZz4GjO9xC0E7tbxm9keB0Lp3/R+y1VjY
vcOICgL8bc5+eNcckYqa4FqRA8z93h8nhrsYP/DyMNBXp4ZUsEfwgNbn5Sj7yB+KJLsvyAkZdXSR
QsjZUtFqxTJZxZVju45wpSHAP8CVAQaJagpFqlKk0Dd4zryS268EELRyMm/xlmCqjV4WHyi8Z7df
2AedWiIM31PXKMghkX6McgT6WJJJsmMgpIDZDvznHoprN1BI0Qr+ZfWUjA3JL35S+CvEiEc6HTEZ
gq6D6OinqtF1w97uROSNRY+1zkfciF24p7rQEkZTBp50D8K648Yw6wUL3/y1D/JkTt4ifMUHs6ym
W2rdUmQjyog4yxRcoBbSWc5V4nja17rxyiFCrUbOyEYsudEZJXV+2CEvw3YxrUv1XKr/zdBj7UyG
xJQzAebAWvk+Y+mWyA+0+CAE6/MGUL3pw/tCNWbyh5ILK8e/K2rL2SAUGY9Vs1u2lkL8pAk6NyBI
vAInHr1nh1USOn0WZprm2KcIRCuUshKvcYftqaDBzK87G88HMOs2fAYesF6y/RF232ZUMTB5uDOh
sdsUCjzUfGJ9e7Xjov1C4+po8Kc1Oyl9bTFono4qltDG2C1ezYRvzG4HOdGFmgVyjAR1npYZFx//
dUjX6XvGSi8ACGfm59LfwJgjOXC/nzJQx8r9+qTfUH0ZtVBoiuuSjtV/dsToiCLJpcNLy/eLqnYp
VkXKJeik800RB5BKZw/I4ytN3XZ24mGeeITwsERKaEjBHXZYPFcpLU+IgU6kSydrrdTEH7JRjwOE
15SxA0teHiABYbRmUD0GndVrGo0OHlfyppxllN6IyGNAjdKAHiG9YOW++v0HTZI54NdG+qbCeVV3
MMMDNIe+e0hz9RT837EFa6AGR8oaNca1pVUNvCXX8tIhhWGPAxdxREsix3ZkxlB0sxeZ1Yq/Ln+h
4L5+SNdz90vYCeF1cswhQkN2OdmOxXkJ6kz5EguhzBEcqNm4W5P0RNAAHPObxUCbktAtvfdy+1/p
/rnht+6f9Z+7uvwrTT0NXcJauWFbu8i08AZrUAmiRQbNH/zC5TBvvqFDXMPTSMrgynGqaYZWtfaI
PIpiKwOGEgC5sTSJiUxg6Td7PBTpudvu6LeibAIPRjMK78PWzkcucEaoe7f+dM2TJ8T4J6ZL7ELR
by4+HhlNUO2XCD1WJU3tNWZ1pgpZp8kTT539Zl+C+vqj7Wmm36SE1NSm3Q3aCQCxb67V+oM/KHOy
e8yjXg1C0NWNn8Jar3kDtDBodnjnThvRbnEGEGifv4zu2D9skhbuh+YQGVcAVbNNUDqw0EP9/S4R
VtUrhLUP//rtUpjI37IpFNlvFwlr7/ZkrGiAMOGAj/F2vU7Do2e3Ytq22ix2DH5P0GOFE2pS951+
eYj/KC8GqP6J/JsQfXjL4VKyL2J48bxKR7IxXPeqnc27FoA8F0RhXC73gSol8nkSL+bfROpoOfOB
FVNjWDBsvcvnhbF7sALMfdpo/ati6f27yQ42DoLMuXUAWfmrg9gl9ju2965E+Qil68hnE4rKN1ju
cutnCpg3IrDdg+WRKjsZhN6FrK9wpdypPXdslKzoqe4t0Xgm7Wg2IOxh5MHK0yW4vL65Ebn+6J38
PWmYHteoulXLJcjTwuF6Iqzd4M8ECYoKD2tad7nfHm0odMxxVHKQAPzGUZq1Xnl9/yQ46a+zlqR8
YlR0PZnNbn60S8fnQVXoblIKRl+T6lG6wNASB8RO1IttCq29WEzQJyN06OV2VhIWWbakVEhh0qcA
zDmFyhvMGrr3Pcfr9bXuyi2Oa2D/nLypFypEiRb3KPUJ5n4891sw5zxNXD01kKSgw1/GwkRspQo7
wWwK4IPzpTPlo5WI1hmJD6j6F9bHOJJPG6cYzu3VXSkEQmFL4KMAxFuPRQ2ad3jfqdVNV7MAmv2p
AWJ7gJdM9y3L5tkiIPz9ffVz3w/W3spiS99nzDgX1MxUo5JNHfdlKefvjyXG0Y2gRML8RZWyFOIg
WiiIFegyHjQ45nZ2kY2vjntPAD5T/H+o70iPpPyxr3kJ0ErY7o73t3ZKQIXLGhINbZlThUOUzMTn
6TkddS48c2XVEvHqlD97EKujSyTlNYJ5Qt43PJJ6c6DJciZ7+cSWiuahmuRXlALkYkTdyXRHIbZn
AQVlgS31KDNOePVZ+fouhmJpWWCSBw36Pxwo1tjtODhaa745s7u3wO01310IyXf9FGkSvCp3sHNp
D0rjdAuRbwRAfEZY9Ig7st12dUcy2vdIzgL1lvgfplEcJHzbW9zmX/OZ3kZwblX6TCNvp9ssM7q9
7/QpC1sOHiLDIdvxWkSo5Mql0FQ6bq2vH9f8Wk0EDQbLDj0yDYUNUWxq0x1P+7shICRjLycq0wkv
pkz5zOT44a+jSTNlPt4vuV0vlOvDgNz0iS+c+jiOHs1UqeAGFWpDjzYo9PwOsiU924AT46Z99dBB
6YPp/NDmbK2PT+MijaMZGlr77qDmAPyl43WGTSuCfgv2dxURN/Oaa5W4VP2wkRzLDa/FAmwQpih7
vxp2owEJd7DKlFS7+hKhU5s73JBf3FvPy6Edkxa1n09TuX4UNwLR9GzK+bcNxAwJwufDlP9OMzjQ
7X+yB/EvfQJ5dVtGupsDx6nEuHJEOdkaLe69/vLGXKQsg63pX8TA7s1QZUkB/IeZ9W+f114iw6Ir
GPFRvx5MFi/j2quSyO9s37J/GQdt4nRQtS24UL4bP3B9cOJ9u3IsL98BwJzRQf4BrWX67SvVmOrV
R6uBJlfrEvRKtNX3QvJ+R+EUXgxPtLk3oeCqaiL9Fyxnoli+Fa6TtPj5bLXljgmyQ1c7MArnzrWA
charjhlY6EeOZB48Mp2fGFp4rFklIVUeC9McXpaBkD8HCrGG6iS5FucwsmEXOa9Vmn8Eq9+KMzET
Fc998usMDgWEB4uiffBS33UjArZ99KRjfAARKbEBqjW86QXfM2D4DylsrSaHE6NOoJJ9cRO7+P7Z
tbiFM9X3WaLpge1sAZG4aZlYer/hnZUxS3whye0P35aEZEk1UpYhTuAOW8XGXoL6amMUEmQM+Eui
w5nxrpmyCp5su4A3xX9HlzJ3WS66JVLSjfomehXSjN01uuo9S6pgzaomsUj9KG2xrt+bMlODYQ8y
BcG2nYrMZdvFfLy+EGQzNl1+XVPl2r5ikrXqu2B34ZPWdNbMnYc2jQ9olPxQ/Dlhe1lT8miKaR80
5UGIH4fdToR5Kdun0OS/yPQ2n9e8/JCgn/9bWuPngzRl+Cu8ohqxCYFSTDtKZ/MUEAJlnF/Ga9fl
q67uinlNPbHkg6ZAojOPIgm5GypdB/wHxPkMy/m8EYJYPPQfyfNHZiJPntvs+4MoLaQXzQmd9dCn
hP3FFUG4vm/ozsGQnkY8mm6AuJUuq5I55SWBeZR/9dwO4XiyWcuqtTIZph2JmhEZ9IiMoC6FH3e8
E5L7VxIOSucv0ColBJJJ7DpENlQf9w0PVRVYGHL2YvaMpdtiNx613bo1LSuGenm5OEd2spuD8CPl
TUsvClltG5pOL2bPUEyS7tm8D/pk0PbRzyA/kYV/icfoOPrz1Y+juf1+UnG3N8X3yml2YFNhDtC+
Ut73G4FvZj7tyn77hQPxhp9qsO2oLRhIkNgolSAphyeVWYPBiVekzC3a1QvFqn0/HHZydWGVjf9k
hlKNFIAdJ/orX57kXUoIYJegbQqjFT2UMt0UzQKAqi3vBuXsJbJdgvZf++3s90FdGcRbDamnPu5V
KggOs8agvNcKwISktWe1v5k7zja0AlBZIGRwRl+lQKXGOq5VgWufyeismMfUG8tlYJBe6Xmp0Wxg
ogCwmFz9IyEnwAdfoHpQl3s4tKy3kLNvAVwR8Xqm4fLf4+I6Z3S3rJK22kD4cckMRdGf9BT/Q6QY
N/A6Gh4kA745ljAIZhTHRdh6lOaDapHPRw6megJKMjm/K1hI7VVkicpBab4RJIyck0CJdi0+8E37
0iyR7Q+sNscR07TPLgdq355PDb4/+nHxHLRB+kBSbqjxBtgZtmAkid6AtJN/NODOMicUKXGYBQT/
05FsTyQ8uMITgvpOve10+EQQUHbk0ODQ+m38EAv49yZkC7qEUAR6wzks+Hri+fj4ygd9iYirAKJp
/eMm2gfge9RyNkPeEmVaNs4Rya1P7cafRuYAVl5zsmDv5g051nfcluQ0NaUEmLsUX8sbqg+71c/R
jDVsdjHa/83rgjIIHKdw5yPGKHeP70pNYnAgWSrBsb4h1Vd19IYbhydotpidUqmgZmMSH+R6QZ3E
ZIzAa5wj+EzHzmSgtNubPr5fkJHfK3tSbq+sv7vmNhvxtJNGzw9rndvHkYgF2+RazpB4ABeziq1i
NctbpmaKyuxSvFXnUboNi8ja0PYTqhFsG2X6mFoE9kSJLOQTbfMwHQRKQQey7AByOngaEPgFiA5n
DbfbcGxnZmlLjwq0U60GLgg0o3JLo16RNWwAK4LUjsImn8OSCUcg3b3iIKL+2Pd57/kfBXaeHr4w
7/dQ75dy8VKrR5riQq+bxnB760RloV7UwXz5bGVBXvu1zlNuEsGHXcJMlpY5o/OgL8jaD8Y6EgjT
+KHK3QqWYWME8hNMXhZ2AvtfBTzEgubwFGXPyPdbtpunmPfBmTtPE1x5kpl0U96hKJA4akNAsGOU
ReY72DOBYIX8PYvcvUVKsxi/yYjdL1D/1RW/FpnI5GXkNn2muIVt/3AcClSvrCFrknNk8Uy87NDV
7ygO0Lxm3Iw9J3W5CNCjCo5U+8R9PYTjmH1xu2HwR4TKI7J6WclyJAiroSq26yLxei52Tvzeng2O
qWS72is/gl5p1EI1m8icRaRRnPjt5AIGDnKphdExhDsVL8fodF7fwnuc6xJKwThd8xqsL8GHqYYJ
v4cX6GuOB4nnAFTCUDxNaFHXQWohUq8gpkHn+cd5sSprHdVJaCP7TuKnP1mfLmLzhrCwLxFe6PTD
Dl6VtpAVJkSCMj2nRyTcPyZi2JP453NePcL7BgrRhSmVaqO3qwOE1mTc66J5vutXPh71Q5tqj7p2
XoJ5/9+EsUwqMivLrEGtLyScFGOvU0LRs5/Dpd785e7idElloOBRkyyz+BUFHIfOaxWcjg9QY7KM
ZMq4aXH7zDIqzVC2tLJdXbplqleNFiTevXEIEnr6SjcrGuGpUm6EZOLG3MD+VH4Z06rvHV2ya94O
9Qy1IyQ3eXavShzEFBsGhgblaQfleDhAxGdn3ZnXfIVrxigAeeazVSJmYEhx/zOYSh65j1rDNSzS
Tb8+cgFNl20CnkoFV0UcW8FYjO6aVJWqn+NmiPHmVqtnKn7JY2NSUMdOaS5MOlDGMJIp/3RRZdCh
YVfv1S8TZpUpZsqru06fCJhmSKTUSM+cN2SIFhISj9Al5wj0h550kbW/hQ4cdTwQ7cIs7r13j35C
CXMe2KYh2O3bwMiAjTB83HhOFU0S+ikjFWK7LTiR8GWzBG7QqrWvrFm+v7IVWdy46R139e9WyuOy
La0VKZFlWc9FHLmhCXEx9LXDL/tgvK+hR4bGc/rSRrbvm3wsW5L0B2GmFbIGHcgBThP6vh15nipc
9xzFt6l4UpwGTFSFwN5lt/gMXnhmJy+cLTVJAqynmX/F4RiKt5rZnoRhQQJXbSoCxZo5/KJnZLcb
dNp5w1D6agHBJB+62nfyBefN3at9/4NNzAmlL0aDpNuqrhBjePaYKwCKS/y6cpw20fCQfW2Y1bT2
MxC2GvxZVxO+0lyrUSI5OCfhPF5zKRyfdM39jygEJAbTMdXJ9lIqd3kfowwoqG88bKIY0nbO/3x9
dY9PjaYVCnXLM9PsKUSHf64FWpYmwHviWYiIJvkHyITSu2nEqBk5yQN0Al5K4DtBaodtMJWHC7s6
eAUiSwPL90BGG5LCMc7gE3JnIKRHoW0ARSKFoQhPZ1RmQPch9VQCX7C0rVdKK7oiO1fTH5fRSbzt
7obbYlZxcwH3rXyYRlgTVjo57UovSMB45zLZNmkQt6Vukv1bZ+O5mQ05eOUZv5IEKnpu3R0YnvhI
u8S2Cn+0Iw5g69OFqUoaoW8zVE860W7dHf3ig7CqwpLHl74bn57FctOXOSHwrjfbXL60xhlx566j
GjmsMkxlLpvEhrevjcP6VfSj+F50Ek3uKOz+PQl7zHbCl5igbukc5qghp/pfL3UAu7R/o152DF4s
BqJQZz2kTNBHvi45KmtOU5eOZL9CiE3F4k3LMATVVkX773JK6tqxB9Mx+fC0qiaqecljq4JAfN52
G6/G5VngBD0BoBQh2RBMZvhmTwU7HhA60Ej0jnXDN9e5Sljxdw1LpBtv3GzR4wi/NKyOsEShOCMB
1eNsT2VNfOfxmgjAFZg0Oxoxrw7ppNLoraZt7gYlDTUSM8/3BV/rf48cq+r+G95q7dBoPBINI700
RRxYJmwdJm+gZs1eTEDpKng8FRnIEZp4RwcnFmjdmM+oDrW5QmfeMcnMfDsRIB0fnL5iKu6mpHDM
B562N0G+AC9V/6irbkFo6+mFfsy6nwf2+SA+AxHrLBJLuzRIbEjWDZ6ghqegndxcde2hMXN2jVZA
ug3AJPhwHCn6i8ew8G9/JYBTIt4MswJ7VzN8KlsxZtrtHvLHAM7QRNbUwCAG1kHS8+zc1wMGevJV
QYwLdZIw/UljkQY2s/FX11c1P7//AHxoHREhXi7QXja4mAeZQ+qloIhVdPVsrFx0YgnZAjqYGstL
/+4IHvC15fxVyqZjRQ/v3iZmk9x+XaOgySh74ZM0lXFdBzw+tRW56USaSDKZPw/vWbVteoCNPQQ9
vhNUa8btYiJ/XN1gd56l6fk4PFutnXfS7G4t81Q7lq90Z80BsIc+LyS8+eJ5wmnE57ITU5dCBcQX
nuJuwNqMp009wYPAlBJ/yuf5qFQwfKhAlLuU9cHAk2dwo8pV+SxB0a6heC5mBV2yhdOMsJsc38Gt
yU/1fXpdI4kDMedcJKiMwR7/FRtiKkpBjX6zkX67sInaocle4t47Ak8iHvJtjO0fyU7tTlVIZIui
I9x5w0xzYvLB51OWfwSO2tC9CiG6jZto/8nv9E797KcrEXZiqiVcUYCI0fMDTLpfCc1HgljqD1GS
OHCJE4jK1NCOerB6ixbZZegrriu2TNnGFoGiU6h4U6blxTW6YYzEjNrF5CRgScv80p3dVLgG9WSt
FJdvmqchZYGKKcvgzMiCRWhNWce2Ovq3mNov2s+Q7H0nDIbkCyvbe5cen6IRRYBSZs64Imcdrb5D
QAf8udX8sBnmjaqGDpfswamXDXj9V3c8Ti27laZ9YYrki3Xu+mBrw3FDodin9WdOQ4qwQ2bGRv/c
4jwjBh5t/7uPPcqasLegRTFZAG8CZ4M9C93p2s70s/4YdoSIvrgtm2ntqN3B5RDoFkNiKATifi2K
JIOlEkx0xLV2JonwGOKpIxApPIi+7PQSb2298ZqReH1LE+eOJKM55fcyyoj2N5qKVTmYTlPi2dgK
gAju1f28uC1FG0aMZxI5Xqdz8ytAw/AqV2bOB3/lIKf4B6hOlgv/jnwvTo5zX0j+jkaABmpcuXnG
e2HO/IGZaKyfr4IPd4+pvBE+bzzXCgCSRtpgONIxbnC1w7B/XAvq3pyE7OTFqmXyLOJXA0GoJBDD
sxYKdsl3aySz8Uc2xheL+Nu1ImtYHoyRjiBkNZ2fANsQawd1nO2SVJRsXg8ncKMdnwPMJPcex/No
HYDdtH/dq/LWxDyBwrM1OmqFfs/9rszhSWLpok15SkDineUjArU/MB1zmRIVTzJR1kRIPduO/usS
BDN0Jd+HDecBmlzerr1TfOHmyb98eaULtvGPIP+KxLjX7rtOFf7J+AIrQKZTf5Rm27d/+CoVZdU+
ZTLepkRkHITern1C9XEbOlnNwVKOYKThNlQ1y2bBWp5I7WLub4aoN4rk2B+3Bku7ppk+aW62YVQr
fp+x+K6Jo3MZcOqh8Lw7iLnqzTOXkq5J5kuWIsqiEyDecABdlLicBZaPBvZhW/8FQR6cSOT8s08L
uHGTUyUCmdrJV6SksrrNJJhGMEcueUVRKHoif51XhUedH48Ayb8YXkWnwugkGoWe5wSRfE6+H+pE
eKku4f4Loi/gqh7L9s3cKjjPJUYiuSF4lZvk3RzbfUDPCF67F2+EeoTXkDIomJnAzXidW94MukNK
D4C6GU3otYPe/hZoRtjbG2hfX2H0wCQADVzu22BD5IA2f/ibQMDoiVmJDxaBAahJmDHkx9dJEY/+
wXBLS0MxUQSe7w7jIHaXFRA7JLrjtbTtPO+q1LiudEB+beAXDpBQ9FWNZZRE+/vgWjMqus3unYAv
2VjaE0cAiMPTiJM2AJ1r8Ln0VfDu7KxQhsoXsCsXTiHiK+6K1MQ8NnHBIfW7qsFDS6Ja4msDQV8Y
mM3p4KifWYXhe48K36PMNm7kAmY43sGKEhu8R1bSNp7944UPNxYydn4wuLi3qbMybAAn6yL8qGJp
yTrqNHA3zVyDynWRcd3Z9i5rT2/S2um99I9JAQqBSzh87697whzDZpSEcrt31M7U7rVFRpIy9aP0
iDR5IebqCfzSD7wuJRoU4XiqF4P8uOdbHvUKF06lBZOYdHMXAoJ75HUxD+ixaJ5r76wb+N7GwAI0
ctZer1cJwbs0Bot1AFasQ+unvHhbJQvVtgcoaDX6tVlEY4hu1IKbWwAoR0xbzhjLBNl1hfhaJcp4
P/Td99hOu17WjT9sCKigQurj0KpvzFSovsR+Zk2KwvP4YBTnbvuHdW92RcCPacKs0wNbur3WtfqJ
2rKggh8JPfjR9wYMRYXe9ZP8xDspvXlTvUf1J9zgxR4mtucnudNL9mqyqBM0ElZw7hZjBun04aK/
+UaBzoaSPtNsWS1E+0F6gI9s26W8TmeSWwKwcvjEKc1Nmzz8yVSFhp1HpwiIOTw+YCPgvnfXIQ3D
0o1nFBOVvUeWSIAnxHONaDj8wVGxXqwh5rUcwfmfNCqHIlp261BQfwXlLwn2geQ8lEVB+OsgJScg
GfTr67M10zSQ6zFsS6XWTGKSoFpPhOlQf7wb7foFMfKrk6BRtTi7k2GNU7ie7xXatWgh/jkxw7hm
bHIn/34sEJ+V3VY0v24AP2FeZJrQVTX5IUi0aBGy/6dERzL2vBvze2HJpd+a/0Y12IowLREWkuaY
nmKGhM1+PMTiTicT3+Kr2tkYM90Au6LVlisphZXfRCjSuYmZm2HKD5+sHepMxq2kyfQPu1/wK8UE
qk972QTslmvrfXIP+x7g/U3OwgauRWGGm6txZRzoKRIdttMnZ0mJs0aCly/cqpcU4PeR+xnMPITb
ebtWspcULfgevMm+8h2IRC+xO1isDycR9C7IqW6vU4sNikOw4SxEv5O///0JYyQiyby+ibxjpCoP
zxjzcgnvs3ABNgjtTBF5rwxoOjjkuLJ8umIeVlu9URvpoGfA8pk/eiAjJkhhSx2P0TPTyzgynRVs
Xp+jXA+jGgtKXeqr+EOfnlFCi8DBTSpOYFAUkQgjMwO7v+lcpRQ5L9y0czsgPK9WhkevuKPMrKKh
YOiHZK9Ntce2hZfernq69CXO8AdiZ6m2ZeUUaO9J3u8kmGIzYS7iiaGhYQqClb/4ujS9p74S+IK7
M/2IXolhzwC00Wl82PGEVJPSEYrJ4m+gSmEy0Kpg0eHUmsotihyOlKhU5PtIMOPoO6xsaLzYwIk3
wgteAbYEBIKvVmSdm3xc8Ppfq10hTF/M5E75mJttp/HYbOCGrv0pU2Z61vNogkZnZeutCzsbso/w
f7rEueiR6QhDndRzAVbq3bw/dqmalhbNA5g7NVts1FRbyR9DlqufTnMyHdVnOsZdFnIfEobf+F4y
i66oYZGX9QxHu48wNAov+AbnZqEZZAwZQaws1sIZtOaf2LdBywtUoi4wM1mpybjMLH07ao22c1+2
QF5tm5rLLKZ3Ll7/PvqrxfweGxetoVxyPeU5J2Abv0FjqNTDUFy8ynYLZWNDVjaVfyyCDMMscSvF
AeyzE51/rEVd9rf2MDgXzyrCCEoYtd0o4+lYrCot1b300LfOw1D21bXkYIKUCEel4FRrwXXcAylB
egJVnfcubyoSEqRdtgsgRBM1EouM9rZRAFJi+HVE0kz1NFfT2XxVGodMb0a8QS4jKwknXTqD8ADg
WetFIKsBNubTAj2oBlFcYxW0hTGYQ7rUzCh9tg4VCLkj/eUSsDOdgq3MQg8sYI/D1e9s/GZqCm2U
0Gqc0TfTjXP8U+nOgib7uB4ID0Ad5Pcy1UyHUThoJ0yTOffzelYEbF75UGgDvoazeJlJr+o4ZAz4
1cwViUrmXmse4OJFZHwJ8MYAvMWb4qYAZdD1PATJqVOzjh0VGQn7o96iIIqGjHvmjU2UiTu+mYd9
SeWXD8rGbWGOboCI6o35kxCgzrXsFdvCi+B7Wef6vZXTIEcOvnLQecqn7wfNdlpq47m3sacNo+Wm
laUJuTsFA690ALUiv06IhDzrUZuRJg/aNuSN5d8XfoWggq8tFWpxQs10wYfdincIv2ihlr+VxpRd
iuU2D3wEgpOWEMK4lgpSM3IKMcIdTyRt2B9bouhGxPSyHesxZas/yMIt6nuwpTNkbqTGKRXK1dKq
ustGADhbjqDB/NzpzO73qJyr5JlFDd4CKVIVJrG9kltq/6PnaYfjoiCIqaU1n3QcmVX9RpM9Ky8O
jRKF7NYg0khURfgO7Ym4lrXAYww8rJ4zMkwsZ7VY2MNNbsCOuSMC5mCx2dgckTzMnMLOJNNPn6MV
7Yyrr4VVP477uehYJsrBzfc7YuOwRfJlxeY2s+WGuJiXDJxADYtFefDrYKsq309bNdpRjgRgf1M4
1dnOpZpZDFEjZBUf9VaIOyeXt2vbTSdrOaerMNCpTdTsx3B7gxFwtuVtX2sWkvf+IRTlWQdFjhPD
Igx/N1Gmk0DozzhXQZLfmh4L6AuEiszrtRMgTF8QDY4TFjxQ4juRzCK/TOKqqklYT6UPGCIXkP3l
jF7W8K10zM/hjsybOavMHnFRTMKHtq0Udotkf7ZSdSYuT015usTVAwVt7n9R1FXkiTVIxH11gOcr
diN0THzTEPd2cG19/Y7xkugZhZ0rB3gEtCYG5CrAE8/NFmDqunu2sjVxa2Mx+IZ7AIwfs77cDI/+
+wXvYmDHK9xDfTnkprway7hvmWoVQVXuYeYY02CS9MVXlBn/KFv1P3F+Y8h1jC9rQbYZxYFRW9s/
x+RnuouYRsPi5paN9XZmq1GtLM2Ji36b1lDDOuLIfky68nLCSqVUYFqITP3HWyYRVyE/wICoZDcE
oHpN02QvTf9H1uMRz0QqiZHUP3wdhTpErqNlVqiAaFHCKDJmcqDhyrPMfrcej0PqFxWTCgJpy4mU
iN0y0G9sKb9ogWtDRad8zSiARPzVz3XJWM09/9mTd6Xg8rnbddgJwFlDZDtrKJQC0zDjH0lzSZis
e246pcpN3pxPy34RgvgVe6i6xtw8EcT8AzPHjmOcozou5AbDE6WyvQfAlDDouHHStPkWaFwA9xom
sYGmaFB93l3r/F26Wppd+CuToQRn8fQ7zsVmG4YBdBrZVstSg4vnsVc0IQlyPIryqXP+bgp5p3DL
PKrcIWvlodI1HiaWjZCoIz03zh4pcJ74B8EG5RZJmzPNC7HbIzW6L+iKZOhE/6cyWJDayrzVsdZR
BnNFqQwavHA5ZSKEtv+QwuNJcAoVBnr6Sxve3Fu6/4sLDI0aHIzZsJzfjMENOmY8TxrEO/LTLXIy
1sc1gVozh8qTJjEdmU42f2Dn0CoQpLLeRsv83L2IlxL/tfsZledQjxiHliP/ZMSWpHMcMmh6O1zH
Fkv3YWPUCNvKWzzKnRUqgloa8cknBUumgNKRGQRUqaFmwCIRukXeBGY4pZlSCndzXMAK1qnx2GM0
3re08IEgjvtp6WpAxw5k8DdVSx5ClZCM+jCSYJIsdu40W3V+2cXAvuRNcJTe9d2Fr38p4Eh5UA/B
+wbZMo/xGrLbfM2Y5pbDdn8MF7FbNWom0k+M8ejNHpwwlNK9ahn+1JJWgvJZFwE+C2asRgCc45at
u6T6IHsc922DBIzSdMuxXEUYNpHNPsuRLY/qHHNFCRChwLK/ThDj0Wqr5GaNV3gYSuAupT3F8FQ/
rjsbbv2ttzdMDWT0YIHdQOUurKjAX5dqAVxuan4LxLb/dD3wZvY3hU931LMbdQb6AElFrVALpnzd
NapWDXp1+DCupudOyT+dc5CXad1xLUPZzrs83XV706/PuEXwhQbmbZyBDNvaZ5IA/lKl1z/aie4j
T9s7LCp8u6kmW3nxNKLVTWeS7psbBu0hnT52eXzSoF575N9n8RLE3UumoPTsYOJoWvqBKxcApjUn
L6ucBeAVy8CBqpuUZP5Tc/AHTHDcc0xyzMu9dIuwaveo73nAR2TVaSHyEphnOFqCEliJN5Tnt4Gj
r/+Q2KSgU8UiQSxhohiuba10MNPw4Q2PHOgqU6KI0Pj66RrRBUPqXmquTVqu+B1WT1yLNgQMPRbG
T7a+ATP2OFx/uruG24v43tAHpLdFcEHkz5GLIhjO11D2wbM1+pJ7NQOq30GO0B2yhcB+rw9JX7XQ
ZGZfI3GAEG9LrJPbQwLEbf5b+n36PUqJo8Ug4JksgHL1C9BSgpfsgF2pJfwI24XX1sOrI4UhmRrr
eHpCPYIaiDV7rSfv4G0QvMn7cqYsd9TFhfqKnKadSVyD0ts2utLJnjurC7e2IZLKupjQjPM+XD2h
uc+CB+IvbXUXRHdtaKxRnEMMcEj2/8EqfG6InqPrk/N2xjKflJlH+2dLhfC6rpzlvCSBChPHCiYi
vQhZ4wx9SkZN7ijMAmXV8p47ffpyRAo/1iU0kjR6VqKT5Jeiwm4/gtEuIPvEdDq5xbUu6bLK6U3E
oTkVYHpsJBINPHAncxw/IOPKV2ZpdC4OhkS082GL9vMWdPRTGeh+qCHYyxzznKb+7dS6LeSVdCin
Ugm6ziPp1LuOdReDrrxyt34PtBcQUojG9hRE6jiCP+Ey7FSEqynpEGi2Tagke3T/EnAtc/NsdibC
kYrQd0rZaJHJBZH6ZFJtvPy6IIaujLnG+OdcLBIkE6gw7TLRKcd8ObNfcqgtgiCfzg/GE8jW3ulm
njXZNkoEKMHiM1ZTYV1Lt8fLIvO1FtrexjGjGVgohOKb+xpRG24J9J/5F7rza9y4ismwsQ1n2oxL
3VQryqh+gMm+fDSts+0EsvRag89fBH9vj7VHmsvhnZWI4nBPFtu0zVdUZmTgTsWbRRqTlOL5c/5Q
gvLeP+HC9CWS+oA55Ap+57SmIopYBxzlvGjeCw2UqRqGleWY9DTRwehPEchU0XPMFxoAvqsEqcpX
eHGnqa9N6le9gnmJXdb58YB6LdC4R46lgoFB7Ced78TlGKwANp5tnSwqDyN86IWxTvW5EDeYoMES
8lm6pqz+Z70a8LvwoywQDCvC/d5SlPSZUE2U0wts1InpN0QnCiwvDHX65xWDVuVBAu7uTlHcPK3c
6BEtQ55Sbz4xvgsGBgdvQF9rbZwBVYMdw73ARQ7B9iDTMCLcUVSz9FJ/FqJLTJL+cA/QuIuvtqb+
DXyJLIys7ueUGrsH+ksXfF++ROEgAO6B0yPng9fVaWNew64Z5bEkyFq+6tGLUWKrw/J398+hgf9g
DtEWewBmUMGujYqBpR8LwUwqA+aupHtz6IiVx2zWJejYD+HFig94H96240UV0TTgM6VyyLYxi/BY
9geEsuwfSlQpvQL/NMl0eI1oeoWbM/J0R8YSiWMIXf83DRxsplSe7iYfRiN9L5i73QfFoDn6Iqm6
o2Uqwir1XDmO6fxVUNZmGmq6Qu+xoHoXLgiAElNivy42jC9kBdHEtf5bl8MG+Ku/7z6k+KMYZwQN
3N+DAr+Y+fMXRQQP3dsa7N9RV9wFGqOzzIhPgmTwAYdiY3GSw14uEP7oZn5V6/GWpSzPv9dvfjbr
ZG4MczeaUyvcDlj968dQ87XJ9bnvpnIi1x+DtHYTw6R7jr+jli3GtnYfZWuOfsv0dO3S5QUAucXk
/+CN8bSu/PcOq1pqxCwLxPbLR55Hi6XBTB/H82NFitOvzetbSyQxI0XWSc9Sl6TJNeUnGU8NkKBP
hoEOJUmjuFRftZoK57zSOfPm5w6PEDbRpRcPIOwc6CaUrofBKdQjlKxbxusjoS5DTkapbuWBfL74
6zd+smtzk6f8cw6LORSMcemISzqpMoTGbCUrJng087Aklr1LyJkYdRdfDnTvnHEum+UCweBUT/xc
PQtkmwnxl+4znDoVOsSKqvmEtWm/vQt6PUv84FvnxAypPe2pkR3hAp2Zv18TpuPJvgSbB09hoVU0
A4veE4J1jcNLGn/N2sM6ET09fJ/V9VcUBdP2FoJVjYATLbStlVRSXM7x3+J8T2cm6QtoYEROkmUI
qt6hoovvxW6/rnkBzYfYD1R4qhhbPqyVFQDJkuLptUl5ChCcHhkrzvpEkkwrDpQ1VQUtl+YMjXmB
6TBK+P3E164RNCJpu48CVDcoOy/+X5IjD72SK0nJ0wkJ2JzGSXvyTp75hSR7mV4dPxGVpojS3whX
ECUbTiYl4GSXUZeayJtCpdn7AJHMhyFRqyTqLvhCamAhOYXdNKfeZrQ6fxJIZ+FjFCYAOEc12+cJ
mvm/gOqz5MrFMvlQfdF+XPkQMn5sS4k4g0Dg0q9PvvhDsNyR+9MxR7TTP55LsgPog6Qto2yX9t1T
rfs6OWA8A3MDN1IdSLvbHymxKYjJrDNhlD+raOJoP2pCIp8fjZwWwShKCp5VarbB7qmmZCluWk3/
xms/0/DGg0tyzsFWgPeIhX9O2W+4wiWanNJhWPJLO/RZFFWhbDD6V5FkuS2ERykHyXbS0UIWaZip
smHAJ4lFLUc2ViniqhL1RGHWdhM78hcBEBjE3kXC07ORmRGQOY8DW1M8pvmK5OcmWY/RXJaiC3RN
dT8CAjKF9/dCLRzQndIkZZuWy/BbJxDeGBmefVnGvrCXSH8PkxzLonYhORhxcdAMFDNoH14Xjip4
7ycIk+PgPwMab0TaGc4cTfSl/PE9jlKrIMlZ31GJrc3oFEgIWe6/9X/+6jiDxGA9UTD0MJ1fJ5b5
lg7B5sNJEewHc+vcLl6P0s0JkIxMtnlr+NkyMgyOF7wqTy+OoF6/lvyw5NFqvwBtzuBWmb4wDd1a
4JpFZy2J76zfibUD1BdnrFl0eQNa9+ANKmv3wqOhLS+OItzHU+Tundsx6NzVxojqtSVd3fajkjP6
JTkBYfxD5ncVIE92keIEtJQFRgSty6jJFURT678RsPy7iR89TMIWpCc8/RLl5hdTv+glDFxxE9sw
Pb1pOirAYqvb/ijPAuayQuOhwalgerF0hG6TGsYxZ7KYkqRDxp0HTqHfOvPqiMahPXzqPIQ/xt1f
Q1LesjcuveeSK02YOn35WBpWkSitYGVm9t+EoecAODhvWFn0j/n2YRTmKqKwAuCiuSQT516e1kVl
kmVd262eRsV8PFSPSfqgppWWTosqHc1LW9GQ9kmCJw2wzH0PJWayTugRMcR72SjBACtF8xPL3LGm
pxMs0poThQGaUJi26/OBu1G7apIn2vPzT4eCfdai32k3DRHH2OY5p1VMNZRA5g8hvMthPstLw/KJ
pYintu1I6K7C/hMSkJua4mJL2kwPmXX/WV7jEeu5Glrg2bZW1PSgoYccjPqSJuaBUPUQ36IhKItU
DVLgCLjdWgDKKAXg/NgQ4IK3MJsmB33z+LSefkeCe/IJzTmP6UKoqqD+pyrEMAI5xZD3mmpL4BK+
0s8ONmpGaiQHj03nzgoQPFH3e/Ucv7BBanzmVgXuZJrIR8JVT9YEHys/aoFkJ9wdZCHHiZZHEk5x
R6dTMHpizkqn5wxD5EPQKZuo7boMCVd4hfN/5HwNEuF7Ro81uczURAX2M6XuACIOPQdyDvFSKtsA
Fwf9zEkH7TMYDVTk88uOfO68ixVhD1udRzxfnobrHQRQPEvBelCIlhDaTK3stOabo94wAeIdVOl8
jFst3oDmLHOIDORqEiTtrc/sQ5ncXYNTj9j7EomFBPCX/4RYETjDjoSWBJ3tWIy3/5SmyUy5R3GX
lUpNKG1t/LYQKHa/ew0h8sHmRkoRfCTPaHgb1iOesi52vxpzKL1Zqu9ffy1jEor4jXNDBnUuvS3v
Najf/DwqlhFK97sOdgC//dsJ6VHr+LDeYgksMSITG3ShGaJmBeyQmu3C3mJKKsflLcvn39i6fRTr
efMRF8+tut1HGhefaXb5xZuJApmQDS9zMCW8qVMt5iLCjye2MJWhRyFjHFIUlGG3xZ5+BH7UVMCf
41uldwjI/LLvGc4tdX3o+R2mX7w3RqiWN5MV57Ne3d0vq/5exs1i+Zob7OyyP5EaIaV1tKkl57KL
2AZ1QuHWQnFddKivG3uG3ed+pTdKR4Lnb5+3dQaBX90pksjSgwM6kfJdkzsn9U1aPQjMFRp1HeSz
tmnUWZVY2Oo1ubyfqNzFBupnZsdWGfRPFCinGv2QEsvWUGO4fMEcSP9uGOdgqKOB45Kz2w76FoJm
dcnLEayGJ6XpHzJgUymit1FuksaNeYdSYmbxK5Y6+o84M9f8zSBCmDpfPMA1LQ8pLeZ9BEEqstl1
HpuuSoLf2Ta6RdK9l13mXpNrXTZvXt1kAqDqCZIbTgPUDRwnNs+lE+dtw5JxEEgWQibtY+y4ZbD7
g96iZEtRH+XKcxltjgkOqJR6Z2GEvlDHrbjOaclFZ9X5bl2W6Il+ImgnSXnNH0e4pLq9yf/NN53g
1kEK8AU+bJOPOgFh6zTY+OnwFx56TrGj4onUWUy+hAvsr1s58izoroRmmJrEPKkJFPyzGK2k+oyY
DQ52pbsydxnE2sWoH9DkmvcOqblpeCIVXKzv1qgh7//hL9LZaloC09CQU2two9S9gn5QjwMhfFxK
4/ieq3rHoqC7cA6jbOwm/tcAXvl+tjdAnic1dhGiBN/ZsRqjMT1bpA7wn78DaNQ4GBs3JkB7L0R4
fbkst9FG0vtWtiULfS/oeS+zHIjBICqoOHpFnpLlJtWFvzRS6SYJPiaSzgWpbc85CI68ScdZZLpI
nuqPUYDtmCBULbjYkxmtK7oLRGW9XgWDOricjnaJXq5yH7WmTX7gZhWznRa7HdbZvHcqe6oLDdvY
gOPQr6t36ZVWL832Joqk7Db8TKqkhkTjLdKrmt4ESAYW518uhHNmRUeXGAPe0nMDWlK97jFFafzv
VIB5344+SBotzpykfZWvfGn06wkUcnbFE12sYlbg6LzLOJqXHqDqShD2wzYCrqi/8KtG/4CePKwq
6yj7RwGkekqePtsDTNcjkZFSRLfCo4G6XQnSjZ725WKsjbesIHFuvvtmDXK0jXbIBnJeX9Y22B2D
U1f17eiP/asLvtu18AxzLUw2YHgqIQEeOcvFRWMxMdkpxlx/v61/KjO/4DbAMn7vU1jhcSO6Nk80
rIR6XV4OUbsQ1j8Et3/nJueq/kwLuMNFzhZ/94JMec0jPqn5OKPiyBuD8m+jRmM9jqvwO2wc5HhI
US398IsomFhwE6vSpAZhlizk/IF2XYE7JzuxBUH3XdmMEsXxZypsCXOR5/AC1YU5p4lR0se0mxQz
mSxvyGxjQixGY0xHewgExSXZxcjVOh38x9oNtXE/7McI02Wal/0kbDA783YwTODoeJYp6ho8d1/2
LeJzbvfaVvRafiuaOQdAQWeW3Olr+ZuXWFAOLzNeRr6SnkrBLA0ltTS9vnSmRHO9qNH4cbjmxOd1
kLK3XGI/lPyJwv4yP4NwiJCFdITT7IFMYPBdKpIVtNA3w+fdpRTDWqEECCJLQJbA5qCQdtUG7vV4
jeKXKLzVjLEgEtZ47iX6wo9wPYj4cKbxHd1Ed96EW7NBoP5G948ztyStpDvsU5Qf2MSsn8L8U0KT
K0p5sIaNdY7QYdspaZoVdMGzQLaruTRyWzrQlFu+AxoVsMgOBM5grEfxR+F8PMWMBSuLxh71+vtE
woIn+hq60YsJyAldtx7s8Qy7w+WiZ4Fcj1ckdah6qDtFOYG/DFQc5HDTpLSjAQPCQH2M1M45J3NK
aS2Fcbws/KFV1Zruq/4crsIhroIsvSeisOdTLdtOpbok1iGBGCMzZChu8ZkGch9IIIaax/z+wsHA
t/Sz2wYhD2URSMGGbZkG0Qofb4kBU6g3eMEt5AYw64gvA8b+oiCNUSu6YKkZHWmt0q2Nu4nhA0cz
NviPbsSiOmeA1i2d9vjZCF6bNp67NPoKQgiJDVHXXuzOG6yIE0y6ltKtQC7wGJxbBG7CAmR0v/eH
+s+2Cjx4eqc5UYxL5/beIiBjqcB0hCTLZsSCw0B76ifhzAK9PrnqKsLj9IVwm10VaDugIHkIGeWV
G6Q0GjbRhPl874Uc3JhGyhx4UnNKY8t6B8D2oVPMYyNTgs1tUuhIsqAyp6/FnLf9HA+h9dSaBKsV
e3x1q5sOnxIOxUjXXUc3jlqP1ZlJPjqR33ZrKDvxLvHg1N/gkpc57GyehvQdtdgtMr7S4N1svymi
NfpbtwRfYMcbbqMUQTV/OGPLElNxTEmgS9S6S4G8i1DaZ2+/jpZKAJ6UDzZHFewbR3KYyOv/28WA
kn2kYHi7ZSb6Vck0srUsyiMMPXHC0A6bNHId4WcOFmH3NwPGNLLqjCQj2Qw3OWoNePZYDj8ROo2j
ZyRCcOegN2Cgr2RgSyt+uuiQnaO2ahFiD1sbU4irQwYYC0dPNaWg9u3mkuddGVi8MYdeJ7NdN+d+
rkUFDnUX3S1XsNfl5Kt0LJNkPjNPWyh8LSbmxzRs0cdSGHSdhhQbJSiGTLRx4//stDroJTrz0g8T
IRtb9oyGh9NLlP6pRq2+NBAcdflwKSev9iAUNvlhYdm8xYs91mUjchB0fZ6IkJ6f3v0QXq9kcjVz
bg7VeQz0RmxfFcYSL8gpM5nDJIhlqESDv2e5lG/Yfsor3orvCugXR/bIXF05L9p+SrDMc9E9LpEg
MAQbZQdk1SbK4KBmlbBdi6OhWCBHOqNquFLY5XWXD/NFBxnxEyc5pC7cpP8USSeFzlkygjRKfwVG
mjPXOeVO3l0NFBXmNkeW4lDOyoE+5ChlfdFBoP7qjsMB4ZXcQ+CYG0oTXyF2AEmfNfMMaEG8oNt/
0AwUYsOl6YybxRNnPhWT2o9DR8Yt+A0XYqOGwYLC1adbuCNrKCVCkjHaaD4N0sMnnk8TJBQ9arGu
lO8h1ru6W7CZktAK5Xo9xTmA51tgaTvKQMOTTrQNgAtmDL6lYMoCXgIXbaAgjcawEDekOtTcTKKf
wBMJ564S6bOYw5IYO5nHC5/Oy8sfS3J9clgllWehtpVcUjzM+WzvaAp3yy0Lfwk5GvXUQaTA7dnH
AtRbbmWicCSGhceBZ+cr3u0lf7FOOmZ52mmaIUyJsE2uecD/21Fa7+9z6VWctOAI48g4cmIWMolX
QOFsbGQefBvF5RqZSMjF8J4KDmbr4BdWkijOsZLVZZ9yB0tLdnvpLj0PNLdrlXjfJ4qsYPA+WtDL
QwWK27LolVaHixpFUsWgR4XdCoQ4PN7wrNqROA7OYTG/MpxVQVsCumSXZ0HB8Nv5zdDvQAPyxB6x
AYGnNYZSH6VLUijVm6Lp8+pdaEeRT+GUXbvxP8OO8uWPVZu2IuONNm3BGHgH4Q9BhmjlJIE5E1vl
rivo1jUTBiXgCVSxw0WnoYjG/j0Zr9v2bfYS8lnMwOr2fD+1GGDSqDEwBY7gotI/xSFbe1RwpP8v
Xu2hoHRelMaqiaYw1Y1gHkq3dEHMWnqeqOjHaFHRJSPuWbjC/1K0USQ/HLb5YJ3M9of80S74xal8
rr8EBZrP9dAqSi3jfa9x4WpiW/ezKhNIvUFM7JhNNlYyCUqK+kBeLhBeIQOFLd8yLXvuP6OfD3i2
U675CwdSxQ2M03ilL8kbyiwzUUEP8o28VLNlH5T2/EMS33vg+wbrO8waxk192Nh/fKgaGwmii/Ip
mIT7tShG+SQP1Sz0EZLbeQ8luUcmOaFWt/sVhkFSmFL268ijzKpkOjzzhfn+lca++gEnuTkQlAXe
NtG5CtJk5GAXTzckivd54FYHaka1AVRJyKkHeCAcXRwtj5SmGmstrUspau1lNWIt+VtiZtb7bJjk
IfQSsWl81/WN8ewRjmqWFruFyLN6vtc8jff9RrHkB9BubAemJnWkfQwqeXaGXfxV8e6oqdkXjQYE
eTH0CWP9HheagIlvTNEgieNseIAi8DHy5jStKBZIu6A0jbfQcFUmrNb6ojc5eQKs1NIUW0+X38Nr
6zrZ7VnZZWTiVThhbY76Z4y5Dwgbdp8VEsx7L3otnrOnK3sIjBj0ZYECTYyacSdEiEk2itl3QynN
2xmA8agAxk4Um0dkIM6XCg65u+BwuhcdhtmWX1FN8+C91gu2qio7/hSkof955BjyTYQHW22i5Epp
KFhaL51lCL+O2iz36obL36YS+bZTiuA2cQURiL4sZyt5L6hu0hm12xu4beuv0wDTiadzsNPecLbh
84XnoDIdYpI1Fji+vC1OClHAtE1Z4+fQLMeI3KM0uYt69HHGe9swMHKfBF9s+ClZOBuB5uGBWAhl
6Y8VIrfRKjynUqV15sW7kYT98vCViQg0YU4f8lpEHiCRfaY/nNOf8kUzP+Hb8+ZeXNnggKdeE+Q0
yApdWuXv1EWMBRu5Ml4aRKH4KHuXU+9sygYXj1Qjr2gCenUZqtFCE6Yh0Ait78xjj++/NdG5bkyI
PgqGbhGsA1jYftPlgVF7TyqXyKoL6b10rBg90RhmNaEq/aoZIXDEGohpQoVpKZUlg7+0m6zDvI9W
FTJLtdsHnqDZGpWNtQq4qFQg0QTecRfLHM7cfwZAPB/lorp7HCFSkf91CUjJNZq6nRaAvhZPayLx
UNrHO7v2msu3j6V7EH9ZJp5fT6ksPYjat9lEopShpDf2ZeoNcHVEKOU6OUiVIuflyWu0vGEi4yRc
KQwBU5jwFitOcy0TLAk7PhuTwk0eog/EDcqyxtWnGEPr/iYh6CMtX36ryTtj5D4SDoIEpG9mncrS
3bJ1ujxfiTKVe+lmY4ys3JK+lGcI+1NFMvkts9rsdHQWXwwUis5FOKZXHi6HUvhK8ZabbBv5hnBt
tZkToKcbrQuK5al8Bn45ajEYIDiAq2oHLAWu1ZDSt/Mbk3Wv5X7DZhN4rNg/iZybRHVACvh81sQG
yh62PPlN4ef42rnVwbwf+72a2JSkc9OFJuQHAlL9yp+FX7ZX/oAdMSBM0owXM6Uih/pcFe58qgWt
YvTzHrJo15pB71X9NkOk9/LS3cnEFuC4XGtdLSU/Z8Dbt1wpWMMmBdjbMuWUQRxhvaFirXxTk52C
COo4ptIUZ8Gzh3xFo1oGX8obuVGbY0KrIAClbQBsYvebIjJ0S1/TKS6K1AHrsyojTwYh2SDMeoUe
nZZe4djKxH/JsUvMNf8/6znPyg6E82E1dfTPUiDYzfBQ1bE/iX/J4Blt2AcVKg3iz2kqmbrWvFV/
s2Kpcg0PTx35KHtGI1liF+CBfRtgLm4qX01z9EXykdVzpGNm6ABLpcCv89m0upJaskli4M+VzkXA
PnXQoKQ/SnVfHpEWQBso7fSzy5WwH0EXr2QS2MGMtFya+CCCBQWa41uV6K73Q26o0tHPv3lDa/F4
Z7f2YDjmmVm7++tFw7EyyszLYRRjDzjWgW10vvc9LbidFri28o/CevIDgeN96BxSYXSzfahN+Rsu
O/SyZcfJu92o+USD+0mXoUDdn0ebdmJ1vC6LnG/3ISSD/ccbBEWKFvwDZK1cXaScsaPBswm7VLh9
PPK2PrlCVjtr1Q6mY077+t9pmo+wW9lZ3sk6cw0MkdHPfJzikr9/cXdTYZZtiT0FphcflSiqRtKt
UqQvDCcMHX/U2ILw04aju8bLLCASdU2ydI6ixU+H0FuM2QwpNOobWlPxehzmccMDuX1eMe7b+U7g
quXZC2LCtyL41OKJ1RrUkRm0R1zhSnaihIY6Shp8m+4u6rAuSHIpFBrVWnXcMvIMrV+VKFq0ggv4
C4Tfh2dtTKsnOJ+cFIsWqBel7Mqnnk/sNyltF9JNUW/odul1gpE1bCbO/LmoxKzdhXIkTarZwyz9
ABFLcGQrqNG5/LT0FzQY0PEPxQ7DtlzZC7j/x1xzC8j/mI48KXfXZMiYCqjh1CiVNMk7YPM220tH
aZ7wTC3ZcTXBk8CDv4jOxUoUb2XMVW+ajBXr/p8T+xxy/eYK1ZRmclOP7G5U/U9PJJRRS3BTqDXR
/pomdkkk88opH3jW4QpXpIPpehgnh0vqEZb9/3+xBetgBbmufCjNwaGnVlDbHuA31QMraSA7ScUX
eSd+VmrT7C+zwMk6nRG5tX660TsaJLN7SruDWLHHPtXbFOiGmDJWOFobg92EKXI98ajFbT3MUO/i
QV92YbwqSn3PnOTZ9+rSdcny9kX066O9DFiVSZnKzWAIekSwPdVNJ5cABNGoLik7YkQ65d0euep0
CF7TKoJ3RlkvZyMHiBKFRvAo6ldSsMXaDzhdbxdFwHi58/6jX7aGisec5JVP4OxDVaIzXM2WRTGu
NImkIOwLMrPXc/IQgNlGw9cACCpnar0P5miIqHkr6AHqSoeH6h30aocH8ksDooVAvxieqo6orbTZ
VNHGmbFwWQDwIOpYX1Kkyr7uHvTqutOXA3wPYa/jHZgPkH+HWOk7VjZTvZ3MzB0J+SCfcC/OuAQd
v0TAqtrKa0xE72OfNQcnF9gTe0nhMvZhCUX4OigK0+NZrjBYAcsHwI1wtAWUZpXVPibnoWRYr99B
noLAh3j2EC2E80IhE5aSv8GkXNJWrApdytGg0B91xLhdjkZJtfK5tN+Id+8iYU6FHYG9o5d3bAWd
E1kYBOFS4WUlCzh419++XW83kSEmICx9we4DMabPQvkts7uYpAw9/VaYE+sMkG9XS+0XwXUd/gCh
KKmlnChUjj6opwhTHIzELPb+0PlNlJcbDNxv64EjvFdbFYZtJ1AOuJtcTjTHhjSRbKEOQexWXwDN
OM/PLEQvU64n8onj7bhtIvA209KWneqzHpGpn3okgP+PyPIAji6o+myJOqIx1rDyAEL6wqpFWVgy
og7nx6M9AUhUN+A6a+YsoQ7orrlZZKAHuD2tbJ22hcljbOlDcEFLdVUHbnDgGABbpqyj0zgqBjon
ITDI0dyf4onmutwjOi/Tl9krP22klmpAIgcnHVEln/4mCQ2+5bDWfFFXSajLH3gIrI+3pRRKNE7Z
XP2w3VnLcGtQ3bpHQ6LHxUUX+A6AxLAvS4kN0zCuHB3RyFzJC9aSoK6MIRhvcGUhvSKpmqVcrNNh
HbJI1N/VGIpY/GEZRL6Z2TFHjeMXQLLweR358aFHNXi5RFd/QEXZetVgc8uk4EvhRtFlQmoSWPM2
68x939jeyMabhf+S/4xFs4zO5y3XByBfzlRy/5vHb6waR0mg2/jO9Oi07157ME2kPh+6Wolo4ZxE
YSLV3kRuHjGyz1ruHZdLlcqBEnMyuU97VmgATmE6OFP+YbtmqTZhEIqr4WUcmx4QqyZqyNe1uGbo
8K4Dyq9do6Hdj71H2kBPrxbvfgSRQ7oWMiosZahGCvHYIuXUbRfYpvsWiFALofGf+Fno3EsNBEZF
NMKwgLv157crC1vUIRYkGRl8cWRFpgvebvmgF1K0iTbakKt8n6ZNiR+lyHazM+bSCEmNcT+V892n
K/lttkYL6fx6esHgTFHMhEXHJflMr+0kWxFCsDBnp7KTL/fg32BK3iN+O3N1R4calxvhTmwFtevv
cIb8tl7idOsP3GX+HYRCu62SRMR8Mk9n5ryulUtx2IC4H+MNBGjXiyypLeKPCMD0oNDjEzw+sMQR
ku9HHJd/j4pjrYPjRNteh/pqTDZCiXOIp9j9uij/5C405TdCdL511SOF8gZGAeCb0oxuNHumVYsm
tD5S56abLBB0ti7TTb/YtaRGq5T2vUmQBMpUDVuKthoROysT6Uo24gTfLovR4km0dULLUN+DaIcQ
9Us78SXJhlmYrpSG2ySEbOakCeuhLhDMq5+DyvDzC4YFHMVw9sjuuOGtRLV9cjw2bWztTl5FKwFD
fQr44hQWcHLPmzqi+5MSGY9uGgNLbVsyXH8delUyPuDQwdBJo8fXNRMzw/NI1I7WIfliR8asQtjE
5QhWuZg2P2j3zMoZpEi/Qb34rbm4IdMbbQrtCUgsyCeuLkPnw1DiDltC2iUdCZNzKceEu32GwPxI
cvRRMp7HB2A8WrUyd3d/yRx1GR3Svr0Nnl/NGevQaxFfsHo5HuK6/yKQnD+tUOM1tIEbPyhixj4e
hd3MiErDAviR8cOl/N4gLKedPfzVJ914/i/h2NSJaU5YY2r6hcUuKZ2VMjMmGFBFdkmnp85mVIHL
wLWOCY7ddD4Q+PwV0Pd+OZDFGpqGb8yekUkVFV3JRNwgdT/MfDXRpqZgNzF2eHUwffgsZu5QZrab
/kkonJs/pdBO5QwSsHtFuzHXCFi0Z/ZwEGHbwzuabyoMAsm3bAKqrKesbTthwAMdIiNXhdAFSF+t
QuGfgKFrbGmGPDay+ymbsXTugP94Phe0zxnz0GEX5u8PUSzTQ+vvSaUpg25HnPQvcYZlFkRTNz0p
LQMhIkv3creCZ0sMvwm6n1R+NgUT1KNi1rgOmPTpfZy1OchINzt59aX6qWDPL/fYY+9nliFVghQW
ftGMxojWTwB4DrqJV4glXBDuXzKJ/h1qVry6rH7yYgQR89bP3d9P8K/yFbD8D+ucrkMl5X6osAmH
mZ0ZctSka160/JxyRFwHv49aH8mu6Yslg8mxDEwr/l4RdBObMlf9L6ilimqV/lF3f9a6T7JsGLQD
pL0rf1ekw+vcLpF8ji5K7l5EgrEjHsm0TN8IjMJBJ7qwcvTkO4QQe3txOqJelVnlsWgkwHJd84KQ
4hNdbZp/OVHUGrGFOwoGjvszO7QyrIb6hTCME9h7e8ujoQY7Na+5//bBU80yqYbepSpDsvlGR3RT
7HOjU5gsIwn6Tg8M9jDrn0yNoe75HGjZ33OzDPw8+SejoEhAR/lEthx4WsedAf7oSzwDWiwbCjpD
gNeCa+r+L/D45r+jk5Q5Rg3Go3+9H+SzkN2Hbx19n9NNBeSssZt+qNSs97OxSBzc2fEodzDw+tN9
bQ3ynoMseXQNw/EBYSrllo1EQhMkOIDiydCowL3b8DY5dlfTEOHHraiF8Bb+5KrP+O4snyP1DMJ4
YoI67uN6SogZdhj30e4bZelO1Lnwf7sGABcJ9Z5butsFORjtGzILxnSlSTk4Ghvz+Q1lsvqnfe+b
f+UdW1oDaANHSK+UUwG3vwDlsn/yVz9XPQiXRPNb35Gr++COLZK4ZKTYAHOF/yifLNjMNEm7m2Rh
qxt7Is4tNsqZzewCddA845gCLYdg3M1vfPDA0CjmUKt1w1rTBL5dkNC+T1xKCfzpRhdGvW3Y2GZu
tOq37vk/foufMyGyG93G/W4ULbOGG3BsRHEhLLimcizicRzBOhuYzfhYC4nsg7KbQFuqXLpi0IoJ
65RUz+4FJMmXWEHD7aoRAUUZWcp0d8wMqiLoVId42HplNJvyvdBS+EnaU7F0VI6kYGsw/88WnIQc
2vE/Vhl+qqJnSbmZcYeYNZMKhWbotT7+ZcbJ/cOHyWK83416OwnoVrnArlUhy7H3LY408dL93I9z
PDoRvbt52Cwm1550JKS3xc8VErsBziXmZamK2K3VMNSjDkOv34zb8QnG0ozotE4PODiUptEWWM9w
EvLVi+Y2kWL8q3TSWqhU5m2W0z33R2Qq0HESVoDlooiPaHvTO5DJX27nSmjtHSW4CLv/hbPElPcn
XbIRtwvqeKTsCgcaG/zYuyOXgs8bDQhDaun7pwTPR68kRFp6VhZ41vzyRdKKzpkQS7iQ9lWd2L3A
1SXs28oewJb6boEjPg4A48xIfB0VoqY7cPefKRx9cZGbGvY7rMwZ15+vokbnUgKyeutcom4A6KKp
Ni7/xHkWU5Z+8+AqLNmZwFg2Vd9uyS/7H6GSl3cSxd5xM4ecNVHQRQgiT1dqq0lcK9Rq/yH0HQeJ
/axYepClGjvaxrsUzw0zlCSghQwgg1zqjN2QYXX5nkJjO0i6/v+kfBAR/92GFEyuctaPw0wPFQsx
urbQMjHFSaNmfy6waRgq4OobSk2xhE6GzhavMS3YNhKdLRmLS6l3BMmo7VjnuKfrjcdmkNYRcRRF
Mh6dc+nMMaH2NEjglGdccG40IbLjDA+YhAlHBMalpSCKlePcx3CI82VDXWoC4jfRUo45JZ3tUes/
VEqn0YIVJX2XNwcT6WAqNAl05CSUJWqGfo4QKvHy3bX11NSjXL8Wbgn1tv9G1oanCdDHMhbq7QwB
K/jUN6Jw2NW6CW15g22ZZRDzDPEJie1WQuNSJdXBMg6hsVJJ4GQA7SNox0piRV59Xs6bFJlli8F/
5aP5s33WSfUDTPjeNDJ6Q2HCePgSWk2giJCeZeFUe9I9H+UWAeWaV8F6/YKG2llJYmGH+gjHuE+Q
0X+rRcFkV/Kz2vXqR+43jJ0XuF/1m4wZrHDAdErsFvNeu93mJx7x1/K6Dnwj9d+XlyrNbNHlK8bJ
jhr+8IthdKulbFhngOQM94/EH8MljFFnxVEuyaX8GkCHLtg2P7KkBF1NkYKbGm4QiSgpYo4U8AQ4
pQGNWoSZDZPgom/pymlEZ4iBkljQTkw9iYsrhgIkDosachlRqubAKosvrJQQyaDsatoRuOqpqWb6
UpJUexVCHoiM3LtXzMXdpC1p92YQC3tF0mkmroqQ/m0fh/d5CCSXADeO6RaF5LoIP83EWIrTmDMa
xtLfedsXcgmuWX0hf5TW1OYvvXRWkkdNAl9sgCCBT7316IjlrpBU1APlPqJWotfQjiWlPCJWOJVd
gaCJDkHEMwg/cmG8J+28sv3TNRM1YtIjT7L/YXPoGcFOFtiL13xtcDjIgikbq41kAWvtVVtPVY44
qIZvWQTPnxjF6eVjzD4/bQJaLtxg37EhgITQYRreQyrxmrHeNviexhEEgHoAh/mwAoruFgpECssA
tWVJGFdE6PFZ6XJeevqWmIQgLeGiAT/QmRHRbSXQNctPYzHSfosWlNUNguNgXEAY7J61flaru/QX
PpaRJyNcon/gOtcYpZOjrHWduyw/1lJYCt2CKZF+5Sf/zKqnQPCjCmmLBW+eG8CfuRkSWo3Alidv
yvb7WphNM0RYAcs5UvGlgz0S6zOgfTq6rnbVwLhqEA45yYsO5vQXnruivwrKq8i85en5sE8G7hY9
ck1s/oq2pZ2Rl3ysCgosqH2uvrBJWmb+rR14rF19vjhOru7kqHzEnhV8ccfmSC1BDcxvONlIBUtf
oJlzx7x0AvhAZmRbmIz5g0heJKas3rO4z+aCqZMJF2tN02okU3/3IEKibjG3y0wQQIsXqwLY+Aou
5uU3mKOY/N3kG3A2ZEA09vIQnXlVgWiwfAey/cHdWdV9aHSP0MCBjHOzDLiz2ZdKFYRJfygyzyl1
Qz03pknyHmzrMwbwXLNkRhngp6QSGHbCtmlB21e4V/0bu29vphy0idYGXJTlGJLdgxOgnpFQ2f7w
dj8mBMRBTRn9PHMjQvnw5XpSpGolPcoMJWtwQzy9wZvQJR7daW0A6BZNQG35kTnRbN7kmyk1UDz3
Lv1GaJlFp2Ll1j5oRQb9sW63mnKNKejTuG8pio+QjuGrqL3UylqXF1w+zwjLJ5jUvDiUBaDsqB2F
KFKS22nKAxQylh7WESujPQjJzgQ2jdVEFvgh3ZnltSCH7/tBir9s7744vePMhOH1LKyVC5g7taPn
ekunS2+R2Aj2GLeSkVknfQFf7TwjnUHEfGBRXct5Mqmh0grtIJKsNAUBlQStIPaMKya7eHpD2t0r
xkulTyELSzXwtvj/Izr6onP8db9IKOGfNf7vzMjbO1NcoV9k9CP5IrUl+tkZMYC4wiB57yZq36Mk
iGy+oktaFhmodQ8LK8cxPZCeDtbLVrJB3UzDVE4aBKtTcujX2ObwsUQTAajLpiMfm21JVzkdTewg
WJFTyagBB+X/DhlAq5YLPYtaMlrPyeFtDgKNeggKzHYArsRrsm8YaYRJwKa3TQ+AW6KvroTrQU5R
PjVeWUyRexoH9AkN3ayCM77xHmWwZ2nZlvuNvmbK9+ZGULc4lhx96hjSjmmvXNtLu6F1gUROKXOC
Z7U5/1kOVEPEhzXdGDDSxXR6wKZsBIV6+2VamLt8VXzaT2mcCwkQNANh0RR06pX9/cSx5T358tDX
sfgqxi9c+fOTly39Igb5R1ZYNnFaUtUyk6osqSC4kSYBi0/lpaCrN4NS2mmvxgzZntIk0OErfWaD
nMDVE1HOmtpOax1t29/zuanDT9+fQeMwHvnOk3BN686f+vegGym1gWRKFugVThHxP6a2y+RxEe7X
oFYgvRWsnWU7xh/H51FDDqDLbWiOqlrOfq7s7JQjd9iHZPYbm/Jsb1FesYJMphBsaNWyc4ZVW4QU
dlyyi+j6GS3w+AwkxSEVTNxCbgYS2NT//PjKRVQKKNtAKF7Hm0kXe+2qfWE3HH7YmCQ8qRld7wTd
3rJ6qpl0Bs+aG4dF8YKTcM/N+J7a7MegNo4hi8iyW4d0Fkogm8FUTgHFzZDv4wVJYwxE8ssDMc+B
KwaVjunqYP2fnNrRLN3eUqScyzLiNIjS74r3PpRwfro/qEPbPGEJhSrvSo29vmhdYdKcboFWnWRm
z3TALPTR6YocaWseYPla6Jpaposni0FUbuepILgjIg6AAcEUhG8r6KIjrj/HvQJ4B58Q+YEen8wr
esfZz/2iIH1yco8EVijlTGvxbXyKazUFmnWWjqvgHMn/DWfiU6HvaJ1kGy1cC65kE5hvK64pLSpz
JCYVM4gg2Za2qY758wsxDMENAGIm7wvJDZ1EqfRKH4XhjvqcKqCXJRXZMtO57Pe4Iyx6fF6nm6R5
/Qpnhm/oczAyyZj+zW3ijt24J47rUnqEhuO8W8zjgLruqQJoQ4daAUMFPx94g3dEwQ/xu/1lW0Qz
JGbe1WaEa7/K9rxDLce2Y6j7/iUChtQjevFzfBMsmWb5u40e2KQGfe/HEzgkatbWBZWnIbORXcMU
P85o+enJRAu81XSjaOijiMe9FzA1e2784/TQsg77cB6Jj/yntZeMG9aKpEpMZNjad6p6ASWJ/DzD
YdyvTj0k+gY40MZot4rqYqga+uYZ2/KAytumkpqJgC2ZdX4K5jowreUksnSz7ts56+x8XI7Qjuul
5K0rWetRwC9C0PLTJkWU/LZvwaQ5T0vbr/xh9h2jzhQ6+sHtfb9f9YKw0nhMve3rsfBaviwyNVPb
03dkuYvVvL/LelmjSI8Jd6i01Qeh/QbTtvFNnvhg+CEjPUQ2rWkjKxNDdUmRXgJ+QcQS/TsrHrph
xWiDo7uoFcxYng3T5F1utdDXZTqkxAWCXEB8fEdH++k4MDKgvOtZGTp4HkKKC54qlTzPgnpq2GVg
K9iWf21tAeIuvdHmnP/GF/r5H9jb+d2YP2Hf5W2a6mr4+r89TxQiQkgJxxlbvVXlt+3z1nJdU2yM
hW3HQ6NsVt7SIC18Dvfyft2/wLJByVAf9ZiyrUJ3M73MLCWVGckxC5LIQECqM4NMsvAM5h+OY1I/
VTxYIW5AqBwvfeMYaWQT15kE2nYJjcSQebCQBwjNxYCMUjVUdpEJ0O0aU/PyTYOEDr5oazFSZsYs
I76BqxvuJsnQsPrpB4hQ2XwPZnTZuZLcxpv9GvnFEdiCFzXbKTAfELpysj/Q9xk/4FndwePICCg8
NO8STM1w6qd4ggNUk8EcyW/7ZA8xkj9kwf9ozIvSP+3Nr2X1gDAjN1zgdrAggoFjA0F3eURQ/BuR
O4VPlxLnKQ3Lj9YjyRzp/44AGGZj4zuxzJknNl6r6lUxxHkx9p+ZjP/Gr1/KE3Ul82CAPQX8Nmbh
3U44qAn0xATzxDsvRnfO3di2EhTtLNrGPRBClJ+bwXD2EUJXPWCyn4sZsFc5ZT6j4K9j3CtJJclE
A8PNg4K3yZEtXgerjFzsQmYzTmoFkz0852OjiLIAG68dMSg6tsbhLDyD4O7Mo1hxL1ZPChOduplq
J8hR6AZrNwU897trND8z8xsFOnq1Cb1OYQ3VDQOq16wh4WsM5xR49yRc15avkWNi+lzWDoQz8ehc
yTxaLg7tUiE62t8WyjDJP/qAKlmlPIuVcpH6x85LH6VKg62E8E6pXbwlqefFJ3zf8nupYD9RLRP1
2RNH4e+gAYsDoRuTcmmmE4M6xOAcjcJbUQihPgf2mOPArrh0Bxr2gKa5hWMPlOmttZ3aXTQko8N0
7U5X1pJSA1WGUgN9NM8g7BLj4kQ/XEVZ9SOaEAypU+U8usVpig998viVJaGmhEJkK7uyD5LaX8WE
Nh0VBaK/HYDNVKb1IghP4fiEyoYXWzI63er1XGFGOk5WINNa8un3z+BnH/y9ZgPgJkwiHzKgJtHt
NP0jxynwD2ng022V/J79QHZnZA1tD2y80Hs6jPs5ZAzw30+NRjb1VFszOb0EWXvqK+AOm0E+bLbp
KHXGUwlkWjpdfQYI+H3cvDMrcUdx0x2/+SLIq+6nJePvdVC71jxntnX2M7m1hjXkYR4/T2N/1+0Z
ZTbcLJWZKiIkXMDWuisBVVvgFlbSeXbJOu2Hs1186szpZK4HZZR6bb67jhXbM377L9kgirJFdVyi
RJERzXcic5j2mXIM2BYqBLasM4mu/J6QU6FdPJnr/zTbyMdEOgqaNeXRax30pges1drpKg0p0dWn
Y9QmUswgyvcyNCijE8gutvKfKiePsRwha5W+qhtDSYFE+v3WVFjhUtUj7vmNuvZsfMVqHn6pGeCG
PESYtjk5N11a1vY8u/c0xcbu841Cm35DJrgR1ih246RI/JQx4eSGH3o5aaFvq8V3LHJMqMJP0A1n
RDqnVovyaLTJPlhHm6CNWRl2K5yQ/boqA2MqvVGiazH0gA/qGyRsoAtAdl2cY6Ojsv4j0WmdMGVA
u14zA76OKVdJSuJBk4pUI9B1KHaYdqxJJpw8XWaC3znLBvXB7C1R+5mp3RML4dKZ1SHBWB+541Wq
jI990pVj9G5VqKwNTxx56LGHo9pyPNof7YJ0TYIVOIgggFcJfcJCAMXYxGKSCA045GjDJR4KH5+z
4Y2elgCRcF2uuFOgi4L6sX7wv9ntYjWLDTAjHj50wsG9iacmEU0hdnRm7y/Wlz+qPcubW3LwGcZE
1pZpHRXtpXrgbF67cGhCH2qRsAmLcvmae1ef1AsO6d+zn9pTHjCgPrmfvQqVOjUAPxGZw8e4ojKE
BgeagkowecDNf3pvTQrij/xlDZwOQV+Q7qYE4PIzl8Z2CQOSRpXWofmKS+PI3Wxx3LjqO1rkrCFd
oM9+KsLQVay52G+0GSvWZFGAmWMYhH68TAYuH+JNYZYz0TrzPI9fUu94JciRa2RUEOs1RR2DzATR
qrI63FGA8nHieeHy23fvVwzRO7mcaMNHJTgIQiOyLEAL8FOT57YvPwVwsWCOr3/4RPLCSGz46zqy
tp3/a1d+AVwJirUtICMLQVv4lmXZo3JYht6L1kkElPDwcCUyV3N3elOTJ+N+w2Brmu2HzX28Qc8z
lBpwtVcwoCnU87PWSEF/pBkcrI9HIP2V0d4pOr71HR0CBHXgZ2hXY6vDd0/jgMnhisXrlDka/Aah
gi1Lab7xXSUAPE8rghRNtZT08BiUsCFvGe2UsC16amncI+7/Bkew2WQ77DoG/FJmeDsVOV3RoGRU
0ohkqI5FH5RmjkTZZCT/nouRBH2DJjaxE71ENR3Hu7ZyU0H1mAZJBcQ22jlvpIqlMFwj6zJ90JzZ
67fR4ZHinuvznWIejRGUBzbTr9yc96kW4h6K0ysKFWTVIH7rc1sFD23ExxX3JymOzHudhkYL8EnG
9iA88Zgxb6JEVyAGqN1jn3ZliCIjeT2b+PyKGRDoCsQPpjoVKBmJQm03r3amjFvQLuVahwnvDMbR
SjWIRFd5VzlLHOSLWerSLIWK9jlmFRTAeuOwDmKYPZaolIAot1SpxLmYL9O1EKh7nJOtMND5ipsx
ZvhT/EgwoCcRrXuSp/C8KUMzK1PwH+7XSwmqjOu74DYBuvURtl0BYB1fhS7vBNaS2Qg0pq2oMejU
OyPys9rosrytGRs1iK29P/LOykHVBDyG3uiI3AujSOYHIwben89Ly52CFgKSv9UjuOaRX2nvn0p0
k3TRIHppPKFq1B/KnwNseocuU7JV9jLeTmv3g3anR0FFD8m1KrLNi8kFMxxgFqyPaGAXL7GVTJDf
S5IU37IZj7tajDfWuKA3UN3HGVTwESKD9iJn3318XRSl7zTQDd/VyGyhLP4/gp+iu50XGGTksqMl
1EgOu+6SJdVpF+yKARza/LwxUkktBqHVWP20o/dre0T3RLp6pt8tksUBayb5zMlxs+13pk0kssRs
BZ02/uiRaptcYdPtasTBNZnC3/c+d2sAqkbqxBm6JT2ZIdlID8iDJFITQiTKLEyAVzVDw4fq7LMB
9BNLYFSMasExo7vqpHAeXSWhtgdhwUiPX05782vx7JMt2/iRUzZ7NjaeaspJwfwoKoDJ/efdwmy1
wuKCaSSHyldWgXVZu+ld2SPFAm0k/IxnGQibMozM7jqiqJimMhhGo3KTcmVIJjje7yX1faL32Dlr
h5uIssYStWT3i0tMyviTTEgCj5vx4vjiZT0NgtcgutJCcs5IfS24cgWsD6SsUJVS/jyoe3dA8BMK
B00TQTewnchrKXh0nBGqAPJcNdVO7g3MUQmgvIwe3xVPZW6n7JhBdwGIAGGROzHH4e4x2PIrrfsN
u498RHvhXmDoPFa4amcqRNmM/ocepoFkzWdxaSdbQjortFEZos5QmGDuyKpAxrTjDa4Y62fPWG58
mkfuA8R4AO8+jIHgURNLusROWn0WjpRMblZnCEPL8qxjhL4umwoHlP15/a5cwv3YC5yk+SKLn5m5
E2pkZlg6L0R94J4dKGbJDdXdF97Jd+r4dx7a0z5QyfXTSP2xmfZPzPcDGSUV1aFj3Hy1bnjl/ds4
8LvU9/guaK7pOcgKrGzHwyPkfDIU+SAD289r9/qSuGWXsPnnOu1Hu1CEkoeVkWtLX10igr0pt+SJ
rhListv0GrF+n/ZM0yQO4+mPCIxeyqyI10iQxhz5z0FlzPa0QVRxj9XGYcKTe38Jbpq7jT8j4A+V
EuMqJrgu4hVbReTad5lJvXLx1AH+wDvrD8LV21eMPeKW7pjWl7OI/060sQrWR2cSIUN7zEGysfvP
d91RLd/5iCkr7exvZt11AHLwwH1p7PQRkok+Dti6kJF/PGqsXeB0lXLjphrbUAIFZcHfrQe88ZEb
R7DNhd9vE7ty8NvcalVrBDHRyJNwhv2zuvh8zMVCBKUwBPLZjUmkzy8U2+0tWBf8PAaArpO5ImeN
eeh09pdx8gp0ry/KVPTqa2a4x2cO3e8VQsNoE3WsHmYF/vSacKAPTkI3MOxjLRD2mh2TREzRZV0K
jvYGkv3rIxiyV1YW7sKedDpjwk+ImvHjAtldTFD3kuzfpPLK+0D9KqGsKwrradgM/uAyjjfqVHlH
CQtDedLVJLD39VZ6vw7it584dkEX5uXI+050xY961vJliLEbo9K0LMnqak6xIvwyPh8+BY5c8qKV
i2ZKlJPSmRhr9+2luP+/02bdlRcxjY/vbGngL7L59fKBSQm+7Oa3/yfFVoB0cDzkXiwg/xzUSap1
S3IoZAZZxwdEao3cJekW+a9XpjWT+M1jhYWEr8qbyEf1OGM5jLKKpl51TVHJ4Um0+bCZeJbkG5Qq
9qa4KVEMPjJyrwRMV56VB4dQIxWngVBSMo16XnfhWNlbzlwOjoeZPvzo5YDpfejJq3xBNsFesHPU
hzwQculTNVKunSfHIyBhY6GRrQCk5q/HpVoYGxMiBiGpSZ5l8qvfyNaPUOGBV7jyFSSxnK4UJ+k2
aVeFRMeKZb5api+sx8lXYejr4P8FX9zg/si5uFARzWSkso6aPBp60nj7UJuSc7qTHIdixQciUsRr
yxwwx63Dhb2tDMO0r+R/ZKR7IS7Oubmd35vH91emLo36WDTeYaPhPOB1nXag7jlwf+kJcfZGmr0X
EUkPwQFKJCsFB62eoEvgjZyHA1/OY/1X6l4aeM5xbHayFFv8/5Qk/1US28snKrw2YSVblLyoagcN
PIrUcYyoxr+KlaOZ1GmppUXfFLW34G8GOo6fE2o8m0lP9gFd/fj6u0wSL0CTP6QUNknb5CrFGDf4
gYZNdVcgmzt3/tejKvCNaVhox+YiId3ypzRr/FlmCRO+oo4VVJhz2s7ttfr9wK6apz+YsuDoB1gH
Sxi22JncQpNEdllLGUzZi3lRxy5L/1qeL9mwTWkeXoqr76xFiKEdWJspgnsQS4LTJapZkmCm744E
qNpj3CNuEcQ7IG9iQMRR/d/64DsSxmpD27ddt2G48X4SRk7R/1VY6Ucp2TBxfodBzlrUObt2E23J
sbmej+PuWf7e1UCMczQcHuVDPiKgfYBtx4WuYkNs+VG/0emSGSBN8xm/nH5adL4jJPqJ6XqLRcg3
2MykCYDg7PZ59i1crT0o1v/ydzk6ASMGmY/rDjxbiB86cYTyEwBx+qq+MNE2p+aBEwWlIo9aRSR0
miwOhmTdmJFwHmZDQ0aFgj8O7ULoDd5iiABoXasN38oPl4eXXaQl+BAJePFYW3HNkJu4GB3yZijl
YKX38SEoS93NRO9zEVNAzgdpYR4q7e8MXvuxehE1S29Tpnli7Vr3YEGkms58rMZFPxT5zuiOXZ3i
TTOOUfSx720vrDOsCJVlgiVHnMz/ftFC+bZ7IQCedJhuwyltBUZZgfJ5Cdo84O5UopeXEapc/DBT
wi59tNMjo5YEn+XNqybMQIvUSZm6sWEOLmXe3Cauzj0DVRPCefnXHNrL5v9NLggQmQixIg9F5W8d
guQ/euBQoj6viLZFo8gBIzuNlQsNngKg8BSq4bzGdLdl6R65ZDjICiA93ERnbL4FUOenNI8/Fpft
W/1jXPVvs5CPvuxkLxKs6c6Uexu2mRWSU1z8rBB/wtCvz0x29cobwLvpoiTOXXtSUiGniB33z2FB
ttR0rzqsMTVNbDIUHs7lGyoH7r+8zV6+g+gjWPLQXj6ET6WKhHZr+0HRDcY8I8pJTNRZSkaiTCwE
duh5jEtmNUwcMc6aJHvqPvfqlRPnOM0/sfM0+Yv4+h7CBFbVfh+D+peepB03zq3sCPbyORApmOem
CzblOYlpJfDb1YnwzauGs+irYpTyslyTlYlDsDTViWvipkrXlTXe90iXuDTGt6fdSCO1DD473zIF
gSmJ8S2p91ZG/h+tgXs1L75ga32UPQC8PFDTa4CuzBop2k9hSXd0uRgRt57N+9UvDrEk4d/KEjgc
q0zzh/hJnWONhEbjWv8wxw9ZH0y3xJbt//UWy7Vl8DuNwLDAl8wtEIbyr9Ze/5GPck1oPe0bR7ge
6JGTjLLfskOFuVpk3kZZglQD/q36ty4k+sxNDJzGkzT0Z44ykx1zIaUoWrbCKMga61k+Lh8+hd/N
NSnItsKyLdgdpg2ahInnO+3BR7G4864ApGB3elSiJ3YdsUn6PS8IeExyeuOEDfn2KPrBzXxnIIMw
mywlyF7jtPhn5dHmfV2phHUpnw42ckp9DetB5ywY+7lFWtzpXiqcZ5CbDmvR6XGVOq06T7qCoMI1
wj45AEF8Y1bcm4cmLLM2PAefYwYje8IXYDsGufCcAdUt5tMdZ9jxuCI4rJ/ELxeHgaGrI5ZAe1F8
0VitD4lVxoQozwpFz+z2koNapldTMa8wGce4sOHJwtB9mTU75PbBAQSxkKIJqLjAHLCH23zU9RPd
ghw7aGc15WKem3i7+dG8QOwxqoavtRPVhCpfleKvdFC1KcyeBu/Mi005+bxHj1qXfqbCdCmkIb2D
3dmKy3J6mFPdQImXcgH1yQbxNNGVABPrsFlyd75isjZk70qRwfzT4DDK/dYePF+rA21m/Wn49KY/
jJP3OJgwfLqQA+h92G7aQPtHY8b5kKERHEygnqenhA+BxrDj7WJQDJtz3SEofiry/mhe9R4QAkrn
jC8n5UNbt7/hpwj2kpPIcOOSeonW6CxJGtORFoUibggSe+0woswYhJ7iY42B2vAPm6MuaTHBZ9Ja
c+tz8z/eb3zQIpGxHsyI7ny1wrkxvoXRnMcRp9EFRzBlq/kFheH+jEDtfdYT0ZnZ0tJIpw/gBWpy
uPeSGosjN2R+gkUE5/SaEAeVuBXW9DzvEYENrsfoehs7zk5aiXAajf3HkgY2ZD6586T2BiK33LcT
B130Nvp9hQm6PfRRXGmCCVW3pazqSWn7UEpQRnHEWsM70kORB8wmUKSYaKVMmeK+nkOV8r67F6pr
qWV++TM+85ccwoThK6lE2x9ACH1vd4zA4Uzr2fLtcRLZ+WC3RVsTW5I6JvWKQjdJgA9KhlAjt2x7
Ib/c4jI5VPDGmvU1JOd4w01ZTypSVkPiWTmynDyY7qeiwYIdaRq2hXQzn5kv7WUUn4Pq0Wewudvz
4PmetP1LG3VtK3DYaIlaf5tCU9E1/Le4F8zXLHNpl/Sd9z6/pj/wNQ/7WcR2poT/S0aftgljQttn
xJsp+ihb87PE7A/9NLEAJsLPXhsjwrUfpOGUZHmb+WmKMgTDtGEBAB2UDMPy5NgiddIxVFN7QxBx
1rAPTevu3R6LDczDE0J6HRjsjzu+1q89HamMQVjUsc6w6fpmhAi4MkfobpyjtwicdfKANla//BMg
RtZKrAB7VmFGQaOpqa0jbz9nnIcP3A/8+LV8794NDnRUgezj34FPbT/vLW+P7XnfbrX6aXwrPkhf
8Kp4qTXUdYViwmhbsZ2jT0LD43rdip4AKGFNy5TxAZg2pharQHZkHJl3qrv3vQKRO4b7lXpL0Yhu
U7d2u+5eTCGXaEimkFmRwxd2i4novtbhMhEkKl0Jtc8t2Z+IpRBejUR8I08wXYFGyWGJ7hVjbwQs
2R3tPNS07wSrFvk//a131EF+VtapYM1t1EzSH7NrlAdhY1jJwvsrnK8zMiNZLDwo3IS6sCn6NdYN
n4kPBFMGRkTsjrZhNEZG/DSjm+zg8eWnFQa/OBKifODHPI78menPe9YOj54Bsx10uPglqdYO0xak
dxgiqsKK/rU5zcm8qQ8CSETXl2yT3F/Usfcebeevf7YJALuWFr8C7jQtERSZrvdfvwgTnjKSRQc7
QGIy24CUMFxTZitdCOcTMzq29ZrC6YisX7Bd29y2XwpRtKchLBE8pcH83hJjFugPfRjP+IlA4RdR
VcxVPZrF4R1CBKi+jA31bU7l2WbnGJPIvsvh8kztlllYvApjGx7/6DZLCsBZRedmT6m3UtBJMHpL
l+AWBWMes99J+Qrf879rxGW0jlz0HQQuL8hF7VPAGuboVe12gMIDgAl1F43zaEhd5dNnaKyLZm9n
JeWPUNsSVmgPR72yNjRMaTDOMcz7J4tA8Bxjouie5nj9W8me0uPhH0CdVdB11XfcjY+dzPkVkzsZ
43+KDZtYOYK8ytjo2lLVKMBrko/VTj2r98WN4Bx/IQTKPHH9k3jvKZQDB1vi4ToPWxhjJ78Epwnd
egpu+vORlDjpcwvsYRAoehy6TZPXEXx2A8qSl4YMuW2rXinSUVHW1A99jk+se9TI3glk48h3VekP
IUrv+k0XEdL35uTWYflxy1tA76t1foTr0z2WMkzKBHBLmG+zJWcUURxCZfVlDaPwXRt1JJAe3j44
6FScd0RUSzs9zxUXWTQ1cORGLm4LkztszPXe560gOaPwq1MfuwNZBpBrL/h0OIiFCtVZC3M4M29+
PNqxvgdhFGZZPY9X8BRlI9jHjOzcCag0HmccT6BZFg0dHIhx4lt7hr7JC8cXNgA9fc3zQDgSqMSK
Y+8UeZjRknmg18dIOAqQjwbySsmXIUrEKrCa0LNcvnhdrltwiM5oz4ir5c1MRjw6L74EXqpi/sxB
xhlDh3pnYDvwmqgiM5T1mXqBtaR07gfSAZTFoDhvHCJjkMMYRcisBHelw/f619RNH9bB+oWl630d
xK7tmTc96IjJPza5Y4mstnlBe92NJniQntIoVNcRo/GDLqSmhfayizrNNgSUXmzuDnpZ55JEvEzS
KGoU+nuyRcdlf6kxIyD8w8ti436w/DSppn4fO8RLckKQPRU2DD53pe1XoGyuikb4Tij3tzd9PFVm
ENZWeJ3SFdk+2/iX8ZTIr8NNK/jtiMWCoyXr53iLy2cefDEdD2mPWmpncnAVCQF9QLr1aKzTdRoQ
qAol1xQg5mOHepZ6GsCo7vwPRUOiJQf2Z9vMiOv5+b98J8eeQHeYFr6a9w4VWpWZqT5/wLkMGkxu
+lSoDNT94U2bK7Gzb8CqgFCAL4JH2N7v1gZjn6Y9XZTJwR3uCW4hqBVwsPbfI8tOPK+BW2Op99Os
5HIZ6D2gvBylUMwXXIBVHroY1BsRs+YVA1ci0/vzCkdTajdp4BSv49iZaIfDQeU0A72Q1/r1xRl5
B8QCN1DFgm8OjkX6V/rELHfQs+iCE1OoyFxI9stGYzNszSh/CFoCkIgpgkaV0674H/LC+/so7feA
sOm103JEoS5Y5lmczYFXnadEn7/iVXSSdlmS7bzJxo7gaPCZQJ1ha+cD2/+Xd9J6aHPzO74ik+Z0
KgJm5CBh/X1gKGTYJMEKgURQFrSiaNTI3jnHQ9wSWn4OMipz2XupCxm9t9bp/opDM+NjCKtseF4h
S9WhWA3bRJtexd9+D2HoWOA5opcezfftr/rp2khN/X2qG+u9UR1jkaQyKJA23aUAHj/EXi5DuWvn
C5uZWQ/J4VNutyMRkz8K24JUs1CcfCsl1BXqDsoHgf69nSAgX46qsQCeGLCGVitsoc/e4CHP+Sqi
VFip/E1fm+aajAZt3SUsgwEqQTQ0Y1D9oEDUvUOA29SdPmDyBjTteyf5naWGnBUH1pP+oR5VBhgi
/H3TDbS20VyQOvZqR3jPTf/5ef0fqrdyj83NV1c/iTpb1LhtVGhKQCRthaJ8NuJZmgWQHNtLtq1N
G3K703Uuo+UWW6h4dUzEU5Jg+JGjQ0soYAhX+KGU75RwowYMiKaGudJR/basPP7aCgP3yShMNIUn
M7P5oYDV+3bKS75Uo6CvM4sZN6HWazz8GVpaA+V0FzEzqXmdj7cN1K/z32NhBFSsETJaj/zIJjir
omH0QjlJPSFTQ0vKKaoh0g+bLRo+xdHTuQSXlFO2uQxxE9f2HjnU/9A9BqZk9kDm+0l4JGUrIRKU
kJLzZrOPcjWB51clDQbR4sdkvDwI4k4CU1eMsDpAuaj63gVq8aQCAquxqMKsyp0pnH6jAU1v2Rkb
flDNYR3DgCENSKCNaMqJLt9YGLd7YTKO1Q9N/BXin0B71ZAQe6ULilJCylSIMNyTbfW+hV0sOHwx
W5Jlv0lclDxEJcVc6VejSWLxiaD1qhNCP4j3Kc6Eg2wTpO5bAcgTeLTVtemOV+0w/cFUcns46XYa
kL4W0CnXRieaL8SP+2sG5toWXgi+Guh20khHe36hTfV7VmL6mUpQPWoXhhuQuzcI+mk/VqlOXSvR
zgY/2FWAy5PAtpwZhZ5TLdL1gRZy1zdVvQy79/JDL5seWEXUsO/g8wZ7kDqRxyvYS0Y9xLZDU9OP
DkppJekWVsbLNcH1phVCGPC/u3ijuVyDbA4ADo4tlA3FYWzeBSP+rCXsgwsMbjodb1mFnr549YmH
Y/2yggyBqe1ui9QDZ+Xh04g4I0xwdMb9u3AoOJOPmvl+mUfjJ5qjg2nkJ5iA1vab4oUIravjo0oU
Aq2jjT8R83Bdc0Uw0ugzKw8US3GoI2DF3goOOjPLL9bC3sO7Gn5SMue7ci+7b3vdJnTfAFPxaFad
Hggvl5eN3RUyt6QGZEQ/nQQLoCBp/pHW71HVLpjS6NhwvR6kCMQFHU61L7F+O8TvdoQB337gcdSK
OPtVURnSxEgwhojGxqe+jxa4idVWuGjNTjflJ9hF2QZhsFH8TQMGqnzdJxGo2E75uLs4G4j7gREZ
mPiOx1XLjMZ+bafALgB2Y0ftVx8sbeSUYdxxWUHJ1cacZG60QelnZySGTU8muECi2aCahYFjV6Qx
f+72zHQnYB9s7Rm8NR4WgbgCy66Nv21wglhmyFaQmmxwEVvLdp3pHDIWVvgsvTx8rgqmYmRTShzW
Pp8C7ia3EiRTeRVsjlIS6pYgqzjcxOr2svFcY6fxuZrWqXbrsiNh6Ckj/KbE9F/71AipS1U7IONR
i3xBN0faw6ZGNtyg4qlAtOCeJpzGxywkcnLTxdxwuPrw7WBUrS29Abrp7fC6zoDzyGbVFzI9vn+y
uTb8J+ljEoPZ2Ya6UGLoPG3yONDxp2rCoFaZnl+YqzS3RAaG/hl+6RtI0p6cFcvrZ6iVrO4OBK3l
BmQ+7EONp9a7u9UOHgArzIf0gS/oqdwjF+TFTaRuD03hi7UWRmVt8HiJ2yroFMsSUAmc7Qu02uAl
8eQYITEHkwrEFoiorfH8cr9PfGUnGQ9kxtOF3IeaVIOgP2nPyUUBIQ+OjNEpFO3oZkQjV1JyQfrT
Sd0rPaMhBLFswwd7PmiUlQJd71t6hLsJ5WRDGLiTFXFS+/e6+DhpoRuptDv2Ua9XXw/OuV2xqJb4
ul6h3HphaQ7rjZZgNzyp9Iyl/F2PZPhGWSuolX01U3AAANVP8YwiRht1X0CfTgow3yjK7Cg6ZKUa
LYS3065pH5oyDjYj7+IUTGN6okKpSFTAnOO0CDIXQ1fY78ka9/xFTplTSDPtmVytFNJfKKNkslkH
bY3qWIclP0Yx1/4Wdb85BnGhG0XdESGMA1c0+PU//KTBfaj264bDJ8Fzd21abFE0Ax6v4A1BHPB6
zKca5hTg2HZBnu36XCytXxBMm8esSHrk9H65QPy6FGGd7+2JaVulfTzYzfipocj60LCXPNSzF9KC
7dqEPLE8gSQaTAijxfJNUTFe2VCTm0VMQabJc5UTPrtj7aSCojxvYw6XcRxRKuHf039Dwf6xxWQb
d4eW0VfdFZkdhpqNtmABa3XkFr1mmFJgfksCBcbrBOh7koZy0s+HDAkQmc/+/F/glpNV/YKslxia
h9pqnJBy5uUsTDqcouvO/Nzkg5Hzp9NHWzj0bFp+0I8sJNIbMBHKkh3fJ0FxCmhLtkFdkh3DZqci
VgTrotBewIlDyUcgv0sOKsd5pQSIGLylf4ito9LTxrIcbGyJY7uE2KPVqGHt1yaby6cCid4oNAB+
L6hu5NIFC5YTObT44a8HhO1knd+bhcgidxGC1j+TzXBe+tepb947ABAEIt5jg3/0it/k8966cJtE
jEAfFjIJfi5ls9RHPl8F3rDKHoTRuGvfpDKqy3AEC2wkgWZCL2ePN+VJxCPbzXxhDy1J/FqXnjOF
ZpMZGLkbvypltWHDioBBEGsyNkmu6udyph+9WPst4ug5srw+D8XLoOM6kzPEnphRxEkymV6cs6hP
+qf+P57D1LF9ofDr2R/KMUZAzxqck96jjxByuOdwJz5jqf0ZBlcwAhW6QIWJfN24mx51ZnAX7aEo
nMt/JZ3/tBQe87hgWUJe3ZHQF9tSrzQ0LgFTmroG3e1t5eK8+0F5XR2WAaFQnhwIY2dWROJXWGWz
m07xzvIGWJIOwchfWNeollKda8UB5jY9wzqlDfgBvx3TiveObd6tvYdU5G8YGU6sBVwRDNCpan8l
w0o4amQU2YRohtYHPVrm0EM9XuET2awbBjRvkTAqPBkZC6QVKUeHrhi0EnVx1IzRNfWlD+oAeym5
T43neeOqu11HRLCBVX9mBQgPsAi0fW4sGOAk43a19TaBTbE+mazMq1z1+0+G6u4a9H+3rsJqTOBP
/BuMjo/FKE23bFAZXg1K1qhVp7lg0s5Ouzhoar75Oz3VbNJYjVSQFkahFUU8oNFpDLY18MVr41Tp
PoZEXQw4JL6+D55pBhVtYuJOhMC9AIKgkZen5qOKYA7bIcYfxKNg1Iz3f2ajw9eG8r9QXwk+5ac+
UNp7Ly7Hov5by22aU6trTlZ3yRzR3JJDndoLEr4Cn5HcKfky+CXiy8Xb33dzqKTIJTEOPFMKdzgA
t25N7zhnlR6Xsn3L9IJezC0yP5ZrSbntdiVuP0BO8K3cvGQTTAF5uAlbRqa+votI0I7Fvh46yEk/
2isaF7sVDUnwwrRLdJcXhgy21hMu9R2ajxAecYK+6nDHsBSksZD+Xi70IHXJzJFxAXJVatR9bA66
RSBCGZDBAeue/iyeb3PgRY9lGHNLToptRwfoYjYmpP0rf7Iaz2/N76lYclveNO+z/XuXUA3fampO
2DqHk3IOeOZ00aEd1NNr71BhAtA7YMHeOxYWx0txIZTx7p69oWyLZ4H1uvhmKa1QI/QBuNY7K3N2
ZG5UdcQocFFekm/v0KyEjFlaxjM9ZpxLpStrbmexK++XxQxNgiImeyoaT5Ou3jzo8seJAjpVNBqe
qthsaR7t5o+mOcSK2PC2bY8wj1zwNLQUcaQz6ibHcHqdObNaSrjGy0ji8EEHw42J1dcHbfHUwnHn
kAyCFY0aKHbkRTqAk3NsehxsSZoUYgavryXaJXmzcDeaLcmJsC9MvqFf7Tr+7pm8Lgq5NSjM5MX1
eozdhDig5euN8RmYWpCl7oe2InViTUUCpIdgSlnylSAsoo2iNO46vgI2BSFFwYv9MBSUHkj3rkLL
e9lWy9dZl2X780iIC6i7PMX3ylVNGqQH5oI0OtczMj7wWl3B5CNjMGwjT/BX1Q6Ws3N3qrDYAbAs
cfhYxZAFeVkMl3Y1HOI+9+gTZ5ddI18FtnMiagxnQmQbuRVRCeVZPFSrk25mvn7X+UhVot4me77Y
MF8RPRzkgdKWEcp4bgSJhWQ3DlrG5O2nMz4TUmH5DATXxXZ+tdBdXTUnaz0LD0H5OXCcjOLoO1Kp
ozjqJArgsx4uI/Khqqwx6rsY8qZWlH+Vm6gjkZuY4MEMM/VE5DMgO8RjAUsr4eUvLYghWh/0g3eU
CYl5oSKsdBHjlqzYecup2dRTAHwLqwZs1N5+zeL63fiFWy6CM0iDVmedMHAe3AnR68LUE+eUSrrB
WW5cUkmmyVCBsrsJgZWj15wn1cCFDOPR5uEcp65E2EVG8B5OKABN7oHeFsp0cXRJ00EcWiZj4TVA
g1meLipnTQS5yVSBjDI1QsEKp8wpbOjpYNmYHCfe7UWbDhYFZhCDrt6vOy73jiZRdqhyYPqz8wvv
2yeuXqvW+dPfK9ebBEnop9PWTbfx2Z25nE9LDR4QFuV6jp0e3eYes6wZN8wncU9DazUwVVH5Pl8v
Q/1ISIYmIHH8SOnxlu+wi7qzwEx1oBbGD0DwHpdGOjulL8SApMxQETnESscgbWl/QfiaN53Naf6I
ag3DRMxyefajXDmuc8nJB7YVhSGoX9ddQGiejcXQtT4/ha0KcHj8EGgi9HUuQi4pB5tt5xSg+4+E
6z/mUr3+IP7ywU2Nt5YQ6RqOeeo/V1RD4DymCxpCoha7GmbLrMGPYIM7VDwKKfRbFX7m7sZyUAR/
jYeayRGseDZ2V71FpL2v08EfmmX1vx3hg5IEkDjvDzL+7O1BQAkqKHbBanRAfospAUzLBS7bykFC
ahGL88O/9Em1QXAzOr5GpcIxE+74ywlMzvfAqbHQX2z7zSZJ83v58T3xspTzeH6DvtahXK/5ACTB
1fm/pYJeJqVbE/RSy8Zch5R+Z1Otdv1L7/g+hFXfipFQ+lY18oGpSKLOzQjzj4Vv2jpRUasdFHoS
T/HvZoHnB2rGr7slUpyRehMzv5Wd9fnJA/neB5++Qt986ALrRyBCSRz50PoiTmOiYn3zHYSodGaG
YuBn0xl7rNICXiDGRt84vI7PTH8oNV+cFoZxDEq5EDmsvKZdv2nwromd7SDMwv6lJjLKQyOTtuOy
DBzq7dj/7L4yj68RqhXckNGLKHBqMfd43xlH9CXyG9275Rze9eNpQ+HSDHPUM6+pjRw961cgfQQ4
LwYcIDQ4sgYX0TAzD95Ob28wDtHuCbF4lJK0lbQu/mJJv9fTIP7/UaBEwaS/JxCgAIH01DjZOY3v
jbLOWusQNEJd5K3bfA6X3akq6xhcD2rCptrATJTcvK3xjvSBMnIJgJjBQ4sGP747peXmVkivOkh3
2kWTAZ/DgHH3Dyn4BiEcIMsEphFqfELAB3qvs9TaFsTtsdsCZkt7qSsteDTz4iVh6d2r/Djv0SF+
iSjiSsVLhTURrDUS97Sxsy3y2SezbdUX5u7c8XsEWLSdMBRW0yVR8yBkY9/OPOYFR3uwpbgqRYgS
CUGSTA82kmIO+ZmlyesUYcp8txWhEwq69OqCqpLLYpBf0LEKQlwzvLVD1AVjbPZPPPt5Ygg/E1rs
5LngFIzN+Im+uK5iGJ+1FGHRZgVKs5gEjVjiMuJQzqUOkD/79xbnmRxuePlCSS0zRG0tSpVPDHe1
XV+8RRwRmiI7jmsH8IX5fhpPgMOUrOBG8BXsr1cpDfFIuyZ3RgirFdj1Pq3SnoXGtXc95HMkGsBr
ZALpC/XEYig33ScXC+BYsCkyI8OFtL9OTQ7rK6xbb7TO6Za+lJ31Wmhpr7WIxbpz9gRCqd7D29t6
edEVhC2au42QdEFBrClMoeoL7KGUd5iPCK6bDouAK5gP6K4C6lIdhW/G0DAVaivVRlrViQlcc3lj
isGhrfNrM9O0HcfJt6ALUjdQRLVxH0BqVBMKKoDMOCMPtHWsh3246eU7KJZ/vXbZsJO20ewFzKYA
LVBE7NPLzQQ6Eel7OBaeHZN2G2qMMZSIfUmqx2SR3J+Nn7SeV3oRnHyy6JJ8tgIpn2gUSp3Hslsa
XVHtM7D6gt6FWTOWtsGDL734kDC73NLWYRdqYUydHi616CwVGZGplk8MPVqOnncMX2416pGOfzt5
XvWt1bXafrj6Z5UHUsS4UwBoDuqOLz2K91fJcY/nVfG80VphKbtNpmxWGULYvPh7zR4SIiyxltxA
OKuOwK7FkcpPKdRm+9rrLWecUZVZLFUvTEn/8ImsBvwL+GtADGCRXH03Jt9UApVu2s0IeRqkRVm2
XpqP8B14ODyv8Zps04JJil6RGxZUOQz0btY5Z7an46CgTDVqXSgKpKOZTeOVrUDsfP+1cgorrNde
FVijct5L+wG5HYXsUPdjgjP+pUzwYgUdHIvFx7PofZBTHIUse7OeS/DTZ0J8bx6jrd/uJBogSfWD
zSWdyTaNvB7vbPYImIvz/ZgVlLgBdCMJV758B85NGO/xiTTyckpLDIlz+IytwIEQzbBIBV1ft8kb
5SW9QyUThVok/zfWUIojCRFkvImCJ4FNopS6I7zwcYMoihmwyXrmmHsPkmbG5snO2byxtFMajByx
koRQ6jDBSkVxt0TANYGISh+D9P8g8dQMV6njm3/SMdrjJGwDGl52cOqTvQBu/kGdmuY8JEYD3+ch
jDpIncQqMbajiLcPXWLIxMsgfewA3RvtPyMCUCIRg3spFNwE1CgPCriWHmCYcYOhx8m6105XwICs
E+4T6CKnIfnkxFOM5B/xjTOC2OJfNxuj36nVjTFrmLAl3vHbqPwHdWW5kta22+ijCGXUNFHM906z
LSS6q/B6WCHPH6rETP+hZBLvKnIQ91uxvIpJhADFXdYyxp29+cNrhQIrJHnBATuPAMd77EbBX4Qi
tBZn9intYoD4JyLp+Qr1j9DaAxenBqLdsS7FPvL4m11qb1fJqhR9a0xo7gyN+7GzGGxgIpz4D9Sl
oZBG6b3v5gfpEoBZeObVBVNdGt9bxPWNaQJ96UqDcED9z0XayAtAeT9DJQ9BTsD0yES7Toq9SgGu
VcL7/oybixmOhVP1Tf53AZHwVJ/hOB3tSlWsEj7cR+EihuTbcYmsr4THsj0iOnCYMvl2uPGgcJt+
ORMNPcx+YSsKFUHpoTi7My9f4IGOlQmHEo5zl3T/763mKJN05h6D35tUCz03hW1iQe/gLN21hVaa
fe/9+mtZLC/z7MyiHcf/oYCWA9SOm1Y/Yq05EN7fEgskiOTTNYGtdqxqpnvJz/bmjWDbvJL1Usx9
wAyH4apsLthFJNpqPapVOoESb9/DCqGUeAmVMMbBUbepFsuIFzuJ76V/BK4mPFeTJn068vPrk3Ni
O20ncUjzkWID2ThCpBWulWkqSIyKObXiHEyEaOQOOB2LwaVAi04lKUVoWKI9/5S1/zyAiKs4wfxf
cZ2U/wNZHweQv1WnNHRb5dE9cOIElWhIYRwg5cdYK0BOUS6C0UDSe+SZE8wjCvzqdlcOKjZrSfaE
sk9visa14evy/+cSAZdy5jjPNxYtitdiQ+laLmUuUeMJ516bb/Kd843Ype8dyDbxavCgHavoWb1p
vegKqf1g2OSRPNtxX7/jBdVrcCIQhlYSK3d3CP3GjPabt67ykBhWBidAjo3ybTcXD3O18CzzmTD3
OOkh/MKgGWpmqFVV8B7j+2kiK2HkbZNbTMAesPNA350fMYJ1PBBra3Xd3FfC8JgS/B/MEAj0vCkA
vn5J16SzJ8cZhf8ldUk40dSqO0+92n6QPiiMb/qOTXuEb0ScyI32ImL5Tf+ESBf+OWP3DAnjAYE4
WzzsUM8B8pRGWbfLZxTnxB5x41bmL17i2+GLVUj6kVZ+ABQqOhFeeITX7eouB57oW1ku7CIs5wDO
rsGpK9h5MDau9jruOmz/P6oxna3MDt2AMRTQ1/+yC13iOODTIU8TDwcFxg9UQHmrd51N2KURerlC
q8C0wI1wbayxEGSp4Uj1cSoQ5m4BsOgLxZ5SrW1ztryDNdclSwaOJIkgtS4dayfHFaPCRL/MjhI7
fLaTZb+Xp54E6yZ/3katXn/4kBuZRPvb0v/7BpczOCAjaQpLZtup/rw+/lZHQs6dug0U3tRUUlkd
0KhVgI8BMvV8wvJwxjwOilzRCIHgiQ7arDjkXJh/a5+SCJkJHaPZ2VRc8br9RIt3P5f3WG2b+yGL
9IXtgPt7Oo91w5OWf9YmhyvioerSs6ERGIrpdOrU5Tgv7lTHu7FWQO+FaFzgVKON6omVEC5C8Axy
/inyuQQgmmRSfgaROvqcCuAtymn6uCRmzNFnSAbFRmzJ7X6mFnHxMnDsPHttLSlFp61mbMwidG4Q
fn43H/s1vA6BDd5rJfQzVxOEcLTnFwd2rs01mZiNGJ7kRvZ6KjcPzaREwqc33gYdGhxwRpAEW086
Ww3X02UMt3kuUXOCEoeGr9c2+mgVLHir8YPlfT/DOKYBJDyDNxMwfbU3VNA1joodKJsY8jmN7JbU
9fjiuNZkghZRrqSn/c4DlrXCKajFhICbep4l96hN18gVzFw5dTBViPSa9+ENYNcjVUD+TrX52nyP
mvsmb6C7Cus3R7XWKIAMYHPJMfJSlHzw/Y0vHPcyfSYELE8wrJqI9rtTd0I86QwRCIbqw1gyfNnj
kuSkUcaN5bsHqwRMYGeveP3Kwxa5oJNfW7wCpEACY2NpdzX8BGMKxSdNrCBAwfbQkED6dO1vogX8
Hxj9fzwC0um71D7cFeGcsygDepMIgU8ZYfjMMgMoPjmCkBTNcppXS/oZyjjIWFAahEy+BSIp+DRo
2VpABvewVqdfwYZzoaxs67ak4hQbXDCi+W6VlT492mevyeb6FKYrxmlS+iaLNaGXWSKRPAdGYkIM
IaF8ELC0RaUeL0NYcaThb89hS6dQ4d3lldiZYNP4twnaV65IONMLDDMJC2lvQlQd3iB9YPZOGOkY
l5Ids6jceZxTs76M/xdF3Wg24dvahQ6gZV93wA93FMER0rlib8lAlpPELeo2LuXWErxVyA3k2eCE
FyfiGaOctKifjjM4DxOHtql5+tRyFhzZaI4TIUzO3b1+qX3yW0nKSF2BQWLFzd9ZgaRW99K6HYnV
TlZiyksGi8qBhRwbnixCvrWr0TKTg/TKjuK/05DSC1aZTFoY9naaZjrNNu3CRXWhTBPp57SaHEdJ
9G8HKKOX7GZt3pMeDmlJzrBbnfKUUvBSVE9mQLSfulm6qDd03cEkli+/Q7yMLyAZ4PiaRHiUE0kR
vqM9x4UuQHsupqX3HYYyLQzWFR28yuzmqaMeGC3IYAu5eEKckfm2qGid16COM9MGj76vR1adAArc
q9/6cti0Qa5gfi2XALuW+k3QT6q6xnFUmXqqWR4lz/UC9f/KV0q11TS41XgukgsLIN0r1EkrxNpo
wuBVUDTw+Sv0RRPv76zVqhWgJHaeao5li6o63LPl7rVTNb3gNlM/ARjoQYMgg50UgivgWkzBxdzr
7T5nqaWFzJ2lTWos86q8clfiUbIFZFvzvvvWJkbj0tS2iINLXu9BREvB3zl33RxX/kzwKj5UJCsp
GIBhSgOW0WMOEXF3Nl6Sa1mU/wy3ry72ElkGOL6Mx+dh1MjkOn1puIfr6LEvXQNdG2ZmjC5yRi11
YOrZOVS5fWle2jEiM6n4VFJeXtCKyusbhTys15bapfGAOBhVsEZWi9GiVZoIX0K/w7Kb1M74lGN+
/zpQwJlC2107fqzhgCkwAIF/+cqd+pDe6r/WY+NV+MSF0/+Cd99zE+nTV3YrEBQtvRxHnPKvSD8/
yV+jUGHiw8BhF+PGh+e+MoWsLYQs8ykJFzLcOMhjznEHRctuKBetbIYweuOTg+7MUOeWnFPACsXB
JkucR6XWEbpvEd2YONfgVa0tp2VR/u2lM7iXwjoTdVLLSG8di9YeCsAF8fKdfu9VBRGxmneXaZxm
rWVFwCpwvmfHaZGZi4Zkda3FfdY0fin6yu3IVGN/8sAftBL2VpHSq1RpvtOobXd9AMvcMC4VYkYw
KIvzlpVFzXKPAOt6URXQ7YCRAAF0EVHslsLVtTMpM40bWECPXm5BG8A9UW0x6crtrGOTEv9yr+ZB
did7MosW3K8ZIPL53mxas7MpXxgAXNaYdwi0rBcioLvUvm0EGDHcEtL/TradYKtj6aygkxNYdH+k
Zx3PNESUwUhhyr3O8tqX5AVH46YZh1Ee9G4QRJuhHj9bmeDj4W62Pycj8hq82DH/uqFEcGP1QADW
pARal/ijckyjpunFfYivg+XqmliewFipq/RriwdZisn362VDwZLyLsyA8ITCxRsXCaIKt474X4cq
/CMCxW/9Hlg44VIB1sjqrrC08dFU/o/W5i92NnLyBtozlhsxNDD22eyryZbx3+vNR8Gq6Et+7wVR
aqYtzhWQnlKuaENhymw/x0N4pfwjiSVeQCcZTCwVsCEEZ3vyPZ9S0enjj/HxJMv2q0K8CFgA9NP3
F/sUOL/XDFaxKDT02nQonsyqc2sjd7Tyv1KtZG7iB3HxzS7QO5tX//FPqquDD3N67nedy8QyxHyT
GEIc553L5GdZWa+oW4RvKSd5DHJNZkrMLmhz2Uy0jfT32+o8FA7ct9HdggKUFwh0110uS/z/WuQp
2iLlVRGqE829VZ1Emp18aZP98jRtJDjIveqIZigKdPjJPkzqiIUYnarsJvXiuAety32nxuJQSYz+
TeLXQnzUt3VGKDcoCwfPOSisdpj863R3KZoynipk+umoJzlyzVsR1X2AoRQbvSj0V3v+JisIqRuc
kzLZhO3eu1hajihqpuLyM1bYLwBUA/+lRET7b/HaonS6Wk7uNj5AiX+Loiv/TIGVhwudhWrEOw8N
4kKwlZncnEmBvJJLZ2cS+mDbS+AyTSFRW07bTcKbOv+YBKWqMl0IQ4T+SGt0wPn7Kr16y6so1b5U
oQrhILPW/RrSaFsi/z/1L3y/kfppH68z4pJTdXPgcTGfBGqcWmLp59K1p2uIKqSGfddYMJNKIIqs
trfYNx2gTEC9x1n086p/6quq5uMd+qwPT1UKK1hpqy8XfvC6JAqaWM4i5R6FBbRzQJSr37fkej5S
5YddPWkxoQrNExIITsO1pmwnoKay19J0lrN25BQe9aIUmjPYGPRmToz3GbW0BewfJSNtAWZh0WF7
EZpyez43Q4kkJebF13fwTtr1gmHi+fN84cR7Yz8eekv/lbyN1WS5OdyRmtcydNxqZ54ftJ/DQrRM
9q+TVOGuMU6Djawi3yar5U4zFad/idHxVsvBAhuGnGw3UWZqqe9AF9ITWrhn9iR39Y+41+2KVxHl
H5z3A+JfVj+YUE2nCVJAkYa2sSSc//VhGTf8RddS4IKmPgkydpDELfpy1uVYmN+/x1yoBThVYprR
pBRwmYrT3v56gfZV+1b39NXoIvCA+3QCujxmDU57KTJDHcjB8RsbwXymMeWgliyHWi+jhM8MlGhu
f2zSfe8/heWXY8yDhxBL+xvE1LElreD5BSjQ4g31bDWkIW8hnzd/x0uV+bZ2NmM4T8Z9Iw0NlsCx
jWlDuBbZ+XVPRT3SF/wtVrpG8oapTz4hI2o01q0+a/3HRCta/TsBCZViOo6wTBFgevJklsDWkE3N
HEQPzPpWOCBbDSyBDv5/NXMnYm/psMvqRV56VWm8VppUNBMGeaiJhM0Ox/SxLDu9qjBpKmkbXjyt
EytOWQf8WOZzitI4gXO1uBb+Gau2td7IRJ9d5QH4YO8iy4HueJJwqF2K7E5eTBzEfpjt1f8v9mtB
JJPc+apyRMuEAbcQC/UQ8cuHZluSuUytYjqCjRieIqCuGmfuIo6D0uZgtKvWGRu2gVzDE0l/pHEI
26iWfTTQHL5EnpiA8++yRRox1uPPvwd82441+eLGldIA8RTfS+pxa29EquRwGWz2VctsD8cf7daj
rqMcfkpgUVEWRCRaaZ0uLDqvfsPnXhm312oiC/K55cDPpy6ON6EjNnbOdlpjxk53iKeIsQK9IWCD
kmsGqFW3qnSXyDi/IseL+CpoPfPrfUSJi/Tkji6AWDUJO+uU0Xoie5tFfgCn1B6T5qE+XqR+hCYA
P1cLiouDmMrnnDN2M8AhSmDeFdQrLfPS1IIG2jSMuT35w20QMetGtY2GgAHYpEkDE8fe8gSH1aSn
As6GZ9KLf8eWxCtXrQBMIaJovkY5ZyJCXbvjteaVEhQnIel39ujXPjRTTE7osxHLaRUS0xC+CZ2d
uwes8mCEq5Int6KhcVDOWUxHF0i30doIz09WOZXF34/vAjZwQLuWwziZdGxRO4syoMzMBpYTAnth
NK2e68AgwdNgLESKocvXQDxuWis3xGB1LW9LETq26MbjfcB1sO7XSgo1busDobkem7EJ7CumR0/e
k56BHEirVAg+nYEezQ4TyThAsoDADk3CCb0aZHZ1xyw74PDJsl5WOG0vX2iMSPckmCzUk7nOHSFo
tg+1+7mB5T7jFGKB2qq+a12GhjqNvbNM2US/+jTnWnUjSJ6QcDgpIA9YoW1erfABYF3bFs9Rxor3
McJ9QEpD8ub7mvCRTGdIs5J+ork6VYKe2JQEAnZzYyLqTWZyeDquP/yRIaKrlHQwZfThC/tp8PgK
OMH/WIL3kxR2s07BOvZdGmxOV0Ylsr4FPcqA56sHwfQExtdZYPWS41t6Rv4D4P2UjBNfptQBror3
aCGwGW6gtKNbbE2JF81HoROQeVExZfbX8xlFhmMOmONK8MDi0kWV1ikNgFR/6PM+bWpGNf9r6d7d
9DsJesH1dL+Jrm2tLoIWf5zXKE9XA0U+bAA0l0bJEEmA+HXIuB6Zvq+znFf0BHiwwSIHYurFgAyc
RPwdYBQo+vYLrdSTJOE5pirVRHV0/ppK+OsF3hS9KkeC3NOdWJXoIIQjqa17mwhPTqG8SaoAb7Tl
5SCaNuKnaDSD+ASgc/2SY0abpUXgj7Z71bc8F1EsrIYuZsmLd287AH25AFpbbl3vQVLVRgfHjb6L
UxumxXcXEoIpJ3kJu7EWMnOlMEbgwo9C5L00seiDTvOF+s4lhO2wcfdWsF5+rDHJbNr4ObFHPVYJ
eJtnemvfqRv6yqIU0DrpiFQdAddUzwon+f8R76WZHUofiVJI4RRg6DtAjRTT+APbpdBIU9STJbNW
LzPX3uplEk4xlj+ebfEJAZTUlTh3CPeNAmVr/Wm0xD0JpzJLY5kl5u840p6QpPfxhLXdbWYOhyni
MCMiUHs62qPlOdNptNUqVIottU1DqwID/bUxbPVt+ip9Qz8aOJP0ksVl8Yfk/RjWWVmuOG2Wx+as
uAjHC0lEZFUfJ5oRNBj7+HboNIu9y+vvXyi7o/yEEJgKaUgUP6iPOO70/w9cS6SXVNFn43NsbzVz
v5ezMekgqxGO8n+s+9eb6XEyDz1zhhS2ZfqTBXtT8gyx9fBflmcEO/a9FimTMnBfX4it/0LQNin8
HF6Rj/K5s0Lj5/A4+33h8reNmsDj4VoFWVMFL/awGuYBE9n7zR/dnyMibHln3OewLwLLSVnJqXMt
efLvFzgElBleescYn9hI/+R8gYFdIcndPHdJyfuChwS942/bbg98q4W5fWBOgIVsnEGmhx3u5vHr
d5QJkYtCvmQbWofvgoYP5y5Gb65nZN/a2UnBt14Vjy5ra47jqsWs0gsm5ENFD9A+V305NxEsMRKG
RRXt6W7L5hUUtcNQVdnThg5FYw6qSmxMyrupqCYOtxDWgz77ckci+mNU23RxGo1Tnndeiu0wpKKt
kW84ikaa3LcahhErQHeT4yzC/cBl7JyQrdn6mLpobZEoLO1OvAWqQWKVetSGxVLcSGIT6hlEYgNP
k49e+ariJR37RBDlryIFs56UaRQr7v4RPEp+Kdpd8SOSz3z5ThSRnCRhsA2TNMSBHHOwT9vFl7Mn
a3bSk99hQLi8oiyIwlvZOK5iSg7YKEcFHtI8zfAFfGaCHcl1BxAcGdjkm45WvsX5/FmYXWA1A/8+
Fv+3wUvYxfbrXzLxV5JkuQYcysdo1hZM8Nqp/ryA7Xh0kPZ2IVK7Rop5XQBtnlIxwwqWvlhvfAnc
YUyxIxRN7fUy+h9bZeQTBOkfVafPOVgu1fsygvViyt22kE4BvaH7h71Vm0j9RwHIAP6BcjCc8/Pu
6o5Sz4MblaJ0gVNJmabFJa+FPOrTcAgZet5Pzy+YhZLtHPkv/snBQnJfaishedyqYQOPHrxAoq4X
5RJrLGO/TuDWkJFRg2+tk5N3yvR6M3VeCOY4yrqapEGq5EdLQae9r3kzw5eCHRoMMRIQGILGOkK9
/cAREic+yESKmgg6/W+8bINNisdl3ka3ZekA8qMXYaP299QlZ2D05af3VBJvjKZF8ySwWYATy7e/
uvMzzYxqstsC8g/AMUp+wHQfEbxxSe2js7JA5r6zOTI5O2okl3249UAfKGPDjjtIjBN/jjSRSZzF
8xG66oF2Rt5fWeFDjkEmu8a/mq5ES5qHEFrtq39E6943F+iy3DUEwKE02UEt8oUvMWkeWBdVWdM9
ZVC8GeUXNHxOgODtnD0DqXEcuVIvcn+wfd01DpRmMXZGC55Uf12PkklHDnN/dQlMkGhrb5vl3Jjr
vpxymLMz3EiBI9Nk6EtaYos0YNeDG/3QY+yi1TMKr7BvtC9M8WTfTc8Y55cF7CEh7IU8BKYHDjYG
IVBrKCRJYjes7VHKnMmBeTFPfjgtUdVf98uPkgBvKW0QiyKkIrmHkMsOFR1chN8ym1lhozGboo0m
fKVEZOJH8vKuLdQTh9TPSq7S4EB0hiN1KbQ6+B2Y24T+wCOHT+QVZERp6tueFE7Xr2IXALzk37Io
CfbDwE76YvTAWQHrU7FhwGYOahTJMBBnPD4YAV314IkYY9H+j0eMUm3LRaX6w8cPClpX81j4Xt+Z
bi7nLgPfO67h5a1VmmH4AhAT1/TlcKm2EhplOIMRpmxbLdizA+l+bbghxzSdLMJdTVoYNdc34rrG
bDXp7xjwlkYb4TJ0TZWk7sxIw2HPAVBzVPXuZv6pZI0MBXGp4HXGRP+zrF2uzrIfEk8BSbShQe3y
kTXWrmQoDP6LTFf5oZ/45LJHWA/B7j7rqH4Qz/PVJTMH7V70gaRkvcb7kR8WLI05d9lZB5l57tiB
BdfoQ10fOy+I7stCc4jFyYueT6rWdv3p5IlynbESmIEVN0hT+Q+yjgVqk4VZdjlBXZkeD7b+zVG9
QZ6NTBUsBSFGm3CnMQDvHoZj+S6fLpi0Jyvq012P0AW7yih6DZugOQqt4a5SjykzsGAaOFm5RBuS
sW7P9Q9+KtAXQN/Ms4sx3B9vEIr/XHxeidYB4rMBe276Vrk0G/2En0hqY05yFJ64xbzbzm4KEXPo
jXBInp7LLKEDSr0cEBS+V04+iQvNGA8brybFQAqS0WXWRG7yVGKfpMVFvAh60tEClSSMR0qyks1M
CvNZUpv54IDsRIrsx8i8VzN+OlR//s0614h5+4ZSPa5X6/fM40FlqzzIM4qtaOt/sVRgURen5WgR
ZX6q66maVj5SdhC/CSa9SPSaO7CXBotdlTxP7mG7ZScD42L8WssQmo9vI6sAhtOVEb7pJlHk50FV
7DgVMyWLfdDxh4qSuATteCp0E2NygdQCcSH1tf5P3CbkVZyMWtRoAbA2rrNyUAknAP4O8YvYR4ok
3YGpxayh1EgTQ6HJwihRjS7XXhxZJfdYuE5LA+0k08W1dqGdnRMiZCuu0AqMWbSlWMvGhN0f48V3
xloAso8AIEgxLLuVN/MvOJlFev4Zq81rWNRjybU+LtT/jrnEIXB/J1FkqBxd9gXeEsetWuJEespj
gPDJn5HpwTf4+60JEz3iSWQFFgBRWsdykkQgEKQj7am7K5pUliHZgvSxc7JPJsx0t3QG7wVRHhmp
cT6TdrF0ilc0UYwlN7IyHxuKaqf6IOsfKwTHl3CLTCyHtqfIlujoLYZ8RUHYqwdU/qJn5auRauOp
Io+JRXjxaS6SYePWLmh5Z7AtT8DZpRjckznEgZ2YAHlPd/QvJsWrdr36dZ2oeMKEWoY4Lko2dNGG
XFpKAUJzvXBv4pEtazNQfB0ZHZCzbJmwnMx8PqiOnVK/DcsNVHA0sO7iXZ/b+h9Kv+721IeN7JX9
TD6rZj3osnS1xt5syriV9G2Ebg5pB3WmOmhUox5v1tTL6e1EDYVlWAueg5TZZPiduNflmq4BGjCL
kCnhC5joa9BAxpOqgjRlJAwa52Y/I2puqDHtGnjNzAA6r7MT40eiIu/VFUcP6A8rJlumlrvzgbZF
ujvcECQDCQCphX1VWjr2Wc3N6LliGZpcWX2JnqBycOqP7gRVPfR30dPbk292HGPAn9LbTfBoguHP
+5Vf3E0bfBV9XI+WdNqTgQnp/QjCe8mjrz7Wr7fpmKoRVkax8eU7xRBZ/ahNIe9xybCpR94NcvhD
FqgfSsJ+LoPN1TRUgjd5irFP92KFuorysac+hK5y6Xa59Rvpj4tzWjCA3iX8ZWpcrSIzLD/9JNzr
YPwVu/BQKtQ6MeSUq+p5p89RJiVzDEEIN6/doF/9Nx2EFT8XZR+e5jEG5EuwgJdy6hjGcTMyIZWs
PG4QtdKyXCqPAEuLqRu92BZ4K8P/Z8S790s92rgNSDg4VDn+IBn9GnB/Vpl74EatEySGzVU6xumr
hMlE+CoUuhs5IuieCAsfYjKajnF0DsTGKC/6za/DFbgTTlEPAawV8LrpKukEuV6PKN/li+AlJbSX
OM+zdC0mJSghcp4gXjsbSd9TYbTlBT5pEAFlWdvoH5dbfvk49rzznXLy+IPRHKNbqik+umoZnu+u
9OyBw12VycwTE40yIf2snWqQL5elP6MMOQEOiWVZa4lUSHxytNJDBxLxWr//AtWksBT9XP8BkwvZ
8u+iB4nTXJEkfmttDr7Rkq7ezoGQ4LF+m6BPtbhw2mVzbRaYvGTJUXbugeMC+UiCf7MSbMGY7mii
pd1OeEjKmSvUexrMGiZVphipvf2ahm8bkLmus5X5nZWUxjsT8nDZHsU1yjq5AmccXStgnaH9RNzj
ARx84OFak+hH53axLliqMYIQkKDKWK4XDiEp26jUM7KOoC7ne/bEwKVZCzkSFS5LOlUISdlMyZ+K
mWKgqYf1csgcpUWmEm84NGNRbZryCrR4xagUX8tSdfaXTtkvTtyxV9OokKNX+4l2GzrxN6hUqz4N
0tOG90fbm4+QJdDc/JlBcLOc7Y3eLl91/vXBLFIfIphL79T8auqSJva0bFsCdBQfqUnjgEdl/Ghv
kbwh/6GQTC7dg0f9hwEG+9Cah4umkCNxdWhDa67cB4uerMHcpxbOlqCAP/bSJmEsKD0JgYOz+WBn
2WnK1z9avd+4C20X0hGnXQr9aJhCdXdU8YPEsXcOGOcT71bBB1h7w+djYBQy52hfmNVOdl4SD4Nf
CAFa0KMl3b+mV2eOEjBDvZP8Z/vdqY4VeoxTomPg88qLlS7gDNHXauaPGCJRry1H3hHL3FZxGuDo
DFGikeI1H4gaIm14/x5HNhRHCeo8S33ny6NHbbIRMAe9oPQP4EChyZkeI9M/mwJibSXfNvH+M2FN
saJYopx64DjZhfzBHVzB3ZqMTLi5rEMmxuTr3rXlmoavkvqse2L5PvkgUCqkYVrPMyo95JfHdPCF
S2F3MVGWmWRcEVqu5wZOJenFqEL+ulkbeOyYsue9YANGRNAN5bLmmHD1cWas9uVURS4SWvTRb+IT
pmHBLfOm0Ttwuq2iLVDtz1C7fl4eqfs751jXsqEhT/vNG+OKepUCI5ONRTk9RswyzvK+lVyy/Qmd
1jHJjlUAkFp2hHCojskUQZqH4AuVlRN4lJ/xuLFZnR4N7/ByVNjVJB8uC6WEFHci9yuFAmJMN5mJ
uyY1BmQL02HNcfKlinIJUW7nWTXJfGJxd4dDRRxNxD2ZZz00F0h3/8x3BxE97DX5k8iYPoMYS3Et
DuVlvo9S2/FZRTLtfr7Rp3YlxzU4EfCS14oDq4PIjzYSbuiZxiD/3LxsmwrbuysP7Kbw7D9wmtyn
nSdX7xAasBTXhrPSgfH4MxqGGpDXeR7z5abHoajpLR/Rk+pMHeCDNtXqZBLCBQCbZZi5pE5VUz+0
OREXpejGvJLu9S28IihclLHhLcGpAsEBRp838A946YSdniBFW6wDiInBm9+NR6//aObK6Ddj/NAL
lkPAlOtOjjJh41WsnlZ9rPPBJg3MdiL4emgHtCZnlyZw2xRrO75bldjIbgyGV3avh+PMLMytU4nn
Nd2UuByBlmBhZcRTIWIVaRG/YN0ScAkc09f5dqCjFH7KP3tE1RT2BVIrcbf6UpMYo/b0n5xY3V6Q
44oAkodu3hw03F3WVvYXEWkt9Nyr/DL7Ll7F/0V71NtCGDX0LVZibk9jQkkFMxdWoOUjCB7B+UfT
UOtBURMqa00tVqKiszP+wfQ00Pf1x3yMQlXNhnvnarKIgb7h3Kr9geCl5raH3tUYixgSW+cOlWyE
h9vRM6iNr8wA4WS62FXsY4Z89Gc4d1ws1qMmiAYsAWjznOv+rwiB80bvdaFNU9nV+6Hx9cLjk80r
/bmNW+yclWyYRaBKDUWAx31R+nG8K+hyRhgh99qm6gv6MkPBAqcN1FfbKIvhjb1+y2XLY7Hg+LnH
fDfX5PVjwUSDFaRpAcwfWdJXxhUXmfPMFMcX3pVWvIQGj6s517lzsh/JJFQQovrwfSfW0czEKwO3
jHBrpAHmdEcC6+WJNezrXM/oCtOMEo+yQmpzB45TYXAICHG1mh5fBpP76A0JgiydyWCB9Rob0PUA
9trGFSrE2W3C3hDj7K9JcOu9UjYTX4eAb+uXeRLGiOHZRashY4Te6lZVTpk9RKUffXuEsstsCJVR
i65yErUT9ojTRNr5733qyC9ZOt4FDWjVXxwRV14F/kWQcuJtjBjs+t+GVX3ntGJefLmz8Q4w3JpD
dbnBSFPMrotRgMkTsRM5wK3bVXsuaJypeVzbEISL6m/9yfdT09/TkT2XoeaPHHY1W3gdrGLXsGnz
WuOGIbYhgpU8yrVWR1ZQkaCFeMKeA9ICVvpKaEWwlqtfQxRdNzDvFPjGE3IjgLqGnVSd646o1K9I
48wQc5u3oMfpeJtNRQGrQzT783YLmZdxCXD1yQ2eH3DNtrtYzkwKmstRF9xJFb+O5+RGVdMSil3o
swdd8BJul1jsPOXX1h/U8afn7Bpc89D5UkiVXE38Bl7fjYyvb9F/O5qkni2n9L702d2SEMiSNsh6
rcDN2Jw7CVxFrMOAo7cE3X6fWWd7ajXNydizW7bc/+pMAFeTQsXbSSFx6+4mXevoq3lnZJ1g7XJE
C77+mjm5fgw05E/w6cvIqh2c4VcXCWI8Fh0ZACUt4QobMFhIgZrFASKlPEmFsT11E37Hlvce0e4e
HHsDTaPJudWdU1ERHQN6M2LjExud5T6qVuYCsgyKxUTqKb5hvagVx15kSmMfpzb2BYiev6arF3qt
cWOmksUh0++TLynfIwgNPukgkcV7xw/av83Qat879lxQJ6iI0euDwjdyy4Upoux/YTGtJvjr3hnw
78k4xsdJQOyCNMdCRdMP3zNRhoJMaX3PsHs4i5e52JXOZUVKaVbTHPpk0eWYUd4LGf1ngv9GwSyh
a0T2Rqp74DFESI9zvcEvDN7EjdXU0Nk+ZAmV3dn62PRa5mvGa0R0PSi1ETg4Tlfo60y4db3kSPMq
2OJXusHFI3/vfgjwzWJCjouKo8tfkt6ZfZ0xDBZnzBwHgah4IjjLZ4kCACRssrVSJC3AAyX6w6nj
kjNvu1ttdLfJ4aq6HTU58Y+/Ftlg4RSVZ8ucZTunwj7WENEzDXB+E7fdQAA1oTIsWovT2suXEI2v
PTbeRJ2//ZAO8akd69LF9F6Ps5U8ZM3QDuqSB50z73+rQ5LDExe+D+agiCvix5KqNE9zeCueMO55
C+w8JQg5nCdH8pFBv0BlD6HRRBAZfUzt/d2kzTSq5FAca1wBQuIyqRN2biMoZTbMN87nAqxG7u1F
Dcbuq4GCZLNyk6aYXH+U8EPeQjyx5rFgYKX93ZACeNrS0j2L6Cj6dal0iMMXsuUDkdjn6ry2LOI2
Nx+/XR7EO+V4VmUOpjRDKju0neRxqzJyUmgowy52bt+w2Jk8P1gIi9EZdwKDZbTmQkGlKJK2d86z
MKvhssPwuyNeCRIY8pDUMAPsPq9hMLGCejhHKc+vWxMMXtQ9zEzrZ4WUenfMQ176oltgvHmv3bmV
nmUFTtm8H3/twhvcvZbRxvd1P1tpbADlXj8Ljv2ZYxAprnGd4sFE4vkjHt2Jtwb7ncBkMXu3NH5i
xP8RINVMBev2wpNESlGdPQcs+NbTR/myF/UsngSdCDW2CON9CVRLW8U8kkhgdKOiJ8XnmMFOcs2J
acl2NZfjz3fgmc09QqgvVDwYMs9ysVGLB3F5jV024aXL5/Kkyj5CB0GECZjXIKdm7b7dbWiJ7oY8
QEIQOIt8zs8XIL5awNU12QM1exAt8bINscujMTTDj2R6/IWEmcP/w2+/141AAV3A60/HkFEo+wRJ
eBdBI2iKLaPDfhNYOw0JgalVIEmYH8Zb12cKr0udvRLVSksBQIfA57TOEA1MW8FtvkH0GXfrPWBq
86IS2LTEYdBSbQs4nG3YFUgC3+/REpCc6KHZPawz4QcBERNDku59yVkN0kTB2YadXNqSyG3sCGCF
u5BUpHJ5Az8VgPKu+z83e6OCgYvGAI/hvfjeJh4BlQgDZc5YnJWHKkbqdp+GRPCl0YO4K0BZnZnX
s7FKsKCMdBZP96T8DziC8iPv85xpCSKcgrmSxHgN/rma+tyECNuPDpbqloqokhBYNoC0GEbUEzeF
JRot5vaHsppNvyOs0+ZdKT45qZk2oFHc1twFaxPSvAW3o3pvXi4twwQalA+cqT+W+zP60ViS831e
tuLijqm6RCichF8hSGN4/DvTwvGZVcTrhO9A0sLNZYNYtUdAsEduNLgqk9MOUdcP6svciyc4/wMP
w5CLMUYsX0aigTE8TKZbW+hqn8y2iXoAkUCKmPl/uy0dckwYRO2txUTd+ga438FBroItO1GH6vWe
ERqLDmSBOLWk6Dq+yan0n/TQg4vF6fnfiC+ItVmglEHR94rHn6LvMOq44WOEQXn2OvxK3/irR5uE
oQS133I6FWstUTdTZYgJA4gnpz8gUFZOrEQxzvF+s2lDXB4019395vl0a8nUuE9Thudm8og/3U+Z
SfV7Ooayvs4nY8ABoe1G4iiAJ7pmb1YICoCE7/+jjy2291/tLZUGDHGiNEtnDmWBaUx0gchBXAt2
zw5aFNIkw5MvNz+s9u1kXvG6t9ZWXt+8XrZyCIwe+oopbOpLyJ//F9wZN+iVhL0hcQNi4AHakTEL
f0zMRObmPdqubUXd1fdB/6ya/DJ9OMcCmo0h5mLnc0/Gghcb7yYCMD9tfP3vDG/oPsb2WKoQAUQx
UyHbEtk3zLb9PEyGzkxF6j9Fg/XybefMGupeYmhB4uoRRin8qZfXYNG8gUaSOh05uvd1niKiiZrM
j92ho0oNljdFqpTDnM6Fjwj1bdRvEtezQc/WdyVyazsS/itzxyqMpKuvIZJsS656uhDCGfSYdX5/
MyRIkTaE3w5y3+ysa7QqB8Z7tumUExJO+o+Ekulu9PGAsy8y8M5FKuINqKxqavpd9nZraQAd2vz2
P1sO9ablHFfQYIomR7mq31l7pQdfKB9M7Yhlgcve1pLpgqbNVICiF0I6EC3CN9QH0Yg+cjRSgDvk
DCdiLm85rHN4gR/IN2uxWMazAR6vhuO/X+HpJd6TVmMLk8p/xfWyn5AduflsYjRlVE3C6sn8NZfj
ST1rZmoMdQPF12IYMMhYQ29l8uSAKrIUN19lVLlJ3aORKvAiizUJLqGDTxWAbRN1cYnieYSN2jdo
Aowtu0j+TlkjuinAsTrdtcMCAy88vFpvPmgQ7yGGS+wzS9Kpo3TbIsHreENblzhkCyCBEmTlwwcf
cyhQhowdmuCkxfDH1SF+q9Mdiuznl26zqcW3lNavQQ5GCHXOiW+4iXoLV0U2OeMdd3XIWPVUyRrj
YWJmxowyYLPMBbpiugf5W+DzoKfN/JWdmvgxWbo3uvynaw6dHrycRirhC1D4oi0eYtJaGAY8nf58
3uNn+GRiy8++sG2Z31D/+DAAuX7bXRfkNQgyHH9VAwmC6gzVbG5p4wLCtaA/EA5cF8lt1oyrH93Q
4OoXDVExSOjSVi85BYnU3lLir77RXOU8+s4itEyEZi0VH35sNC82agpKxpVz3w8rap84CDrwrwQo
OiNPPaopnbOlnqZuHq95itOM/au4XzF7sKFkMMKa7LJZ7KWPDj/NJWOd9WxcvwF4nkskafDSrjBG
KbLxp8BC0zeMR/4jUZW4HZ8loEP0vvpPenDH4Ze9l8i5JDMi+ZzLR3n2GaZHri2BWroBvQE4gSoo
ee5EUOZXvtNEn9lJPNiHsoavHnzZMZqZUT7+qTAP8JPcofDw7+WxqVgXgZDEkUZYTT/G9fPtvK45
+NVJRYFvdKr2sRT3a5N396ko8F/UK8X4M1zLn48uCralLUjPQbZzvLBXkfUAPFQrDqzmD8bM6XIl
j6Pq3OA4cHHw1+zx/pS83YxB47augKB5ZUm14NnfeeNkhUkuCf+GrWWoZmNEdbLB5aYh7qb2tjEC
Npb+Q7XhUxyjEF20+D7rDtAdSBRALTJ9fcmXQpforx36q1dZnU4mnMOKNv2Xu/nOuGh2qFan88Lz
7+Ap61zx/SG2uMF9SV55CVe6Me/LQGnky9cbAey01qsIVc4IU3j5Tjlogx/kAmzsKRsZCsoB3RTE
KPl7eOCNIUMQBmFR+fqMSeimlcb2Ka1rHdRJGaXIAhU3J+hT+8PZl5MPlVHFSwb7dg45Eir9MruS
IHE1SdpqqiIgqrZd6LkClc3umYhfeHH7RT1TMUxvBi4WsQMJDPkvowxaqGPUv12cmQhXvOF5BEgt
fMNz4JJlyQKLiP9pH6jKdCUmtttCZeaPChEz0TG5HUzEgRYhkIsm24IF0O9pl0smwuXsB9o9Qp9f
vMBN9Y/2Is15G5F6QaqeCki7jyyx8iQ8OCFajFMaZKzlMb2q/q37yNHTNuRH9xaNaxNIKtew2vRD
qB1OcEXjcHGsmYifyizNN4SmZgyZxEevudcrXXOZjzYVbfwuGBEKJdziH8KPp+O5xNKbFaFCAQwf
ZXOD50Ezvw2vIeYPtRmqPut3sTt+gwdRWTJzO/3wC64IjXJm7JZ3gUUL90Z9bnQ/W3Mp77jwZhDO
+gXnkzM6Ih0zPjmCX1C8eWzlIfwL4K8FdQLc6N8BocTlJdkFuyrxBirHpAKkcKxn/QIc54A8mrA/
gB7YVPTiDNCb183exEaF4hmODQ/Sx+FTgS/z3l8Q9GyUr1X9vvMJnsIHC/YIzCa+K70MuBQElcYX
Lnr1h4XqgPkb+WBFwrxCuCKgHv/634pIhsWVVGRthpC2ko6A8dl9DQoBvr+/xqGOQTD8UNMQQEdR
rpVP9kbgCSwBDXLL3d0bAcPvn1WLt0j56YeqPVX5iZcfRVw/+u1RjKSkPPBMlNMlaokjmZ7ud+U6
bDou3VmJ8LoBamYfaendUextLbiUl/+wD/JBGp6bF6+wdZq5hvWgoCU4FfDKGwYFI+oCdaX5YoqN
4wsRDUc71B9V7BTeUoou2CGY+T2QVYEAYtgam1iEu4J6tDmXJPKfXWFVb2YhgUIjlACFUvRax9iU
w0kvQp7OX8IDBaQww7tC3wVq0NprARyAl22TSUPftGFTrNp6N/e480/NcSPCVFx/M8Qs4nKlIDZt
IDGMm/EkCxO65R2H9WfpbQkqRg2HyIzoXng87ONz9Q3ZLKYrhnqhCGSXUMrdBW/efUgFYm8i4pD/
vCHXEeVVws/7bN+FiPQsruvHym7iOdYTivBqPtl2x4eNO++TZQa45+rOFtnNRaCk8KzDDaeHybCO
m/wYK9L70OyuqzNhf3Okx878rUNzOFkXhj5ApqEYWbXujGAWdLZz+5FrntXTsfGCEwRMYP5tl8Et
Ywb30aVy20hpq90sZ6Spg5CFvT/Ctc+LwbW6XR4L+e/t6oZVHdr0vd6GUYBgexz5Tqs+6XUV2oDl
O7Ku9pTa8OD3wnlZe0iaiX/9Y03uvKoArBlRSAHR9epmNAePQZbOFjbrppY2zdqjNfPK6M5XoCQp
u8KiPqEmwxATBGdYBjFj5RWrxsHjB8iR5/BsKNYm0RmAGVGD39rKHslW3qZ7JJ9Ky1p2KYM0ZO7g
nrU8d/HGsev0aTooWNdJA2raCu5MlRXXyz+GyBmVdVDSM3IgmQ8CKv34VCKgNbPeOpbXMgUfvwG4
qOIgRorLXeHcIHmopt0FJQYH+Vr+XIAHxNnKoK6xqqv0aD7mcKb2AYe5XP0Qb8dQyMgEGIPKg4H0
VwU7Fqa3gk/UQsdzIX6+5hLtm7l9yVyFkBbTjtaeSJySxiYOP+K1XFRFrljppWEQtZHDqEdd+yCv
b1HbqwgsAili254fi4JlTl5fVZb1lRLK36SJVCL9UGFl/+6zLTSqmv7yYElJlKeZfzyRs1gdGb3A
o4jSZneZcU8Tw7KG9ZEAYmvXV8ZW9C6lSqN3evJXn02bZR6TvmwzCYKd8SdAAjwLN8PIJKBsdeDh
poFiXENDp0pEdDjOfqZBuPkJ2/ZuSs14MXRpyposPzBbSxkc/ikL2MqNem09OYXiHMG6E9/YDpPo
CkrLHLxLZ+c1BYZz+ut7Wb2MrIbumjRYr+CJQqSsdC6JfhAfvOv9yM/dQeq3CMxyx1G21ywVjcXu
AYqY084edxkMUCWeZEkzXlVeG1Tn/bmr+M/QueXcwecwHiIDB9/5yovZXmpnVGov23yPlYjukTHK
7gf+q+a9A1d20TBq/QTp3KRtF/sFMNwLblXlXu5pB+q7BuNz7xg0IV6uRwFe8i3RH1t0uyAhS54X
yszO0JSDgBofWWAOqF7rUUq0Xndi4yl7KVb7Rx86oZuqgbxhItxQ12FjVh5viEoZcSUKZgHe/eth
HTC0zPOt33ZekcsJMGlZC07jPdc6YRzhpuDIv7qJBTWnSJF21WSpVhHrrIGmkiiDnUPmV/Ge8sqZ
w6JEuY7iBsiNVJ+99CvHi7llMPmjZZ7iVRani0QG/ozmylHJ4EAW4hhY78R/XmMfwOX+9OlZfEy1
NnMkH0xSTaWzgYEXAeGmfNHTZx55zPeQPCBeGOMsgWocu+OZoikk7g7HX3ss45esPxqISKQy1opE
ofN9XFnN+/ZmOkkOG+xIBRk3q9LQ3s/X3VsMj7lHvjzsNm5qLrl68BJX3pWR6QuGsHm4k3ENDXNE
S0GsmxZY0tUavK1If3mLqllVTm7xsbVVZdhroxkp8aIv20lyu7YQFGH1/F1QjhDy9FCqHgN+I9EA
zIRCWXz66Kxz4anKSTeMzUX+ZcZQh01s7uqcBxAnLhhWHK2N+4EnoV609479MidFsqyV3LV/DhiW
VPktZY78QZjFKoGLjmHRc+RQUuNc1sAEgFbjCuEJmPEz8Ysc9q2BsGSMYakS8X4Qdp1uxamYeomW
fzB7sM9t3FbBgqptlzIEW+e9QL34M3W2S0a2ISUsDflvi5rLDfJEa4RtM+gsvbFBqWhA6OwQg7ND
t8p/ih9ETTJ/7F6H03lxh79gF6r6HNDDqHs/ZPpJyLYjJEhF6GIYPVt1LA4Xax3avCIUxBnCgo/2
tTOGJJ+N7+86o6iGVZFXokxWiTIbeENRqqLv3PF7ayAt44JF86NW+j6pl8IEWCm7KFvbkscQeH2G
TAhlJH8EFhh0ISOez0CSxYjx1XV4FAJHGSVE31pq1AXTnBpVZK8SCLALFnCd0fdD5EBaYVv63p2S
lP1ujC4mXjR8ql6Cfb0FxOFm4dR2YrfHfI6nebcTnuacmwrpPs+57f0dpiFNkZgV0gEPGqJ/qgum
f0i9eyAX/8R3JqdFiv6jDDIsXxwwuRxGxlkJx5mFAxBD4tkfpbHXw3HQUDxOqQsEaBgPmwCCjA/j
IYm02keinTaVXJ49V5ZEfuUoNDeKGg7s+ecidn6vqhfISDBEtVIBt1jDGqC2WRkWdFLFS/l3g5Zm
FbSjkuCaeZf7yeg1/blU4/vs4myPgRztL7TfQCwRyOvlnLKm2h/dz8ygOOw+/GN9Orl9RjRwxLji
fYmR1it+xmz+tZgT9S1nExHQMA50wZcJZoYZowu6Ve0JPzlC+nf9ePBICrffCxV01e9ixbZcg+Ex
1VaLMF7bl+laZNRPygXUflb5CSNBOCRa79yFwq1LfCzGK8qGH+s4yqqqzOJxexoeVAbMs92Gf8dn
LiaL08EF4GLSBXYEa0kyOpvtluGyzfCNzgliFkcSFBRUrKwrjmstk6iD3+/STYT+7q6WTsD7S7Lp
dO89NuoPgAKzvNoYb6m8Q+lwdx6hnHCjfl0FbkDb23A1CVxj4w2rm1Zl6iXuObTi1hqgWSVKxXFj
afz8Y75K9Qm5DhBCdQQqZdqIzCEvqwbpDsf016dQzgt7ka57+jYZFUCR1SSCjwxhEDv9yaOanQ2q
lWEXMyfLQDPGAOza8Gk7UOOttVJZlT3ki6pBbwjZ2RAfyjumIt1jkjqB2Bh/iNgqqm1iw3Ows2rN
72d2Dyy2OJ+bRPMmAbZTCzvGMfwNHv6scCQimhhGDkC3WJecFSIYvAohFJvR48n4vB3fHPZVfapm
rTVJGoEI/BatMPYVENPDJDZSPSDYEIz4sZVM66+cX5r4nWrGv1IXCWw5WXD4XME++d6PvfSsvNNc
LdEhEZ7LjsIeuYMl5Ud6NhTpl4nZwrxNxh2wAwh1qf0jNISuTeje9VabYxFXXuiaBKQO7/cJZU9c
oDpBl3BJwiULjnq0G2wz+88BMo0c1DcaHeGIZr8W+9b+Z4muorKXirT3L12fSTZwItbNH9MTFHvG
F18KLqbLe0zzIWd+udavTlkErFz2bnoEN6YXEw30yBGwHr8IavihDJbGnTK19qURberPjp943Mbm
BYCD4UGUfr91fIn2XqfvNRn+HMICbARETUkUaG2mgG4+adnBn3Xo0ZCLOARehQMp9k92hjPwJkQW
7FMp9cE8pFacSOO8fvIE+/5O2XiXghP91ugvsDFJMF234u250N74Y+Uh7Lq2hDlQoz3WmHV7tSxA
c+o8CV1AkbnQYOj0LNfq0lO0cQn2deiYZf5+HtfcIdf+ktM2/TvU9OTesUWi9dJkO9XHvZoQkKDJ
AdRKoAcmt98OUya872uycySu6JJxiO+IUyJhsJLr+xiHayVUzkq+iG+YwtkK9MLec5TGbqBmbuyC
0/CEPVU0XizohCVUxclN9zoUoY1f6b77tIHuYL+11QMWh9Lf1EaJbNrz9ATkZMNl/Yc6VqYC3o64
SKhpWer34O8jzBWRZwdUZ04xgT4kwQmAQr9gj2oZGNNQn2uidaE3n67bcTzYswJ4PATK/nFHaIEY
OiP+1dRTDXsu/llEI339b38+jAWQp4qcChVGqavBi9XlpN6oeJ7NJkrQENRGzBX31vl59TgF+WhK
TfBsU++3JT04uFhzpp+PaWt0gjV07K/c/wh66wStZyP0WExROYAvacRMHZvSc7JTVwyZKeqNXAwG
zJBUTdSdXqDiAQfCXPHNRfg0anAcxTcO0nivrVQPLHdh6+pOZQf+wXSJrptzaW2QEkdUhO9pvdW9
spPBf/SmYmrzOLDIz/VjQqmuaYdUUd0d7xXjgXQY6rv90UpawRVJPkrFn2koaa7oQK2RXoYh6HsV
xZ7bmPMHmau6YxfK5wQb1Gls4gmmoHrW895kiI5yzY4cd1y89cWNdrlwZ1+/nv0E9K3AbqYLrgzp
6erj3xo2LyupyzVcC1H2pk7Vsjb7j/rkSGfgJyh0j+NmuSGdRXQJBGtNq/uu6hYodK9yT8Fm1AVr
lHU5i20LaTqO+jFprqpputpxvpirD/sAzKDGdYypiSApiHU3AsLIUj0kYL1CbYSSZq53Fsk/9ui1
7dCUUB+P3YxeekrBcgDPJArnrUPP0F/Aw7Lmr1ws6P/TBR1nu+xUhfMhr8zimnEU18bLDPJ//owt
cx03FwFZ4rgXCLf01Fk6mnIgN8r/DHdiH4v9hH9vZ2ftJh6NHBt8HYSq0otrXbhrH6jth32AA45p
d4GXt7nQO2ZqbPhZtUUz47j/YIMoZjcjxz4N85E57SJ4ikd64zu98F91xSWRCqoWb05u3NZ6fsye
3PS4ZXAhccWd8OukRJwaRqt+G3TcDZHfB1aM6orhbnjgLr3rAVGe8Bpt/MkGw/AZ3oBgsl0+Ekkz
FaX6GL9LpGQjAqi+Gf3syLpT9LIsX4YT3NcUWNQiEud2uviMm7HjGox1DXhIdWc2xEZ0tmzxjJmR
KJAVvwM4s1D77Q0Zh5YkLYiP4mz4k9H9NgNDBQgu/gW87viN6FCIaVLA6TJcVatedvmSxJ9qzG+K
L1ejVZKqyaxDR6bV/a+Q/7hzTthNzs57DH04ngL2dZSJJHDGr7VGjG0AJ3VfcmqxrRO6ojWeceu2
YKx4Jx0trQFNoGQuZ5sOCkx5YDbjZ93Fa2W85c0fAhNSoDy1Hpp7x2X7E2sR2LAxfuk7wZJCWFB2
A/CWlzl9s+UttTK37oXlvPCoTK4PWydntbc52dwWGmaZ4EbvZLWaRmPK6+22lcbaM0SAusnpBgNA
5dR3PKbOr6rgrqj1fo04z2mdALUpnkio/xC08x5U7tSzvFku/vJNDfyM8hH3STT2U92+9z5gzQev
Xm8aDRIrsJ9NRT1ckJgE6juQalNq2Ci9M3RUtw8KR/Hui4KKR+VeMOpaj1rWuzygoseDPGX535yh
GCRY4qi+POrqC/suZWtdi+R1d7ySB4rmjVUXizkfMNGs2OtvtcOCBTeP/Ob+WR9qeVyhhc//Xihk
/QcyVxQyeOLZj5npDBex/oVi2Bzq6JTuGHSGHn9GEEpcmZiV5e9Zah0wHj3yv4JxEX/YISYmx7YG
xpGYoTYhOyf+pvMehQWzKd5u4NYvwpHJG64t48CteqJl8YfMBXgKvIa1QBaTU8OO1dhMgzjkVqeP
FIXp/eDNaizRhU5AORT+x44BX8cN+lsSiF1Qh0yc6+85q6C5Jch98gEQrXO9KlpQom1kWINN3hgF
Y1OqA1tMBjvKX61e/Os0grJV03oyDsCKtqgPVutEAYlfrqu8xTe0aS6b0iC9DzwaU8kDUclOJO0E
gFDyrh1Eyl2+DH4pF9L/qUxjVt+3iHdXEClaP8eM+D8hwdZpNXbS5ZNoVzw1H2YWnZHgLdBB2pnZ
4s0UVvxTs9SWoapSk2SZU55jPbVXMqRK0MB7/KfjRdiWzj4nvNoSvQHno7gy0iXol2MD0SNF+TNx
hoDWWPEwp+d5ODJKVnK74fSVvE6ciz1jvHyvT9fpdD8trVQS4Rdghld2TRSZNrCOIC19mVd/H1aa
ro+UMVh+UIpPc/qdqMOmr9+jKYrR1cXkkM+soWyXAaTkD2c0iZcg7n78CK5iMd4iGfifYdYW9oSz
BxkUIQeE8PfKsfThxwVMlP2cBcNNJ0z48r+Ih7fdr+DGNcCA4P6aIYNr4DItdppkxL3LQmb67ehZ
jWP3d6fWDPNR5RydrUIyL9jTKa58CU7otRs+Wm3QMjbkmEnd+nV9c/Q0Ks4Dfcyc67pO6NP1yLa4
b0mkRvDExjMksCfqhycxSIZU0ZeVYEvFxy7Flhj6KawAsZ9bknFYXrBDkyt0FKffsB34SIAlnIaY
PsvRrLwuldapZ967kKek4aeKJsW8OkyrTaka6jhIpquNZQpKWKX/f6UAL++1LGZ6F7e0f3TK2A9d
ybyCj+UsPk626FPw2cU05QQFkkS/3mbEm8OSWSURW/qbZxnP/fmczOMVtOBB7Obwur7rfmBYFz76
VwnZ2ItRQmqhskB7jZ1PPkfimCeOTmafXb3Unxu7pyiFtQ4cPZmtx5uaAyYuRHYcxO12EI8rYtrS
TZkuNyvP5pBqQfjjTof0bxFPv396IzX42cGXN+jWFXOCMhmvmBbYrFq5cq8AQS9RVC+TbHttAu1d
ES0TFW3sKFNUBn+CF25gcFoVBfxTMDDwCicuqjSFrUD7toaPIB+rXuj1lTS8TWVbopbFrlNp5qRc
JvLlh03wjLepgHtyrqEwa6+kfhBSkEm0gt3Z+zd/zNL9Jht0kTn1du8irGTqvOPsKYRBAs366Ldq
KB2isixTKIPjLR7PUBzyn5CxVy8tvHWTLMmK52kfGQVb0i+HevmZc9ByQ7cl7yrUwSrrA48N46Tj
rcQMsCHxb5iAOAyBYc8LGWVQEaqHsvFCmwAuaERjx0GGQGE1UWNvq6vd2JVVk9xfUoir8afkqM18
PFyXnuGqVMU3BqTR5tX+EL+MSGpW7KqffDENR31eN+D/oM0IDmgoa+RjBWQQJ09rEkvZwC6tULW/
f3IbTwfozQMfW5Q5OovcUZ67rnBarjuiqPoTLsPFAKcP5G3nyxIWZ/7SJRHf9cGCcZVEhGvenAnl
hDH9OWg1kM+4jQP7m9qs2qKKAgKNLaWEDHKJrtMy855xrfOXTBGbKOujEEkh3NiTrkJGoE7HVc2j
7EtB04ORDj4EsrUNhBRB5DF0p7GZXl+ACr/Smj3izhGB4huvrIetP6hptIFp7DSU6dbZZb+XIJov
uNcJnL9Y2ADACL6WAkPW+HE7XepC6uLFFDGC9/6cIUOkqKdcrVYLzYaVM7UcZAZk++YHBXbJmk2A
cM8CMz1eQTxYaOsIsQR49TBZxdw2ABtupfYGcmaVBkmiz7fY6zc8r++B2agIiBd2famEgamFM07D
5ug1HHXWvx8bfxMaB5EDL+yosASqmw5UzBZQeNxuCKCZxX5EGpSFtLpCQpsQhH20fNlkb4uh5acr
TbkAyOoXeeRHYwmACtxuqC0EJntkg0fbxipQ3ekzWmpGMt7H3hncNhEOLOudifoaA9PKwzp/Vgkp
xJrvrAXHuxUoz9QdcONOSZQ5Kb/wzopApD0CIN4NUhDheyi9uoM+Zt8PYqyOHleCsT+HTwxbci2B
Q5ddNxk36sbGCO6mS6GVEZEnvo5FnbeJBOGW8VUpeOFg0bIxHWmHTldBel9zEN5L/9iHva9k3DIa
wyrUtOv8OfPLEa8n+tM+kqew9h39cbBWf3XDbRnCtaOOMCpcuern40bBmMthi85j63BVpFZDTg3i
9tSfeQV7/clsVveYZrBfWGz4uYbqkCiu1dEDRJ9K9vNg3gi80kuCGOUKU2VrxBeSy+AKniX7a1/4
YXEtEzowab5GMY88r+c0lVHAQoslKlfnm1DbOH1iNwero6DZhPYBQ4NQcRZFF9kZbot8eevoBLsR
Yzp4jZjn9g9vWFGtD8z9VYBmDnOk/6sfP2fze5itwsqrkv0eDPqW+j8umxRySMH0Ie1aJ47cVtyW
H3dJRBhknm8Pf1tzYNkRDWzE+kjZWbhaGiTlv88vioI+25dIfA0lxUlgDDakrbBdelSlaFNp972/
p0UV3ylVCOEZiqwnPcTP/jSAUdpNfQfHRZxxgFegc+hd7xR63nVZRD9dFbkVUe5zffWTLUQOzVW6
u3ZSAEnVMt0/T03ezVQFmGySc5tjCQD/o6qyK0fXk6+hEfyOXyFbcnsSOM6yUD8r3ISTHHicXLsM
EX6RzqEOwgHA/B/10iDMIM8MLssZlExHZeXCqrVMDg5lvrMSBywkyQjIzpsAm55Fc0RbefnGifFT
U9CSmBPfF6ZU/Gn889WPoWnJVBfCLYB7JuKXEunOVYMVkVmu/mSKVDELcoKOVq7G0PWGeOatFj78
ANgPoWNuXGwK+ZHrLqYRgZnoqjkcrcXEYU2Qe+Nz7WpUo3vOLVALdU2zcOjq757pcdkJzIe+Jrdb
MgIGErinLz0+VQrr48zjQnjriw733rE5f3JJxfM/9L7ZV3URP2q7Ncwte/wvfAk3lE9V47f3MdV7
D3G/kEpIv9KOvgTD2VPFz0Ml87znt+wDhgZ4XWg3EgLiZfD+y1jNyPky67mIPg0ZDY6XobAyMg1t
r2iZxVAY0FOnyqYcsazuxCAB7SV3aJbDNlQds6Rstr5MzSXoQK9BbtE7khtDAGnDQilRTDPnRBHp
s2wNQiZZiCh+kb/Aat+cnsnpSW2MSa9w7zexCYgz8vz8gGKNGBBHjb8TIwv7Ia9F/6fcTfYRJgDE
h3dNn5yJwBpuR32FV5ZnoZpcFgjfVXYSxDwkA1LKKaOUfxkozVbc+uFU+ltW4P1ooHdVhD331W6g
gzDO92ji7fp4RwH3qDQN/6mFJu08SrlPz58hD4bkDm2U5c3kEFxEzlVDIR82UTZGL0mT3zbY/OZb
vmBTqsxMQaeos+YTkMdXLOKMnnlLlGP4Bm38h8CRBJt61RnRkMPqu6xdEIWQ0WMdGQws4iws+BJK
Q3NukuD3ubYteJkjt7zJd6QUB4G/pFfFTH9alBpvrbfbqvGqMw6Z1Zogs2GqFOi1GeWu/z6HHCSz
zWl6hXl6H3/Kl9xtRWR3MkFzKggGNVseSoWF34vAlu3TBTcrN0jgtmGA5ospt0log8KeqiYHld29
fIHxtCxu/lXeRhTjeBX0+Y7czCjRyKT2Ab94o0o7uwoWtJ71t+wQYQB65AzTlaRIKCrPN9XdiWYl
5kXVZCLnXnz9FMj6jklV8UfsmvVzWk+uufiS+g8+95UhX4O7Iv3V88QSLNE2CIhw+nuCGgx0dFue
KcjJlLF2InC+rabqc8Kt35rwVWBZElEJIGOofGlaAd0uPMk6Di+UTGG+KPNu7xVnIBKMjGEf+R/8
9a36+yxrjL4KKmZRP/fVbmLy3vwntBSkl+/dKsau+PsntU2qc+Rdaz7v3cv8DTl4ixJA3d3n8DHr
uK/Qk/a1UW+RmhH2LqJhlwe3Lq/0SwTQN0GqKd0jH1B3Ad/vpEyg+1Bm91pmSSlrhreLyEs4kkx1
g7NfiuG+YQqs5e4szIT145VRak1O6DvUtj6VY3LlUCeJPsvOm520VPaY6AhwxS2k7cdXu39EqwEA
rIqJJZpDyRytsXxwcrKprt6+McVtfhv1eZopvgtYTeMYt1h6KjpddncuIEQuJhQxDspCheu9Rpzt
aGM+Cqazq5K+GBeoSmCWNhJs+kqBLfAM1yWsKytL1oDoT/PfghU21+v2STOMUIPRq1CnSCdQ0jTr
EozZh0oiako8TsiSjwDXaACX7gYjrg1nKz1F+jT7mzCPlnkXgXBMUEJS1gK9+Eb0G7Xl+0mRPiwW
mt22OtRUBVIOQLTW+ZMwYwKgxQIpwBwD4tLCM03eWCpSllQkzRNmkyVktr1SLZWkmj4sX2HaZkK4
T/q5eXPfkC/WLqfiHA8ivaYswoMi4s4IRhks0ydR0UJrX8A0ia6PaBmdOoO1bFNCf9z4oE0wVCpA
fOc5ccdT4LSoJnzbOoe52q8jldFZ8nbZXFLFWczG2XIxUtlE+vm3myIqZVuXa0Sd1cqzIfr43wIV
Xx9gArLjprMi2qBvr0z5hlAKouNISsb2p1MpdHfbVHkICa/iOmB/oRh/fy4wVBskiRzduFSblpwd
fk5TOTe5ja0sJ8ycacfwcZPHnJ55p/SHC8oqHrlKwlsljEjUSM2zIiQQBeldy3+kMGygQdbiuog0
vl7vVMM7ZnS/2GBJnc65NvLetPCSQ94vjXbwfgbwvNzh45GVvHSipAQHLMGjltooUMjgwKQOZTTn
hnp/qDVpcNr1CamdHwt4thjljta7wsmOvU4mQEs5HEIWCvi5wsFK4N2SPJkg2Rx93486CPjh1xGp
amm36uSP/+cOUYDbuahWdDtSpmAvY3Z1jxnscBLztgmc7vefv82s8mQ7c9qvDvglicmMtxfRI5le
YoS2RPclBC8DvCwF/bQkytt9sxH7D0dWQJrD5hwyniR08akqbduAGmZVzTZcskHtFph8fV6Rq1Oc
L0AU4qJnt6mraZyIGuPknGSzBIcqUNIc5CMHnpMcsygTw1Y1vSeSr53zrOKhOj8tJQSEkYibt4yA
b5L7HSUOwiLVVW58ad7x3Jm1RM2n704cPXmTy08qhHaAhinFWI9CowIy8nPGdTE3pGZch60cd2r6
57qK9eLE0mqxCOtQL8pwLSQ2wuGHdEQeFzds56enw9ZuEDmniWk1lS7x4ar856ehuXW1661nOOLX
UMi4CH1otoMUBfPW1WMRXMJHVZt2flMf4xSMfAxFEANo0M/r++9s45oJs3+aRrawNtVxFIke6AtZ
6Ey4tQD7VKHPMCJ/vOgcmRHDNGmirm5fMEhi0w+pxw2vZL3lR/9qZnNpe8+MGuVRGF729XYUEQ2j
iTiagSt7+gu7GYcWS/QmVU05KpavIjGLy/+w9C+1f8Nys2B524hfuUsipRTF023uGk0KjeXgNzGw
296UWGSzdQDbGoAdQZE7ilvNffY5xZFLfnzYlwQZKN941pnF6RG5mBlYEbJSFKiIO9cf4inHM4Bz
mOgVtTICyRIj5ydfajUiDfBgjX6Wfqmdsa8ekfzwpqygsqRMMNh/OGE7R1q3E6emljFhwvftLeQh
BBz37lXuzz4iVjGKXGdY5fTIgRdIutzwEdIwXpOmdvt0phXLKBYWGiUJPvohzVVy4d9U+DT70Iok
oNrGaQZhC/u7z1G3o3Kmyat6sAi92yyVVXncGXA9Rf7DKgEEdqKCMv9Ej+ERPAbx7ffkKdSCoCyK
4M11d1JBWJphSVvLEsCDrd9SSJt9+YGZbRJDLHdFdFqWq3EPLyzp9bg0bz0h6nFkYsRxaLyKr4lx
Dwno/nyRqPEgTdqPnmpdnPNoyL2IbD/TymAY5I6Ka6GkWxMxppQHfODgp4OIsJeE8W8SWzucifGK
cP+Mfo8zoH3sHAY6mGNfu19fR+AXK++VtJMZi6T2Pt3Qobw+NvElzzk44oZ59KVZNM31TL16Hmhf
+neQflgguXLl7smc9OXeer7aKn2w+uJfmifC1K08gdyvwuUPMBVGL6Y78wY6VAb61Skcj24D6vWK
BbJvBEbhNcYwIekRT2w3Hieyy8eYlGUclgYSM+L8lvqz98MKLRhfAnsF4Pw2sLnCbrLl8oGqzds/
WrTxlexdglzFOgy8l3VdSEmWo74s+RsxV68RgQtdwWnuGMT5E8uzUYOQkipYO1Yq5wKpOL7prLn3
PIv1/VJzmQXhSKfhO+ziJt5zkGR13o8t26TOXwCsQrA0Rz9oZKjCaYwQibbWMNo4bLXJxIIbWZrV
1jvL3ctuZWcPnOPrryxuVxHSiD5FDDw0UVmrDkUR9x75z4GID41NjFnHXpYGPaGzPxaKHw+4OzKz
6AP+TDG2N0x01ARJGXfyAW3wdWI6Td9EdR/sI9le1a5MyL2I4QzBuX40QtLJ9rJH9q9fQ0bGogfI
fZ6vztLfFQHoy71iTM+iiW1+8ZO3d/Zmej/Jgkwn89Myp9ypB46NoZsahNdrXUuoMafpyNcnQm/0
twJTr9xoDiZnWv1i4gU++cRZB3eHvgTJWkFHYAlgwQXj3Q+KK5P6DLg2HevItSgNMO6kT+yRVqoY
RUoHtVvUlr8I8EtVHXunz3aCWYK1Vqb+NQ7tBEa+7+X1faCLNbpDsQDaCeaUHlnRbbbz8X9Fga5P
t3GqqXybmTmORHUjVQw/mtyapScSIUTpmSF15n8eHm76WvKJyVXhnQLVaFAeuuUwa0yx4I689ir9
r/HTdMqem/ZjtkfA9HbbB/BNYGQrKSAwcZ/EHDFVY75zFljZliVTisLlLy3OmH3ogT0LbQW2l3rz
q23JIxXj4uQzOVXnwJI1he7vHd/YczrSNNPcigSheu+56j8BpnQSigEIRefdbwrsgvA3XFuWlmVM
SvAT75BnPqqKsJcC4zz+GaU2GjmKEYGe5PDingXyWm8vIARRYHpJmlWiX+owjBilijRRhQt6rw8P
dooJI2mUCtyG7pjPIjtJq0F2zgAuKCkhz4S9NbdUl8Y0XpWMduFzUcqqs+RHQmxsbLAw5hTTVpmR
4VTH3JmSNAwDo92GXfn+VDfAAd2JMXGZB4aoiZim/MqMh8FuBdSmRLXxS7NM4kQvrfRciwpTLMMr
5qpH5PPlgaC9zwNa1cwB2VTXZ/BbUK6IrZkFejfZdDf3KgDgZZJN/pdL5EqWXS2HK+/xBWEpYo74
pjCsIPVuV1EtMy5zV6Kuc6Z1mQc2p5GrtyBtoMQ4UlJ/wUUof6TvTCUC2Ka16jsThAVbJI37gOfP
xNjYgqZOuLbQ22yX9DOdfQu2DKbdwhLX6w/L3qdsQryDB0qQA2+H8MS1AZdb+KP3xfAPH/XARAdO
ln2OtBfEzw3dGQdplp+gssMVbjFOkEAQZ8ugU1w3SlaMNlpXv4JKLI0nWGODPHBZ6G87mz6V43kM
TS9azc0Q9Bjf8MxSqfcTygJLRPM2wxGbwGoaDqZc46RI/w/YquMfOQnw2p2cYLxe2neeoafCFa4z
iN5fVbit9S+tSw2ldq4B14dgmCniqSTRitMG2HnK6mcgNyKXh3YXCL6nZErOBZAvSo9e3WdGuT8H
Xn+I5NHk2+OPM4XEP8T/2VZFBPqGzQBTuyBpr0ZS01Oy1Ox1TKDbeAjeVl68UOzPWEWBpW6WPnfb
wkrQ7B0A5uKnuT25ghSDiYertvJ6CwbgRw+Xn7xRKYjy8z0WA2ZmFmUiLIaiQdnYNYKmsInqGs5A
SaGQw17fz921S8LSZs6ynTqEmhZKOv30p+oSSWqB0mWK/tDjvUIJ4N8BIbX+C+hyoPdiHrp3GY10
x9lJm7Etbhc9MnhV3dP2EDWRQ70xH54oA3y5Mu2s964y7xnMrr+NBSHhryfWqLTfCHazsfIKD4DH
wmKRl9nvdHGl+zTQQ4gmuJPauanEHH7XJxq4aeTiFqqW0pT6vb3iN7FsJVmyU+xtlCIBsF9UJOtw
2ytm0DQ9PyixbtQgP68b5uRvxU+9nby+zaAv6B/UdQSShIBeAekAe2Mf+Ae7lsJn+Tuh3NKEwnGH
wTRvQ4CjwcgyzsQwRe/C81pkPZYotbwuWAZc6IVCnTNhNqjLLMQOKHqg06qlmPsIEVMvLGzp+IEy
IHv0YS/LISYVgIUmqTn6+QmsiwhFfAJ6V724rQzsVHhKa4E9AYFuRjn8D5mDvWr/h59FyjqsET6j
Jo6DpqUtgRElRu68NU6kEAM+AjpbFEEi3vIQNPCFdzQ94Xp4CzM/RR1gEgw/xAoyW0GlGSmz08P/
HAcqa/V9erz+Ic1EZfJtx4IbJE0YKTyRRai1/BqC8oeJhcaEDV2byhiWNJ03TJ0q0fqSxWyNNxlO
5SiW0nY6AaVdTfW/M1/uDiHv0/sjkSAEl6kwFGPmJe7SuiTVafAQ97VSYfrnTs86XEBlPPf/ddYS
3phcZL0iFBMLVEMOH2bYJwoFYM6P7DFjezMuc68NrUsnel+LMluEWiWA+xBr8EJ8fq7W7WFW+xpo
DC3aZSnDyW710+06NwoVPLPdygwnJ1LefwQBKGqXN3L+YSMdHCgfD2Z4it6gzSOapuaoiudgFqXX
gIA09R4y2dhIYwZWjXOY8sj0/Qim+c2Dv0FkNl8xd3dd9+FN2Qf+k3kO9WeXhEfxr/puIqo2MhoQ
UB5mUUrNJiHr+zRvrEvfNQyBPSGdRDdYa8MUyg1lhUFk6wwF5q5LbRfoybqg7tp2sa37cW4T8C1w
p9MQBMR9CbDIgbEkAfv4tAYTg7cnhewa05JhodgeFjJwv+SJ6cXfycNrzVHGk/43j0EbahIrscat
wkz//fnyTEtTNgPT/5GNVCpZ55CajaNXydw5qb4UYCPE5bAkKWdND/ECEIZMjQ73g8FSsCyMGol9
zhiqmM9d/FxWteXQrw0jTpdVsR5k9ffmpguCK48wgrw9khbp4VXWhsFQDesoOJbBR3lmV1fx79Wv
15b+A0UY1YYPRxbD0nSaNO5gjbKdaLvaWG/bXwrzWp66rTlv7MCYgCNxIoo9EjdfrgX/I/Ui8hb7
W5YYS7Q9G3twEgWo4Vzg7oWtJPaPq9VqKLbT5TMf8rlt/c+WVi5RtGk30MVdUC3N/tavtYFW8ygS
vZg8cNsQDSYPHQo/w8reUjQLFQnyGWVgNVvW7iehrRAWTN68OLP9Y7WBopioBwy2AP/HTa0Zz3+x
FVQeL4jX5OlbmQErvfEx5Q2MnlKX+VWlNESrB+av9l+Vv7I8CbrEZln+qHqlE+ETnd/IlMh4xcVl
4THmCTLx3CqXzo0EzcDv50VWjCvLdoIsuwoT1eK1KkCsKGox2TdmVB1+04mDOAVS1X6XH5Dp3SX3
ASiLRMKotj1nvKjywxSjej7foSl9/p3YZO2v469FHZeuxTSKEjvLKJhkK9gA5ccMc6yPL415tm5M
cAxpwE+2y9KVWGzwHvr7ErfgZYc6Mx/9h1aU4dOuo5NW5VgpMeC0NBai5EgqBw7y65RP3NyAz7jo
fwYiW7XH6upFR0VPj0bvidCxNlHquSYtBqZ0oG/Y6NSNDwRitjvqt8Z+xWKU4kzX56VDHiY8PmIB
2GTZwt2VBh9tEZqOhQJTpGNNcdLMUZpGEDTjlJNfY1ZBxA2a0iX4krjz2Baeb8ZnN5VqBsSnrMK9
ioZA3P8egQX3yDtG1AIFyrj60aljhvZNmSiwk2ymxiYlDoq1tnhkSepb4nykRWGywU2JZerQW6Fd
uv5rRYYdnoS5V57URrchM4ZE2NdW95qv+2okazByQCsqh+1ufB0tHqvC4iqEnHaiTAQ+rxRwm8wF
sZfrTGwQ4H5b3iaRIb2/QuS50Pk57G0P4lk6BTJ8OcYVCpK49EFWyjg+rGXEhZLqa9edd9csQtHu
MSbYVDvV2NN/11CaQHDAkIz1LVQmqL3yZO5vJ+Q52FRuQNzlTx41LJ81t5uwPKFLlXf5G3lubicg
dQjln5GDW4gnF5hnTZqoXUTYrZn6oJ2eNBCTeOtbNJ84RwnPbxs29ozTd0hPQOQvrCDubGAWN+yF
8169a4w6jIFl6TOwAByV8uLkIkqrlgk+EirCbJYH0rkgaF20t1hc8UTAU+FSCsKif4ff6qv2a0gI
5LVLJ6iAyPdlW1+YgzDSduR0JVq2lh44peAoxAbKzjLlEFwNfovStUCKHLgN2cTA78X4zRMezTCL
9yV38iI5EpQ6CLT/dQB7D+qwLuozqIn975lmpJKKC3Kpwo8YOI7ESnWUtM8jZgvo9jOKDYVXlsTy
Hl8/KfTT454JizvG/DBgxRpCdQe6vl0ezvvtErXZ9iuaEWEZKEiJVPSXBrDkUcVkEkTI+FDAwlCq
zfKmRPlCF8C4ew5MkxNo1+1qm+tnNtl1o4ifcfg4GGl2HN5DxJ/FHlsmr1wAu1ypv5aIfrQOUa38
+cmkXujPzgoozmJkL8lvLNWVOQ+L/BpttN5dEu0MNWa833j1B/+Mp8iFtD046PUMQkohjFUKVTpz
bihbWHyirlHFLn15U4uTGxCTlD3TvhEyWYi1HvRa9TqUt47fwotGJigrncWz+BIR3bHkgmS2h+ZU
BWgoHFmwWkbiNxpa4jWANDl7dspbHZ6jeh6G883v7Zat15RaxfD0zLLaqSWMEdiu/iWhR2ajVRQO
Ywh6x43oiehQL5l8gUbOkGnwgTZ+0SWmlARggkVy093+5ZnV+PjsSw4RYeb6+nxifOBVnNiecwXo
2R7Ki8/Ad16vdqJJZPYr29Je9TSNX/OZeB945zQ+uXi3WuthwPlx9aoiJCzuPjcbR6RznTFWO+rl
wPnRkiiEhJMdP72FDzfA67vcmGcEf22mqXREQIgbKwuIH98dPOEllflUZuZ7WKeJDTnKSThsrTR9
nE8ESfOmHmWZcywHfug/WsBWD5v8phKpwGeBHW9YoA3IXfLLZv2f+gamFsefNBspHXtM2jEPJ25S
oPmTK5sve+UdOuhAOTHT5V3Vf8HebAmdzDnCrxvrlYyPVDeKe4y7SzUZmOO1e4nNNGsXooBRn+qB
EzRQ3BKTPJcjm/g9KVVrv4V2mnghexUcFkcbnBAVZfnvCYL2xHdQXj8McsAojX3+VxsVebPDRwU7
gnkQCPZuJN2HTG39FU2qX8zdacifxl9EJpPLIGp3uOGyyPKNyFRmsn08TKf/DXF9KCy0ddMUjw3z
xiEA3zAz3afaxpIzc4KnU8BzlPQe4P2fMpMqpshAvt+IPySSkDPJnfzHL+3kKeThDcC8n7MPxqaK
JHee5MqmBBxMAyTevGNCa5x1BfhvG6a8ICfmgE4MYa85VHzoLKwGzncJTJMWd2UCbb3Ege2bnpxs
aKfSFeyWqkK9rmfX31Tqx7fvPrMm+kIU7f5MEsmWXvQ4mm6391Eac0RqfPwO5znetLWesp2bQTH5
TRQAaZfmqXdYjvcD/rIYXB4LS7cYh43cJikg8dX1ey8vhFgH5DuUx847nbfUNjIx4edmBIn2AcGN
wcsxNAefES+Tob6/IAytzzKaKdUMuPSRmygBjl0NHU93Rx54uAJtnANynNiXf62Lfj0CKNxEPVas
/ae14Gaiqb4Tdsh+JpRT+iT00/o1p5ynFLaW2KOC+O7+DuJT8GTjjws0Po50IbxuGCafFa+LN9Dw
n1/xV/IaLaSAdFC7DTtLRzKz+AarRSbviUDUdT9waUxn0f6clQoR6mFjyMCxU2bR713lcyyc8XW7
nmUHaYuKyEVLmRLyS3aecLqk34vuWNoxRMcdUWSe4mqkeof7zx+FPui150YrQMOImnGEdFAKmHOF
G/5xn8COAqLpl1UgeMRgCA5+G0xsmL7v4BuHJIDuSJnkPxzZbqm8hCJXcQLhpqwsBHWBkC9XF2Dq
2kalwfmTbmDZhlKlm//2x6AlcoBBw5JdzXkzTZZVXGVW+QjZxWlYpEBfkdJrkX0dqotzOEkKJX5J
mQ+JSHf5uxSP45uahGHUKHmkeLrMjaFnkPQ3BWoPOxJKCCz5awZAEOox0YGGceLmzHIpZwlaNS3j
tu6Ue68xDTh+Gj+Xc9siWNFtVO1nscUegf2ZCSUt5GwM6NDOUevdPVpmVTB4zyGXxh/xIPoQ7OGl
ceylRjONmZPrDJWGk6YbD0dmxirzb7x9xX7sYr3HM91fBpAV7m0TuwwEbVUabWm4XAHdAuyuAASn
BNtPPL6ZPAJ5E6yPmC0s8rMbPMU287FPTc7WEn6zkcVA6rn1M1FcERm1iCEfEkkB5u2T2jv+vK7n
kQ4m2FmmC63SxcCMXMRsqpY/+hSO8gW7qIW/PpP+eCcGep9GOb2dnMPp4QpyOuKG5nvdacYG8aKt
plLthV+87miqqGlgZMluJCT1psOXGsLBUXfW12gChk+5GW4ubHUB16W+Jn/s8r2jlGfxXwy16IK+
JfxYs3s5Ct6R13MWlv903GDlj1xwKkdjWkuTpvV1zpzcNUBtK8L0O6qQWHKeffaoMRZ9EOuqcAAd
C7yVF6Q3byyESmFjKpY0Ibo3Mew2D+JVMPPExmNFxqAMpJ5VUgyAyC2HAlfL8y12o9TqYoQc1+jd
jukVHM7p4QMBWg11JqOXFoWImqBHeRKr1mYQEc+7MwuXh5gSV0jlJmCLK1sjoNUTU/aSCkhfvAHg
iOCGiB6JKJezyb7DR1B6Np4ZgQItVxzRyT6HciqynFKvmtd7LxtZDT5np2sXzSPmHDobgjrkK92j
+2UZnFtaSoELt+GDppsuzORNPabEz4Mc9OUFdwuffdxsLSIBeTpLAJPNBS58YgsyvWSikyq6NaBL
YYfqws8vGP/prOKjljU9wemXszT6rel2oKlM7nSHC1hV6Lql7Dyqfbt4XvUCa0itMhrevJ7KFk4s
mCi6Houh4LiPVUsBOyKwoA+bdU9PCoMLoMadM9bsweDvShwxAE3fz2t4iNlIfiD2/k+TdcF7PU8t
G0dPMLk41bf/myANwua4ilpicdKaSJadeSMsswShHGYruaVr8SqiOBQJOwVmKFvq3I8WF4O09S4F
jrgT+mEjOnnmeLHZhmiXwQ4nmZOCSxTELY8IqBYUWGSJ7efbDrmJFO7w/4tlp0EWRZN16mtzjrqo
5d2P3I2wxceYsURZhua5eBbxH/V1WLld2VVUEUbI7vJua18wtLrflahX0+xi9Bcbo5rwb3S5WXnH
/3NGBb+FtXioMr7EM4LH86JFhxe97PEXHw59T3Ra6DUMpjfmqCbYuKlRN250kEL7Y25/M6yTn12X
igPw72Uj5DhuTtMgbmkqRHG3zNO9w+jQmh3tsOc6qytW0zFGD/cHUTCCxcZghe65KPTkqSHkkkWM
HE7BGjggTWa3D3H7RZgu5tozHG98+cWPXsPA3nUsGKv5V+Jv4j3JmPWB+Uk1Xlfn7PjEWKGtIeW9
ief7iuZiNvnP1YU5jKB/IpgVOhskn+kJNjAKJuIwVdwW21chgr/GvWeWsL+8grPg1EncvW1nDxW/
NgpJR8dj/poVdnyko0rhPVqeYn7Ov1Ipzlqhlhc4Ax+tX/a5AOnfd5TVekBP6VhxOCxdotXrftTb
H1OJqDAl9b9cOaaSxH0OvvpImBAQAZhaKgTAdTbDsRuDx9kmx2KbunHEMu8dZs0iycqCl4fo30M/
FqvNf7/Nz8KXeBmqZmud6pw7Wix/rMCIMWicNA3Qbij4GFCgIENQdPJ5L95VAEW/MWOxsY/txV2+
dxIkpWYvfeG/6BLSr6AVXO17bsqOehBuVVxTK3lWhAarznqyYtp08YHwWqXJ781GWDG3OT9PqGpf
KnpgpRQccYg52nyZum7oP2M13NMGl4Jrkuwm01cShNXk8sLGyBBt3FrImSuZH5Au0EaCWU/rkn9c
lieRGbudGFjszEPa2sXnIk0lNWrluRGVC/e4309O/qGxgCLV6ldBLBz26CRixIGJ7QmKYUa7nxoH
twg97pmudWNMDp+3oTA0cP70Ejj49a1p7K6mod5qjBXTgFiXqsnjNDnkKLDsa3CLPZQTegcizj0V
UGYp7FNyIn5FHt5abzG8sQ23OW6GarRQgR1XqtgkcW2g/DmDav7D8ESPPDEiL+cLadIXRic2fIQe
ZVGOKe++3YmyPv/GdCiT779sg+6X2+nU/FkmEz4ww+hBmnKMZ9dfk1TBFHzCpPfbzNTCy+1If0fT
oHWIR5tcFLfjDlPkv0+utFgCnXX8PRMbfwcv4M17ssRDNGb1g0X3e2uzL949OWcQT0dVNShW0QCP
hRYv/JkZwTifqXzb3LcZxtRQ3G2xaBtewl/b1zTp9hyjGPwUDLNS0o+93lwXqY3GK3PCAhI1CHW7
/snlGEO2TJ5nqHWQ8Suv4g3RpJW5YHNmNqUxSvcd/2W4kvE0/QFMrRzOrDKTM6eRTRi/WucH9TPw
wtP1zq6mUMu8S8z9PYLYDAgilVB5LWl5/4DPaKH2CtcZ18OZs1oaBJ69uDiMRIajQyH4JHzyYRBZ
8QuBkNKmolm3RydpMQnhzEtmVty5abimI7Z/UnbjAZFO8m5KYIxTDhkTDbf2WsxbGIqRKpQ8SALj
O/BbBBo1vHnWWxCuVWF7eUd4TXt4rlimChVBSHpfw9RSiytGibp7wAzcn/Kbof93w7fRkF8Ad/wZ
rRxnETIlgoRqjGsALPRB78eUYT0fLLUFvsmxjrQulnJzGaQM+cpg9/kyIdHYp6gA0Z7Q4HZVD5Gl
Z+VnYGFgxKx3OLyLqvEt/tvKfpmiwgs/sXHxiiyuQC80SEFoPytwpIj0uSG6XT7l7GkgQrmJAkl3
6nMKAuxpozB3Xk1du16/1Q1BMy+2+NSdHYntOHUHmBzZFAk5yp4Tg2B0sz1ZULh3ICs+l7KJQ8nO
yItXdDinhfJXVla9iWvy+Qsi8B6TkJ/W1smNOfG8TkUg1QtcPPVWMPMUGgBzIVkIxHE5qtcz3XeH
6WJ0kHLBpFY0Tz4ima5tqxgHQtJa6gWEFCIe/ccmREeyYWeZDyrt1qr1Ti6b3ovLkkSP8d6OJIms
RpQJrwVVFSWxtyaDtZYIYFAfgtgDt+2Efm0eQav0t0WEXuq3+SCGhz5ku28bjY/+1zAHF1lkq9m2
h8bZOgbI1VAZEpJCMdjp9wz7navzDloXe9YjMBirLi+iEQAwxNOkIbyvFa62NPbdurSv0Rexx3Nb
vYU6M21as1wfEmrxKn/pXWxO425yISy5+xevr7fyVH12XOkqNeNaZ42KgSVGvEdF4kwGDKhLSf3C
SkKAXCwufCdM/TFpunR4316BFH1+6D7rQjX+BuRmVcfK+6PqNAr9PH9lco9Iyt5Z3m8eUSievYr9
MGc3/K38EcYctKRvA7ooi9hFAcfsbNm1sk3kGc1bZXRoVi1LeNUF8XceFFQoqXNKu7rwLWGwmGCh
Pu+nMlUCJD0bxwTtrQTS5KkZpUnWbbGaYglotyCE+Wy53Lg91NTeIiwWtzERzr1NqJsb7f/0SXJ3
shoN0/E8PdpywGgFJGWmfVF9zQRye/p68Dlk0G+6+91lrnXhRIp+xcT8tWyb2uBQG3aNBY9TQBZa
2RK00eFdn9fs7opNDVQN+AAT4IM+23XE+WF6HAVeYPbhAJvE0jUOj1bvQjuMQpZ1z/JovV66Lqe4
JVAxioFVXXYyutu+ZcFJddb+A3j64+cdVVF5WO/AzwlRK7v/dnt799BwvuPVP8XzKlHIZ5ZfKwgR
30h4FkR4meqLp9aYldJw3QpBFo4BpfAu/iXeJ5BLncLxQJSz9QTRoB2/1p+lKHuOvOBGV+GAMAD0
nFeZasMnqVqH/izG2b4EYzv1VLW6du/WctUPZ08sbGguUrF0lbrH6E+zkALiH0wFURS0HQdynKxJ
V7kQrYSISd/u9LzyrR6zWbHYrbsVrSbRvaizwpGkvAsD/RoHpOBvqnZf1mAapHIWYE3r3wMEluxU
bkI2zuVdkwm7opV/TVDxlOcJB18VFazFo2Tyfpb8xOvLbyk7ZZIC7VlzszgwF+kb/+B2wkb0MdyY
ioR7KdpXKdlbFXLodLyRUtJjthaGMGWJ7HagE2uaJ61Yem2PRwoB6wmfPRmGyhpWVQ9H37+JsO4r
kBw4TPAZH61mJip/DoynEi0oh2qvBDUvZAVSxbLv9qdIYXiOWxs1MSgAMLxOfIoK9M2qikEqL+sJ
hAh/JxN6VnT0jdiibnm8gtLvKbYcIjHBK9NWF9huigEAVsXgV031tyx0BjWnhDhPQgPM1V5Gl2YV
XLrYllQ8w1ANwS7J5jNPRDMxJw+VdZ7v/dQPzmrgLCqEiL9geIebE3c0NuKiDGYQ6bgL3vhw3PJl
LuYQvBgg/uTZPFkfhFXvKIGeLMcHsxxRcwPviGkbvEvr1km3kYJ7kTlEDYFfSjv08doH6DjIdzND
cfbPvdpwPIzPVpTwbjh9L1osz9CmoeRkPTfVaGstSZKS3a47rX9NpMxpTQS0SPwW1Ivr2swjDW7R
ZwpC593I3ur/49R0606JsnhLQb3LNkDmBuu9rqlqQ0NYvC9lE5PAlA48VeV5gDmZ8wBwfnjmQgcO
HbgSdlHBWbgxY8sNQVGg3rycpE+FVLNGhgVLezIR4si0+aGNcJi7wEyXJ3f3eSSs1O0PUdkx1tfW
6gNkMbvLUdBAdk2Qhb+GAbbDUDZG6MLwnO824WV9FfUT1Hm3auttQw8fQ5YfSx7zdBDCbWJNs0Z+
aphI0usUrSMeJA2z9PXVOhJjWFYzQ8TOHIISTkFwzeRfHbF9D//yNjNjT43QcX1DP2jLfJHO7klV
HiKwKMX/adX8ciIGIvCH+pG33w2YMU2ohPyQZvdRVz7jncUi1pKDb+nnkr+fL2BEaFyuktJcfEfU
98u9nuOgC9CG0WP0pf9sEhU5HMoY3N9Zg9wLtxGRi106bMA8CzQlLCN7xoGUp2sQwwtrMuCBTpQt
/CHZwi+h0X8W4AO/r5vYv80JwT5U7Qsn3aYOHT/3RjkIuJAqqbW/9uEsiYCAPSb1HGM7vDfvJZy3
dNM9ZnY+MceJVwmixoNNtG6OIv+D0SkNgAeYem9N5/8UNvNauyuNCQzQhriTN31G2nlZqsoFrWSK
74bID+lRcBgtdDAaZHrpDreoUL5HRge4lgaJbhw0qS7b0oCrjX1JZTFNQ5DC6c/DQH051oJzkFhE
yd5Q96zDZjhmszIZYPUeoHCoiIv9VuACQg3n8s+I0yp3Lib8qqf9vzYudJToyLyyIVBZOXtTyXcL
sy5jnECkXYUlWWeotdNdYlafoghF1dPayxYszuUBXy+V82ECQWgvSJYVWT5hVI2OhLBUFMGBoC3C
o8D0bfGeQVVOk0qVEH3E1Q7TldYMQbJ8rPhL3fQiunD973G9Q4zE6JAYgkKIUT19j/JUI6FA4ac1
mcYyfUuDv15IcT7V8cddcFvlmI4wpnKEpcfEw5gX6gyvbo3f2GmbcmRy4sLqhriJX+rtw3kn1U55
NPf+NrJi7sdRapR+aSgYFweExRErsrBsEEdWLsNJxBDdGW9LgEwsfovUm9rAe3npjd1c2DfTYOn4
SA8xSo3HXFOWxLzigc+ko5hFTrmxTpFPT5R02IdHHV0e7ifkZZhWODX4yfT+HNXB30n/rlwJqpKC
g/KTDLlKDEQJZ61aRv2rEL2VypUZDZoLdMagSmozlJgeT6c8+gU+L6Pcj3ZblJuMl3kCbrPAdmJm
OGEZ9bZAjaxLNPQOkRHHp4UNSR58422uIIZeW9dRYNQkXVAbR28IgsSZc8krdxt5BZwZsHhsC4Xy
1+JQxAkGJVf5KE4rEwppNcZf0QUYeojbue9EIISIMvsGy9Cc8g0e1DITALi/8KKCs+GakPOJzBW4
s+ZufeXaEBHXF79KhHNvRH9W0MRs8bHUrWNSUUu2DV2It/LiqXk31in3iyzQ3YeX03JpStlivP2C
pZk2HwWbHpqcjFuRnzbcsDeMIX5h3ee6xOHDr41DsP/E/DWQrhWjySTbLBcGOGnZ/9eTYGV74+Zr
N0YF0ANnf2Ju1R8cAYifVNKoHC8Ll/0e5jZYbMskdxq+qvCgdb2yiAEAyOHKKlMg2wBQLdoaKUej
Z6wgwp2ktA1oCIQZfGJZKwO+uoC2+cidPXxVXVir+o7gsxnlyCISeB9/YhAIiIqE1xB772OhQOVR
3SERRCMVhzlOso8YMCmN6enO9sQ7SVbPA9nQsP/XInJ48p3DJxQOTY1A7HCBqcMssuXwp7cywDxL
TZCaB5PZOInBVgD0DmvDnCK5c/tcPcQ97LSs/Z300nkXUPAj5Gn4xmF2nJGzTq6BcpuhNoLN4TuS
XM9MUHbTnE/6gDz6k7R9EcP+sgSIruAXbYxk+FGKaBg/lrYNq4Il0gjGPLRBUVr551ZlXB1my5b2
ob2ifu+x3tBFd3jh5ENLHB+Mgd++138Tonh5TIYL40DHPM1PGJbepmluzfnrIAb/3n9REjulUewF
zniNknRg+x/dTQgq973ocuYWQy0qTzzi9P0tHJzhg4fd7jBGIrHV2cpO8+uMtXivBjuuEUqT1q5J
a9GeIgXgiNroFHt1VoVTdLaDZtvALNnb1mRQoXrs2HibGbyDIvIoUN2ruvF2GOEOCysPrDA8EndU
No4Sw+aX6cVgLhrJChAPEExn0Xn//MvfhfRAx5EGxq8icOdjZtsrwxLt8gmBnvittLwhVQr+DS15
IDBAOJr4PHZZiKF8RkpcRd4hDW2CD0SAZK4yY0CZ4ckJk+Rg5CLGT43gmm/hty4umsKicIWSIND2
vSuo19uapvja7ER2MtENjFm5o8lhZFQTqBTpbMBeqDWnV+bhucrnqqX2dTvk8NuN9rke/v2eNyGN
uGA9iLNtHL3ZBRUA1JjKc/vMO6mslreOkJc+z2p3o4yBvY+bPtfEblatgExvbwvw0+oi7wwm5wpq
fwsyz4RdiuHbl7nhlvtYTBXwsRq1gdYZO8ba803hXlv6pWutdIKP0SRTE315GiUr6x3T0IUDXb0D
kCcIKb8CIbc6POLbAby0EowjkLDthK0L8AQficGg/d6gPz3xfzrgnqeTL9otHkAvyyGMZa3GXWb+
mYl8xcc+AeJO7roSQAZHjKn+iYj1wPkl4tK5L7zadfOY4xMVCobbAsk0B1ZBT0GzRWQR4lO48ECu
rO3jDNZOXlMm5WFjQnxqoYd1PR/DY+6wmPjsAEJe9iQrcXV/CbaZ5Ub3ZqFWAeCsxzkb+PRPrOfp
kHhpWCzf2nOJXfuBlq/oET1x/lEE+LLIwcPoCtIlgMNbX4P2QEkyd62Ei3Wz9QHk1oJwqrvTIvLd
34bAwUgtHnVjvo3VVQ9YFCSW3rWgSsz/puPiwtnZdBgtx3G8nGLxyl0flhFXfvCjo5y5A+invumo
9wGdIpPbQcSpZ3v7ZUDx8cY7pXTOYig1cJEpy3WKHUJgSkwLExrKPRKF7EuT9lURwtBOwG9KfkkO
z5Hdw6O9GWlODD8XhTSzLahi5/AN1FZ0VCdT+m2kvrLvQ23imqyWb9pdJSF+45CE8t7Mztpao1NI
kEomxINIpKwkoV0ZF1Qik2ISOUQ9DsJKzQAaA3JwlHWxWOJNeIDdFPqDzfTIJ3tA8C/ym1eQNmrJ
2N+IgtgosT07TgE9QgAcyBGyI8SPW5mtvffO6aBblnq7VJQKbuKpfvUfdIoBVulcHvyJShGwP75N
z3qsQFXfez4ERWA3+BwuzryQngli9KpwA88R5n/o1I8gdufQzWIs8vVWgN075CpLXGEdhWqObupz
/USoNZulqNXd2CCN31IgIvabqMVRMrh4wXtkfg1DNVZ5nGZJjlXsTTlnjpj3YQad7AahJ4aLwiqw
YhTPvI9/w7RIMX/H2vMnMLoxwrnfGiPQwqIYGnmAHaqva7i/qLKUmI7PRAOtCw9Q2Pm0gNLfD4bE
19e6FNMAN7Osc155sqtGy6MeOUvwI30BFKX8rFZIxP0QvgNWsW6wPTPjSksD3OH+P6DKeA061p7G
REyi4Xax8nq3x2IPldYpPSNM4O8bBdmLRfNjQmw+JMZpNN9oBFrZ+QFI9/bgZwhM+9kJDw2Un78z
7u8tqDTrz5Xq9sXvkHz9oJwGXvdBKDVxH+qh3eUtGiDzal2/R/2FNPXbsnX82U2JlLvwcd0GmvsX
ms2Y+k15viM4gRD4JIUQGbDGBf0dODbMcKY5sw2eTzdV9nrw9SDZDC5dexrUgZyJUg4fp6Z8Jk5F
7GlxhSzLuIvHbDEsZqSMwV4xqXCqOBQDLfKo/1f0mh0RtPT3sLwU1zZzJfY4So1ZSd62g5/ByEdH
Ug6kCs7BBhZpnmyN9igs5BgwQlCmng5raupZo+ALh98ZuanY4Cg+BxoOEXpdE+Jlj/WXzCTZzK3K
gl80/zNokmivzsQvRFe3xYLwHI9aTqAEQZCH7WFhPbV6yQKphDufWVDBUUHqOfEbkXbRCqzYjp0g
tL7u2U17ozQAsQNIeHrFwXx9HIQioAhqKZ76lD/wy4j/MWoT04mz4RoZmCEoA7UtH4zsZvlNW6at
WmIKw65bBOpTUfX/R2xFkFRz76AjiAz35ykYgWSaayrWT7SYH1MvqWITzCYHYboA43M29LPHYzQ3
dFHuXRy+5aWnZmAfMIXin9+CmmYgdTOn4ncQx1nAY82psDhdJ3otFnAY2/Py6wljNpnolIKVaeMn
Dpcm1D6tSV0JFGc9i5+zGA2+0Uc5RGho+op9OFE3WiTScvJr+4V9HyEpFJdbXaxYuW9C2372DjDb
jylMTGQr3AieSlXiGqmJZiSMfrmEqp2CnOh6py6puOaWZDGHW5Wn96ndAoPVjsyyIpbevBLkdYpH
xW4hWgM7AoSoyP3YTWkMGPvb17lMJ2i3DsK7o6CR75hHZUXqa0KSWiNUw5AnKDl9ptTZ5gjcvSZH
q+cqSL4jjwcOXkMGZC9R6GQR8N8gvalQsao4qbbJWscrXGih1jlO4xP4QkGR/DlUA/H8T2hJe/Dp
CpFjNfJPv5szhbQMKGk32ORJM1H8+7q7J0p8cd9Vo4QyIPJ9tD/hNaw/BX4WpvlRsgFSPvNpndWk
gfgMkbMs6BeiuOTquax5qvMddIZ0InYHKLhYQIw/HWaHBZv8123jacXThpGqsidI1f/IKb1oyg/e
Cl7rJacCgOWMtX+CHUcSvs53NjcqXqs5l9Dh3crMSYSy4edQf4D9MdUALV/t9LUdpZKJI12yqAxC
EkKcB6Y4woYKrWkSq0JFFSv5qzHR58sDshX2vxwA5mSyRJB7mTFvw/XKbaapGZoa/UieanpNh9xi
fewJOyrdEBrft8SmdTBljQ1Vpi4EQFS6Toxu0FmnwImgX0vYM6PA6fYevas9MltJRF/UaSKuKZMq
opCnCF9QknbKh5AMjcsHQAl0YH8sV627nDmZBvXMLaHrXWfRt/r2FutVNiGmqaJiYF/+FtKCwHj9
/ntFOHXEYO0r5AVdwn/KwYERoJiW4WBry3Nf60PRb3Bbt6Vjq3iJ6hg8xLeRAklIN/PoGPwEO749
7XXBvTdf9xe0Co2oisNZTwBvwHUTLilTADzNfD7QNR/CBjQN3bTXgMcnpjm+VUOBz8mLa/tVjDCf
vRyNLoXk7Lzu18G91Nyp7aBllHULSOPJZWLUB7XEnocQdkl7JK+BAe7vm6TgjF1UBfILhAqYL9WA
CT+myFaoMWkrbuYVeGlu5Ejej55tluosAH+kxtEo9r++LQ3Wfrc22vH15IP5a1d72tF9QjEOzbtW
+J6jR6+1b1SzCNjb3HlMh/ESk0ZAeJwWNp3MpnoEoTbBBuBAa47mY4Y2y3UWwFIsUIJ5wimZLA0j
mDKPI5w5D5vR4ukB8wj1+LikiECSIOeYDac6ExoaHwS3gq1QyLLCbjmzIzNf8+pM1xokLWlhnpfS
VmDFAYqWQ1BTn3wj50ynkec/cdllUfBPyEbODp4H7ACwE+R5EyJcr7g2sAuFITR2/N5xwzD/w1tc
YzSCr1xhl+TXD8SJUfZb//RZys+QaszUyidT7659WJhaOs0KC9FzDKdcK75la6HztNFtX91QfzqR
hpfOBDCpn11F/qV+X9/1SJoSCUs0eu1jMym978hoNt/hvfIB5s5S2UJnWt192IvvxMkAMw5lPkDg
c+aEa0JwpV+8BLIVObZtcnU/JaWOqPa7N7BivO+S89QhtzVy5wxY+ozrBRaCIZVzXaxbb032YFTC
1DjBMgojW0QfwvDVrk4KQ1QpSIPf+Abbm+YBV8Lvw09NvoL/iCdyfsUnvuucoFgzHvD3niGuzRr4
mCVfRrZG1bBQA+VE96/e2vWySmf3sjKpn7E4CBhh4KSdevkw/40SEKYsUcFmjZzA1EP6dlFSHlYE
gGdunwoQJIDPOB6cUHz8EyHonTRLdkkbXWCnXuH0kVjr68RMASACrJfe7lQ9fV4eQhrHt/7qDmuq
cJcyIZyDjOHBtt4x77ESW9tnrv8D4X2vRW8eeucB0ktvBG0CVa8HpInEUDxsUgh+cTW5xUAvMQLQ
/8WjLPGsBlr/RelgQHz1H4zNncxiseK9Iedd95T5bC++mgG40DAXyXc+ge2WgF+N1rtGgOFs8jV2
rxt3s7X1w1oWJy29wnph1eHYLFtvXC25Ul919eR5hAvilPTQPQZjnCTmW+RJ9tH2hMEmoIl3WDQy
8oYeA6jiXKj2q+0s7jghk2N5v8jL8KNTUD9KxpzfXEErbo2ZYIDhXYDPgjjy3qX0IzYG/lXEjBx+
WUXGk/D61ubKIrAWitNZEjTz2FrUoynBgnlY3q3L8ba5E4oLySwzOmEKUXsQihH0U24mvwrNE7Ah
YMV7G4VTFJIoTDUUGXxpxEC4WFdIaclejQxVg2voqbEI7GflhLCB2SwaOiC5F8Lyf8NggqnJhNeh
D7r1bSiGHIgNmTrMG3ICkRiz9MaKl3CJjjsKDk+2115rRHJ2uZSOhw3rz8tcHURs6AY7DtxivNnY
+o8GDbSjMXZL+fdvPd5a+Nu/LyarrIK0O10TXt4KLaa4fPT3i8f9KOaEn548z9gJI97HQspoMTJH
E0IgppCghmjPqBL3EVZTFslVnEzb/V+A5jDTEHLy4h19OpjGVz45e4eCu6ZMRcQUk2DvVa5Wc5+p
FOt+GIY1NgsBKBTKMz5JJCAFz+FU2BnWRYuhv5VaERns7jKZEi+ZITpNTK15voNDgLiN8Q2fz/K/
X92vHecQYbt2i/Wr8KJ6uKYkR6ljwx6MAyrj4BRmp7Vx9QoDxDGy2DmQu59nhbc18HKg4t2xy4AK
lEpMBzUWynA4WrjZUv7/5HMTypzeP5sEObleF9TUflPCC51PuYhWbdMuuennr7BrAcENqDhnX938
XJZg4izqzrTDbfFE8yZFUdbx3RSQQ4DudBqV2EnGBGWaq9VkdfZE/cHtZGL21+YcYRCe/SEWL0sx
ZT5QQAwxEVVi3C/kfpkVbk075j1WpnRV0rw4mhmoE9dH3np1u1IaXNsujPLYNZ72XWMikNZc48wF
mLbkGY5mJcn4vH9kTnhUJWxdDfbTBf5KwHQybFEjyVjjvtanDCXulmWYiD/AWibcq2aP9/qFtHa/
pWS/Zsmu3ZEGo9ABHRI9HCAJ7KZ7dDsxDgR/Kv50avVF2k+LJVw3Hdim+1iZQZnjwMuUL0lWm1mO
dTkClsIpm3dgtS6v3RAy5CDxt4AxqpCyaqP06XEceeXiVqnsXWB4tRJpj10YDE57cX9BpRH/CfpF
A3ughucSSwXpVZbus/YJBeI7KVz+t1pJm/99zY6LSa9/K7+6ivDdfRU28Lg3svBgU+ZQeSXv4MNf
2jCdNUXlY2UqRCLDmWoZ5x7qG9SKl+RK4KXZcZSadozmyDBFucoXNw/vgbBkkFvMDqbkpx7YfOyw
cY+hRM99hl9zk6c+7KwSl3TAY4NoRx7A1CvaL9dhYDfGz2XvFPwZOhHbX1zlXISDZTF8HFErw5o/
7pCb71mR/De97u77QGBRPy8+FqdbAd7u/pOVNx28XCGxsGfDS1Pt0/PRndlAlobFfVmpxTRuPvxL
B3XoN9Z18CZXAHFtmB4QD/KULbKxZ1Z/FKdAhwIs8RWZO3Kx8kDFZXo3/rK0XIU1gCbieMWxirUy
8fATQxyYNoKo2oyNw3SC2CarWMmABPlIMvyPMexi2hLnPYh2SdUWUvlyjzP2hJLV87jr4XSHU0CN
80Y4hyzy+m0Zee7WPXwKnZAyqxUpWM2wzwmE/Ev7mcBC0ft1q+ft2rv7hMnH5Ch8iBxhXXig73p7
RYrb10Al6G774qvWWVoNnreaHLbHbBDRdOOCioFFinSKfp1WNokkr3jy9bhLQuQL40XciPfvmIN3
5nRRJuZIqXFmsIqw1RF6hIqOkuSNHnw0IxNQg75OxzkHPgw4LO5+VHfgpRUtfnmWl1ndCwBDazWq
TDe5S/YJKlOAB44CD0uHYZ1p0Ti7nsdUM5i7QKH5ikjSWZUBEOELzwfMV35z4Yi58q3DGLGhCBgS
5bVlIe/IlxeXiDbmDx9XZgv9sYpzohN4WgWbuSDunM6+fTiVxmN3VejI3WlzNm9sZ7mUJQ5yDFI0
+AEYntcwx6skJIhGxorFRqe5i7UYkAIYF60kud8ACXfq5R3Nv6u1g6IkWLgmN+rNycTp6gARaoqe
2GbRb3ioqw4VtRNyUNakep3FYXZmoASmr7s2ItSdpTxZwQxB5TSHN/xyXabEaW4ke7NUBKyuPh6J
0GD+eQybtMcU6WFGgSL0q43Vvu+ToeyrSTighGFr0bqwZ50e68OJJ12wRPN9t5SEyk+gVrhPgVnL
92iGytl6KcxJYayDk2Yza6LMJq2yd6o/QFRI2CRNJuykYG2kezY/dJLg8hu7uCuGxzGGMjLPvwge
u2lUowvUMCfAB4Uv9fmSY3o92OSRYpfdUGOqTMkl3zTDV4oraPyQNicZ0WFh9UdutmT+4NpSZqNU
ks2kzIBwpZ1eWhh3dtObJv2QZkvogfaYRf0eIZILBV1fs/l2H1EU8Q2T/8oBRTo/lrla20j5xnRv
dp+hXmoEHewxxCRps1LgDSKduoUpt/p1x7cznHaQsF6oXaZ72l52leysq1b+IuxymauKes/+OJiW
tLQhnUEvXko1pu/bI3jvMI6npV0T2KaWqIar5fz3WyRzSPVyCMVqAMjZ5IwCn0w85c4uVStjjt3K
IVN8VvRO1K1G7Uq6AdpeS5bOp3PEAkJe4captaGGZjPEek2BDHIiu4sLe1ILb0J++V4XcylpnrVG
rHrg2A3+nnYT1rmBgsiOZEuTnLUGMA/zgYfrADT59jvU+qI+uhm3z/s0jrnjuIjhqQvE15jsMiDg
dnVPgJjGUUr5yHFL0PkulIS580iu/gq20YadOaC5kWADaTxzy3b3t6gjxFa6AFJi9V0J0H36E4R3
g8peC1Mdyayj3bdYcJfFssuUNYwZqiGM0aTaDerwLEPd+RF5SWT8CRjfQ7Miu3xzGBEZ4cDwXiET
AmD2xTmYkEa1qNL/pwnKn5ByvRf44FPDEvFXwi4HxOUbLanHrbSL48/wPx/KkQtiCUYpZKkeuqvc
89zA0fjblVymf7FK4ex22jwuBQInHeDTmXzRZHYUdckK2biZA4nmT1T2OTYqboJJzTfAjvjlJTEW
YeA2M0TMrq9nHeyPSq0WqLmGcqBF813IkaFjtnKpf7W4+MnqPwJCsmUXmZfOhsqfdfjdZvP1cnJc
qf9EU8tggKZfJAhzGe+3FxZFDZx+KVR/a7oc+pi4wC6CtLFBrDIlOFpIHCfFCiqrCDlQ//Q3RLTp
P6+x0h6ibCDDDrWpngBAwUQxu2YdS+z30hm0jfkVkz8TLyTGHvH9E5gYogYzm7WqGxmJ2BOiD5Ax
GNPKLiEN1njw3EVA2zqfhgW76qkwwHAp++/K4V9/utwuA0Uk16u9gu1U9QOhScyvHiNky4m4AWZ5
3G9oCeGOhiwkqqK1JlXrug9Osycyg6vy69kzIcUHcXjFTtwsCOwpkfYlnw1mtxOYUQR+LbtzTcG7
WT1SN6u1Ii/l8XYFv/nogo7IMpVG5qtYBFfAJEzsuSDbUVA6m/mZas7WBuoinWwmT1mw+6O0DRa1
FTze2wk8FbtzZjx7Fb1Diir474zpHv9wzph+NkH+EqOrSrIPgxt7WrjbnNV/gDl1w3LNr7Q9caa1
h/vAQ1ubvv5gE8H6ydpIN9nYct2uR6XVnWBYN0scHKgGnU61fGhYJZFr95qzMVjMySawQ5s/ZVuu
+vMbb4ExO4U/EZuq9PjYeoMGMee6JYAjYzorveG75GDaPYLtcGUbR9LaCOj859aTxavwZHTrxvcZ
+Sm2ODyqYXKg8kXObNE0+Awckzuez0I5dl9yIdj1XuKvqMV7h2+Av+a2mIGBr4S9mK4pm3B/XMXX
iyWnO1u1LlBBGx0D2rUv2phvGQ1pHYLZa7Yzyy5k560Rc7imJNArodLmX69QYkZGv8sFlPHBCNeZ
CBkCbXFg/PXWav4dWGaFKVhYZusE7tkACkgW069KKFWub8/KOE3VFaX0MTlL4nUWCczpgSFA85lZ
TIlc787pOxUzIIWbhN9/uLv53iihlV4cuqXtpl6SaBfC4UHW49+Ef0tMzA2IFiJTbqkE8gCeOomi
j1RdzUxxiBI+quSxKc4A4LtiwRwYJ7YLlCdpr+6HR/yxbpxgHIWC/GZoJUSzUq1sBGKWGGg8UzA5
oBGNpuJovLLMA+Yk37eLv1HYhhwqQQwvJXnmWHOx2iI8NEYyb+yXkwpECnQqC6J+qv/UP7CYwsJX
oIUfXfXkk83s9AKvLEBuI1xKgoqz8j5fDcfhHeFwT9jjQmxK+m9NIXycUVld+7UQJPffGkHEH85h
M0/I+Y7oWlHP/WUGSkaPTh8X04azc2YIW5GgIiLtUytmOf93G/XTrrYbql9xmI8e0ZdHGJbb7txg
uxOXlsmD6kM0Pli7CXB4RgGU0WPlSEqEreuUxepkw5bD/xlqkjlOMa+GtlJfagXedMbc47TCoqfu
aaEgZi58xhNlL2EqQLLDTGX7o0wcJPgCH186ghAc+BCAbQGiOnKtPad2cGRAUp1wrI5SNboRrndV
y4Qy34BFnhrCakbwel1OviSaf8fC6dAcrMwQdK6leSqK47fHM6NPeDfuGc/k3V4p3f+TVNmuEZxd
U5SluIY8DfxXhgH97zSHOamDSjF8E7xDx7nCgyzV3fgpWF3TbDeNRGtBSQ+yndnQm2USr8K12T7p
QnciYcs212UjGGi5D2/UyJ3gyC9EGm4eC91ZTurRVhSJHJDVinsKy0PgAIDIYbX6WHLPgR7bXiMz
+hxC+gWvUajZyUKsOz6RHU7wVWyvVUqCYTBPPR9+hiY6PbPWc+AOHJaATo4ihGssY1smx1OXUkO3
SHHZIcSv4XNhNjEqV2kGCAAuBnKa4EtbaB9jgh7jHnUp5qDzJuBHOtoaVEIlV8ta3q9+JeNzwgV/
7yKYcmh4lPfNsKElMtf1SKHgaKwD5DKeb4rjbSBWDgsCDabEBmwBxcMzLR0c6xoLI68ZEkOWem/E
851hzNBsjaJczWWARqR7BdmGimGcBvzv8QsmMzO49LQ0jKoHebOzQi8d91ubeF6j+bTZ0Yi6v/Ot
w1uyZ+lXVbrHOwp3huS5ij4YQgMTr7R6/c5BTzEby8LX6E7rZ6rC9oIB8eAHtfsFfd2EcAoc9Rsh
T3iFa4/dEXit822HuBct/iD/HKDaiyNpY00LFqNdU2jirdu65UVU64quu1JTj4osY/CiHsdmpPcg
W/xJw9J0iIh5GHMBMVzPWrvFxqJx09XtOqpHkwBZaEUWUgml9s5njD+7hYo1WT3RNGVeBwO8VVXt
Dd7ylsGEbZraiKYb8037l2CKaeV4CBTE3kL6ypVrD9B6tOZFpiAjpsVWdpHWy/PB4CAbs6wHA7xV
58XETKrUd0N6SFjzwIvtN03otcYl2SMUvt05wEkCidlwaC6VHlkUMpGI1/mIDixkI5VQ9LY1ynvA
KDEEjpssU8isS96dHOQPx0DYzKvJwdlbgaaEmCkjB/BdB1AosI+v40nlCcuJ4FQQlmCO1ijUVF7x
bO4yKYsYBH3fbp+s45Zdewbz/oD77ZIv4m1fw3oxVlcb1mih7bsXcjAUCi4UI3+YABQ4R/Jth+SE
yvDrGljlka/28HLW3XZ3c3DQ8pX/vbRBB5KsHyie034clbeL0mFGoshHMxQEd9rVP6EqDQ4pTd19
NpFqTZRDhrl/o87glwvu7wsjuECXZ1P1RiHhMqcTsVnUVcpqDJaYcM0sS+sQc+lsRWN8Z4/eqS8x
M3n3eLt/ievIcpt7sS/MCFVR3Gv5spqfwgvgji86HaXtklqBTE/pDNrFCyZuUaes7zASklKPbnfe
aJxJqktapNva9kRahuiGqLJjUI6AVtM8Xuangeid5b3YntQZORk4qs6B6jBbYmsvgc7bdKnhkxf+
OWN92HwNtPT4K747JwoK8Xyuf6DM/MAd3o2xuk2RhoXCY42HsuWUUcc7IQna5xN9bHZLTjcaHvpw
+sOXro6pdTX4DhcQIYXYPuJChKKgKmFQ++1dOzHp2et6tV1d8DsnwhmULMoebh2wknLo5C1/Y5YZ
HGNItr7ot2odbdqxcUstUgAXrBsj64xIGsL/WX+2J1hNFcT9msaGpjoPgC2sVp7yDErdVvEcdVjZ
tHNu+mr+znBhO+NSeHKRkokQXEWp8nE+2itWwcqQ6VH26cs1Y4Yt/1Rs3VeZLIuhwVJGWbzUl4sh
0Ndlx40S+3rUnlgJD/+KGC91B0D9/n7QSLZ8ueu28aU6zNq6lVd1Ri7WXSozWqkzykTQjUCt3d1A
5OGVstPnkIP2OlKILFGEHRelYnl2OW5FdEhwWa5ZnAJbCRXqGv2dUQumX5o10TOpkiY/8LbzBOzM
KBhMFCeNNPNfLB53DNf2uOHMceWlZdoa8a20w1gIOQMOTYCoPSk0RjKp0b9yMudfJ0K68axnFwuu
jkun2PmRo2Qqz0d5LItpI71V3sQaWgawo7s3xCy64O/zVfGT27QTuY8O6m6wO3xzHX6xguCspYdZ
sKtnjmHcSxZoZag2ELyC7i965ZKVP4TYkQZ9ACP6r31lgrBi6PWIK6EOoMv75iWfiZzRWl4izck7
te7fueB897NU2RH57GEt17G76F2B3bgnMViZ9pFHiUnyd5W+t2PRvYvtp2ac9vda27Tu21028DZ3
2zxwVMBZBwcZWYha8VGFDrM/+TdJy4B8utiYrqzCvkb2//CzgAUXjtn6sO5QXcICGoadt9tNB8h1
jKQAIEm4JOyiXAZvZ+ISYJ7cYSaUEP3x5HagXgG7Q4udc7H9uDvLfEJSBkmoTVfCsIl0p+5U5vvv
m2hgMjKPhC3izGpmz1PVnJkpfnbmW2Z8RPWXz3Q2wZA9QzmyIw8U/Ub81R3cPVMCoyAlMP/UH+Tv
F2i2T2/PLqvJFw0mnR06SRZ2Z3yYbX7Y6pCIu1NCFbrJGtyOkjfIw8tcStZZqf6MCb+jTtzeTtVA
slOQhkVEf129bmx7OuCA33xWvREcw4B5cp9+vIYE3Mo+xEpSzrWIMyvn6w+BdRNPVEXimuObuS5v
GXBwYxD8WLolSwJQDzOH4CTzW0pAoCvZhz3mOIhlyPZkgkewVeSMs2QBJfzIoHm7iVR22NbeIFQ7
A70ILd8GjD5LMgVn15Dgh1mCKDpT1FiOn5W1QlwENuxZ85ogCFTmfl+rXbVVnzyWzvdXtplo1QpP
cYRreYWyqEGRxWd0s2fOwSxdTJBq8EoktXAn9mHwN7Pm6lToZ9CJlPsfP/VfsgUd7X1XZvPk13mw
OGr7TsGwXgrPqVPz67r9/+h87Zjr3n8CV6pARrNs1tO3J2qCP9QPr/l2CU0t/9hIXmrApnbcaD3c
VZFB9DQy3QeLuAqb/4RLzC0x2ffSc3ffn8h7Z5Ncv5q2vwjZnuw2Lqw0Ii0qd3XvvcjjopYygrc+
uxDMU5J4T8ceK4furqOpX7mIhkPAkzZupLN1vfsTC2DT0+aGOXEgmKtLBmk+QvGBIMmsfXk1wNy8
mv5N6h/pdEYsLeVa7OsG6QGg16Lj7WFUxycBKXqV5MWtuihWcpDPiR+9EHaONdagS1pziqhICJsg
KGbi2vPl+m9j4Axqb/fxcLIjomOKhqoQ7iqCs2XJs9bFXJ1QQW6njvsm9t7Cwoakm6y+gTFTezCA
JrIq1k4tS9GjthDYvFQazvoGU/QJC0WYng6c/mtmWy6PVgJeKqR5f5qtaIBiwR1Dpl+3hSid91vw
dcg+H4kcyJbWZ5QL5lVKz1pALnZITnHNBYJwFNud/JcIOdeQZbGQrGkjJItzJLMPkwnMLv4xZZI1
XTQBxPUu5Jdokplqdnpzff0uwCQDiho/pFdko1KsMc+xqqGlm2JK24C6+MINf8VycQh8c2Ox50pl
TozzY4+e81ZAMrr5oeAb6TZGX8F75WcPdJLiLRf6MfThA2z5wdCZJhi2XFwFkft9xvzGrtRbDz/z
mq1yaq+nn9WG/eD2I8ZBHN/F0AQ9Cag/nr/AEl3Jxq2dZxL7AeITGwBVFkm82RyhUbd9tMPO9e9y
AkJEu+eDOFxfUS8fqVUo6xqyE6SuQlVcF0i40rLTwcMiHE/7Z8M1PxvGYcabF4vY1+VIKDiXVaS8
myF660dLY29I4vwJF9YqnzV8pRT6Mgct4o1kCTs27pR96ZiVKjc/6hIb2NsQ4iYQD9ChS7g/3MXX
78SXJykbM9kzjfgMhNGvfKle0eKkR1QjFWq2WWutKhB+/aggGF18NPwvlRv/6LXviP+oI6+DPbo9
8bCDcRrzy3Kxt5E4xil+v6eWOW2UGlWUhF5rXJF2siHeo95C07TVzmtIcfSZhCYPACa4+uzEjJaB
oR+AG/n8Frn06x76NNT3rE15s3bUooQuldr4JVmW0Jz7maUgZycPrqEeY7WaR4ScScZ9lVcHpUwh
LTVWVkxbTSu2B7biS617eYa4Y2EQiTzGpG2cm+wUkLs89Yjg6WvpImVNFF24+O3RH4XzuW5ah2su
6tWFAbYRbmN0kApc8C+GnECY8ypVrtqf6UECPw2p/iV051bUv9Tu5/sNonu/ifoHlzJqE7A/9Fvn
bwXs2crP2wkQhW6HkSY6DoXcpVgNfmQ8QaDRf9ZqlEaOkEcRVeuvCNeFJoKj+ZnM5YJ7BZbzXHkY
v3Wh+LARg4Nr+YUxJeyE/hw0x/3FTFS3EOEhIPSFfmgJhn1w5yGUYdt5+GUriTa7cDSLnRhE/E0L
ZctRg4GCzEDne5yTOEg5/OVTzxxeTKz2OqpgK18mWOWG3Gg3qGrb6heKvwHxzaO0Wjr1EkgPx3qd
FblB8dNTXA88ILhvg0zaMXegYzW9QIJ1Gc1gKD/y13YVRfEG/mkWLfwF45dn+hIxF3OOUrDfm+xz
1vF4RjAjNgRZy7VkhLbdAfGXwpCZGaLNgkiWjtmLfzgaEA1JZO+xZ/S/3HGZbYLIvCFMzOnjCtPq
JaQxH5Cmmu4sSLjQf4CgTJNUaAJ7Wmn5DCmluIZPq4ds+pmZqVlOu7gFBpWUUkOV1r/xsuV4CvMn
JFJ0Fkv/h4efUR89aRrLsMQ4/YVoUN37pgH6twh4RsGccL8fH/vl81NSPWpH6wTPYX4arglDE6dz
dazXXEds0bBLDHK73BW45y/fyleFxG0BapRw7ZRaTQgoJsr83AFr7GHEVo0TWXBRPppFjIse4RR4
uJyjlcMqEeypYhRmk9BguC5hjEZG1rKoj2QNt+3CVWYsyvXHUmlRWTyCx+gMpSb4N06FGX3gJ8k1
wSYioPwtzXqUuAaEhUWGWkV3zoqLXjJQQEI6zKfzyh5o7qluE1XYp/QUlFYU2lkkGD5OrY56S3y7
RbZdX7a3o9bsVU285oTGYK8Hi7klGi/XaHWLGhTaEOeSjMTHzLBccvXRtfPBkf1AnG3JwnWSsmhE
4b3IwCLjvlKPnX18tNLWpSBw1aZ16kzXxYbCQzQOo1fB+w5AioQUA5PCS92VIEYFrfSS3xJGbcE/
X/9LayIMEPMv7zeYhpeqxZYXbFbD60tkR01+F24N3bXIzyZTZf/9ACKIuSwmeOEbWToSl/q0PGv8
EcL7qTqdnhTjcJQK3+S0J2ObYmh+pIkaIdq5ow8K4q3ftU/VPGkTKtUgkV0mj13nhKxoT2jFuPFg
Hk97x3MVWkGJjbABas4l8z7SgmEUdLAJnoBjBEjO1N1a7BDOYEqgQ8UoPYH/K0L9zk1sygtWtISQ
EcGL0nNvUv9Xd5SZVyKbNcqwZWEmDHV3ZAXwitb5npvpvkPAtK/RJbhHYgYmyBlfIF+bX6pQASSG
aW6Bhn9T+Mgu2V4TVOnpNwoGLG1x8XyjFRayMeYg9xDMYKULMdoIfagbzctcBrj8VhEzVOn2PW5V
B31Y2KfW5nqcEZoU9r3UCs+eMshBcMomOo8cNjwMnFxOalozRMGPLRfWfdwCdswaPDKJAon0odQk
elx2QEB+T8vrcFpyt/KBsDWbdc+r7oDG/U3u0Y3do0ioNUfuT4DI/kNZboVELOg1lCx/Dc0DBMUD
FM9wXE6TXGonCb8AfPvBOas9fQdJYMY+fMN2P5dENk+T3Nbn7iMXvtMZqPryE+YOUnJrfh1fJ1LJ
snGuVhQNy5M0c7yvwOv2QJ1byw0g36IBYMjs26k8z6GB2R3cHm/3UDRbEGVYKKWD3U8m6XCtyjQq
av9q8RIZIuGc5DE/Bze+93suHT/2lVjQ0QTGfT7F6BN+djvJ8SzxYM5ht7U9YUsf61bE+cey4eva
uHchzt5Yt3ymJX+YaC+QAFtZ0HeQE0CFtJGyUmpPpCOnIHu0tt1/M3OeqjB3iTK/a5Ai8RDcDL8a
EUNj9g8hynvsF2R07NUHG2wmkf9UpKbBptYJK9i0bcIDhBwD68ryYbd2QpjqrLjiY9vsPDK+NItj
x+SilRhQOYQpTc4zDtDLvS53WG/O7ttvV1Ny6UT9jxPnKO9yRu6743KVz9uKbEbP47S+w0gAh6MU
hIqIV+p5RY2rRHV5N8lg7JXLjKnZOxLxmX0hw75AsQBgjkqWwlzw5VgQUbcxY+YdUfxEuDOA9qRX
ELbF6X+FqfJMg/8YSLcMEmPJc6mAjR5o761bKG6vspAR5QRGU7c9g9Gz3ob8IjjyOE5iv8BlHNW1
d/v/NYtIrPp9949OgZlTNIt9Md6+wTsQJGtJBLUIh5VqZTLO5yn0esKFXsQL+/c1BeA78OWg8H4V
6aqTq5Puln0mnDwIiBOgj6lIbGTUdk7zImuRfSkPfZnnYI2z8g7FpZghK4dE5Rd45YTok0oFzx/t
bTRw2pVsV9cv3VjGmriGRNmdomh8xJHFzTvJ+y+KbhWDtSFqVG0zmgxjN/o8DDL1hzaDCrIwlC0J
suwTi228MfbS3sTGyjhlr4WJ4d1Q0f0ct9Pn81fyzSSoYDw1UnmpSvI4bPMj80R8ewl+oHBheYIp
UXjN77MsEl9ifqpQtRxO+YmDZNlgrNy9uV1IyFlTCLRVo7YbRGuivS2uqszL9Ns8u+A/4xugP/at
/xWg9wuu62yRBXNZowaTU67NF7NicTfOBnGWJUttYKqkGRJJUHDcw2Ra/mrXa9Vq78jFQvSIjSGN
xJyU3yHllR4gX6Sxc1p4mxHc0j1MoMkYHnXZuEUEVvQakTazIvbKLtacrTswrqtaUSOEsx5+Sjvx
4l2IgakagCbUkJopszSP5bRf61pKi44pCdNZyqMLbZIGjJiXQbVglB6bNXIE82i4XS6aejCJQhIt
ZmUjUR29Vbz62e1+xQnylXLV9frjLuk8LrNAbnFe0jA4E9jZiztKhIG81iLCfSd+Goa4NMckqixP
rdMjd3Y2nnI7ByVARiwETGJIa7I8naMjALa/nQSNrgwkIzcuYBIlBlpA0ObvcHhHLmOLvoYZ3bfx
0HNr6ar968Ni4zgwohRs5cYcf4j6Xf9WZq/zqqyg7+6vEMxpFgwbu6rx6d5558ixN5senr1ZwUje
7BgCVvwoaUp41xKyrTD/JY6fYxtFhZsI/UWTZxpWpdpkSpzTPorQ4DhdZGM3l/eXmHjA9jsvHqOA
TTin7c/eSBbitNfib6SzSuLPSTF2qcl5qjNs5AH3VKYIK7tZOg0c14IkpgDNEpQ6XpCbE6YRYoJP
323mh9/6GA3RYj+yRNlpalbvEFCsOxxkUx7kVFyqxcsWw8hGo4j05EJFymkQcQlfhgSZRZTWwwfB
aGgKX1mJ4jpP6943AaXIk/a9aPhfQWIVlMOpGgp2d2vGND2U7Edp1soRH8TwrN4Do3Kk8VjoV5a3
mPkY8eCd+NoZhGSN+T6XNaD9Bw8pwiWUzEledcUGmnbHNR2I4e/KEu+LBAxhWECyXQ0wfl3FNThL
MnI0vGvLfy6uSnWjo1h8TV9cpFp+VDef8zXY8FKaEfUNXdyR34dVZrBW2pt/LOYYM/0WJrvuPhNR
Rm3Ta/+fgLM8gI3QK91WQuc73IngHoZLOwFkcXUWFEEynYWBDknU+RpJ+CWKCXj8NTROG0bkoolG
X5sVnt9afAsnBSga4q2OgHfN2GXDlAYeWGpgeKUVfuBy2COW1Rgxsb53S/kkggRQHIktv5E3V/pd
pdHX5yOnRFJM/thNv0CPtbmJ3R6YyLKSvuyWBSP3iPwt11/IeaojrbFHJmPgFAT2OJsMv8o8FRWO
wUxyyg4acT6RSIcr/9Mo5sZHJijA/mSmHmH6lVfUKIe2x5YQ+jiRH1vBVbubxYsYTX8yytinJUvw
SzjIAL4BMWUFpezP+BHwffnpSwMLORKQpuZlMK5x/uRpdZKdNnZ28BWqNTB7eJT2LUj4XGZTTvTZ
F89LyhF80/S4LeJ/OcCZxPm5sx2HhKx8oVRcfIg1xGWF767zy5OyKHByGtnm86IFLg/TtrNXkG6Q
hH2ywmolA+EhLCdmKepVwXrxuvkqQjuuqoW1TMMgEiknDyouS6dt3aHIqemCpIF9VpaHeVsP+A2q
J9x1mMYNMMttIaM2wGPb1i1ONok/nZA62yGqd9/8SXJkHm8uitUMTfxKdIgp+5jUqoIZC1N8tUdp
tI+TmwZheb1n9wOzNVNMFHlChiK/YhO/RWIZZZFtQ+WTyeQSLP/F9i0OfrIrEsp77x/kEYnQ8584
CBs1l4bRG5he8/ZF2eUAnIQPoJjPqvxSVqEsFRYgCMo8WG0kks5wNs714AW3z2Y2t91HRrOfH+7o
9mY/2TGZoOSuZu9aydn59Ne/8ce4jjEjDEjD5hmo5aM4iNXXNLBu+GvPy+Hh0AJ4P9y65izxE8PG
BI8DtbhsOHp/E1k0rWSjUTqtiOvrTUjkNYZW0AE8m0gIq5vVmtdJSym1nETJQkaza0iaSc/a225Y
Moxmjvbd1FfXDK0daUmr3fxbBLeuI9QrS2ENhSOt+wWXFJqdGJBiyyY9zHFPrdM/sQY7sMD9lg9h
PqPajoupcTGS7Gloc0SZIJ75dDHmD0wc+mi/fp6ddV+5vlZMOSY86Xz8PkMNKRYxmnQ3bR5L8iqc
gYTzMCph20zy2MWRX+JSKkupa1ANIssA54nuxrpk/k1iEwbFksaL0KUQB9p3ybVJp/8Qp8KP/mP8
RsaVGdaC0zsMeyGv0oXQo1Bc2O8kP6j+eBCf9RCQKOwSRGFYThDMPyMR+5gnnmSE4n6v0wjguqnn
YF0fJqlhqqjwkUdMpjFTzb4izGWE447EcrUZ/132eC6ByEOq1iSBU7lt9e/5awFndHKIrKZaQIpW
E30h2iXPbY94IfsRybpQB2jngxY5DrOkmQKqfszNWey4n7BYzKVQsQoCoR2/DfQfE72tLt+xEvpE
ssepFe0GbgMFVM2dZAlpEBvKAg8s+xH54Ie5ipjK0wNJdfA4f04oaiquiZSEGkwaM0tVQrIx1q4V
2pVzIQ/gYDhAk2KnE50TH5xuX47RUMLiy1bPko0meZ0crRV0NxoE7c+xKpMwcQ4QRV9VGrT8oOip
FxfhIG3qnPGqPd8FdL1odTZaogiwzPGu/p1BLqH7M2ZVXdueVHYntxFzFoj9S7pXISzQmZ00tdAl
aYC5dLm+5eg5rE2OEmn7s/VHlcEHCDpbyAOEPUUmy8eGf4bR9kQbVQe2O9xDRrNftE8PGEEGajAs
KVOsuNYEIg0gIb9fcIhYXv6f6b6awxrqpYisS99iomaAUZOG4pvAnfzYG6b1YIOOGYYKibsrAHya
/PGljo++VvMhGs0asFFXJY0UAy4a4U5DG7QSWgD0fMmjRcbMpvae74qVGMctrnR0rWVscGCjJ/Gb
xGgT5LsYgt+fWai5H0BMBOib3YPlyfNDF0PRKGSUqiOdBAbcOM7ZHvfxgzbloVpAPb0LxzXuAJ9c
IaT5PKHrV56lu1lQFRjpIa1Am356qRM13tKTQQV38R4dM8XyctQyOwj0JkNsnJ9AHSn8yIKW+ARk
g2wRe1n7JbalgWaTJ8TpirD0dan5JU4C2wwT+II/JpTSl4kG5H9XzndAq8wpX9xI3p8w58aiRJVW
43YTfsaM+ci3JLpjxJKTqq79dGuGxNqoH3qAqj1nsPV0svbh316smTZABnnluGKp6dSRUv4bcHnM
3H2i3Q/LInqJjnbhSpDK68C7UxZUKaWwDKpZ0DYdeHwlPlzavUArZ9wmL64p8MQdMy/v1sVx55I0
0lFjj21XcC4MZWhP+bBuMMlpdz1oqBG8/j7bt1tJt8WDhEhgW0YWQ/myxvJO10TBJNWdEvHPl9CT
q17Yq7DsAHFpgm0iUCgQWRInQhwgR72CPOxACMyGLxKOSSXPSHqsuZyYM5of2N9Boiqt+y5qtg64
bgq+hwhDOoW21uteU2Q6VRtyFIon5XTM/iC0YfG90Oly+nFFPqrnE9A34Zan+SwEHZyR95A6oV0C
WtsU/dwgKe/6cEEp7XVXJvAJCaxxMY7pI9EFDO3cEJQE5QeBDOkC2FKXrDjEyJjJ5obs9Eh0rkJm
Q10YhTlQ/aw+K0x85zeBucy6ALIMFCbot9enlq6LdKKfPslYaXTk/qtbxGUQQzDHIc1otpOn3Et/
0gBion8k+SSBlrZ33mLHXPr2pUPBSLCSjBy+sdFN7IsSz4ddER9zIltDntrDrxNHIF4Z6juBzzD3
SvoGkkbLQWP6EfEnh/PMEw2cnjfYiwVb25OmsDqhcZSMzWHuXNDx1rpWBeQ/xTv1fncg7U8Mq3sZ
j+yhgRwZZXsvFjBWnEMoj7kEZnyT8frx+JDsDgiabT3dBXIhxSI4u9VRmoKAt9hSZmGiiFkSbb3g
vbw/2o89xBDlTdhBjSgIRZJAoiYFcavMtZm1NH69ecDKlPzqj63gK9gKWpWBsw0LIfmU0u6Tg8PK
lCpUCQKLoUIBCLY+eRcMYi0dF06zaXO05jLv+biACzM7uDl80MaNb2hfjq12MhDmiH6vwgGHmi8+
/5rGmGzGh7dhGGNv68/6jT3hM1vIYjlLnLq4pk+tDfOUMmnZNPUosj7J/bB+6kMAj42izuW3WdTL
PNc2U7NedEQhKRt9402n3lIJYEgpcEqzrRQlviQnjA3dqIC1IJ2Gt5BFFYEfkuc7wHkUrg8KteNW
SZ92VtnZQaVSfn9XiJYUST1vKzt0IwHww542JCKXvoepPglTa+x+h96G+9VRIat4KG7AXxn/ReV4
ypGZjXaT5hvFL4q/nEZLu7tjDzFPRPxHNzeqGp/LGcLIgJNhrxRMiFZNDrwJCBCULfA9ffZNVqzn
nZKzTRzIB3bf4ybZwQKB+gpT1yGo+XdQi3ePJakVBPXJanwHiH8zvHXgo2OJ5GnOeqdIh28GnZVS
n/ynL5Ou+8n3Ecw2pdbsfaP+q+FS3jcwhBXLJVkflx0Cf8PqRwwA5NgdMtUT5d6pwWLryZri4wCC
00fMU3fOvU/9TLJ6eQ7iXXCw8vRBEQUVA4aC5fFmoEdfWmLQxnrKCx69WVwTbEFXR0gmIXEt8AiA
ogGXEDeD0r3mbjLegIO2eNIPUPuUX2X39466QxnxW1vswgvvHN6ANTSeoO9o2RVrdXxL2gTWEhDh
piD+vOfJot0j+I47QytI37byquO4LsdxXLvWvw4a7h5WO675AstIuYMspjamBJRaAG+8clT2g52L
XL2DnSc3ke2BD4/ZSqPlb4Tfw3Q0UzD4u1jRJQ6lVAiPGnVXaKk3yj5ngp+f5kFjLPmx8ZT2XZ+X
n9aeV3H4xYYM+E0FEMRvVQchRIy8/tU8QcOxIYHBIi8luO9J6BTmcVU3nZrjCIySf2Vk02pXAxYK
s2zKCCCRLZzs2nZyT51aK/XCK+4NGyx9H8upVf7cCz+yLNUm43mUvK+05J3uZONH4XxEIbzaIPyp
WTWytvJrN83YTmiqkeYrtB68EHy6FpxPaVfM5xt5Gm9grUU1xAn/WOnE5Vf81SA8RB69SbXXYKy+
2o3vJqBDhjAYRDQDVNaK3CfHnOH9kbV3Yt/TPYMavC5WCw7QvMjCc6htcNCLCZxRD0TORDBEcB6J
PeY7QbrIu0cVAe2ZXr4xRVXa/CNWywVUkvd/zmLkzWt4ojFr0CsR8kIgH6WEVpBd/4TLF4YPtcNz
CsZVZy6KpbPnH13n6ZFu4qib0tviTn3Yd+2t3jZeCamTtK+G5/ZRix+CjlTaLDr3F3anUNnLkBrd
2HeimIfDG+OnpB/oLRyBtiGPkN9eLjTcPcea3OfTO0h3sNX/v+eA60rj+Y71un0gh8lfc5f5yICF
PGi8n+lVSxSBv4xd3sSPeDdGZ4smxWSruFzLXhTeJvKdxdfFGlt4YEUV/TCstalcshS2/JTFmrtN
Dz4OpCbhFFne4WQuIVJvWphAuEYvmwaNXJtYduA8qNTBhXEGYX7kABPlThffrKWd8c3TkhZ//+J0
qyNwAjyuUhCpVtrgAT+xoNhWPpPHZTegH9LJhNmuTj0Ltj/zQ1ATPkk++H/Nz/EToiO2kGv8F8yU
b+rrk3TrwWjhNPdzSd5cbBmtnRVXwINFbH850d7okI7L+fcKwHVibmNfxtmsf1fCnvAM51aNGIZ+
HDwWD57Eurw1ASKYzk30hCijpif10SXG0V8edQ0X39TL9JlRNPIde8uomnIQJn8ry7a0QbavWRFx
r3ECKJqOZ39iSnqjvQGTPTgUDKk3dWbv0M9pWsbNT18Bryc3Iy92eQ/uPNjmzEZ2rNPYHDydx62f
/+2Kex0A+GbdYzxPuuVFn+6aknHjif4NjICwgXTw0ADwiy7MxJ2rgdNr1ofbftZEj7ejx7Yk48Jt
WtnqlgnxoOMoGG9Q5x4Vmmq+dJ1gFa1L51FUAqaaPEjNvw37dXGKNTYYT+BuumGroGKOYobf+SVw
WbeW3R89V378kpjEkRcL/Z8DjPBdTPxgOfEfZrplY2ekgruefxVm3zKHj+whFu1ALglnN8Jwo//F
UY+fxr5iguf/yENcdVvy13doMPopKPs3op1ZYe40FuZaQrvfl2Ri6pCouqcihQuTh1V9l8T1ggKq
YMH/2QIseLppWbkHmizMaW14QlSTv3euHvBLW25RdhTfYKC3WyqTQPiwHW5t1xDgk+PnQFTvxajq
+Eg5yF2ztGCxV8jqr3VsGDhoY6c4fWsoz0hsSzl0UpAE6wia+D5pNMfEsTkwwiwBrLmodSbwS7gR
wPUrbD/wpLMx9/mABBL6q+/lQEab7TpskRIC3TW8H8/dTSv+WigU9DpAVHFmRpY+218PfBUQIKrB
tC7Krebj4QInTm3KHOJAPIIb5kXwntJGlQETjlJ+07UMvnYMOdD0dHyvtOf4HFIbcsSLx8/QJzDC
Xog/09WKzSI3SWXxxV9K1qzVIdo+BFNABU8Hox6ifE2JlA35V6sKCR7niI4Nb2ceZk9Aq82sx+HK
FffcBapBVqVsUAhcZOq5PUJPTNdCTW79RqXHkNkz+4xwYmo0Pepn8M0myHlclwnxmw4m1yLP3Tay
PNHxnsdV92iFBTM8VIbO8odzJABA++FodkozLu5Mqeo6hMz4f8rWX6MuC6zqV4ky9M81CyLv/C67
2vCQKvEkPNbXodD8xPpRnPyREUiKzjdd4vPQ+1HSC+DaDDyT7dRBRdvHyETd6d0xALzwxMwK2PHX
c+z5qYJYYQqM8ycnfF8z8+rVqudf0o2vnUT5WwCZKFx1LH5pLX6OE7MQ+a74rbFmc8odIZRm3x+v
peYDUFq87qZrBLh4FdXRmJ8iObiSOX0BKnEg30iKNyU7ypGbf+BI129UeFUCTyfPFxyQgcBLSVJj
g1QGBre+szWzNyRwQ8doaa4fpsnHovLJNxAVOPL7fTJGejJL51P78Hkb4wI+t4hGtCRfagFb/xHo
sy/u6jEVdJeHfNvlEYJaBN6s7Qz4NfVyzcU8BMVSv4g/7RXf1hStNcZCoA5tBUW2q1YKY38gUcKo
T2v2PSYAS4RazJXnNQpEallW5RK+nTw7HK4OTBkhvSMhnb63T57rqIMFC/t0AsIIEJGZmCo5j+11
AN5pFkW0qEXz43i1tIDoowqzn6eem9M9nDIcfVEF9Mkqn9WY6rS61H/IlOL+YsJ2KUNqCtxDhdPU
j3KHPZaPqLUfp1teeY0WlIiX+hqG7vO/V31RObxCkMG6/FDviRN3RpOvm9z5eol6Vbf0Jc8dP7yx
DrkcfhMts7Wq92QcEou3XDZedN6d3U1uiMM1JvMim2iih55bMmMjQ7yAdSQAX3ZMipTg51W2/OdP
1lJwucX9bS7qxoe8ZvD/Qv3ottluqhAURBfok4Q1Td/QYKfqhoLhVVkpKSSF+eqD9QrgjxyYRXO/
qOywj5y+fIZyUe7AtMjqATuVB97aLgG30uc3XSlta2PVEjJbC7xQ9IJLbsxba8ACYyxOuLkGZ2yB
m5HQMGZzbbzKXV+mbH0JGwzuFDYbRDcKP+dEk+00KHO2AYtXhDrbXN6KxwadJCoDshOwiSDYDSNC
lJdDoe8X0ccT8CMxSLuyl24HC8kAFuART0JzoFuR366pByx2VzuMp5h1IHcwrQ6qhFKdO835ZdOE
319bGtfOD84giDiiZhFRsJP1Cr/gLxQTAtLjUyKsdhSbQDM0R0/O0C7VwM2ANqHuYNWrMhVB6NuF
y0j8PE539vnvB48LGB/oAr7cNuGk883QQb2FhBELnKWdFLL9ufy1lhdgN25tIHNhhAfQXGNXJRHT
1aeuNTEQgP/w0Qmlojc8euhu65m/K2uWWhoEa36YcQAvWHyOTDAKMBO0A575YDrWFI+qkG2FfABK
dbZG71pph/yIfToxc9kY0ScwMQnaZALJL3aUibJWiyQIBEkbtbe7xh1XnC/W3SlXc9hq/n9Q3ZYc
fnDNXIfUWdsTx/EAE6YqgoJhWDf26o1wjpqMtW87exQePo7/8m/F6KbEo9ijoZHYFxOrRaWUQXuD
jXn3RbBPNaAMJJhWakalLj8/UH+sxX9d+83U5rpt67HDSApBds/jyWs7Ng3lsYllW0eN11ZgKO+D
VXHlNmop8BRiI0QBma7AB4CLYWzU4NY5yz3IME3+pNW0EbL9oFKxFb60u6v57EFEINAyNeWIUng8
0yavT4sIRIFiVRSJDAh27hNDMX+iW+zkq7TpoSGM4JvNDZcXEVJXroYTSOpZb/zNQx+1oBW6ywHD
DngPtLI/bpHarENFFt+mKgIorW7k1ysuRuhwxClycljFPs7vXWQTsVh7AU1pIk/WlYtbTZcN2xvs
ryV1Yl61BgTjagFWhfyTHe9KIQvXcbVqpdwZJDq5c+/r1HnCVmdjuGCCMD6qiU1v9AX+dh+gDjbx
qBMIwSpNvSkfi4fMXC6jKnGfB0Nvy6x7euDJ5uNSZheYFjyCuNyUmKoFyGLHTwIf7U6P0Pnqj+3m
UiSy9t2jA/Nyat8Zc8h4XwEZs3u2EkiT+oiF8+/nn0+qg0UNcjurMF2wIB80jvggDcQm6vNOLjub
IeC6dW2uCzuxIutcRZJwFK/3ryrjaaExjcFQxoyJjaN3y0ooiWNK2AgDZXh/71fJF4XF4aa7VPoO
wxZJhLPAkuC0Ru8pYNiVRSe6f8uIlqZxVXTCt7Qv0d58f4CteZVx8AZ7kdnQGF8PWSWRAt0Ka631
xcY5k4YBO07rVze1l6Gcd4Me0xOkQS4Bo8fdyz6wMBgGh54GrQuJ6AZbMiChSdIoPofFqAWVx5iE
jym0ur4dy6TS4Zd4blCLB/FqwX9RU9Jz1foS/R2uorXriifH1jFWqvXyTtyIAZJ0+5YPKXfbtzwS
6z0yk80+2/XZ5r+eqrkKod6r5tUf+HzMuQD05+FFrpox/icn7UEPvl5d6lVNVS1K6yzKGq1OEpjg
lDCcjgxxG/s67tUlxPS/Z/A1VC0Wyuyz/N3jGZZFzisZyTeEgBFVBRrpFwEmFMilVPgJDeLRKH70
bS/PBWOFnmcVuYwEv6k2WiXPSaLQ328ZeaCZ/AgFLt1BYu6cklURZ8pvYnAy5vM51UE4pnPYWDA5
o7c5rJyv7rH4ILyZrQUdcY9Vpk1mep5ZQpDApENPRqv2fuPZGq7z4071Zi/ZJlLT5pJoVLVktzwm
9dYP0RKSXxNLGM1bc/f0SrByzqMx5kvPhDxFPeRZiP7/yilvNPeWN4KcCq2xbIMZGCfETyMtB0ee
9g2ZxksgHFbaj6+Aji3nHlz9p6UF1gY9nNGPh8iw1X9Rhv6V/Pc0M00GkMio+cK/b5gwOrCzkd/w
k3GHkNCn15DL6SREt153VzQSpe0vdgFl9WLTtWZvCJvqeEwcZZZC/14Gxt67D3cURCI3IxDTMuOr
U1o0WtnkE5I3Twsp/l2DXpYD9GRfryhBLp9nL2rE5b76WVxGCL0fSRJ94g5l9PpDZZaUQPebK8zY
YeGrDQlguQX2D65IncSo6OHGHez6IaB2XL5HnSg1vdViWSU8M8EliTc1xNbl2nDGBf5kWICY4onE
WSP0mthS/GQSdtDuJ9X0jfO4w1WgXopYpnNkYAQeMJnNsKYrlFnzZkRw/LW2+eOli/O+bctVK7yJ
PMeN9Y2jlQkdvMAFJvOwq7owOw0m5T6bCsQWpw2Ys+TqJ82/B658aS/GFc/PUgroti2HPr4SEk/g
km61V1dyXBH6/KX9vHyrhZukgd9YNKKoC1aPkdVZVsTvsHfooQb3BXv4v8nJkTX43yaFJHVBqB44
ozCkSkOPguX2sihQaK+HBrWV13uRO3E8uUoh4fz3NDJ9m3OXSbAW6r2L+/P6xAkaIZZxuHSFEJ28
3ObJmt5a8PyGDg+MscWvMhr5qC5xVKmHBh5kNTEUjTZjDZZUOhLitgdzEwWeSMSrshXlp+SvedJO
KiNxlxuOWkXgPgicdyUcuKy/2uds954k+avkUdqdSzwYC5o/iwMhB2wp7xB3ehmRvjF8BkqbhIQK
EW/FiE7DeOh/XzvLZSvQCTdJQSzJRzutG1hpz3RDkgD/0OlGi2adXzeWmetdkSvAlYXS8B03767q
DcWF0hn8x8BGcRxFTjiTxyyVKR+Zbg4+RSwiXmaRMKMXcMqwJ7oBiFk1iPI29/qOxRYdzE0vYjBM
L0v9RiWYY4YlBban5cjuS6+jCAlr2RPArvI1B8b2plHp8wJgBMIHKdKhNbRYH1YTcKKhk09rNQwD
0GFtBd5NC9UszFCeBwM8IRGlKE7SV82v8Dco3C9vmV39gOYLtC8un/8+UGdFKv/VU7lhiL2Rfg9R
ZOytuyZdW3spAYlLuPG/oS/PxVO0OpcXtHZ97jDcp75ct+sjkPfNJotlHPBpjQhD+7/JJsFvP8hp
Kj2Nn92AKZqD2CPaj/+kKphxYB1Jg+iuqrD4PZ6uV3iejdA5L6CwhhT8b8yFiGNqnIihGcOJMGiK
lZm6Zb+/M+6gUoggLk0jnNRpKijHPUqKlOqWpLpTI8Q0/JP/MtT9qJG8NVCNltyPW47k3O+xlDyx
bOji7Jae2IMTnpQInKE5p7JAM0jgnenqNuso0CoQDIVLMcvrZxDvZRWnqagAi4KH89DDYwUgtmqe
jyT4Dnc4rEwx98mT1qjvjfqHYGEPsNhEGLGyIerlhuJHWDGB42imAuq1Zsqk6DNWjFFH16YaSR4/
EVfaevBPuTp6RVGC+bi2eCeJfYCApfx7s1ZwnoaCMjeJqTzgLnS0ROI7b9b1bO5gMNKM6STuz23u
Y4olTXmkzmXUIiPa2il9VWu7T+q06sE7VL5z4T6Bx5HlhQY0ZnpuQ9SVPR58uq+jVubCzWXk/7W3
haqJu1YLm6B9O/3GKTCPwgQec6QlrCDCYryi231FLYMRZ8qxmZ2tMy4v8G86B65N0tDFCovMygId
nBzmOtJSdsg42gXYD1o5+tmar33QkpZuIKqDgLZFjvKNkZQW210c6YxT5ydRqPAZ91BFEKDYCJId
rInVmNyHXiw7rDcpyrKlr8k/l8dbo9Mvt5r2rfI5sD9fAyqwTIq1IlDoMk+a+4/8I7/RhsNAhHBN
A6EKHp2Xzapgh9WP14s118dZ8///jJM6OCuOIEOmusmOdd/97sEr+P5oObtI5z+M1vLDx7RVk5Av
J6laayBM4532qxr3K0e/P1Ll4IPh8WVxYm7aCDxmBcB2O/gOhS66GO7iJWspBKcT+eWD5/o5CNRq
04T8drHN7JE+hehu78F9KI3OcM3ASQxKahhcWCUNWZNL56xcRcIK17cbZg/OoU6wv3D5WxDscfiq
LNGmQ9Y8VhzGVhCRk/SF310QQmkdLs5ZiiYCIyxTJqQcmuf1o0s8cYOXnLxX2CO+5w5CLNMwym8V
hu57gRrhLR0WOPsQEtVqpL/FgeKVZjXkRCgQlhHrOZF0HI1zQH7fYuUY3rncXBuelyiu/NHDc137
TnFcymanF2sNcsIF9mIqWE7zO0yPOg3vpiVhMJog9/N+zx6Pzyt8DsplSp3SyP/OBxSIK5/FmVAt
yU3c6QdLnWy5JSUYrn3/AV5MuhDsik98RzeV4mNwzztEPV2Ul+h+xNAxdJ9+C5Sihv9evS6IEGOq
aB3+UKO1j5tZuZDuughkpGGBcErI961hB7umMocN+72UvkpvElfYykeWg+htjZdwYky0x6HIG//+
9vdARCfY42hg7sifQjWP5K8bn+1tZpsuUofWKyQoWUSd7yJICYG3BYi7BYl8GS08rfnjh1hWKNny
eLWWRkUdBjXHBl8HW/nWc0u0QcNOzPeryhtmf2uxjlQVW9kaIeqGzYEhn0+xQGDDqz50ZhRwDEOr
Lid9u1gKBNUAqhUJMxdLkDGy0psJt5xU9r+Zdfm8LJQUQZDDUfsCOvrtCdSLQdDl/IVyyRw6nqrh
0/8XTDsHOXnMJXOUoZCZNw4guxuhwspZ5Os+04lQVa7vAFTd0nGNdaxG5DfoXVPpHBE2dqN2EjdH
ppPZ3Jv7NWoqE/qFmAB3W9YHKx/ybq3C6QAtH3l3X8g7fBQHmiVDpUw4Btw1GBStT8M7vAb4Que3
0LeARKJ3nTKmM1/8OJ3zotJBy9dZSzJpH7Y/tS6d2WvdcPnvjPzxSGzb5qp0rFcB+oFI67xpoAoh
VsHpGn05tMaxMlXYti6aboP4ZLJP9ZKc4hf+HoWe/1d5gKNkmO8P+r6ezzeA97AXgVduFk2QLkEE
QSax4T1lujzPK4oyyNm8oPWWFROedjzlU1wEIRaOVxIyAhvg+MhtnNPS7IoFCI3eIAbTdNJbGVXm
2cI6/joo6PBNsfFp9V4xrJqYFzWGczRlbZJa/KTkpLCsIWaKTkNfzHs4KQOE/x/zzNEgnwUaqqfR
Q6zS1qqg/Nvww32XVtHpUenRqAAr9u8+VO5Jly2O8zXNTEWVr3Gmyim06sMfBNUDv3jzyEMzrcdH
tH9EV7dWgnLfT8+TJ3sg2oUSPjREusBJZ0tV9gi21G7GQlfMygzBknk9AQaejWadyx68Fi6X4ME3
Oo6mPb4sgQH9m3f7rRbh24iGvvpZXx4J7nYdqvxd3UwdKQHySPpvyOJPAI6nYo9c6O2vXqcMz0F4
XkWTTWZTxVzkLGVvRuSzRKrH4ANSwqHbqPP83yDWEJxd/UkrjoFERVe33e9+OHW0ywZm6rFC4m8j
pCSKr3IZ/dJj17S162ButYvCrBqsuh21W4cDYYWn4lMxMTkQH6XO08vR5WGnS1vchfoUHEp73XvE
EFEF+vgFuFxVCO+EMDQoPsJTMxFvVVhSI8fZRsVXi9+p9xJc+E9csx24EHKxoFvs6BjZLv5w4BWj
wZqJriZj22O8VBMfRzQFjJC5iy5KapckzCrJhN75qZRPApFka1CxK684Gc7jipQMMTeO/fGYYNdx
ifyDBXfQFb40kzVJ4X9GjgCc7ihcYWWDIXw3nPKzW7UaadgGGK238t3jjXL6XxMrfQrPXp/j6zXu
hVRCV4nVvoUa2M4ORXySea5V0GtKbXX24FyLqs6iK4BpGRm5lyxks/CPtkOTofrlRn5E48zLTgFY
mWODPVbI7lDy8nRImdnQOp5XvRWMRNAAUM7s5rL1dajdo0hGIEFUPmLpixRWdyQw6qWGUsCYrsVm
vp5Y51IOgXRG8caxl7CpIh/tdymSLsO3MxU4vE+wEDqfg0e3RBQtd0HIQiLL6HYYMD338OIu3k1L
p5iuFn2PMQBBatV+PURDu9wRLh4MgvmBIJRTu/1SolOLrdV3f3PUBhqWjjFUqg/aUu0fIYHmdEuz
2XkZuWX2NghDYYvkN3L1dwGCiGhqgC7rKBXvBPfnpJ4M16WQdBco92FNiN1akAp52GIhQGprStWY
5E8um9Lbo9lYfkOHLb7YsYuyJLaSDEQQLnEXH5pLmk+A48C64Jlg4Yas0D7eJVOW8X8bTF4B9YN3
uUUmymHATqRS4f88IAss473cjaqylf6BFFPWL09THKBV9wb3hor4DSyCSczVOHnwEQC4P2XoPYwh
MhQfuYM14cajpdfNChuywuhYh6humbcsvRGOO7J/WcjzhPUBUJPIFRHfvmeRp0lfuXjHRb6TVVCZ
T3p1/b4yuJFWwn3lY3rakNLUy5qa+3T4Gkip8j+2qpwoW2ERL2qe+zMYQce1pE0gt0iTtCh5at1q
YlGsvFgnd9FWykZExFzs7WVbbCDgsJBtIU3WHQAoMqLTTLjGAqu6G9/RVhl7vd0H6iXeBXixBcIR
Q0YGp5YdMJU2NH3n72NWKjGssbR5PT4T5EyfQAxrqswUevNZVUys5VmekoPygRbA4G5pN9ghNSlS
zlVGEUIzdZDcgM4LQlDiOotOzIPjzgCvm1Upsmnvi6FJEsY6YvvNzQVbfYjsjwzEW+CMAP0upB+4
crbGzKijagTT84rDDOv6Pnu0D3+/WrLh71ejHaWmwN5ki1q2vx6nCO+9f1yQfzxF61S5bHAoID6t
dyDmuh4fgRAlciZYKFJehLLBZkvqMovNtFOGNNZC3O9xsG7+DTEJsuZRQRM1J0TODUladZSM/Od9
ZultbndqdfLx7iQduwXjJnan/FwscYq8m7I5MzCS4838P+5P2h02RrEtXsB3RrJsMfqLU/mt5rTJ
5Ln/k7JKofU7nfApLvPzp3EUvU2XoYyxl0CHJbatrcwI5ofQ78SHRgLaLvH4278VnRZDBq3tSdnD
gI625jX8K67HICnXJB8rU6R6QTJNQMYbfQkkDm7Wt1RzGq6NpJbjrccYkGdNxKp1pOBtL9ZtQqbO
3UgA5oGSh3aIb+TaUetdoDv3X9/CrzSogVYIUWVy3RTU+zCPwtvw8gcCZD5O91yn/OGeKqdbZB7W
NPfh3Yil66GCfUPjqMX8JEwT1LEF+Ct7Su6KdrEqHaov7pYdx5KCHTJBwDzaa8AmrBtEg+mTPtxM
u/HJLr04ei7ZHc4/Ktxx9DCX72/Aw44pxSJb8Yh4vzMEYlMoEPUznf0rai8koR0jpNB1ASNO5C2V
0tPeWLwkl2kdRTht89EgWSgwylXIOwliyFTGLryYR88g93QiX3cVkxRFVFylyU1OGcgxcJ7n4vzG
QUOhTP9rhnfyVtxf/9FP80hDz0jyrpSjHnYkcFfPT+C4bmHLFf+owYYg6TUyBVZqlCkhlZKXOBBE
tfk4xvWE1H282ofQKvvYs/4YclslMpo0VbfOQIfeC/A8O/dO2fYN0F1H2nUm1059HFEt+E5VasVZ
MnOs4Ey+7mv8jtL9GgVYUX/5/k/3dkSTEhlIJf7lUhJW8XYXhzTyK4+iElkl9y7bwRdJOyfw5CqD
/81fbaSN/Jglcj/IwMJwIcak5m5yvyayq+sfEZbfKsmqlPNqnPLWXDbwNlL3dgeI0htUcI6AGPIh
lbWiyK79B0AqDcd6S0l07B6CdyI4ENUdyn591+hlFQq9bxCkfSGuxQr7v9dOkTFPmHARD9eExDGW
35U5VaeoFQTWMb5zz7Qr9/+P1Q4uAuxVdBYszeXm90yowE8bnBbyJM/mGXoP42lISNbI9eKZgUu3
1zZleOUjDDk3fpXUf5nmp6RKCuuw+Tr7UBh1yUEnHyfwXhTGewWAv3mF/jNf1JI3wbFVDKquCnPW
zPcTkpY2xPUsN1PyeIDsdkAbWk2rUAtu/+pdP/zaH9bMeN1TRYJwP1PhMkA6G7LyFwaAXLCHTHN2
Ur/I9H2mKpapuzZU2oSvE9OxJyXr97BWlzBE3e7ZVi0GD6JU3nVOcwbk6d4DIFEGRSjTnIyCrq8c
z44/uC5BJj25x5zV7SbX5uPEPfnHTeDVpOfB/UhvM4Fq4t8Vyja0tjOH9LZtIr1qLEUO3NZVYq6I
NJLyAlFv7MIDYO8ZWqktRgSZCBfoj3g1Ql7icf2B7feDVgqb/NyWnRfu7e/o6gf/s2FPL/Cx9CYO
6336JSG8YqMuAF2SgbgcmLMS1BAuY6zxGL8W4+e/tsKAuyH5kvWnyoK3bxJsa84aZeDGVeyweKN1
fnooI6RBDWOAzWneNJiQJOSQ7exW+MvAYFu1bth3uNBkymq5qk2OwO/08XeJ867b6jIW+MQBEw1g
FTtjg03uzHpgYGKUDr804wCQDGi+K54V3U1DiJD2HPpEI/QMSuhpL4MB8psUHXZvT2vP5+xsAWDZ
wh9/B1m9jFyCtKrnfhfoI3PRc0z5hNHX6TZgOvXrpUaMgB96Mw5tSUwrwIVj1bW5X7bs1KFnTAC/
5aXTYd94n4ZlGNLysAF5OU0in7gjsIfZKnjAyFRVcCs+8go8x355V4mYaswVQ8hHSm0ClI03J5QF
zZSisYnH8LsCAaLR3nFjOxTdAcktwfIT543VNe/El6YnC1pVFj03WxfHnr7pdnUNbxtd5NXoeDO2
6GeUdtwCoalEOzbSjRlNUjKQYylRxB0zl99uturF0Q+y75TSwNS/QNO3jj4XO3FoW67aYOMUEI3U
/GEuhS0WUr5bK/joreABZ3W6QLCmC23FdJKNOpoDGSvNg9PIKBdY9UEbmlLXB7evKV3t7JtUp4DM
46MaGDAlCAo8d8RWBoK7p6I+8h4rtnSpV/VBJfCgcUipU+itt9gAdNDy497RsoQ71r0j6q9LBNW0
XwVBB5tXaDMhtAziA0pQ1u0JizYvLMNImY95Tg+GE3q7ZKzwF4ATa0FcaR4am3LzGvJhJMmtZ4Uy
CeKiZTJU4FbWtfcYvkZGtbJTJk4HSjEQGAmm/nHc1WB+qADp3AmljWKicdIInZssqegM7wWG3qwj
6isinha2wkuIhK3aOb0BFNAkrNZghIDpJ0Umg+qNnNuoly+1MtrALEyT2MFH49ELqzhpY0Bb82T5
RpY+/NEc6mgRNdu+d4f4wXFtEsML/rStlqIU8GSvndFGpVnivUV5spREPm0LWpCt9IZ3BIShsTbh
rZPPjcUQ4+UarP9w6WPQEpHUZGhaiFCJ38QWI3Hmy4hk1h371PZy09wVDQefdnFAxBpdiOIwDTpa
aiJyv7xvfMWQPIcHl6sQK/r7Wasa+8ra1b/TuDid6H7OnbyNPzonaTVG/d61jA7/kaX9Rs2O7/bW
I4WkT+3Q1EImV0yJS33C9OhQ5UEz3am9acjeik4x6PE0gdq8y0ljK5HMarrksOIEDPKT1EQnPRGy
LCSHjRN0Zl0g7IFjDxq48E/sIzW9Rt4ysPcK7PJSFoxSTQBR1qI9TinlR6Ju0FJzrPqhtqazf4Wi
Ftm49F2dxaGT2bpImza3+z33WHj7N1J26oy5Q8xHi01YV2NfngRAQLeQR5nLflNfpmItDBHCZGnA
TuRdN59/RXz3wn65fcBi9OgQn7RvBK7aX+0JjOZGesDbcPjYgsKoQ+EaKgHNrApC2KZEJHypgD+O
byEbUskkvevwSRoFJoOdrprwl6ziFpRNauYNjAph+B7ougTGNs8NcLndJz30ngejaLKNWq42JW0A
w2bMnqjGkQ2vEarEUsVcKcbP5OPhxTSqgVyTf7b62mrLwvabUYuNr6WGrJjB3FjSSzG98a3n66Aj
UeTCHgizIrQPCskaDvVuNMoSec+jWrtzNzIf4hylPWF6a7R0PBTgx0UsbBdOfBiN59c0bUR8jFtL
lbNBNGAkVkjwRz61T6dnfzdxLBpfz2/bc1cbQIDnmQze4qlUwZD0Z7tnLrY118L4W+Wks6zdzrY3
2nUOMTXQUjhFhlVik5z01ffjl8E8vyvQYDGvFlW0ctxXiczg8UesWHGiIiIdOLTvVBM/GrRED7hB
dqhyfwQY4OWvxfwtOIYSryLPpZe7lN5avdOO+LNBNxsK9+suKvPtXBx4tF1Zrm0SRr+RkygQE5b9
l9FViRPXPRBC9ZtZCv2n350iumLCFU5IfWZsSU04lYR0nuR1ECzuWXVV4jf0OgI3X7CR+mew6QJZ
mcedX1sUO4T4gsjvhZk+f7UBIQmItEeW4YisGa0ZRJS5MVVSqEkkv4UfjRx9jGINCSNoJ2EGwWvh
sNRDkqRE+0hvJkY/Dj8fce4zrjWqH703Zfy5Wfdfw2FbpSA4zsgEY4C8p9JKixBXLxJZ10XUj99H
o58RhDyi/Lxgs7jLW0UwcsL0OStKRkEOXBjAQXo6yhegmJXW7T/EftJd5oEk4iA53PjkZFnAOQ0M
buKsZULGg1D1hG17usKOqRJKv8JJogiiUubom3O5E8NUIimSAPTNwo6X83P9iIY9pu/iiQKXUC+0
9At1U1u/Z85A2ENa1COYQKdLPvzc878HvdNpJmcxXDlXsGEHgVAf6jQJhBvd9WeZFHgcmQIrZU5a
4g+BD58sLi4twQxk3sonfWttvpJrevCjm1Ebr49uOX5kZA3CA23LRoEhwkaBx/5YXQAveEkjnGcj
dYzoJqO99kVTtyXYtxQU3QKiet+m2rWqutkx70ahqH5w5b2gdJkCdmxUSnK26e5K/0EWZ+gptuds
Ug3Co/W6iYnJdYVe0a2DdjRyCBigLmGdXcpwJMCfagqGf8PoxuOmUS0s37ShaJTSS8atVeVvRwF0
GsguFmKStzcQRyfiJhKLgvYwMX6+QI+h76LGpN72qxE0Zu5Ea0G7MJxY7nKD0tlyE62raMS3h9Rx
/zd2pbj/s3zffWGlURRIYNF0zgoQESQ9QWAZaaOKQRhp8wTmKyHiol45ptpbgAK6XFhN16cvrtJP
Vt396lSrCL3NqSTLme+GMo/yvKVmUobn/L920KVLsf1kZx3sBo/ugbeIoRNYxOAoScqKZ16v3LWj
IAdrMSY+STZp12XJd99yxa3wUhTkfKY8MH5IM+n890ZN9zPoFMj9JgAPcXSJcvdrCL7vW0GEIvxc
SxuB5KIEKFoO2Grk3jEMf3Hq6M2c9cp/4mw6ChRrCAwVVOz9VI6mTSEjYZ/Ms2l1nvdrbcZD6Yn5
l4msXB6LW8x63Xj/scZG6Zjq/pLxFdxCIvfrCZHgchs6EVswTzoXUyNuznuMPuqDT3mwKyeJEauE
I8hIW98/OtMy+qthXWZTxz37uV/vycQJ/j93Z8Nyov3mKK6eAhrQjcDSR0tfnoxra72rC0dSh4uX
Y2bwuqNWBh3qouevB/KdgS3iU6DGMrp4epCG6NZqq0UbCSOdNp+7DtM+xmJeQ5VNns+G29Af2+iX
cp2VNudu5zZEN39pLyP2nlqo6r4uRAMqK5TztJxyyFqLfnLNTa+qABviiQx1u9kQDnqzT/7elKW7
Y2ey8nbvSXdaB9b6Ok7oP5AUQzIqzfgsmOyDLCYPw6rqSXbWGqAMdQgONEbRBaukjSwHARgIAYgt
7eefbEF+IJx+KE5tkuVK5j2ZIQtqwxZizxlakKXV+zPhQ2PVMpgcgZK012S3Rubzx1flbZzLnOgs
LKSg40/yjQnQfONheppirTYlHD89pH1qLfyAKBT7TQEP+d5nwRoKpkDCSYIkbBM8JoINHsiBoglI
muY3VSg1fa+H/mBc/AfCd0zH0hmMQo1oH8C2COoIq5AFjO7tKpYGb2PbB4/035oDz5RYgOCnTYz1
A2P/VbXnEub4whufGR0zEgshJZzGJwsPpexQjF8LMlDlmwKCYEpfEhs0AUptYZ3jQYA0S4s9kaiY
Qm3AnO4P3aSC/du2OfT4/VTiRDbA0KRysaLZAu3u+MteOrFHFTHaXInTzkXvlSlV1Im6KkDU9EGA
ixIlH02zxdusuLXXtmQpCtaj0HDVmxrrpbx94xbThoj5uXupXwz7XicnTval9FxEMiZ2mzVI6k2T
RCVzDTh82qH73xZyYGzMAmpzcIKPmR0eqrsbr5zs77xHaIqlP9rEu25zb/eTlZkru7Q11+PaQqzf
t2Thd7Cb8wEayZSDDvq6SquYgMCYPyAudr4EbeEmBeEAHxTv0SZQ1uvfoAtmodmlBH5OmNMNAzKZ
MTY9kmej4OyCtFarUXJ7P/RtyddipT3fMsLBhGbPBMfAsZv7WrcjrRdesDZCAIkBHD5KWfsyv9Mb
mBEfBKc5ctH5mLbXeie7uTQSqLovbbSbJvkh8F8pQSo+yf/QV3rzlflCRAYUEjL0qPnOuT+66AKP
w0FnH5lK+sxNnBHT5XYc8NngbkxjeRAHzITd+HLakPpadvpplTQjQxVMHWUtcwM/xA97m9TUZnbG
LiD97+tbfUwQyCrNWWpQwXeIabtCEvuQC7nKBGP+8GFjfIXMv3g6qrelaqmvdzht4iAlJQgqvvO8
VygQ1KxWHalS6lSPouOmIlygH8/92MdqFVlf1wD0QcvbHUUnMSBZDZii4ImqYPTPFXQsgHcFeIow
XbDS1dmJoKzsQaX221UxajwN8qpd4jCnF8MVsX7NR2kHSwSDbMRO6KaEQbvYR1hEGK8zO2IqLDJf
tI3xZzDc98RKzBzkmoO9DXAIf/anrxg4NkcNhe14MbAAhF7NRas8g/hluftwKM8m4BVpObWoZYK3
BZb4x1fCQc9ze9nWJ21EKw59cpIZYNt6DaH723KxXY5zC5cVRmopKyp8An/FlmX/v0POj2luTtm8
K4N+I4WTgHe2zrjltpyDobpNyhisT6QCw6Qo/My2X60eyclGwflNZHypXSYQ0krBnBp4AERXEIZE
jHt9O2sakqjfTi58gSb9f2pk8N9N76yR9d4NtTVWmBx8EO1SkbIwiAb8pukerBowvD7eF1Tsf6zU
5J41FX1Jlx+BXb8Tla6/Oe4FW2nWrmrFVZIt1u99Wy7I9W4V+D0C7u3xVYl6YcgAs2eIQk+jNfnK
jxiG+XS6uR0mTXDd+vTtHU4L38fEhRQSDH3/eR8x5/vW7FSi2gtO4ioo4dYwIzh5VopgDzDntPno
x4hGGx7AZqvQ9QP5rRa7+dV375PSSQpB1V8B/94uyS+FlZQE0z2/UKs0w3/K6j2eYGY+257XNmE4
CH59EFgIwfP0xdcRpY7VMsWZWsNayZactawM8CbKIH2evrQ7cDjoqVpea2k75OA25a86LLfVLoqD
zXcP/fVMHY4xAkawSR4k6TzMG0yy9/sP55XZWDURKUVbNKgKxCYuT2TILtckuvVVoUWfDNs78A3U
d+tc6z8QNINE+7hBRQqnWGK2mkz32qQPCi8tRZscj1hELbTxTGLErARs7mv7Ks+kJktCG4r/1TdJ
8NQ86ugPM7kqlDW4E2hBJUgvzF5sa06Ntf8VVNdQz6VOrqfxsg2dnUZ/WPBLGFsrO3hdakUPiV/F
bR6+5z2yo8+qjfwxQhkF1IK/7uHwgOGifJhXJM+9CU9KJWpnnYjvU9GYNNvVsbYsDFAITFlt20xv
2jdJachWW32/uslncJF/rAsbcPxvwtHUhawIbkAbmfA2LkI41SlXK2+F79F0FFm9oNEKojPTxj3M
ngBS2ib34zXFFu/W1OA792gkmJM71csKG3u0H8brmq/UxuLVHQ8Dn487agTATngyZLyu4FZO2zX4
MZN9Ql+lONUcS6b7V5fVhp178CkuceF7URWT3C9RAdL73cjk858llDXxH191MUaqRzfaproSjx3u
JMTst4bQrHKhUtCWnzgL2uZLfmXFBXB5MuBupnz6i+h8GQT5kGDwPPmX5Hr7U1tXqbi1dpbZ8amK
kPrkwLKmTO/HM5OKfNGoLy3HngsXXvG0afX46gfFox+K0/hLGL4ZlxEr7bB0vH+Ljipompjvx2Kv
7ohSQi+6qCPmQy3pvr/2pbJoRmX6bHB7YtB7SHbcLRf/w3L/WaxldURDoYoOSQJSLOUjh1AWVQ8X
2TVNQyauxWbKzO143p+pdqUVzL0TGnWglX0J3pkUD9mgEoxmQjP9QS7ID5dmOvgn6z6D7+TN3YCj
GeK/tK28B/ftuWQs+pG7qmGEOPvDr5XsTVVetI3kdMKsCn9gXTRbPT/e2R/qY6liMghOpsSNL0fy
YBZ2x5idTb9GFXDTrrbZx8s34px8AsUQPEG9jEadvPR/4brRZJ5oXs+wfbmsg6xk3rhoowBGF9rd
qlpXLTmlWW3qQIWc/oOV8WPxKP4A5LZgZIKRz8qArBJomtrdY6KK9VX66DY0CFVoRk3qezsPvW6z
1V6quduMQPVOzImGh5suusc03L9oOebGKoYKXJKUCNddjunI2unfGLl3D2nMH5wV1E5yxyWVqFUo
3q7jOwGUDUMFrn1CYF8y0htM4WVrGnEEhiucd4akY60SLsoigd24KLqBXB6n+D9N4/2ml/stE+HB
w+FQiAs+wFwG3NOkOhrJO54KgfC7kQxv2YMUA8qcs6EQbEimkukzncJZ8bsEaXTTXkG5Td+YWNYh
s1dgCeAPRt/SL/+xRzH07xvpE1GIXlQSP83rR/g05/1k/IK41SbrAiju+QWONU913fnbJzu085LM
06tluzJ4RNMr2sixUoG+6hr8soqBPvzJCRemAZNmerd+CYid3hXMHetoKFG1rDkScbe7mgwocszx
AC8fzNEInceuSy+EbIJibx/hx51ilXJOq7g0NGhOEUlF0AcrBw5LMqmgpWYTU8fOPhRjJvovrZAV
ns90rtMoZGlIyPjRWaMu6fcIlAiAqV8yMTQBIHkaft2r074RZeUeuABzLr4AJE8W5pON/BWMlEE6
jkWmmtoRtG08L6+mYN9CZpB9b86/lvNuTxDPiU2c++8/FWDMZFLK1e4ZipERcvmwVxq3Nj/DqjE6
fK8efhJXWQoBN4x1i3n+tlcfvHqfu9uxK7YEtDaIdIcVhm0Hx0pD7RVrtAd+6t4oCPsnDo8lAHHt
hiJRlCXEj9Gp2DHyKFVFXy7G6ba61qO5SJw/GdN7HZZYMw6NiGyDG3EbWn8D5kBA+70p9SyQql7b
RXUUIjed/Lk/rOwhV1Hg4XVmRWL7n5Cv8orSq6ZGq5YduKgk5VLaEaU6K5rDtnuoL+jnsIaqxfRG
D1zmBanUy9kfXk6QNCYQo1AjLBaaAU/1jlYtnH8bxCL+s548IUSeH/b4CPKb/0g0vX5lwa0f9BP0
xveqIZdcafA31LXWYIbRQi4VOvO1IGynwKL5Mi13iHcYHvwosQ7ZzC8vjsghUjGrgYXMqDN51C6f
/i89gH7sLFEIq6Z/sM6H2pXtTj7WWUlSLAJG5cgkJ79rfaVG5jS3PnvtLyl890+RwwHvF3IwoAIO
piZ2sJOu24sNx0eXdWcRE6RUN6mw6zYHA+jjOtSG3esqiYFcrL0Q+7d5nIU4Y1zj5yCK9Wl0y3Qz
OSbBkCBXPFe1Ctr/Mv3jfkYoD67ji02/sxBxrERtpt8MXyfvXMnB1IrvL9wRxR96yFE2EsP0A8IA
A38T4/eRk55ioCzSG2+dgyUWlT04DJnShqfCuI54RtvmFpcUHznyuVPQzwpsfTnT8wrqDksJEAOs
+I7CmrOd5QTN/BsJ5wyJ0J//xPM6hFTS1Z8+c6lkDHvYmDgjPNeBAmUKVST1u20oi9y8V6IWlXWr
5kOS7n0fiSul/MyorlZswFv+HZeYpDE2sldYBStOJF9MBNmfIUcGNygg1yLsYto8S/S4uI+ljxTZ
ZCinmRk44DrHo0swh4TPTS7mjYwIOF0ETUAmWI9qc8+ky4eXUgozIQpwkCznwGhIyF5ybLtP1D30
h5XTMOcjKuRGeFlUvsFUrb1N9RqhYovoBF/HqbDy9GfTqJTDd1C574vAONTf6gsHGesKUPtW7HuQ
jyNKyBNIMARnloMEd/yyAiDRffcj6DOM47a2iszAecM2MdnFkySTgZphWkQ4Zr1rVgYzio1Xivwd
0DnZGwedj5qAkxRQd/KUXQvL+e700gBcunM829eWicF/bXzUf4c6iqXa3QHJ9+T8T031W/RqI2pf
KCu6dmK0DjnpYWq4dh42WWpYmEaG6jNslu+8GcNjOv8uCrqyFliOzL39JjZN0TjZFyeFBu/kjQNa
4+dsYQIxJ0D3QOAP0id7IXJ26LQN8ykbGFDoP9f4okwxxP8PsdR2toUXrgvgyRfjsXhdNw+iO32s
XkGamYtn6cixD8neIo4pyMbb5kkMwgtfR7LQk0NoErpswuDnBRTbAkftK2wZMui0mo91GNUNheql
Y4B6u5sYDsS35LziCH63p5MzDdal9s1zwn/QuaXbS69cXtFUP3uZ17mLA+5yCLIYi+r2gSi8FLAV
FxYOTV8GCDZBbrQhFK/SZj4ufYTEGmm7OrSk/7fc6nuRhVGXBOwdcMS+SOlynhO4yxngUSMzEiQA
DHqrw5kX3weoZBwwHUsg51choELHscwspQY1F+HLQjIamaxcB+C9bihT4flTXhALsIWqWwALSlZj
7ujspQNiu8Fy6mECRurtnZva4zuvRFQGgdfjmkXAtkYpPor2+dOy2v3vh2GC0JgsXss9iGdJjISW
65n0DqDGbU3BwfXJlqYZjiMp/BIQhT1cS+xs2+ALQarzTpCFDzWeTLHrvD1BFd6vCW07wzrkmMoh
u7+jBU6b8OZl734+UFZn+/QD5AVqEbszMCNrMXNVaUdjhgEBGGdub1ol80GLsRCOlIl4ezo+bYK/
Pi6D+B8nOVhzs/LMhu1Yrdo6B/583bbu+WSFQ3RdBTLjG6SMrtjidx7m6kBWP6vGuMQHmRE4P572
C2t/odnmc0l9WrJWpStjONXx5Oa7hMf0wFx4WA3Ddea641gJqLC9USrY1eVZboXlmjh2o9ffQUZ9
7G/GDp9HY0zWeHpsipNaSZIFW++0B8cCi2SbYuP1ul6r+K6boX4OP24kSpHqeDag31Fy0THbRZn2
kwmbm/McC1q8ke8QwSkR5z8OyDSTiM4noRcHqn3UN3FLpzK7ZRhmIuLkT264nlMhZdQUCBvNN09n
gTEaDpyWkGawFY/rLaVTPGVr8VJAV528CE2sTqIPxjpOxUN36YwWcpaxH1J5gNIgw+nTaxd+B5lc
I0qFRbrJJ9iaKZxg05XUSQaHhWzvVuLPu6pZVTicA+sDsVWHqbpkDoqI4twN8jf7RcHd+yR98z9r
xdxj/58IMJ3WSADyih30elkZBEW6qSCsI5+Ot5HxQnD/qRhPpZSlcx+fs9V7U5Shoe+s2HMYs6sb
qnWN8NYbDRRs6oeSFh0ywJZHZmZOaEJNlzGrnlj/g2sAJxPNNcyyWDXU+QSeVC45g/iCMolA0ekw
AsHPoB/XDAiWlw8kuVsL2HCu0lvp1oCIYTU4gBhI/Ai5npgomjcsMKPfAAd3jLKhm+r/ankjYgqB
fEyh1/juH6yupawnjKsWjeG/zFYwcC3RByC9pbaSF4VoYx3c8F7pjkUxfD/DAZTqYAOa+z2GNuqw
UBYR5H0m/SXCLRj6g3Za9RIxWiRz7MSnDiiuqlN4MNi01ZRR+68oHx0Gk0BDoYAvUMFPwCmkxji9
SRbagn9+Oy/ZJynot5r6iTArxysJRbBUbq5figZFw9ZYzHO0qgClJNW6qF2pB/yNFwByvmXFNNFu
w4cNhz7GSvLwmpwF9J6RyqWHrq98S3e/8UlXf60pJW6zlVwKGQbZv9iHOqaQ6SrYEOn+91nIYUtO
7OEBTPqr9RN8Gj8O78M/4MSsCxPJKOP+cFWNv9CsW/2bM1OeIe9GjX52qgPxHdWdSn+bY1znA8q/
fG+3NNqvJutCpQfL+Ps2u5mWednxiHZ1kqNzomxehjytPrE+XPGOili9cCAu6v24VNr6hr9fiPHF
UXyE9PO1hj9Q3tXm5EER2NO7x3eH1BB6Fu39/Av+eV3qLNi86x2aMAu/JH7H1HYFlADN1zQaCqKJ
fQFaB8ta2lCsn74gq/RHmscd3t1e9AJjtRHVndIgY09rsAVH1xbCGGYHRQIODXiPWEDzuL54yZAw
F4z9LamlVj6tJo8m81Y1ZWz2GsgacthzBYzBeRCrVrQDHfdzDaHTwUL7XIHhdi51JvscpNtYodAk
ro4EIVmmoV5G/GHT7UQG04LvW5pwdIKAQ1ldWRA2/VcvbVeN7eiaVMc9c2p/5VazI6MB0CHePM8t
rGFUafJ0SAwFbdTgfDBQG0lWINO+gDBxd0s5n+xODmPAaC+G6NLWEzcJWUDN8vp72wnEK+0YIHbE
hYUbwjiCZ/31/ZiQlIl2hQLJw7TV3HLYJlF/R1yRtdMo5RPz5jDMtT3LV67hAPw4NpNS5OGmJZ90
IOxJVm9m08RIkhJXT4Or/t2SOMi/ZCHGSp8uC8MYNFnwYiOTDNRj1m9lijX9Iffy8nfsRGoeFc50
vtfGYbqFlgGivvPM2lqQ8x4zAo/1lUtgdu9DOYDTaW9x1ExILFNvAkgRFO4fZRt5yva4HY6m6PTm
FRe3s0Rq/OxJmfvKVTtxHQF/I+Ze1qLgFpF9Ez22YlUovgjx6cuBJeXVZoeODlHKTu4BUD37sWp9
d/VbVq2vXfFKpcaJG09jTqytzjuxYJrOjr3CKC9VmfrbUWoWzSt2yl45LnG+/fF+3ILg7EtO3DU4
55uqPm2+Z/Qle8dJZdF1g1rDU5/p2zACB3zkB4kdvLzHMTL33yRq3ozJGLFlo9q2PBECzBz5IJWf
jHsKd2+QUf7pMFRW0LF+WgJlFwuobb6LkKzp0G2+R8TaH+3G4DRbk7NN0/GzXQ/eUaefEgN4wBzi
v/a90GqBHC9cPoG99nTkUwpHb3KAJGhPugmx9rktwRPh5sOC4E/9z0SQehlXzLDpzXAOkVOyINmw
Xg6nbREYZoXm7p5Hr+7OUJuokgOTtWFu4aoW3Wxj2j6xSkI796encXhswxX7zc6eOnuHqBH5z4BZ
T+rsIEjt31IpZ6SWtQJMCNDIhr9wC04GxGiUYmXWspht0HIABOAOZnoFDRBoKm3OaQS0c1UphA+n
KiWK3sU/64AgBSKXJGLHlveU9SJVzkYUws4OTdpEQdBWwX95zYQ/Xic5DOMtTyEqeYCcz0g4sM34
LhzFWC0DttUwpSWP35RiApfQ21+4ljHgNGfxNKSy9Y4h+oIrTunVrwhuUxgv3a/PlqqgqDbYuuvQ
RGrEW0paXkvtvKNHW16bbIEGPTXP9QzEHKHsMwWu7N1hN8h1s1VIzFlIJWuNE2CAIMk/nRF6dDUh
NqFo7lZs6vD8qbI63trS6258xzkEuZZIfMn9gKzNC5WcvlBHtFq+FRWS070ycNqe53oj+YfSlVA7
62ollf4gElsZsd8dew99tRbsHYN0vKZWSml7dXxO5RSOHW3A0AUH9+HAUTtJkw3gbCc4XCOJvx3w
oRgufSn3irCn23NZNMro0V0749EQeqN1BJgj2FCMwt0qYPnjvuurx0juIgcr0KTXyucd7zx+4bTm
Fu04nCsXR8EGNjNxSRtNv9bRtxcvym0xKNQh8rNLh/TqxEY4+P9SEW2yrOpBJbhJyAlwcksjsSFy
HFvMuTKpy4jQH1FvqJZrJpzGsriNRVHj415f+IPEtfEl2V+fAWWGfNWNGl5VnU7wBBWsNWYKwrj4
8XP6PXnYjCpuCEB+GyXlCgfUvzieH3LJypQ8Hbn1/I1dDO+JRt2imiyQhUZ3yQin6J/hAyQSptp4
4vPmALkDrY0mEXNpt638AOJ7WUASCE2IOaPSGdZVe+9tZmovUjhU0bakGFOCGSQk+2s4qcCman/+
r1MYxGusNY2AK+FgaYie6LrBWTk8K6rg8JLmWa6VTvoXgohHaBX1YeQ5XQAmFQdfciPlBkguFf+J
toKJG1Pw1rx0vNGEcZPgn1APYKw4k1Jr3CQnL/j7ke8GiRenQXeHaV6G9ZRJak8ymsjWe6CYHbKz
zzjRtC1qeX0lWf9TWHe2aok9nOlKd8oBPtZzOCHrrmVmHwObylP000sE3cNO58JJ6HwgiFbOYz0Q
vkb59NkXTnI5N2/528aKWj2VxJjgAI/wG/OkxN3dbjkXu3y/WJQ/9YNc7JLSK7EOcJDi2RzdCTsG
lgoqABEujz0MS6zaxivMaT2bzLzJR7ydLkSUDi7ooJEvHHY+BayP7mcAgQ2NV9ZNRGzLteHT74Qa
Kzv9LC4X6FzrzIPLIaGX3jRKRBa9WZBtn9zUlo+rRBdGA2XgpS+rvYNpho1glusYb+PvjbVUPZsi
W7we2MN3E/X3nbjj6woHreB1QvxHiqdxDxeref/OpQpbP7b7W95EM3h73xUVYt+AQj50Kko/dwl3
8Sk/KSIGcULQYZsJd2wXVwegbd0P53Mq6vot8Ciqe8tXq4fw6n76h2g2VPBCBajQ52zvH/Zi0aU7
lVzAcCtL1J+fXzVhsSOjTizjjSoN6mfoL9VGVde24niD2sjPXavaTiN9nAQsKUTm4vzXLF3kWN6M
zYEOBXNbmLH1m6EdP3sRDjirfxWVGSsGPFm+FiU4LYEMRtVSno0bcGJvLhy3U2eJHrHLuB7cqtnh
h6sQjZARekGAnNolfpoP5p7fpC2i4bWRNe4xJgVMRPSS/lOWXj8fZ18IA8G6ARQF6tnxHk6F/BWG
EdleBZD7OFD5ZRH0WRxLXWfK7ezRBcEtFIL2GVIghUAKxhHr4afZWypesHbEPlCu9G4Akkge1ECH
QgTVt6y6o5ZGugmqm/qXqodeRMHlEypzbmRgkSpFa0t/U96e8Et5V83NuN9whv1B2jYijOy2o3uc
ADCxULMs4efPRIfrL8HItseVk8qEwpFN41Fw8tOBvdRC87AALVyS9BhJ2T9O8L8e0metwJ46Gtuh
AUtf756gV5Mcb3/LFTr9y3ukvwQsRdkcbNGjxX2aczpSmR/4qSt5yVV9pcmtpz1vOvan41ZV927H
VEIWMy4iMdscYPzgvMytEcYOxnIBO2DaJ0WOEmA2HAM2g2LV5j5vc/Gpnd1J1hcvR0bYple1dvQm
y60GdbIkmujRzqc4kBwPeUhQiW3z4OQvga33DFPXPxcOnhcRJ7zDnhfVdCBkbgvDEk+ghzjczZDf
rIgOd9BheII7Bf1PyuLA4XMmzIDTRkjDceTXvHk20tmxJCYRVl3Zy0vRI5bMttagc1hh8PGoHLa8
MhQWqSWHNF3jqNJYwrRETK3oHFqcnmcuEr/JFCA6k0juNRvxswWPkii+LW3X5YufRbk+nL5yswdf
WIRSPzW6XO3ORwiro3eB3V1wAJkyDlUvU4mV8k/JXmc9OVEVKwpGG7lOvOscpGimPgF0NROy490M
8XQnGWEwgyuekZ628eOmNt+rYyv/0zwYEydqy0IdCw0jCyrCTm8h7emIfaBpAQjwBMMV/10Oiu02
cW1EVYAIJHKT7+roe7f20sn2EEN2tAZxmFi2yWmNYnl11m0AtH86fa9pdOTciYVfVjNrWosmE62K
1YkYXfdEbYg7vQJyf3CUM8tHWLzz+bE5m5jwrSYfLQYL26ycIf0YYG+V/dPPUS4A3qCENJ6PMZr0
Eq2rlvnF6njcXe+hjPmV1cgnvFooZjdzl0AQWTL1YUNhVyR3mvB56Y2b6Ul96M5drUzQqLd715YT
3phuFNFrXTAgPJ8O1iNWxx6K6SidpqdU/59LJTTM2UuKuFYSM4iixi/02rJUts9o30eeZF8AwQzR
txxMpmHlCi5j3Vitb9ymYeNColv7myinHUUcC+hacpdjLmD45TqpOImW8dECNAI1DXAsJ0n2KMnD
ji6B7D65uMU63l8xfFiq+lfkAfLqd2EdA0FvsMdawpffcjVuAkcX7+5/WiW6A5S2lnHPcPnRO81W
qYQnSeDwvO43TVGJP30XkUJp48vd8Oo3TscI9DrlJhe4xIrFirM8uuJco7Ci3EIcieHvwPEda7WV
uKINCk3i6pplzGckNZJ4bPnfZJQJI41XErg1IkEf3VpIMmKpPcP4QB2fPX+BBFTk3D84zKL0SGu5
yGCP+UzpuGHm9/e5r9y6JDHw+151UhmCljQGzGfNNBoYdu+nE+idIb7NFLQCgbtfmGusWNPtmBkc
QLYH/Vt0t5+G3EiSJAFfMHk9VBm6mjI5xv3mMUylFDM7Hh1UowSr9Jyzq8hTT69H7kWZxlZPxD3E
5649motgUyxdPlxgIYN+5L8LyoBq7gWxgpS1MhkY1rBQL/gUrofTSSgC6eW6IMWWw6nD6n2vWeVx
hk+wr8KYDtoP+SxmOlSAofRpEz4mVxd99Sadi4XE9JaSUpzw+Bxxirj5JaVvFqdQF44bpYhH39Wd
IW1zNmqS8HqzAcynYyMFgg31kqZHttn+FukHN0Ea3jR9v09lapffDFWm64nQdrciGjhjYEm7iJm2
XXzwfZnVtLBzd8Y4ibJx0LifDQxhWv9EeMYr2S+0g9vHPEFqD2IBv1RK1kqp+AV/oOjr3beG0w59
skI2lXiJMeXG+EGtGXep1W0VeCzZ8deFmIo6PSjqYuWu7xWkl0+9J3luoMVm0obW3RUAXYSUfiiW
22gvUzWKd/ivr/L/g94NoJaqf5HMgGwK6B5H7PUYriT7gGA6OlZRLWwA2rkkawSeWsNNHYmskpTz
e3t48Ue9efYwuVGG9J8Ses3OsVh161OR+477ExuKbKrCIaDUxyeT6/1U5F41fD6oDVOBOQs/t+iq
U++EiVKynYf9P9yg/xEBPK8tYTHkKzTeHtG6COFc/mLG2lGstNtKk6cC7I8L1OlEI1CtQNx8ydRh
MtSbkDBRP91e7caNJxIZy9mFK1ARivlfs3CIxAJTbi5RfwxVuz3wzb11d91J4eO3CpD7eqprDg1b
17yAOQ0fH5Be0j17D04OUcPEwz+O92MkwjOrfM3KQAyQ2ZRUIxvf/lS9/xCGbdI7hNhbMW4ItR2M
voou8PovxvdbxbJ2Zpnin18kN9Uk2ThOB/VwIRWNUUXrVWAw9fMmZ4Z1ztNbS2ZrOhSMsCLmiakH
UmdpMd2l7cxIzxjnkCpJiyx7tF3GdRRE5sAZg8YoBFUIIzv8/5qTje++4RZ7PAh/hVLInHlhr1mt
eKPD6eQpVlzuKVnkIou15NDSDm7iXBzoIUMA7R9qQpUMub6a60ac12l/NjxX5M6OcszncL2hiQbH
EWj3Htn+26OBLCtfYO3knbazICh+xPhiqhfMDCiKtx3DirmJaafJXhNuqPLVqqlmnCIyDHjMeGuY
Q0+EqO3fFXXw0TMXvhO0e83mq4V9Dwd0BK4ntmVGX8a2g9Oj1XWO8R+4KjtA6suXTMaWyZgCE3N8
TPJctpA/k3d3u8WpiePX82jyxvruRVebAkskrmJ6bsJXF2ZXKfcbuym+jEf+XFPABMmLTG7QxD2x
TJ3TDpNQoNh5ox0fOmECuLaaagRR44V51CrRQJ7GNDeeCQ0ibxusH20loJmqkFeluAAU4bQBdsXi
481IjhQpabHs9W73K80+QkvvevuT4gtnexT/Z4XiYbLFIeVyOf0xRdB4yOYtUwo3mQQXM0D05cEV
sLbXqHoMNwrrAWOYcqJ1mcW+iZMHqqartfGX6oRB24ElilKpT9AP/bKJBoS4jy4to/rFSvwfS+0q
FMuSr5iHwQ44Cf8GV0rPaQV2u0MOSyzvC1jKdltjuGsEzbkYauX/uizviFxBJ9L5DMBbLVkrUptU
CYK/vibCQPxnjYNrrbtFirE1fcxNHsVm0IHPwH6TnvPfTKlcheAF/PR+xrdTFTPXH0dFqFo4Sv5I
RTXDP/A+quiJCIUoZoPBJCdA50rf7C6qa1Ar+63aQv6B2Zu3jhs8h0rYUjSsPtq53ZMKvCoEdAES
Ii3bTsdn/pPJ0kkSyAcTQJfppYhvi0SkaUHU1PTZzL9RQOZMPdIiMAd9oaNZcw6sb2j5l5K+Rzov
hnDV7p03EG9Z7mbHu88Nmjg/e78ZJL/Gn/3NKiRLX5wfBLPQAXT2M1o8ivpu9Y2FglOFnppz86Up
4S+tDE/5wxfnQhAjRl57ePWGMgBCCYPFx/4C6+eG/pKBBYAJnC+9AlAPhErTJA5rqJzZe+aowQvG
malC7iYG3wrdX2MoQDPa+lWSDWf9SpjFzNEBdxpXC4BpNYcLTnzF/eON3MRu3nsFp/UOb6I7dCXo
gBv3wvOtdNWEElKF3dicT5G1nMf30ie+1bF9oBKzjQYMZb48Ya9mhbeiid3h43Tb0OT7R+6o0qgE
5P0m6l8n4cSk63Npvx7O/hKQq76bgyHWvBSVPzSqTj2lGjmSH6gdJNiekS0fIu2bftexVJhad+y1
d2buoGSg4XWfU1FhZpnp2VFT61YgM30ov52KMt40aru8A55wcQ1TJM3nX1U2bKjju6+z1YU0E6YS
i63mGiU4rtEUhJVTAbkxvmJ4H1ydm4vhOjRWt7Crjm+fVUeJRUBHa06+MD7NR/WGsSDFx7MplUil
389fVn6VMqqlFngRAsLSXmmgpXuU7rRmGAMBTrkBGPOLMJv6pSVoGuJ6y6fFL8ghv50NZz7kxAQd
Mu91vT/7nA7gXsxBje7REyia2xussZn4bysfKFdzX1GmN/WS+vEqwrzjaUt8hqWIMIr4gRUQmthb
R6zRYvtOx1YzOmDElIMPH0Ju7bYd+tfhUzv+5T+zwdxr58if/d5bkpqHpWPM9nIgjolkF4xWMecw
MZ9+5Pm33r7H/pkRkrqGx4ssAXpjWR0GZOMsM699IeWpWpOusuvmW+0ZBJpH9F51jeOHhQa4FkQ4
UIU2kQD+NmblSvfuabdiSpn3o8ghNtXDTUlQH+clnZlk1z97iz9D6kvEycsVNDaYjJKXMVZ2p4VU
4W4EU23UIGmAVKqQ2Ha5Km5WPXTCwEOPHZFDA2N1ugGrEYaj3+MbhfeB0QMlTsUxvJT77MkFzUD5
E3+bBZVJb5Qm53kwAw74tWA04367ubnNz+6Eb5eJECLKtV7VssM2FyWZWmIa8trr6J7BAf2w6fQi
VKPSBQ6sIVLfoj8fb2gjMByGUgaamUtOnrrOp5sWvnrnHHljvDpSTaBJK5CIfnf/jvF7qiUuCfnF
L5n8xFDcxCOspHf6YIYxog1yPFkFPJuiNLsCKfg7te5ZWyUP4+CjwKp5FH5yaBRY0leVCUinRWsx
pkKjr+eukqxb+03Gbf1/ij6FiNGhSozcEU9VX9baLQ/JvwbBaexm/FSOIeEBeelRHKHrW9nwVd0K
E0oa6DJcial8J6D4ExpW2Owj+UWgFSYDiw9DBedD2Sf2Ob6NhRInnRd+JAgYRVDgcIZz0fg0jahV
Kg3TdtfG8AGotJKIs6bvvUY8bbLY3FE4MmWEJWiTGqxmIXIuJFxwrSuQiAhHe5MbZa0v123fApkk
CCLFFcI27a2MI2N8ziqH7MeKnGz5pw04P5BmF7YopIWQLYYTSl3E3cYHKmeO+XhpoJXzMQKjppC6
32v+KzHg/XWjVfMLpbe2jDFEijkFuwn9mnq0uCcbnum/2IEstRdKMTevfu0F7f8pyh58KoYUx9IG
rmBQL0zwdhpbLRsg8fYiyybfg2tcl/XuDmytiCgAEWAxBloKFVAWt6Btd8jBjLxdF+1RCUec57jc
r9l1Cwe8n5EfomxK76MaGAQTBIlDevdK3Ta+y/g8d5UTGO9mHumIcg03IA14ignROEvVGI3Rnf/Y
AE068zMQASZJTC10E1jjIzSlzNKT4SXrTodYD7krNiG7L1CcXiLd0ksMTCBNUxg4hfs9xJu2W3Z0
2wa5rYxANXICKeUNAdaDLtZql78sX6BHCLo0jTy/fl/pNciCa2NUcxkjj14hIPtwHy5cK32pNrqf
8lx362Lbmdw+K5uClHfu75u+QpTCITChKkAY7e+Konx6eivib/cUju0HerH15KaP0z+Lm9+IAMhn
qWTaB7lUaWrmTlibbhbBTupCI++gbKsFXjsSa91x6kAn4nIGN6OGAp7cjxpsasDIgyGG/MlP6/LQ
5rG44I0DlAgtYx2Ak1SCHhrqV+mqOEe3lSceO2pSakh0XpmkZPgzQSiE59B/uek0lQjJjd+3L1fM
OsbnOgpX4Sh8GLdjYt0+6/pjrcD+hXEUcGmN0ervQ6w8zhK4WWyuXULjmqZ0RR+0F0sf3cp2TcYs
/2pYWY5Wxi/1YpetYCEtRhFfOfc3CM7xkke40GCGy/+dFXr7zcpvfU0hNwwShKbOHonMjrB0+oZQ
oVXiWy2B2ix5S2Kc3mvLKCETClifGUxs4jwrtv26yCi83Osn8M0yDbrXVIbkqvyXpzRPkKLJsoMR
9BmmzATiSC4MGO7fAQQjD5NDjYgtrXCapp+Ts18LQ4yedf4GW9oWFPxOwa5DwIGJPCxMpZW6F0qk
rBZlXnTd5v9MiywUxuxf6V6oGLxRzvzjVr8HXHvjXoSbPGkgnbzJYaYJqC49d+38Tq5+4wcbc0tY
yKU56NYhjp6d2TZHYYZjVav4aesuYVdRJ5b02hcvPPo37pPEE79NZL9Oi9RXSp59o+I4MhLE/Sft
/92smmX06UyoWodO/KKDgNRwlbcVfmclVJfnO5g838XIwBSOW/+sV4yTFqyU/j9FHcf4zh5Y1ifA
zfMZ9TBgPp8qX5GbC4v1cEcHYwwR9EssiVRyf39Ymlyg8hlBvSRXfhdymC/ZsAPZDzoQbcWVclqQ
vbAUsbUOS3AWHIHvWmrZoJ9jUOE41bCjUW9JRktVvo9XUAUlnhpO2A03IZwRJiuObdBHiytXEPw3
lsI31xQYATKSOlh1ydesFJ+ZjsaRYfnOmTp9II8lHwIFEYYix28GAZsX+XEKr85ecy32g+bAcRWt
CK/EiO1O48csSDQ6BzIvP7MqRo7MPRhlR6XtLpj2xu9uDDnYVUUaDV27AGV02Th6CpGM7NcizjRP
+uqA57w7FPGSBmT2WmWQDvfCpcEdjanNwhNnQE/+XD5wRff5N3qui8l9cHqALpMwYxX0fngb4yfi
FPO1iucTeVLBnfuuOQTanlxqVpkLybPxnLU0bhnFKI6Q0d4KDkc6HepoHQR4kB9LlOszwP1bg+8E
QRNmw26szdpUsIDp1QW8ErVX/y14orXRUUBY5/3LxGkBOdiJmP/bC5kIADYuwaz2Ug5CI0rQSirn
Zg1vWSvhcQFSkdLvHSi9DpHIPB9xw7bAozstpv5cmcHZBkK2gvzUScwvSEDQYAq00bLbJrJQ8KQU
eFJVuFlAA4eM3/SNKEIoi7l+59PaIeTsZfg/Ppl2sKKCArdhgghvt0DbLGY2oe5SI7rn/wy2LNr0
Xb3Do2nPQY8VQ7oJVBdgWEIv2ZWK5fXAp9I7XrTJBk1YMneXu9Xa+hFLHO4+lDP9JENo+35NhOL2
o9OCqLs7FU3aMEBtO1ZLXNWcyaYAxIO/FwHSFsVI+UZqKMp6GnByPhRTIoyfJ8Vhm7xmvg4SZ2rY
83bOPI47dT4ukqULYe5LwmvZWGj8nKQ3l8Wj8qFR4wp2qm4zzaRBsaNSJer9zY6ZuNS4sc75tCSl
Iqxz9WO5bQ5+XqzzleNaU83sYsuGtqFt3lz1xNk++94NzW644a/bxl4HtKCM1/CJ4hMofAZe8MAa
AO/VsYHn1Vn0xeEnJ8vQDhfnUYYpW0b7dfzPODUGOtJC7cQYYZnUeZ047/rVXXw3yue4fP3hzgiO
Vn2MFiknPHg3WzO0dophFnNt9MUU2ID9DGnZPHIwqjf6dQqDi1mqZ25c4RrdS/kMEQ/ID/nxVLUg
7Fqh/4GBvlC4dYMYmXTM3kJldwhaqiCGo6s8lBu5J2lZlNZ5UvLPiFfCu8+3GT8ASzCXyWD/x1v4
9O+32im9p3F7r+A2zwn84/mCqLI9YK6MDrnSGrQgTATEwStx+p5bOnWlYSYaXQ7S7/S6Zo/myvY4
RX59Px90AYRvMfBsh2AA7cR7cm0dQxFTSKCCYoBQ43u9d+lcGZK9bA4XWmW6QFmdhkoA/2vBRaO7
7tB45Bb7Tqe4VUWU/GzIK2AjgXGFJEPLVIUL98WyBqpapwYJT6Kh9vJy9bJC0BtNwRsTlvODYyDm
wvP+3PqX3ea8Yzs2z5Tin80b2JRfROJ23WEeaSwbRl543yfbQZhGqvejqA0pY2TKCL76uabxw7Th
CFq7vrz7LlTp+Q/KdxZlhMQTQ9VE1/25Eazi54U9hPHx2Z+63ZTzFoxp3rB0i4otwLiAAEgYP5jC
k6UkFBRmYvZYCcaYPdewA7k/3b3RXeqU/KcWcqpaUvCaWiDBdL3k7zhqw0z8DQxSM//dzJalrZ8M
bDyCIcLovKEADzhBP4X+GzP2D3IZdyYggKPEyqclSGJJDTRTpbfgUNTMMmyEJygjcZVBWuoSa/MY
bkVBWPKUAdLSpX/LIk3Fz8tjoX79WGm0TAaeJov0gOfzW/rMxjB12H9eWT3ld2QjYwVr6zjBAnbd
vyjAKaDyZSsnBCvL4G1msmAOPw8OnNKk/mFiYYIp9UiJCffb1c6tarJ25wihGCNKDxn5SZ9xAE3d
mxBYAPBWmqbKDUyOKbS2sMWMm0oI1uBdRwBob44WCAnNYAQ7jOjz95TmjY+YB2Zti8rdK4J2sx9s
GDtwuSre34DTa020ebOXFzDD8KLBEPRuJTa3AkVj0t7/m4qxsx421ZfO1ZjTC/fVhfL6RnKcIEUT
0shaOF53y0ImbiNlCxC0mwavbwpujUh0NrHOA5zlujbY5yF+p+4mV89CkyWah/aqjPVkQmjGDuKM
7PBrcR0jiGf9IZ1371hxeg3lgpgL9krnm3fxHAyEUahFLBVBNfG8phfeTBuAjsjkMPOuh1QMGF0c
FgPtoSujqdweKZhhiV0PXYuvWKL5L7CH20M5afTrgOjFIvcqeAOjhYvRwgblMblniEQ2J8TTg0SY
koYWLiFGbBRLOrgAZYTtVo2KsTktTfL34HWARVYMejwoZ/S8wciTW/GYFunuDCRf6vO3R05NQcxE
BoP1ELzNm1Fgmr1BrP/7sq8lsINjIm+6zNLh8CWXQRWxB3GWXZbN+cjqXSHH10wi9MlI1jeuRaIY
D9ebwIjvaxS75BjBfNAZm96Nbl5Rnx2B8dzzwg4IzuNFKbA6VtQhAR7vu5TcC4Ft1dwP5FLScVFb
i45RjGYQEKAfTCbtLUpAYH/cH2+c1+43eN4kOOm6LHYDb2Pl14N80YGDbQxw0rDG8YL1BOF+QKH6
A4INiIveDS7jyuvOAKk9uKp3hAjJ2H+MykINFuGP9nrHlN2aq9m+53QDSElBVZ7H/2OUFC9Kj6yg
yDl9u7AiXPCgSbr4L3Qh+s9lLFP6EsjuMETWsgTKcypvRkXjyZfIL5iMZEHXDFPJkgZieQ+sIlAo
mCoBNtnARLsNPxBl+PErfXRHJY5fGtbSRBgRvlDc0jEY42xg+BYAi+N+KLU6rIe4pL04rSLIw6f7
ysEUMGNn1ER0+H6FUtfMiwOWJmRG7KrEyC8ayFSJqvK/ClTy06om06wgd/sm3ekgejbVr8U2i7gB
2TDJZB3z1qtuagZtOGgSTYZ8PWqE4im2mqGf2Wja7o5fbl/pEHWMPBZrF1L1dP2vybORh/1zaJSf
84dIrw0OtR+IXOyRVlnDmP4ewfMKD/u6GrWSZDSzJDOus0RL698haViaeJPo8mXOwowc2GjTIF4e
EBs2w6dLPJMemLdeSlhpnFLQwuylSZaXSvQDsAynCvYrDzRLtqJKKNJlV+Lftq44DdHKIV+MqBgo
aiGnBpe4Zh/Fd69dohG/E2A4Qt/HHuGPGrA34qvD2etGKTQfKYU6LXNBz52G5mKC9iA19buMrLKL
1kPXUoK8OwJ2tpJcvjP+DFdvg6mHTvdP2Clq2/x/P1vganxATnREvgh9P6IPI4VgGcou6WdTkztP
82pDTLrVFg7LNttDHHp+qz0FCzcCo3kjVdXX5Yo+oDnLSyegwOFOCYzpanVAfFw7VUCed+2Ym+5J
OPPyJd6oB6VwgQYJgnberJMYA/7uosCvkA3zmFlTkgFuGG85GC2r/YDg301zblcGdfNv79X9FkMx
KOeBMz1lfwYScpLoIgYKMy/KlLWJ/JK+m2bR3UPm9bvZivv3T7WlgF2Z0YEw8uleNZMwbzsnMpuI
LPcPVrmxI9QGgJOTiHB2kPLcn3xMJpn4K8KTh8JOOsaLuOcNnthByvgKrHPUuF5JnAWKTiOfrVcL
P0GsTQWR9dPRnPiMou5Pyd1I7KN8iG2627U5k8OKUC1BOqUY1Jbz42wMnsCIl45UqHYSaWupJ8G0
ks58pUz1UZOVxO/cXChOPEnvTseOqqtBKva2Fn3MzKVlDGdRlGeklW8PQhvO1YuSK9U0iMEBAiwW
ehSM5WfjEmolLxaP+p8RayiWaZ3xmU10+lD5xFoqse3wT8xUjTl1F1hX+NGNCgzGXc/iS2xHZpSI
PD4NMhTAlKl77oZeWGsn5JuI9i6CclNdMoh5jFZZQEdtAjpcOXX8uGK075bNTiKJOSN6kbAO3o51
4fO8BeRGlgAZ/Lh6LOKp/6FgrQmd2zCTLIHvc7VDXZ57QjnMDI8PSlSKOFdAxp8RTE/EGMnoIMvK
qgYmHiPtnDM4VccRpPXmeqef0kk7Kj3awE8Z4dtPif/9hXqDnJ6kRAofUecj78G+ZntIaPJuqFTF
v1T31tlbTMh0GIlml0heDF9tNGG27cFpkq9LnAqjLBtQPJWDcaLN2WBqABueg1E47SqFNk5UlgG+
KVLokNfsw1xwfoyAeXj3DYckzCuaOldwlzICpnwGxZUzs1YlI6K5vGKwPDQFyhzTx+4u0FJP+y43
n5HHCNgAmcWD5gMd575dN9ROS/xZljcp/3FAXWxtj3pGgHYHdwj4FELm0eUCnrBuJAQMr3M8ccPy
8pmQaVyXiesmjsI/yqNxTsFIVyzceNE4mDCFqqJFvlCxcwWpsaGB/gXelFcJsr7FNlSIJNm6bJe7
Lzlmqh7EUfnaezt2wyYiPG1or8TAeN0vi8aDTYPyxGyH+qRcSfHirb/SHoXwW883gdDSl2TN5jCy
GmQYTeZmeQ+xGbkyVIeAhzHyBxsjkJyTcp5Yfgm1h27fzVPY7oqjXpLj4FJkVFwopT1Yo/T5FUs/
e+kdAwCKOj/01A2anq6pwHXrnuUkVg4o3i7KvX9bRc+AkPhpndN8oH94gD5NAkDRnM24pPg4xoDx
C9T+kfzvf6VUIkHeVInFzlUmya4mfCdU/e8LKjNH9JlWmnkYLS7yQ3WQoJHe37x6Ek+DnkD51XeK
fuGYQzi8AWWtl+JFjL1+/ayNHaqZcr6JPlUIZPGxB50uk/GHNjwj1NTB3LD1gOBq4qNgtBJEmUag
DK4ym/xx7n70BCj/p0+fNbTdeAWfvmCsG4zYXNIcXzUQ5cJ651mtIA/h7vsRbLGuLPyWFZXwTYd+
t4QN3evaahg7+NhfqR7hYyUfLhQWm1rvg6/IrLwvAHn1DKD6S2BABIQeFKRRKiZT3prJNWIQSYk4
lVH1uCCNmnHo5ThS5G+c4g/5yKHpS4u1Y9YoT5+InqI9in9sn3iCayFBUXHme/BI1kDk0XDKR3Md
fVvDdbEEXe/B8bE7LwkiCVdgjqMRgL0Oe0scV6am5kjgVy4wOnaMgjbgbRJNLN/Ys5vz7aXSOEW+
mBlu/COyKpOa1XZ7uJe1GXFOInHKxxFEE/Jcp+JggOASe3V4wujsldJpjSCg/8VOCExWk3kIrjWz
tmi0CMoimL5tJBfIBdooBA998aAKJgxoWWDDjcy3n186jDkt4F0Cv5gPxh/+wH+r/KUaJcepntFM
NzTi6CxR3TlNm3pgzjD7J9jcZ0GjyYzPAPOPlWl00caEsKrL2N10KsWvHUdIkP9bJbl+r+boqf8f
Sy47L7sRRJWuObcWZ5nemsccpeLKxUPrQq3Buui3bBiCjPFHpZvjm8Kode74u5Pu7Iuxw7J9D7U2
izAgiGO0zhpkYMM5y9s0TeQrIA31pV3dOyBiCFIpdyOljB4h2WfrGuaPJXYdNMMdfMPT0vEo7kaU
wR8IDkfw01Z/dMELgDLoRcS27nC180jS9j9r5BC+t6ovzGkT2JMzaWFCRr+C1IgkgeEbgjPwvcyQ
byCbojS0zbkILjXzL9owFpNyWvUCno0JVVGJCyxnDh7jln4vdpTSDOvMN6HwePpY4lnSHkxzfpbr
F9abyoTOWk2FFz5gfyiB7db4M7cRZyFxvrjFe9Bb1aGZ2hQ2nD41e68n2r0VAipSPRnQ5PfOHdFC
bUyEONMW3/kSWIWNfF2SUYCmIQZ4aiXbQ+nRURP61ChqiQYknAjWdZR75E07Uo07OF/S03M1oe3y
GqcXTkXRMFBeOz7fvUTJvMac6YV++h+/kLxL4mcxzYWty/Aeq+jspqkKhr17iM/MG3BoLJiN+AzT
KFm3+N3ZSUrUQzT6TGIlkm8K+tVaZyGGlnABSeQz9WeFxQjVgAvLt4SZhjDJddZf8q71dlp/LeAS
tWd+ynAs/+dfQv9JSpcDuMMkCxvam3hlZIRSFm53unrMEezqGeIfjfDxdckZKj8DtGbVRRgShI4v
9lxGpKvXBJmyRGgATsx4aR21cQERP6hpKUeaALj8gwkxx8TxVZXqQbGpQBqfieZIO5SOT7U4nTwg
KbRqnwvVBk9DvxgHGXxdWgyA2oadstY1rQLbPPWNGt0i7+U0x3fvce4PjrBXklFjBV/7D0s8kIkW
FFniFj1m36wjKfgCDydce73WhxFJxKOwNcWh59SCdy+g3rGWr26UjgDIGG2h1MtVBffiZrnJ4up4
ByfxjkDBJxs84J+hAmNodqssz8daM0ct7X10h57VzMbJ6JCe+xXrrHZAHIVTMrYnKb/1I/mB2Vps
c6h2fIhqB3bnPokl8D7vKHYy2Seslyo49rSSWXOJxliPZB/zi2U/7wOcqHkgUe9Rr7ek5W/1C8m4
kuE8iQoasY4uQk1DtBprGqsdKNtRPfLNGfa/BI5Ub9BlY4vaA3XElju/qNO/tmo2RTTUznuwtf1R
JPs/Kgp2WaPnr1daU7NSEwDV7FSsNOzuR6zr0UFE9NS1XL9CjH8/CZnF5AgJdaui5LRT9uZMsFID
sUYbRanuQTBkATD8fqHT3dTmMc/v7Pde+iBGNVROhfiCmbPTRUItDZCv8tlkQ3pbyBEPCntegDIY
CNj/556Z9d/YBUHLXqfm9A1G575XWUqYWkqmmJ14k0JAKDCGQYOC8W7A6MW9qvpC7OyLVXN7BLbC
5hJ4OfI2as90CZI4r2x/HdbBnvECOquV1aGmi4ujXtziR3vzHFoRne2O6plVXaM1DPXimKUPUHjH
Ia9OisHMdXCICzZ1IvXEFtBoBdHkjLrg2V6GraW5Hb218lkDqtKiiglDgKPHBaz9Z3P0Auycd+WA
cMkAr7s0eh7/HjitCdeCfRREw58f+BOTPKvEECtKpFGkA/RceIid1+N5vIAmilSViRwK3BNAQEwm
Y+6bVrJbC0NNziKk4JysZp4UyoMBNDs4ZSFmYAQzTtPBgOD1cW5edtMm1CwOcM5azoy5zSjpG4Oe
GKrqMe9NYHGafNkwfVDlFhm92dY77aCCcpvopvhcQZf8b9uThZwpWmqtG7kzKW63r7OvG1xj3QAp
+B5/04YB7R8/TA7lrEs5681XSEPF084+GHD1dbUJ2CFg6eFfQFCMfSNsktuvyJ486xxes+WYmVJp
qL0PG8yaj9vgoyH0z28J07gz20FYFnjPIv1jm9vUi6tPsfNd6zpk0ZNbF24/TXiYtudKCJILJFss
l2CHfjvmAIog1KKq6nI632iLS+jTQ8IPpa9ftifmTPcJxFEwll+XqRdE0Q83J0H+bXMphRf3yrDZ
koUJDZeF9ZnzfOiL6hB4rlQ+3yDvqmhmP1DvpA2EU7JBqqAcHMCzCpA7Q8F8PtyX9TZWO3YgcbA/
4fncFZqj2MJbTlLAgfSyh5S3mIiFhfZknYWT/w/lOjXYoWhR00Y0+4eE+IYA9zjAWwZi0IJQlPB9
M3yUFm8m31ITsSrJfzUYFCxePwxDfpSfnzDhz652EA4K5M89TMZIpOmyju2xbQp82JxHUeN2DuO6
z3z82QvZIJhLQVAEg7scp5sTRgobk/GxhCk1A8Sc4WO9f1WVvy5SwrY1RUkUATPPAd1bX16NIDWF
ovpOsjtysDAugS+nsY0X4SD/y3o0CqUz294wCbCYPKAy2UbqPHq0FzTEgRa1/bsRCi+H3oRhyOAb
r6zD3aXoKpa90lHdBOVOpRF/Z8eJ2xmhWVRgA19OlWE5MPSrp9dGTvT5ApI7E/ERPY6CCPszgsk/
M5c7UYjCXkf2xmOuDtwxYlJCwPmAYIcWdQVMgzLCdreRkOP+C91M1my/HoWnGUQqG0LiSMt2858i
MGiLJQZ6f6HQNPPTPlijvOnmUbR+fSAwIe4REFyKzMGfHlr5ftR5gDBSnN6uJBR4Gf5MbfeeTrHR
fmFsl1UcGM2zAPCxDJlVzOeEi/7BKKV5U5qEg1F2/Sg1e32/L171rRrFC0OkC8JMfnK7KBrbhqYC
L4PxgUCRNuDqbgz5Kt3NfBMwQ2gDMeogwTSupOBZo1UekffwCWh0BHemypV71/9ew3WVfNzJswg2
gg2S4d7lt02fxk3r1eXvV1K+OZwNxHW1bypeZ2LmEuZrQ5BQm2ZZ+1OJRKQbRQj2uCVQokNPc5DV
pE6XzR8+z9zUuy59argMI8mAdupKXqPFbITTQYDRjO3P2LHwlkK8upKKdvdjlf3sMn172zAAutWj
yYayKGTk2jAJsalkXfljLpfT7hgoFJQDBIyNLhPQ1NWSfQECaZ7Uc2E6GM7+cnu4StIRonuPmyaR
KHhOHShCoRpi3JzAjM4Fzc/uKOZLYB65W1NHXFyAjViTTTrLlr/aRmlxi29wh7HwvsWJkS0Uj7E5
dDW18dnQP1YhZk8rdaomrlwKmZJ3Kxpo752NvL9jYyEEEA5R/uWrwSQtklB5kt0BABu98TeQN0e+
z6TbqL7bPsG0qjjk7zu2QwuNCPOi9MjA6baGD4fg8xHFIhUf/H7n6/uHn28xA1g5a+ad3XiO3a2O
1p2nXlxcTm0UCd+JTq8j9xGgwuTWmkq/iy8OX40cQs+QUzs2Q/gEmDqGH7SdXkCBDuUYqCbTPygF
BtAjsSSwugbY905vwYokSQ0mQ7pGh6jPF61ZIST2vpDUzUEoj5SPA9RzO/FNmTRQPcS8A4IUxoPZ
OQ5yc3CIneKQYWxBRkfqx8wLo55gpLjcej5Ym5xHdtZSCU4ELh58ImYJYyLeYTRyHQRxNfarFjFr
wUoP2HfOEBnFKSYDu+NdsVVziCwgzPE0sV/YOJhswmhBJpnW2kwodwJmldHp5M/lXcQx6b6SZRYn
/FCjCp1lHIEP3GA3ttVlMS5mGKC+KvkOc2RupkgwR/RB4qpo8/1keBugSQt2VIxGWgZXirQORatJ
MMWgW3CCxaGrcYXfjLQr85i9weFXyF79S9QI+K+ZEzM71bwGqR0jMWq7O9bOXbw4ODF76PFZGfMp
Hf7+XbcB1gzk5OJPsX73bp9mAHGugfKQM4AsI7r78Yl6AO38m0P2N/1ZBZlawRlVZgeiKR+d53Mj
XvogF1Fm2VKaZF2dk1xZOXheR7Phqa3fYiHdgxRBx3HLxos88aedMdPXCRFpfdN7YF9mGYGoa4E1
Kv8kGGo85UYUF5rO3EbCuPjxc521QKk1dRkEASMOFd57QVW2kKAHgvn1nOxtsLn1ajqhOPupcvmH
sUPPhkMPa5TAH6VIv2najh+6PbwSOIZBICQIrH4FhcRcAVSk/dcAUZDAbivp8g1TWGMmAARhhQ/m
L7Yw5sVulA+vO9HfuH14atrofBGr2qy5+eQSFx272WxWc17RI5qavU3Dg4Jj8r7gWEnkJ+7LpXeO
+T2F5ZZl4x6tvOPKS1c41V31NQij0ZfkC4YL2bNJJGsR8b74fW6P7BcmbF8nvIAkPB/lfRACeMdM
6axxFBr4Zvj7XHNkye5P8jeb6B6rd2Ji3Ocpk0XcFiDij2P4uJz0OjvaPWTU+x2oCtTETjOmQSeK
I1xX5X44CiAgvKgRefxcXt7F9kXt6pzYy3N9i1GpqYkcdFRCEYUIiBpVTSrhhOgtm5ULT62Bd/wZ
zL8EKBlkk3QUTdb6KnUh9tEWTJ+OxySRLKBTD6YfM/uoekqSyrvj5HPIigBChFpbA2dPJ7Y7gnct
3EX/RzmgMzW1ACh2pZI5ON36SEJoiM5Aw5FVh5bqii1az2wTdq3YF4sURajmSPCiUOS8FrRmBtfh
+W5MU840C5sy+1vyFfF6P8jZ7+SrQZogvEnr0bEF5GjEWjz0TkfRNVZtL1sxch5eutbuRmGJmw3n
VqiHopLzjREAl8XvgjP7yQDpPgh2TBhrcQ6hwYdCtbXk+eQUrQmoSnh0Y5UFPsnq4QGXy2j8O7gc
38ar5oGSLo2d2y3K690rzFcK71gxaX8AXMyobK/q9mxC6F120Npvffa9g5w3LRO8j2sH+ZFFBqu3
3btqQiZF+NM4K7BgUIb35o8U7oVj7MhH8otJRtQSdRhPHGpDUoDDhY/xTNNEaCEA00PyosNPnziu
8E/LFS8BdPyFUhSy8p4CsxqaV7NzKP7ahVF93F36FhnHWHlscAUS160eZllRNCzO/BMG26buWzP+
BXrwu3sXywkMP/o6r7OCq5nUaWWvqwog8VTKLz67bDqOl2AegDd9CU07CNWdlfMNuRJnHR+y8LPr
EYt0R4oWrclMW3L5cQIJKgEY61hSlYgRAJOUgGKxJn/JQzlRu+IG46Q46BI/bhjkjjv6IAogI67A
c3yVzPWxILKZnS0b9ywwmpVb9QFumo9DninLy1ZY7iuxHaATPLVfIzzMyew7N/6ODojA65DrVZbz
yomkeO5yzCqAq6Q/SRv4xtl0MEesdlsKhHVPzWtcqkZtmINJAOuZ23iRe2drwednXzr9KHYftTdK
wEMUuU706gWoZ0WNV5pd3wI6St9gi9LYeRG5EFy13eY3Sq/HCcpQNcM6jUpjScB7cnHxybU1I0Vg
Awzsm0a/fXKriJFJxUfJ+Q9N3iEJjpiSVnK4dATkdZjD3bh8wQZ7+X6mmz9E5Ia34YfmWFft6qw6
H6hMz+BUw2ErauUg1DgRYmJ8nqpQXONvQ2Q49z7IJW4/OwS/MUUiPdn3tihB5+aBwQgwhfACK8nN
Oxhil1BBSwNBgh2zLEpK9djm2R7VsYRRb6RyHj1QJ1Q5cphvhLSJDJlh2ZjrQtRMovZefH3UzAOg
M08eQZMFIYWateSAPE7FCOhmx0g1OPa9+Z8Bz/d7STsJgfITKpD1hTHxd8/DcUvYNCanOZ7eblOY
kH8n97A1RGFCX8BzczQ2POlYa7ZMuOyMowOp/52zS2KBOARFasu3Jy7pwKctp8ceJkf3v9EOTOz1
IPlVGjR9mVT9GUzVwu4LtGzMKZPX9WjBdXrNY3+rhR+rpAbxzc6sKCTaoxZz8FCVtYoLIcehlMSS
w/LDac0w5tqlFUz4DvpWqxVNz5MBmofDdJL8AjzWBjj9chUaHnw9QFDJwiepnrZBsYpOIT1+wc5W
vC8sUBhXxY5IiODVvvPUlJ9tAVLUwIOin8VPk06EfDfLdGncOzenb16mu4Dgfs7zQlzB1cFUiUuD
wjVZgJKG7YB3/xyB8fD/KcoLIEk9s+qt0nksJSq0tchcIpWR+QDBRMUx/oPTSeaKQD8M6UZNctYb
rI9ZIfvNWdPYITPn23INJBzLv+nLLuw/10w68stS69XQhrMxR000K7NXKM00nEscPKPY/Aze3OwO
T1KN1LcYhx0fP72IKYg27VBpYWXepDgbrKLM/Rb4d5ih1qvii7vpQ1nKIoEnI1icFLhDTgLmvprn
RtensSA6mJh+oT+1c4wX1tdac7wjMLXObjaJiKvl4ESt1z36ucf+NtegtR5rsJI1akKwJjT3P/WK
5iOM1DfDeJF5B7cRxAXLdH1lnCANWtaeTlYWV5aYvXoOzDfSFOGCmGZ4Rwbh5CdjLEF0xodc80Nj
jR3kpQJRzHlljRWFfko9QAbD2ib4q2oKSEW0B9kmUy5jHQm4mteWwdBgAgAOE6czE+yj4NqVevbt
Iscc3U2dgb4oGZvxf0JABuc8UWivuGnz227DuObB50U1bm9ep3Gmadb9I515ia0F0l/Asj6LcYnc
HIMjjTfTLhC0nBa1Ha2Js4910xd3NDZgDUDMNPQh5JlezceDGqnili9RyQZkN6bb6PuK1x/yZfXO
maxdZg1Bdnw5oboIrfgfvnWtEA1kiwtlEaWaE097umPShVH7CY0i8rpbv4PiRBzR4Et/Ur6U4GY7
prVdSShD155LkeA7ezD5qRIYz7QczdcVRXqRIM2seR2iDwyviBDS41r2ydj3tAc8wVReuDt8pJxh
S2rXza+EHU7S2BzhwsGrIwnEXQ3bVGRy+6Cy/zB0RaBKZwe+fXsh/dk6eVslXiquIx9HvaZUsj17
FLhhnsunVcwURhGRgoJvKCmsq5GWOIUPeppHP3V/yCPvV1OoOYL4nRKCoDhqkpJKbOxYvz1tSpsd
LC+PkWY0hdSyMzVBdAJKqDVzUbP1BkYsKy1z7/yWUqr22BpNb5VXViqUFF5z5PDy0nt6s9hcWUTK
XzppSA536P/nU2GHvsmomtOT3pQu8LmxtDI12nqwJnzvE8jin/wmz+KJkz+A/B5/IENVbL28IP02
gUjwbFOXkeyMrH3Llw5/2S7SnqdxNkxosig2ZInh9k9vdOYJC4PrO3gmDAHg0nEbnjEyao6Bs970
O6d1U2bc3C/pYTjk5OM7lM9jh9aXMFFdq+u+KY00oJ7HThjp+i5ED0LWAgy7vVBnogiaHGmiAGXS
VW71XVt60MTENRS4yZ87WKTpNZT9J15Pwdqxu7EKGJAgoj1BVUivvRN297d9kGQ1uCpT+ASzTF9t
oiRUFrq60ZwvSLToNL5RdEitrcvAViZ49BJoT7+mwH9HGhSm4qtnxM+78zuuhyoaBa7gBr5dodNe
AZTLW54tTODHuRUQXSrbrwjH5Mb0HQUjWcnGKdYo/E6ZtFG5nkRr2498zwWrUIUeyTtExDkPJdUX
jwaIPiTK1YA2D2FaxSdhoJCGT9CsEWW2OmlFcIFEYmmA2entJuvt5z2WWKcxV9N3Nd6e9PtJOnys
2q2gCL4tQUwlL4GrO++TDnM2z3LVjzUvqdNgpqev90AO49B0wtn1NfGG4/BjaBvb1u+XtMvMYkMr
8iP0+bNJ0bO7FHZ9sVKNQb4iMvhmN7SJDJuorOTjKhHrJ/U1XltmHUJ2g0N7OHLX49J8sNeqmpGZ
2We9EdKB30xt9zDdJwHEDWQx/P4iN6aiRG7ECKQ05GuDlltgfnDp+AvyqibTEK6WaTDlp4yb4n+0
WRD21A4bDkYWr+ErRMC/z7EYVyNynek2HjURDOjdKDph1sOtQqC60rhy+AVD25iiKXHJyejgM5mO
VXjJjtpuYsuHoYfZWPPL8VF0L+oaJvZsQh4xebap2zYR2ZX1UzEbgOKzbLmuAyIpTXCQm09OFugN
0AeNyjIHf/cTz+BIZ2/GDWV+z8Z0TBRW93GBcxI2BZfmM6b3wj6JhrX1J5p82/qEJTlrKX4ZtpwN
Dow0WONCsNrUW440IiBprU6/Pa8Cd2SpXKHvwk3Zo42RDfe9oG10JsXD38/3hzRLFpDZcgJl1mDh
km9XfQksax2/qpv2MBDw5dLYgV5wtbSXuKN9u+xojbXBbjvu6+8UUFbGA75BA3WlWVa7HVIG16p/
WSmoms5R1CWIk2rSRea7avGx+6IR2quRtPs0H+UcCQN0gIRkh2fZtShmgO8KnS8RWfEequay/f1L
wa3n07d8rb3cimvez06HRg3Q/+ihg3CKId1yRfdn/RRUorCjQ9OliA/iLLmm9Ozxf587PVbMKkf4
Fp2GjTfj9ekS0hBtS94cXfZ9CMtfc3Md1qZa/gATFs+1FcQhG2LwtVbTh6oQJTsiZ6y+oYdic4wR
e0aYYJuwHGWU0OInXxZyqn9Y/yKUt7YnezAEzAhIOqEIPm0lo3LeWNsRlzJxn2qNpunlVfEHB+1w
NA6LCblWVZ/lBVca3ZziFiEp1X449ftNNWTmnAqS9yK+PVBOibTN25huIeDtl0ASkKPTZQnJNKOd
yMc+C023wBmMXRhv9MR9/LqXJ/3iKvZMpzPYUP+FTe/yyUBxxw5pSkWpRpjWX7rZXHuoq/A9ZVQA
ymECBl0+qmFnhm5MRt4U8T9Xq9fe3X5lga2OUiJI+9iQpiP15BVZ0okwDIVTq5EhCX3z+c1rOLuM
871LUE9Cr0rScGQjdTRD5ORO2ZRiaHnXmIGuJmQj/iYz4Y7Jw9q4PrYllNfZFuHroDI3f8SOELcX
1TTBziCpxbtbEOxgwmAQYWzbT7wHBwCiPdE608VI6WCitvLVqBPVydVoHTFjioP8viVv8+PBV6+j
iohfmXixyUJIvW+Q86HhpwOZv3VWgpcxofcUT/Dz/Wq2AJnxtN+3BFfqeaTZG1iq8qUcbW/+zqg5
y1HhTnhMoSLfftohZ3nVEDDbcIyiXV/zSYNU2V/ibV7lMlKVAClQGBuvXoj99qYFZkqabVfO20xZ
xQv9SbTEHQSgnT1u4CoSh+LuhQjpYDrdr3YUimXZIyJDqo5E7qnplFosMAzFchjn890HfyRChSDP
IZ118xdiE3jx1sRu0ZCDkcGGe1w4Ln3glVTsbIOQU88avk10fBtK/g1KBzZeO4WLPFP9C+plgbZk
DpFzuS8vkZoIip+2evPXjL8p7hb0f/fs4qzGNzU7lLPnnYXhP15tjVM+TSO/9IczD/Usv4rVDCN/
jYFvCCmiNaI6sywSsxv74aUgqkWYKXEYkEXYq4ENMxbxcs/aEmlmudgdPUq81fkNukoKkXt7Z92i
KEFDRiZG0QQHCZGW9IZwlipfJxWzSZEIHv/Ce1KJXMa9fffQvWECnGdkCmzmcjmESyUK0OIOTXhZ
8k7ipc0RGuLrfFJQ+9o6DOAUBw4JKketT2HNgVfD9/NqV4NVUvUEFd+NCb+NzAqgYGOJj2InhlIu
ejzGqTuxnO9K9d3RQO2uXa9T3F6kEhWkgTKu/HL+1Vr+ptHqFp296adS07avT8Jw0jaroMavskBF
rmvork1YhmabVz60KkeD+F8RQG28yt8KkEaLiyp694xZ1w3uKEaA+3yhAUiRP10hpsO/HBE5dz7K
NTYoqENn2emorG/XyaM3x/vbpIzy+SWN+ImQUNjt+L/PAwijRa90G9DrDY3Twrq8yyms1ik1VQuX
n3ryq9Ji+zv2ipoOGdL24CZQdrSdgHK3aEhr4XHtnsKahwTUy1l1B19ZMLpsGz11/zyyF4DVcsgC
5x7EWCeBpFCFDmnIoXRM0enn4UqJ5vwhxrNKzdQfeXAX3yrPqXmoH1N7k//oEGpTBGF78oPfVebw
0hQXgqWa/nTjJTrjc+L63XCGs25mekfmayK+ZRauZzhWHhje+igLFpRI1tLneN0x/E+HdROa4C4t
ZV/6zmNby93EnDQ43Xrm7okcn7xM8HCcYgqtfbr1UJAyTpN9rurwPpb45bl+6b+O63fqYmaJOqGG
ABRfB1Im8eyjL6a/u7nXfn3fS5B/1QNSbQAO8zAiH3PKvesV9DNp+FteuwymRpvbec1E+kgignlA
KXVLZJWZ3t7qPu3KjZfIatF3dZMMRVDjTseioK2NKJOy8T+0gYvW7ny7TeUecl049sJ5qZeEgHqN
e/LZDpuMMSjrXrmM5qPA73J34Q3fEYB7e+hvX2NuAqrr4IInTg6lylcU6guJFtSPiEXaqdwykuXQ
k/DgQobwui0BjI+34KZg83GpZ3gTX2WSSpU2uLy1+2RNvX876tMaf7XDleB+fAENjr4BcyK0IvMM
oirUFoVMcf6KUhVvQGlY4aKtMEiIoKqSzK4J5exaUfOr86te7R2BSDPwpZYLLZg2dGl9ndJ7hhAm
sPfhPg6z6sGrhztR+yQFxivYzu8kNfGjUcZVCW2leMSdvvXlvm1/IvfCkP9qfVuakV4q0N5XOgh+
h5Y4i26Xy3U6tSYhdtW6Syl/gRKo6q9BmMFElmlHoXWWKEoDMZzZqBy5fjcooWlXbrvdOvvzMNDA
FNZuIj7Ue4rA+ktIqX2V/rFDd4lzimYV2zCAQqDGST/SYFRvS5TCyGkhybNjg3e3m4VxdKBpss4F
N8cdoQewQXPMxLiXgB/ExerVj0RAUfAHuELfrKTHwXxcf7bZwCjnqfO61wgxpfOqWzUlk7QgD+hL
3cmzqiWRe/JCQ+HmE3yyOnymG8Q12IyslsRgpLjHGmpx0pnrsBHcUP+HZKxq4okjDbJBt+2zCD9Q
0gSfQggIPg6ggdD7Woni3fotOr1E1zpB7JzWI5+FxAqhSEsdfMQxhdv6zjNZeyxC7qo/mFCxyZVO
U21RO2xI+24LESUiIo1y+Fe1t5ucjurYEOJeCfyTVf+gpeJdWr25gt0Dndjz5Wz4d+0a5jww6YRg
e0qM6nY6QYx1gZVnCRrE0yvDoYq61tyrUFMVUfJ1zd04Hw3ydyXe7QnGLoOOzngZQzpM/NkqmhI/
ihY2Ag4MGalngboYaMQIPLDyaWdCqSHmhkQQY2sZyDetuZNTKxyunYNIjY5Ig51J8LPjDwJY0S9A
5gYv/p/giz8piaOUziRcwni0LVZB9Vl9ELKS6qyWByIchbsPdIQ9yXkY5jjLycFLlLdq0Xpmf3FI
IHLcCz+GkbAxQGbG0phzv1riogCBXTa3wfCnEtJZg6l85owgMVVTPMXsHXzbiniClAM4DAfOdlA1
RLg+aESN1t/oRSDmqsu7zkMu7/bkfFTNzPAmQyX9lq8dXa6NfIP3y+E9LqGC1kTy0qxGWtEUC1/8
V3sviipR9SWW5QY7wuvQKqwwaUk65a+mwKr8EljK+Ijhw4D2BHcnVjn2SUbAhU+xTyBvYsG7ADTl
esHxuYnRHqkMxNjjOUKnIDhngFo7JXdzyIgh3IWIfLVoESmRMkCHf69rDsejHCarBi6KlDsOqk8c
DpfcqPLuUz671fB9JX1si/ZKTZbZS5NZ5t8MGbqH2h7Rzviyt33nV/sfH1T8ZTZFIokXDPmGOUCi
DVhnQTlGLxfc3ciDiJORF9uaDUk3dmXZMn6RMVpkEf9+wxufuFe05cqhV55Bx3/mHYnYvUbW7fBN
ycaZiT4DxbuRv3y5tSFfEnS1hwYJSvgt4fEWSnqef7MDkDnPWWTIasuz/enSfSTXeeVvBCnsTf5x
bITRJ0ODGnxHvNvRakEN1WA4stLjgB80SycHvvuQvBU1Rj3jv46b6kgsI/vuIJ4eQU5fR2eUuheE
SPWm/u6UxEiQlCjc68r4u5BSVAYyNDX5zZEj0036wyiS8uN2kxi6nnzizNyT1I5lSPxBNfk1AZ9m
bCcsOSWZ4C9eluABaAu4VbYS7Awe5iRCmmNqwOQlxfHoEwDpGNj7JySyVVKxIVf81QQD7XxkyMmS
g8C3qWLVH0S2bqCKw9iTsF/kZg9INuxx1lp1m3uT6adWo+0r5hRrTXsOqsT3+NpHJNVny6FmlSvM
yurx2TMsfwtEjhJH8QDBkku7UnXw+s7DVSXrlEIFe2W16jIH0c8q7QI1unJUV1PKEdMldD64jw7S
pzinIWhKIlQoZGUwE9c8dVL3SKcPTsMmhbgxn5aWYRs/TE0td4HpzCR2KJ9Hdf8Lzf+7BOyPq+AV
6Mbn4jfqYMqeh7Yu0DxdTRBhbZbn2l5Aod+M7f8znt3w+obf+GxUC9obexNKgDabSGRGUUFkj0bq
R4JZ1HPWt8O5g1NYJfPWkfmp6N0tKP21MC7Ns7E2h/md/U/dLcMdguC41AMmgxRSmzKLi75OyJYn
MlUfbwWWdV2yCFls8QhsxujVPUNe2QzZvmoo1MUoiI67ohIqEstXhNDFPjgstja4NE89+t1W4KZm
R7bqhyeNFGBJXRZBYEDfHsvzHEDbNmKCEIBnXNzo+MUS07tmCgKqV8aorXNDdzUnB1vP7d+mYcC7
/sU6hiAEtIWDHgxbOmnHlYrT0eAvhyBxxGGkWGG2I03eDYoK90uT5+i7tc9+RTZC5PX31NCdZh4j
20obFdi5m5oFJapw7VZ1aL+46qmN1JowE8aCClsrH5RvO7pUFDOHbCe/eTisqNAA/+lTLfMQT59G
nk3oxrHZ6PjF7X+6OGWqC7vuKMIS4BrAOQxV5a6Inyk8ON1LWvjPSu8kMBGKuKyqDmgeIJ656grq
PkrSOLjLYQ8gxLOFSYHxWvqFrsAe+f/hG4Fn4PiPBhAW7rM6dJ1yOUDesUEcEhVwtnaw5isj31KY
8t0Qe7Dy5He2Nt4mwBWSEZQ40FAybCOsG1JWcirGhUq7knnaqdGPoUKMtFT/gGoqtqigvSsPub8A
NDtZe90G8lQaxSkR6W6xKMGckrkA076EH2RpenXIrw+fGJCuSUThZrwfeWggfP9LmdI35J3ZZNK2
HrVkWr8QsIFd7k8yc7uhaTDxngZPNGGXKyJakIAuP6anxTUZ+j1MEzfkAB6OGwXDZW+60p6G3L3N
DYwttju4i16Q4Lrhx5pFJ9AxgjFDq1gCb06oPAs6MX/xn1sc2t0Op4vBjKRJqU9re55xsc7tv/VD
dJXXDhFD/tL00gtv9IiGiiPK+IOey8362ulams4bQmOG0rmlt8BHfZf6PvJfIQvjiEzWJSyqmxPY
J05/YwTisKgAEoOeQklqASzft0YfHdwTapjuL+IXn0kuhq1u6COc2M/M+EdgWBZOaZ03XSYnObHu
CUyCOMs7SWZ3vlKxoAfSHDvj58WJZFLBfz0mIIrjlaOH6RxFniOtyhgUigLiZoD/2ERZgZIc9lTz
DAdUco78zIODB+bpuXXJRkBimZIa/QcMhQ4qiy20taWHUWvM5WcYY6AKAZTtQ84a2NQHzCGCQJLZ
DMrrzpAOYs0kpiYYkwuufe6OeY6fT3SVIHs8T8IK3oyRgzkzLQQt6z2FAIJRJGB2adrHPUPbvxDW
9QWLIBotoQQ0M4uBdy/E2M05oLcXjtPukIUSBsyqp4NognQ0sEBDeuoTcH4bz6f7tbj4mPwImpJf
ayIoU8E8H+Y112baa1VmF2qAYzTC4qZgo9ohQCvruToy47hxbX0zzSjm9dgBbCDABCCcaoDNukbj
4Yj67PhpdJnoIGiGxjmYMuTUrICLD0+FCtEW/mJXd7+Vj8GRHByYqRPoXWBejpKwqldSQBwXfI7c
FNXPzdd+GXT2TdxsTl6y+7XNR6Uts3pJfwn8l9rnPUWUrPcIXMUWJNPRkNy0GjhTiCK6l6ukWYiX
ebEPMTf5oFeOgC3yI0sU1K1jn699lHXP2OAeKKuipAvjbXm8/ejygN/cN8Q3Re0G42Q5oEZZo6Fu
hSAfZWNYQbziweCWZEumFSjOw8a96rvr9bcklhuHu81WOR7dS19OTKVn+1bIrXyOo2qGPAsI0lz5
KdmQgnbopbTeYQJ9HuZjRR+yK5GfzmT5reOUC1RPAPvVDozrHcbR0fNmSh5+6k90ZmchMxNF6Tdp
vQYpKyUMOVQhiS9wJK7DhluuozJTb81OVqCFQggQ/VSjBnUr5IH+L8JT9SmVUdel8251Nk3eVcZj
ayl5o0RPFoWQuT5tMNdUR4C6e8VRCL0kRBBNCX/1vS8ZUbLN+8PmrjQH526PEtZZ0fcuirFD6F+2
sKJIuKa9zBg2s8fp0+ZbNPTk37ELn3nFRQUTXM2WpvHAPLI+da1zOOVGZsqsE2UuY+YQvdUlDij4
2S4ymvfWT7TTnpafhQ60Bbf0cO53kJGD8kDUACksGrKU2WFe86+mWWeZ4x7C7wUhghTDG5BNRsVa
Sf+kLhuXf2864f3S9GE91VQYj4mC7E98rzYIAlF3YTJM8D+2FJiXQ0hMhO4MeIryPa9G0CamfP1X
NbOKs9JZYFO6QN3uYQdPmwDtMOni2tMjBRxjnzwauKJzVL6IbtS2t7Sc/olAiZ2XZmZ454eHLa1Q
+q2C8MVkk66IBMqOhW74h6wyJtoIuxRu2WtYnvPG4SbGvWgEogAduYLfMt8lDSb3sRugVLKm+B0i
xkRJG/rsLG6FKWhKCiTs2F7jtdAnp2NLNOgp8HcND6vOGNnc4yDx5TdQ/fxDw+K1qiwR8Z4AHJkt
rNT0aXeIBL2ti/9vEOvkXNNwecWglulNCrBAdpucRf6Z9U2IPvccFLljKSTRMf994Sb3HqXFNTOy
sW6UaiG/Hv36Lnzi0ArXK7BhBRWSKLBhnyIbp4b6ZXzxs/8BW3tjXDPu2HNItQ0Zb/n/4CPxRsSl
yBB/3nIEjqgC6Hsol3Kt0SeAmfiCQJjtmf6a0O/LoZGAmZgc4hWpz0Pg7IWLVBWTC87N17Gm+rVU
L31Q2SQVpmnXcsC+sK24xzFR/6i2DUSfzQHC7l2fcAXQ8KMImXKuQpvZb4y69hn5xzxycaB8pDuy
df9uuii4KDe1iUthKMITkYo+ivtnh9wUdu7BjgSS0XSQv+9nQG3wTF6kP5Qfk81ZXEGr8t4YtV9S
8P8ORmEl1SiUJfSM4aQdNqCUlUNluzhAxeeTrPIMKT/4JggRGyxGclxCkTvONOIG8EAhEnOUmL/6
mZ3yCWFYFLIVxAxPBegKX3IBZhTCSkgle6iMef4+CLV9ibdalnrxbedTVtOMQX0yKC0qv70to7FT
kr/2SaEgxYqbppvi37b9pi4RbJcqsbl9cf3eS3sl7k7s5yiv5dkGdkKG32FDiGoT1nTmyxl6n43s
/iAop1FBR01tNT73S91WK0FrOkO5pcufirBcV2FEZbtG1Xm/1uaMF+ykuOejqV2z04Vc3ojhQ2ke
Okxwg4CaK1mCPYL2DdtLRPwgvzwGE5aarDRTYS3A8nl29Gd3H+z7RXHY6j7br+xJqLup9szcro7c
18kwsse8+IOyDr881Nod5jD4SgFNFzqxbBumyBhJIgAuIo/5mYfrSkPEoO6Q4nD9pYaUOls9GaMM
M+TsaI9PJ2lgXDo2+TGn4HV+WNwuyt3HkVbZckfAIDaxShKpV58/SJC+Z9k095kztOMJIHIwaCTK
vDh/v0A2xku/b1mAGpUaq+MD4hbwYCthQ3WKJT42KLweskAhdlyvzQuKbB+njNt0nUztodKrtppj
Bf2IpMvoixx7O2+Khc9gKVuuYRmNXk+yFVnHGbs5YpSPjuzDBR67tLzqQpz5ZaYjMOF8W8fNUCbs
GjT/MMV9LU+m4VnWmqMQkUm7Q8VtXC4IKLMJ02Tu4HjizpckJDDU3B9f9y/2HUzSoYwpJf5Xx569
bL1lZP/z1umM77PpV+mEwg7k9zhv0u+NTxAAH5RpRq4sJ6ebOqPLgyUR48k+1r4+yh8RsheOMhwN
pDINayee88V5XtuEsA5CZjhAuuq4mnQjyOIZKJBN7+xHoDtP+uAuqHyfUjM8vmWBOD+E+oNrrdGs
OXf4G6bsBf//eSxLS7bttyk1cOxebDvMdcQRUjbra0AamESYaFM1DxhiayMGJ50IxkCvIkJCGmWX
JFfgxB0t0ufWuCrSL/KsgYkcIhYhsZNxv7/eZsUKeth9jNifuU+cg3ICXBhjjzuDq+Gn/IYUXcQW
Vz8hUsHsiUitpUPP5nrUU6scLitCexd6qX3D+8s+Kq0Yi6pcPASL0sDXeVZoGpPd0D4dbMSX2fRy
/CSobKTzF8iiqyPjJz9HoQJTl+0EngaJRoS1ORFsQCcHnspop0LkWfNu0ZwXSUha+b1ZlDLvG8vL
j/AJkjpv4wT/qjfUvaL/yHR+8OkzWyaTLAcSjQUScJJ2aUvcFW6xNz964xrZSU+k1ZD2O6TrXtQ3
KCswo663p+E65NHaupbDBRz+PTd0O16SddhyMz+2gbqDhipeDPGbSYjbUN9GNpfTLzUamc5+TvSP
t+AVU1yd+1rRLqRQUMtj+V2RUBnqjldd4USZo9fiPJHJVPhXIybuD0tw6a/P0c0qnAQVuNNYdtr7
efO/6a12NTqnRWccqnD8LJc/sYkOZVkIsEfVjAUY3Z2CoCL1MKxBCyT4vJaoAM5uPA+95opVOU+j
RKyMulDHF/YFA2+wByU+Vvb8BsDr/mS7Sv+Y4zB0ivHglFjU9U8ziBnnblDSiz/o9BjBgVOOx+PD
piSGZFNbL+4XtbT+t18IdfosvkAqZzd1yZqigdyPbgVBMX89ZnczyvC4DG/5KlbDYuOGIgAWRb8F
LrXT1qeUqHwXO1gdrJYrUuOT5NRcJbBnQKTRsX2ldmpLDg1oi0wrs6GWH0XXqcPkVIE6UjKy26pM
eZH7KcdJr+X1lnbO9y4PXxjoX5/QpMepW26WToHM4+/8ahGRwBc1DGWFhrQmMyB1uoosifkPMXld
8Y2uPfVVTd2CIYhLgIAVOguUsc9wq3Ood0oqLRfsDcUrA+llL8mG8ZAvW8GOQaw5f7aYdxWaJ+y/
on1e9xpJlmIg13N+qNahgZN0RXOvABPwr7wjRGbn2JfwgFVmRd/pEfymxMWkYXbRuHy9g0eBjWuo
LjQPrNoU+kS0UNttAsIk/PKQElxo36a6I/UypJO4OctXPs5mE2Z5G1lYdQ1u6EFHTSxh3Y6e1DA4
v7Wqx+sJbsQDQFAPu2TuIt4pwtmKEgewVYFHnoYWDQHIyISqq1VqWsUpQc3rV43ySWhVASkcM9Pg
wpK56/8fb0GQEIZqmg4nfjdx4/3r8Ex6lki9qIwfyTB3BoGHqtuDWtciuMHvxjsn2fImQd7Vv8yn
RpRx0/FVMMGoaxcS9WNq705b8vqjFNSeCwegxvs8eFuBENsXt9/8hDAIdZfUvZ42A7jVxz60g6/H
GNFx3QseD1aPEUKXFqWNjJv4cAJ4+XOj0mWNSRBAexxoigFnFVhjMZWPKwjumpi4zCC/yvuLg+yS
2wbp+FhrBWmvzyH5sRX8+4fmlzQ9JXyw4YvLv0kfAR4CR/KcFBmWd5gNQDA8hF7mu7cVMDAzNLVZ
18Bs/dYV4ZA/CoAi1P8pE2h6JMCiP/Bt7DCaXJ7dv+Sc71zqQxmZwyNWnB9yZeHn+KNfcjD9bt3Z
v8/9q2rSpz+2dXqQpr/wgRsdxbWU9tLK+k+tcDL8vliLntLZ1yIss64OlD92fnOVgDa8T8VHxysv
HKzfQfdJ9jH86aiEampxKvxeYWwc99mVXejQAtNsr+MoArObUhz4SnvRsMYHAy8G4yljoONbegO9
Q55Oio1MmU/lLEy5RMOv0VykHuoL4v5oeFD3QlpK3HdrMuGxPs3io6IRC0Swq3xDYT+e5ESEHBO0
WN0BE0m7lfFgnLIAv2hXLbCwQiSLDWcUAkBdrSl/LNIAdr4bqu9BM0ncZFLTZzYL/YQI4A3FUTp7
mdSA4MMHUNoGT0S0epx9LnTKTTzB1OaZJVcBRli7J9ed9xp4vyGyj887uY1BFDlgj7fpfbcSq99K
TAB3VQv7OExtjJL784Y87krOhnOCyLnKh6pGkwRb09zTv6XMmEnJrr8Ix8QDyhursObDgAGYXFke
4bNbo0WQJa6/I0VsNuhT6pAeBXgwHopR2jZCnK3vEa4xA839rej0SUEAqmTwCgjnhZ965MnmHvMP
EeTgbGu2uf81k09lQWXc1xanwLBT45bUZ1RYXL22XfTMlfDIHqbnnrhB7fNXYQ3VCXP6/YkxPgne
1HezMo3wK4vA0hwJNrCj0y++hwPv2HN9Y1pvDj0MxznnhCCdDN/V7NyqBdeEWwY8O6FODoKi9yYE
MKWIWJaNgyoEFW/YSQEYOFeL15H6TqfwZsmqYkw/x0p/P1BlbJ2g5DHNmem98sYmWguvoVb7hwLo
Rd9ZrXfu/SpVSTjLuX1LYsVa5XK+C+K3XcXQhSnOcrfJ5MFJLP7UwE0Smf8hpLeyQurAZigOVJaJ
Ilzt0LYRJJvPP03vaSimZfeqp0UaEA/7G2R6vuGTy3DykeXbrf2XBi11d4J3DvSOTSg/3fsBNY1K
ZCI0QEnXzAeVUHMbqJYs7tJazpj9sVlOLogl34bhhdZOyLGwN44Lq1s7nbWPmrnUK0LAWUsmKbu0
7hfj4TODrrqW2yZs2dfTY4mUCAMu/wix+KWX0Lj0tWdnGp3CqVqGiexdIzeMU/6cRhLBkXy7rWnI
xkNZ0DxMlizgy5ZSbIFrbZFQHmG7I4NPvec7vRBFK/odXxjJ5Ioy+Pk4U3+9Nl9gtxcUdijEC/1W
ojiPbcbAyi6PfMF311pNyiGN4iqsIxe4Yv/TTDdVuY2APpSSHDD8bSxlFQrFnrs546VmvloKHPtf
5IQ9opIbOcVaQu58A6muZvVKGvhRuiVwPskG+1gITN6KpV2JcAkURdTktps73LrmbhbRfZe1h/Qo
vDWXR4KeCmhUSl77mgbjq4G+LTtZD/X1+XDn1DS4KlLX9FkpbZl8NRX/r+tenePToCpVar+x9CBn
5fweou59TDYziA4iA7RdGF2dHG5mA6+oeJDKaoHchIwiX9aRlI8zXgEm3+J2ANhtZZ7l0degIeIn
0u81vgKIVn8iqiqbsGZSSsTgSzy6OW0Ex5VXJi3C6gNh0fPbCrm8zKCM0vhQVtKd7LJixvd0EFJP
FXpG2VpHnqc/3LQNMsjV4WghvNY4qDhiNCpzpRqgmecfdtqd22YCyCCuXDC7xMKBTjEUzxO15S/s
GL5x6V0E3Nv/ZJqLVK33AaX9fEcpWLBPAwAN7Jh8yDd5VnGG7HFbcPY04NPKOBCvQ0FUXxXtT1Yf
8IO0AGRw86NTIfucX0ib7GsiS2qw3EZID3Qpuy5nVuu0ikXfHxslqG+JDB21Q4p7s5ojvic43q5l
T+R823JPS/IuWFcbYjJdD6UDldBBElF2d4ckyVDs8ZqFDzxB/NbzdkEWGTsCOdOYD7xK78NgRXZL
GJ7ESEhCn0YyMbBvaqc0bhJyLnp2mEfHL+4nIIZA/hzkhJnqAqptgYrjKrPyPLxcrY8t4Gn0BIkO
ogAgdUzZ4U+oDw/omFAprtbOKjRVORn+CbndSGsCZ68PlnHpR3c6ycu+Q/9xrhaORwTiMlVjYO2t
UZgO+AehzYnPRU4J0fpI2amZS/tTe5pncMnxZYiIQRGJsCk4t5jlx6m1b6QwTEVCZMTrNvQgbdF/
vLphmoVNGUlijuMvZLX8icMwtMJw7vzesmLbce1GX0iHdUMDhSXot4yLOkuxoG94H1Ai92fWptd+
iIvXEMlBOY3ht59zZt/U0e2XYzViYA4wKuKIVccR+84LcremmNlOHtLdPAUJB2a+cEauOYJevqJI
OQNTg4+0ehtQa2hf6V/84YsCFtnymvTg9Syd9CnjBC71uiswsqqVp8v8TtdwxYJb1l7j6F+o4sj/
gm2L52rtdUwKJEiITZ/tdqraoDpoJEThqPk0SPKgIonbw6wUCJVhCAT++t2fY437zbUrBLqqq8lk
eSeTz+hrUYIt8JxFM75qR0WwNX6GC1PXYgxgNPO8D4ff7MjF/Ww9yxo7PagND2DlIAfWbHT0OIlk
E2076clCZFQ7Eu55WkFf5akPYh6WhdWZiJBIqTL0y07wrZGtz2w6UwRNowI8oCeumfpPXUNmyX90
A748tB2gNrgj3oAmZT3cTs59zJUCHwtXrPmSxn8kZE5+nu6/fPUD06MRv9gxyYuJVybAVisRe4Tl
HyeNG9XV8i8HNdf20O5hjmIKrIs/abtyfWrwWJGwzV1KUiKYfmf4ug44zxNbCofW/1Gv3ehAqlpa
XNTf0PiVqdWyDBB1p6YdTN+JdMGLFP4feCmzYIejCAMn3uI4ZVeuQ6dxuTgTCds54FfcCO1tgzDu
BxjH34oTeXfyX7iSCYphspfh3h8NLA9ycKhjH5+KtxWT8PJJwQJTVSF3XQIReZZIZcEy2ko3ZAKT
W3xCXOUrFgf6MoX5k26vaHn5xPfT3GD+PRZEiYC6aA1WVMIGvOsMa56PXk6KcI/KmgLK/eT/EhVB
IYbkdwdzPDKpr0FhcKpVXq/pbW3i5atoE08o+hwkR2REQdM1s5Lhb9mlbaXrGfDLCQ6YMSx23hRU
Lev8yCUSiPbD8HAe0eWePju3QOHkv62g7M1t9PBnu9oIN/7DzRiS+2JtBeEH8yob34pZAEbLlXJp
3pGiC4KG0rzCC47jxF3QO8LZbQaA12SXSide91g92kz+9UzhNlhT3f0hUqTXbGdZztE24B09fDR2
l2MM9MJmMFD2AJtSp4wt27uaRPxDqX5uw9p8lEPgHxM/SWv1FrzpLdl2Efu7XjtKSQVbw9UcIhSl
YSvflMK5Fa859NPoTaUGvBhx+I39zscbBI2WfQPdrsILEs3iHQHvJ5bSzQ2XvoXJB6ZrznPLSRKD
KpXL6mz5ESN4i5op21eJEbIj73BMoeq+PD7/iEVkkfgBJdUfujtbMujxooDU67M59iA5hqFOs6mf
ULKZdGRUm70/x5es4fae3MVbEhDM+NZWprOoZh5ASHByI1fj6IRd3rOyb+f7JYPuXCyapcsxuf+/
P197z+yiuAcdB6h3ZxWISiQFcylnVPvQW8eDAGQSrl5DSJPwIJg4MRgoRN6BQEiY1hl+Ob6Drl5J
a0LVj0PJqpxJvUK9o+gMvWt2fU7CXv66XgCtBELKWUeg/krbtFbApl1ldVGFvEqL42esNkPuJFTv
4hzwA9YNvMpEfmNnZ5BRsT9LkERIaA0hieTooVHxqCYLEJICWTT92ZW+Cjr2zPuhrFhY8gsDhmRH
+jb/3ziQnrTvnhdRJNNDlOypMctKjF2IweHtUg055CslCG334QxrwNvrZ5BA0XAuvCYMckpfv8be
FaAvr4jSDK8eTJooULptUuCj2oZViKbNmsmGkI3n8BuwlkidJyW94IzQvhOFMzeT5VC9HxlFfMyR
ANE9gQXezUIToV/6BgYSoXCSuJbCuIBgaqs8a5MnF9TSG4SYOPWr4B2oPXd5S1RVimoxHqWzfXi9
aqIwQwdBPE4N3CLZSzhOMU9Vn3KAwCqqoI2dnIoqP5gv1H8ASHmDqJolpSI2djFj1nAl5DzLB2ik
1oV3TbyXeP/3TEWP9nmOSja+3RFgGpoEf16pwrKf7xNerWLabLN1lkmMEBpjVi2XDNj8xxV2w13E
9jIeyUVbSu6YDcdI/yR+hFYYFAu4XS/vbW+DudkoT/7lupt2XrvQeuge1qMMFlF2PLMPbb1/GlK9
WFecpfVVzBvQFtBwv7uIEVl4EwkM4Py2OlRSY3aRnR8MPJIcb5ezkGzRGtGxD7GP14EyMaAcmQj/
zRrVFFrJRlW0PpAMWSdu9m5fIcClwX85po5CtYZIGtnlFjl3STUoqY5JZ84Fy1b+7VPbUL8qFYsG
XxVRsWjbi/FwSrNdNteCiUFCIP1ypr/hPQ1PaOecu9+s30e8cxN+mLZAVf2EGNQcYmsQhypHs9jg
tn6NoLmF7+DsLb/ceQRchaXZ/5X2mJVACrNbOK7MEWZ2AymL3fYz5CJwj2O5E+ACFOtHCCofhICt
8ZVlva4q9TsrIeULrLP4OLEHvYF03MTqDKBnCcGKqb2NREnfqfFnct3UPMj9FoQwh71tsNWPNaXf
MJ6y1XOcjwG++OZiIFcZnYh6MZPDFpufp6X6HmahunQek6WJhCOL1PQA6uaQgLxu8YT/lbEB0k8F
x9xpkpHkAvH1w1C8tN6NkDq9cUka5qw/HCCyKiiQG7N3XHNeUppNICsmRqrZs0txynQ3m+wMQ+qq
608ELgDUUrlcqqvhVoCIB6g6GrMuD0wuouHJqOLzaF8L/SnSTTvRaDzPpkpTYPsEVjXRdRuPUCUA
6CE0bqUjNTUaNkflmJNVF/L6xkd6ELJAo+NxSO9rkNPzsmHLkdDJOYEw06HZiUGfGZbeP7s3vjZh
N1oBZvjJBsAYl/Ct3F8ILmEzAGG1/4J/hjXBmVZQZayKKrJhtqYjSx6VfTgu6m30GZw3s9ULkYQV
YnDwMLWbbFd8xGR4whKU8khk37yUFiJKUmoU3q78TqrjS0+AA05MBOlIbEoL/7CcWcxg5ExG3kF5
aikOdv+ilt70fjylmjww7nM4AbvsAxLXRGKLvi7+D6cXUrKyc2LzMHRXQYRryT4S4QNSSimkO8eR
VQnrQ/Gn7FhG+8cRvXjnhF0xmzeAF0GGYvmo6+L7qMRFiy510svCHTLyW9Pio9A3b8vjAxDCFRk2
/xi8fSk9wClxpxHAdb7cdlvGA+bq6w7GkKsrIe0e11K/oNA0I0035cwq8jlSxmGoZSEjXWrYZBca
F13KCTIjEREhoxIeR0vclUOiPdelYMY9wUJ1HuCLc9w7oysafISNdRlp/lqdN0UElZhgZ/gCEpll
N7yGim7cJIQ5E6JI08eP3v9jQbumeuWscRba8HnhKzsDPA0C14CbYkbnjeAzWsnhVuxIl0BJH+CW
2DYL2Ih9NSar1N8/LI+KBjqt+0t1wwf+81GG2wvMpaZuaUZp123UMtQrym52D0IfIMVqYX4stfk0
bnCbcrMvDn/cvpz7urr8S1kBYEBvMfZDBskAS3Yf+2ucKG45NHqUwN6nRXQ/tXyAucdGyxgocmx5
1NIqsaPFbqnMXa49NgR9vGS3HfYYFSSTfcctkJgE+Fnl/7tpNIzCe5n6apiGcnXf6q62CaAXy+Kg
aol8UeLQP/thpdi93JNzc+k2edrw7i+5bLh3p3/gBS/t0rhIF+oGlVkHjo+c22j3ORPbHRP2FJos
ysVmwlhgQbXTx/hjh3uqXDLLFGLKQU26S61zy1IvdpGrbUWOKXzsdylPvytSk+Y6orft8N51YyFh
YaLttxyiBhoanyW1w7FjNMBq/qhR/+UxOvYwOUBhaiCHUACiyLtxTyTXr4SO+B7xvZNNVUQJU/r/
vEsrwK9vk1sdq+fHoZT4zo/2/GV6dHSy2neItnFr3Fu+F7QB7xn3CAOQDp4/OYaJ/TIN/JaHslIk
LlNgOtroMfkLsxtt5TGiPVxNiR1rYH9X7/qCZZsANIhbTcC+SX7AxwVuOymDNMGMxFsCdlTvtdg5
WaINciKAUutQTNCmosocP5X+HSNWa8fhxnYSdCmPVcKjW0/E8Pun+ytP+yIzDW+83WczTcXICqap
lJorrCPRnQOwe+7fbbJL1+38zlWP5Z279cEFVHBQRQaNejXCy99k8SCfxDd+kTnyQiwbf6OykUEx
mr3otZi0iMdRcRcHhYkVRSZQADjc07yc+GlK/d6CUQa2lzoPmbK7JMUkimEiY6fXqSqS+o/yiMA9
ma6RcvDtuZAYO4VZ9+zj7WQqkInDmJ2q6JljIAr7++aK+kkI3+CZ31axXBdqLkHH48Yc282w6YSO
zSSaOAZ4tIdAitZ9y1aoRfiSqpcSJPXH1rQhOV22KBShzQc6JGUJ6sjzxAO0OytIHFKLvu0+zSc4
2N124CYK1DIdNIi2EakCDqUDvo33fZKE9oMDAm3fNpvlp0Gl+ooZifcd5NlHUobHVpx59rU2xFIW
uBF+Aw1h37HnXb2rrwZfMU8i5Vmnx8VrDEgYw/yVEdBsQBh40wEZYzL0uXzTfFYkGX0YX3QvlFtP
RXC4Rp9CzZAIBEKBji5AKNwiwfiEwOOBF2j7vD7ESV04Row4F1b7K6Fd02V1Mf4+EFSV1gb3oBmd
BCmpI9OkrkIY6B8mU1x1lfAxKDLl+DHOVHewclbMfjVQq8f0x7P29cZGUY/ozhM3GYyzY3QwIF92
LxAnshYOZeplzZ7Y8aF/26aBjF1Mcmcxzh5DVR1d3j6AcXSD7eWv+Ynw7HZkK+Ti2Zsl7axDAary
bZtQE3+u4Ydgb5dNQeZ/PXm1cpLfJRLUbbz/nDlMkLGwzqgQkQ60RbYS9mh+8Xz644pPIDkfPT0L
2cwJFV34eKJenYSTLoDEH0q/mQSY1fxTfC+N9tGtBkenKOAT9gFKJzXTf833fFvlC197dqGChVV0
Upts/YnCJIhbI0UBi+KoGFzBvLPiQpJASdYRg/LbcXvUgMR3oOKYMx9QVQQYvr63wgT5rRPgpXqe
xT75X2FrVsnSSoF1Nj2XbXiRle7Q1ggV4DDpNlapSMzNeLBewrS3KBzX/e1AbYoSBXoy86y3bF0I
dMVHrAQX2nwD79T8a0KhlGhjHNyJivXc2dRyxtuiTOdYFKkOHFVxBZGMIp5i1d/ns1YrLTFNL583
ncHCSSkTdVSMnANQE1uE+2eRYFGd9NGVoYyrimxFhDUYTWMFOcUpxnSRmooUL2RvBfTiRs8YWS+7
hfJqWYIhnHud9PfwXLogo6aT7q7+Qd69CX2OcmFHm17XMvvk0kYpL1IF8ZxlqgeeE4fei97r05Dg
i6GvHZv4yvhHiDZH4GB5Y62ka68FRsuk0ANjlqk0t88iZNpd+xFWT3wctGiQd5wb+YqXDK2oyrN0
xjD76JPIFVe1qbxfzcTx4xWcJm0wUNzSfNNAqRDdgtpT92lthRGHbqOzcIsVWzPc8jbwk8qT1RvW
5tDOeqYZfkl2AIb9R32ELJjyEw0Jqq3/oCrFMB3tidWd/gF73TAx7PhX/AIu1nhzhaa9syoI9N8I
RQnjWEzBg4J9Kq9mJMYHwBJTjQghSIEmgdOAkA62Gv/IcunOj/Kh3W7mqP0+rGNMJPAEDFbkN0Lj
TwtB6bucKXextltCX11DF2VkIxzrV7TYn1L/HSbj8ICtP5XTJzs/7X0BCThxx3pUOCKh/RFbZYKw
iagZLDm2g7gGnZeQmzRU3KBSSN3Pmw0Hm2qf83MrHvgofGIzyGgTfFvIuJXrr7kHiuQ9bqnCFDRx
EfN2OJYuXyuA9PxNiLX7+g47tLue1gnCiFfa9+1Q2h292jIdc8osE3AkPUHMxdIHkzQN79blAKby
65YxUNOAmKJ9tswyfD/hM4zQpxF7rLF9eMzl3cRGIqw4S7QCB1r8oanoPYMuUsdq+I2dcciOmjm/
re6BrZRH1hEQQzvaKqSUV7wHIMGM9wukgXvYzzzmiBGbHlCCAoJpawj0t9tLNnB6VztC/Kys72vw
4Tiu28QrIjZnA2j6y6m9YFh6ecuRogM0d5DRi7ohrae5IFA2BsuGdgiCDEjEL7HZBQ1lmBf8mOED
YCqh8rLM0Xrpa+4KxinXCeCl67IfrJJTIcKSdW8I1OqAWnidRcm1G+aDdV3sX/zpaWvWXh7g54Wp
z49vAGvh7pH9/qzMkR03x+31JbALaX64T4rB4LveiRzpMdPvv2zM0hNZ4Gy3HpEqjiy8HsyLj+2V
BesIT1nRs7qaIZ1IsA9zIg7orbgdAEq+Vm3DqRu5sg4Q2JWGdfzBu190BBgd62abcdcp/YdLwrPg
0Knvn0VYdVSSWpqz/r8NM6odMzEBeedOOWCjL3F3WflfV9zDXazRm49bQB6kDVAA8LPNvy28iq9T
knbjiCK2PrOXI8wpeQzm0nFrmuFcNBg/M1AAIUsSGtYw7MLSIMlZ1QeKuIa+4AYa0YAY0WW3oeFb
CZ+pxiSAiEK9XcgdVVC62AxdQG6+0ZafOUzisiWqjC1iEQiwfRfJFm/DsEBiewbfiCcW3do6GDJs
SoahPj5ZdED1SNCySIcdYTp1Vb7G/TY0S9DHAHOo5/A9te0X0lm8awDguwslz5S9hV2QTWmN/Q5a
pUDW3b1wArcFa4PwJpCaVsP3D+iF6JF2FyUw/7gSvoHI5XQuhlcPG8p5gpToz3/fWV4aVzXBLOcK
yJyhevhYrOa2jzXWtcX5zk5t6tA/og/gar+BEBeKxtqS5lu83hA98/RVpUGQ2AFXFoD0PK0Ywm10
xSf453eMU/J3jXk1VOEvUczmmwG4gTIaEREpW7+7wRFEaGcQqC/UbpwSRF1MKmg/RNtgYg6TZ41G
rNUDZi1maN2slJ/PXjXbh4L132TaxHIlDlv3bJRNfw5iOdFI1l+AI6rSRV2wH0odsRolcv80qlbK
agEyHLPiKWmkAMeK7k7TzGCnPL1CeNY1ug4yTnlNaQoW556W6N+TnBafFgboHIXQ65WwovW1yJUB
6IDlkZat5kUfAKjmAmbF4Fvjt2B4THolCB7QaJkQ9lz75/2YjxzcvDVwyN9OX9pvU5lpHLotEPpU
XM9/u/aafD1XrVQ1+YRvGTsqV84kuoT4HPY/SdLB92BT6qf24m/zHT0rI83YIGdWgMHYUWTc+5wN
cTkiNYP2D85N8WFNJNZtXFl+rhlzLIVwgTPQC5jA1yzT10Fqkb/hICn0IOkwMhZ2HEVWA42SmxZi
h49rxhFFz5vFquQ18IlyHcH1u7/oy7AEThEwzrcgHLeRgV3RsHyomCBtzts9rd+lP62HTauPoInG
TT4iSr7SZfAwKRrMaeVP9SdWcQYr9LC8im1MuBGsZQerxSUreXzvALi9p47k9u9NyMxdT2sK4AVD
IRqCj6y7FIoys+OMkDJBsACCmpgm5dktDeR34qmhHXwHcBIOQrlQ5tTtg3ei6a9ImBTxQl2IL2hD
THTxuzw0wCLB++GLBnd4u3xa5EAWTTwDKCGLsgYfJYB55ZZ8VS23weCxWvJDi+5v2ZLt5uDXc4Vi
vozhecQ1rBhDuOqALGp+sIlmoywGpZr3Dl3ec0Q9XbECNmrf8T+12kem/9k4sHNCqykuybot6es3
LXaK7412HFFGNg8RTNeZHSMhJvaHAr51YHesBgbHo1LWI7IOATp9u0K7GwnTG0TmpSJrbe1I3gV3
pMn5HvBlS64yNZ8QWhKWPyxwajWjALaZ1V8mY+t0x72+J8iBAcCH1nH3OE4K3gQc6DACTSJrjXmy
y7gzllQcCgHRV6fzIM+sqN3q5dqmKbEwn5vPKJDyBX3JLPp8UcDCOvJuIWNzrbl/1C2ec443E5sv
GWTdPNPyHYP0jSBV7wer7uBgwT9wo9ieaMJnaG9MQ23bF5DO+VJFUjpzEL4vSB8O7J3+Y2P14dEn
VauAsWDlZooNtS43FsfMmWw17zSfC//5I+il22hu9PJwhpwa2Is2Zap2JrB+ZpWBPomhvJAIzhnE
UN30J3wyBqnH6AWNVrkFP3cF8CnFtS3JQVqAa92DMWzEKONsITa7CD5aq7ArAT0lCJq4ZxHm0Bh0
qEjIQdf8rADw8nq2UkcTZ31jicQmQBV0sraq3xSjMDbdz9cNYvfrQpMPsFwcR7LDIuJTkvtzFJfi
sPZWfeENbEGAETAHrBLEAP0khtfCML03w0AXw8CjhF57ywIidPg7B5g1Kwqww6C85FWjwHwAdO9x
0sRksUKm3lEGEa3AHoclQOZ799GVmX5glNgJXdNGJOyy5kQjtI4MwkpKQay0dRomrhCDp6yuwFSL
yyT/g44VWTeIQdREwr1k205wN1onlzc2Cwa6rr4E3Gf1igFh9ipta68BPAB55b3KLcisnq92Y/S2
BZ3TaAzxEgrhfc2v8oljXY7TtC82qZ+epapnRzHo9dDeQEUlyM21H3V/FYd8MmECwK3mk3f9AkVr
P3CiTh8mhkE55zdFdQjynOVAUhnQ7hY8mdyYoXUqydYqJlmiqRxibfAbC89OkyXXLFCEFB1ushgS
XQaOt6zWlCmxXJqYFtdwVlfxyzspcFdEGEsVR6CMztDtGfgDeys5ytvMtcQWFU8m55Uz6QipSX1t
LgqKVRY8YvIsilx75c7p5WZxyGwSMYqWHuI6G72CqcMBUK6hCf9WG5oyPNNBoKi38TnYbEoJULJT
JvCjF1xH5sdEqtvCcMPkPv6Qpkxu6GICubXqrDDTASHxTgZ/sp70IkoPLWEv+IpETaBMoN4Myejn
hx84MuimDVSzwXExKYxZ+AWphY+NWMV6m+wV9ytlGOU/HFf3CyuDavKW58E/ETou3sR+DyvK83rF
XCfiJYArkoJhHly4cUnHLU7/l3QBX+ODi+EOXwoTnm+HvCsdItMb/Cz7KjP+byl7A6C37hbtbBR4
3HAbAl5/oluLAxJnZGI6G6x4H/HVcwg18KSNz/cQxYFl5u/o0ktE1m9qRbaEwwvbX8+kTc1su78x
artP8Fl+xXBN9S3uFSCju0WtnWaNJFXjoync2wonbKwj145dAKuYLIip3u4shgCzJyfpnxB+0zKg
BHAsDRhPUM9ZMfDLzI6gUXxq1RidQ90IAAs4csO4aIz8QbP6HV4jCCfXrIcsu98p3s+BHXCRNcMZ
cokvShwKbyYJ90HiOTtOGbhChF/vNoUpF7tLaOG86u93U3OtmKmS+fVaM8bmLjv9PYzWcNwgSsrp
4U7BBW8uAkH/W8le4trqg6ZN9Sq15O4neoUxPuumC0aih6bdVZP4odXAt9nZ3Uh4nmPlVfKjGhPe
gZJGlzhXS/241k6/J0RKZVBKCqa9pG4khxBX3h/SN8nrbdpYrlVrS2vCICE/LZJvImUG3BlmAmOJ
FNQeOel4VbK+U6Fae+BTL+9074PKe5CD0e9bIgdlkqX7bFCflwUAynTbvvfIIsJngVpC5DsM+e5l
9s4DA8qDwIBBFyMNKbpUuKUfsuUGiVtdgC9UYrlYPY+xpwW+SrASQ3J9pKh/K2OkNw834XTasGws
AY6BkSYKCUZMlCegGZ+q89GbFxks8USXbrNLM9F52y2NPYI0Gsuu6akw3RPeHwmeX3czT5yczj62
cLnCoQ5/DIsVysGnGShHi9RjswtsdczpqOin3VtXhIdXYIHfCXj4JfrqBZEkm3vsxv3DRmTaSWYu
vaN6T1Q5wWj3KIoedRR1208P4EfyEy5hMKewPPn4Cd9qVgIQ6qwDe6tI61lE4fnoOCOlT9UOw5ek
dQ3dPnScX41ieRyqAbAosd9m539tdbCmwUniwU2jJknHkJtFwt43YAm4S41eXykK4CqA87wAaFW7
coh8C88iEHwIwD/eCLOWIr2oPIaO1VV0A6Q+gZqdXsrqaL3NBBYIjhnPYL3Uz3XJf2TUEsLwWDPc
aB5kV/cpjNgusS9PkcDMrTpUcg6OIqWsVx4YdjdlWJbziVA9nKObpdMVPxApznnuIH2rlEA66uBF
tAd3EuzyYew54muZo+YuCtHuuLh/KcI6zMAy2c6q2ROFZPeR5e3mPaZjgy6Mx6d8JUbhSi1VjTkS
UUoopAqT3U4m/j97BJ4ZpIyGXMxBxLc/MbM1cr1bVZ+gRuWFi7D0EKjYW7i9fYXsYKd0pCoFDLh+
e3o1IpG0R3UZHqOOekIFRzE4+81OIo/pLF5e32EbyvHcsJbUpknwgUBA6fQmSVEu+ZhDn1M8nzO6
TTQIIMKv1Evq+/PvAXsbMHapeD8oNNUGuerlBURq60CiAun5TwcgxSvmMsxlzSh6kyW4rBkGpVUw
96Zjri0khCEZ2JmuhEa48FOeGEs08pS/5F5JOZLfrYK8NVgZn773aLhjrxreYEGkXTEfXja1aVad
Cphes1hqcsfM27auwcLSNdwed5lPs8pHJMqQ/vc+majTqTC72PeNGDohk3lZYr1pQa/KhA5DHBRB
Qx+dPscKrU9/R+BMNHsaFhVIq7UqyiYBVEAIn7T/vXWobgLuNbSZY3fHI4MWucLuG4LlmachBt0d
PY++M0fS/MZkPnSa1NehQ3Y6V8lc/MCcOcgIOXLGD3C93EpTiGf7mHBVeS14qrMaXE1mja+nBrx2
ILInrw/xaqlDlBbJhvJVqcrbyiBKz34DugDCCh5YVjwyECrK4dwXu2/sBQAxJPbuPZy96/YJLyvo
l7DHGku8m7Lz2qTAV8GofYMXpL/JJm+o74B76JKUg4GEGq3nUIsoeqM2GR5e88HWJwjFRHPDXnzQ
+VKgx/fXp393u07rrKP/xZ1cfgGQAwRVfrLiS0aoXSWsLbeAjAWcm02AVm1lZZ802Zpz6tITH/9T
EmRHrH6zkQCm2nX9qLesQ/xq/cZAha+GFjwNN41lXUlW9Pv3gMfZbllpWME2x2htt7pRVB2nAjjG
HbS7zBvPFvkfa7xR+p2jtKbKmyexu50VPijup8X3n5Ege6F3zQykpXnuGhbO9sqiwcivPtRracf6
8fksUUoSxn3K8lCXlmsZQrf/srFryEHlUyX9W40yvpBZzFCnS62nT21Xfo/pxFFm9VN/Yzm+hck6
VQtB7f0OcR8UjiR6dEagYCthtgO43N+5rMa6KcN/iAm32jqfvExYL4bVFulXyy0Y4hiVb2q5E/cw
T7DSaOo7+gMuMoVB5psGXv3RIb6L8iQKk5YRjROC1VsKJK7/OyjPSv7GrieQGSbtOR+2PqnPxjkH
LMiKkXe3v4PP19Hm2qrhf3cd75WXHfh/+Mi07PsG2no0CXDz2leP8Zc+M/K33A1smwgI0DrTbXgx
6FW4VvOfxgvwSjr4qpxZvcnNj7ekJ0tTgxLWG2ZuC+TrHCUqXV0uwvucFLekGx3BcA1oAh1E3TpQ
i86bMfbRLONnera7PBJv4QJjcmpjymVDajJDOIMiDE/Zk27q7deqZOgOOA7S0p+vuYNLgLtmxhSf
KZpXnTYBgfUjPi2CI7XuXAIlwG7AvbR59Yr8oYk74T7ObqTwv+cI9pdbmSN9W/yPeuWtFJflsBzn
zKkGAakGeKTvu6zOpBgf6or9kY+HGVKLF4LdIc2bx6PgbTBhOhWxIKlwGNDe5/BDEOGK318GReFw
v9cqzaMLsq3dWODYcMpy5/+Y4TVrGpoHsaErsp25bse3TY44KyHsIVLVuj6hbHqkmJPQZfKiIsDN
kmEmIMLD5evQ6WqCsbH1w44k1epbSx7kXlXDo4t4VEp02jvhoHvg6i0oF6dNYWuURPdDTe7FN5q1
TTPO1l/WMqxQVRaVRGJrvDToOlowouoUSadihzAnjaX60w2gjMqfPR53GyysoU/PvrgP+QDxU+Fu
37NhoasfmKHMDFzUuPQhDgZ0ZuVnU5rDjetl1Sg2hNQzCDis52WIqu/UnRohspQEGvhAPJgfX+fm
7r7XTt8KF3bxczE6UIWLDOUW0YUANKpAIyffx3JEr1nFbKa0K0UpuoA0ZORcFSHBWI1jlDv11Pk6
GX14G2V1IDq1VAWt4tlowl4dZ5dAOY09bsFC6mw+ZiTcojKgiXg2S3uXp6PDUYlVhR+qGmJCWBA1
v1ZORx7lOA25Gkjf6EBMOcaDGFkodpRz0nENo8oE7fottpPTukM1EX6g4kzUE7qcwqcgwfal9itT
xtbO2jxKkebN45CCsJ02LoigrnAs0OMnbrEnch+f65LgvQU35EhS3Skfkei00DIM9e0+jKgjzru4
il+Pa5BqRpWwXXxvsj/UIlo8PNOwLVkpOMvzly0eheToPOrlsAbzG47IjCj1QReBi53QKsWuOEWx
JrAL5wBfqz2ODS8Dh703eBS2+FQPfJqC2/zSMk65x856q/VT3wzBeQMoXgxEcn8jdCDUAaIM3FbO
zkr6skSlJb45woA+c1251mj62gok1wj8dMiwAwTYf91512T+3rWfPVoPILSl1m3ishTv98HqUndD
wuDLdnb2hwLXE6zO0aPV8QWPvo3I2vVrXuebzGVfHQiSj3FIhJ/oWeZQMD/tXCKaNOhTK/eK0ZIR
9/4M22ZaIrXakCVJTQu7C6/4xA6OSaT6krvceBcjeW/BgKmwYbOxbMwWhD3DdNUXrmOmSBRzX2kq
E9Wzj/uikJMX9ya71PCTAeukzNtP7Q68deV2fzT03Veoy+RRM2VQtiVYssH2XyzaL88kJ+9u4z5d
fOxHAi5baib+dwu+e53IWFp45j0b0XCxNoGqK8RDylu/nBvpaW+duCTXeDgTzVo921l6pxszf8/2
w/XH6ktxYCZcYcvpQuqFnGeABPUM0VUjjE+AD7rbUAZtdyQduhYivEX6H016s04SIk1lhQVtaFhq
kGpLzXmacUbeUQx95wxAWPjMxFhzEpxKpyaEWJ7qeHKBaXIaw9zsu0nXSr1ALSA9L3KwTWb8Xyn2
TW+A/oc3rkeJjJjhW1Tym2sDxgip8BMjvDRLdo948LiL5R2/OvPBwvCUu5+I7g5ValPszmg6RMgB
ZgfGgunp2leOZ4cahVAowgvDSQ5BEncdO9QV2GjpNzSDPJj35z67BYFy6YSyAZFWriNZwcqO/pWs
H4uhVFqx1i4Em3hbLjtIUv7xPMWf+QYnujlD8xJHWcHvt1xBa0j9jXKMAxiC5Nd/cN9mUhFOiM/K
zzPV8qyPMCGemwX9/H8HfdUBuxWIujdzsqpWzlyNhLoxZsMeSserlh1rsQbeJvU1558u4m7cFcJp
gHQHqZEqb8gIWoHDrCb75EwciYHwgHUfPmeUUtWuLB1wtLmQ54442n6XItfd++JcDXue5a8PCLVr
INa8q08JOb1pwNJx5XY2oCxW5iy39oG+SZ4+gKHTk6aVTfeDA5qy9HNBBf5IoeLg7k2V311dWESl
gY7qz9TAIG8mFxUB7DPm+htrGpsvkm21bSLscDF1kS9tgXM6qqX49iBKMoCO5DWPktg5kRYy4n2U
lghC5nKigXyNxNjS0BAb9XRG0mHdbG7sQM3xD1ow2up/2s1TmndBYzDC4t1sWl36yyhxnH3UrtyK
P4O+0dU+g59F5wne30mbk4AzB284SfwGYr8jng1CZbLgpPWkVYezAGNhGgISCXwLARoq6sMP2XdM
rYK8n7PvQzxJK1DmpVzsBqS7/nImwFxqAgPVnmLUfSPZGWDpJvKjdBsBl2FX/cmkQUcgfAom1s4Z
K3cXGrDUOyACQ2Bvhbn0i0wOACr4LMAZuO5yZXYOxRSzwcYwhNDbSMIEyl9rggP75OVXpsmCccAm
hwSOaiBJpSftLS78nc5wQTxOXjIzYjqg06YIjCqp5hovfQNLao5y+Y0c91IkHP2rL51zSq0g6YDC
8eojJTgJ22LmHhqY5grO8a77lrGawdYYRYk2aUeg1ZM7WGr6VF4p2Qg9sxsP8rG31kg+LJG3qDKe
AdfVOA8tPcdA+b3wXAezv/uT0KYc/GV2BtTndm6fQA44tvayehehan+1vZdFwEwWcgXkLI58+rz7
h9MUMm+1voRl3sWpg6jSclUzSR0uoHY60HOA+9NE7IlhJN+4q+ksCmTCYFBS4dZTyiIbc8W2cKVs
xL3g0Rfqj+mu+0UWL1K/m6LUg/liLq0fotAKsHHezZtLgZmTCPP+pyai3sqLhya43Dz91TBrUcY5
OOmwf4tmexMWlAjbVEjJ7bJRJPRHUQd3yrJMohm5iDQEzGdNUrDE2v+b3YOv2KSYN5lPpN9klIwC
2FVW8+a6zcy/cd2g5aDpFnAbli5d8tiKOl7amCXhxEqikghFQEe+R7y0q90u9qmarf00LxT/cjCk
6ZEYg6oS66eDALNGfkMIOUPuC9myJbcM93xgI7rPrEU8+BaI01yvNNzWqUy4quvxV2msSGWlNXPC
+ChW73Lrho79FzFdETNd5tKRSYwMOfgNmVzzypJXfX1M0oiad1p1LlguwXc0cqp/eCvSQFyDj12Z
+DiQudlCTXMIHAQX7H756+/C1W5nPPw4prW/k8hC6RH4j/VdoMvgmXE3i+ll5o1FJx/1w8VSleBp
ABqxAgEub4Fl4OUzUWNNW/DW3A20NF/BFX6+JazFOxrhxExf3vo/sV9a/RO8nWZ/CSNu8eIWLmTe
cb2MogK3mXEkTDF6x4I1JovHIdAYMkCbZNZMkniIDPWVJkbYIPVesXpFIb9LpyxjkB+9ZLwsQloV
Q8YkE1hYrev2ttB2OJeqLi2sLIuIG6AvOqZ25ekcC5Y704EyV/VzbHyzR7Cpx+HJtpu9QZ4u6k5D
FgEHYrKTqLxclIOsRuHe4bngjUgYJN+2z2fm1pyRoILicTVgbyFhR/EMJiHpF6aiOxanofPZ/kQ0
ktcVqt3wGYXdp9ZMvhJFy7hQ9dG96ZUV9Py8FX0Jjn7WR0KZHRPhiHv9B7jIvgn6IzPWBsJvu8bA
aPno742y3grX+PnviurNmUsmksPu25xywFftJxquBBnYTL4W+wl6GSJ/QZRjUAvOMM60+aQGRArn
ofNXHRjZvn3CN5uPsIQi0eM+j6oTgX+v52SjFwFWfJYUEOiJglLm478L24Sgjr9vxEAH8e8A6clR
MsxTPkBuFQbGVO+ou96TRfJVGiat5XHt33h5b9VMb3jYLGx99KmmMCer6OA8nADg4NLZf8vaVp7w
USCiYD61BPeTlOewxWTSx4IMQkVfdYqzsoYnb1qb5cXmX2vcxcAwoaeuTH3hrluphZY6lH3tYiZc
0ECire3+bZWJwcTW7aOULdSMSA0AYtT4n8SEgyJ/v6c5QnWk64wjwSHKpMqooDeEMt7V0XkmbqDf
ZnpjYyIpYOukuanmmVNytzaD/TQPbkibFw70Wd+r5pyH4WCuhhdpqm0XWG6iQqQQvMWOpxo69Z6F
Fl9AL2y/5Mznc9G+7cf7MZn94UpnnCSQYxwjrfPOSEhNjoGYir3frwxA6TOFXNRQKL7HBIvpoamj
SaSLbGJwMl+DwpZ45dT6BlLKsnUh+pLnDsFYGhg2ByTJ9TYm3wcrKj9MpEWX9N1CVdd9m5INu/5l
YvS3BgBsyDRtsCkvUF8tm+q6lxNN+e2IqnJ35oAUljcqBMUqiisonQQSFK/XWQ4HxdLUxzABAqZA
WpmmGiLd7vHUtaYoLp8NXSY+B5xgvRVE78CNmL+yjd3ay6sQG2FbDHS/e1Zc4Y2HVQb7IHpun0WA
PZC44IVXiGzrYzHmvJ1uOC5rUuT0Ccu7Pbx0S4PlaHLLzuf1j676/LHqBKnR/mf4j4CCFznP16YK
0T1KqOCscEdXjOZQWC0wiqOSMa9yENu48s+ELRfCzl9nOr5c8aJPFjn6XMRJqTVXTVjfhX8u14PC
bK1YlhX7cxUkw9PK6Bd47/9QWkKcrHq6dQusdF3w0EiqYadrxbzZ14b+RcjwaGXooThIkGbB3dIB
+RGpjYpmchVn5lZeKiAmJ2zNGBJOVq+osNAdpdRasO7Ud4zEDWYIpiXgqS/tYf2Z4OVuXUCnKz/t
6i2JIpw9GP2HdoF/slhairJfSsEjFkLpj2KHyFUG0ilGOh5S4OlBbenWYDVQ3r9LGV6+5TSkPou7
VsGyV8chkuIBs90oYJEnY6DzLVN2KWyhrHb7h8j1CQpKC6IoSNjGfUzhd8RVmzgLlgoRXwIhhDiQ
05Y5jsO1aNaqG00gcmeSDYmS4SOe7hUMc9vPkKT0oOLP4jTkh8pjrE5wqUDEe79EIqPudv5wgniQ
lQ/QxkJFtzRQL4iFW/2P27jSYV6cYy2Gp0pEJD+s4yRxIqf/K/9882s0jZeBN/H/It0gIm7exOM7
XoX54j5NyZNJTWRjW29yijAOpQOzWH6efffbFtysvfLnk0aZCpwBpp3r7D6Fuuy805OCY/fi+5Gm
1vOIYIhAAxI32R6jYyoq/UhSlfhpAiYMmnrQhMTn0v++MbPcxVUjYnXmdeImGiobKclQ0Wlu5dwB
Imbww5XyQHvXeRU/GewObEHbZHLTqS5wQGAx0FOrTLTcCyYIpHQv6WPWpzfzyXqMlKyuetLIDWHd
tfNtxwFZ8Zh16SdOaN8KgmXvVd7ATItlERK/ibhnTdqQBos3IbnpulCPgGR0fqolqOt9dy+/nBqf
PLwEyXQHiOyMUaKv67lJuQExbqKQQekKjy7SAvM52Kl+jgTswAtGkZ1CgrLNY7U7ynEZZwmT7WJ2
UFWYxS7GDLD46YOzWZobCZnvnPr6wG46ioM6URP7I2up0X4wGCRlakwutgjuJDdWxszQr934Pb2p
EMGtUtdhDHIW2pI0m/IR1llYVbcj7sKNgSVRnqGq+EiM5DSbJymXZQSvSNyiauk99xpbp9129Xug
+F30yftC/L10fZNCaxK9mmrAc6TxmVdNhKsAuygotaEScKeclA/zuD+Jv/ZASwiJTRJVzHyHDYbB
VWS6C8FN4lVGBj00/eJ84gyOteFGYZVfVJ8EymPH6ywiybwE2iH0Lho2kmzUYMOY67N+L5kMSpuI
hjy6Xc3EE++YtWc6oR/e5H/JmBnrpB5l2SRCL/FZdSd57EgGxst70ack3TPC8IVJaRZHwuKvG19e
NcO8qIQhwaxBx19eKUV+bxryBFe1TSIyQFeXu6IBMJxd4EzkPO4FkhOMw8usoNMSgmgesFqOxfnH
R2gVu4lYqS3XX9dqi1QWpthvrSba8JYN9+sHSTKCsEFkUoR3jXFaPJ47qqxWWRFM/U6kRnd0dLIr
hDCDmC04xvNsKgeprPeTcN7bQzTsMQAeyX+MRfgP1VQsZ30N5yCXRDk6E5PE9wMB8RSB8DX+GwUW
myHVvPOfJ4soOHPt+dTotZr8ylT2Ujq6JLgqcoOfhfywZw6+QuUsB7mcZlbrxM2/nhD/L22AvL5u
yOGwIrI9SJzv4KJK5I6l/sTHhDSS2yU8oSP3Suq0fI2B0rJ1npvUqZ+gISis/ftIJeLgmHjT2Mu/
Gkz7m2dn1nKP/5VmDDinBQUAJ93j9nztySMS5RXELOIjI5MU8b+uk1vAKxL1ajEZmglL0hnI3/yv
JM3ILDOzQLVsIEey+vWvup8P4+qPpO9LqldPluLhJQuBfJzd4hwc/jjUjp5vDZD+jiDT5/p8I99W
pKpYuk1hPWfOE9Amp8OY34RWq+HwuvIiqX115iSv4zp5Ibl7D+xZ5I/s8aANrmQXA8I73Ah1d9bj
CTMd+R+jUmUDqrrYd4GJXjoKDHCk0o5lj0ZrAchKbmN7iC0cccHnbunp4I8l1gVc6I86NfEKhvW4
F2BroW8FkxOXdOexLb3QPkmwOrQCRqN53dYTev88PrC1F4qKDd0r1rkSLTqkvGJhnhGdv++mXzZx
OyfJCmDw3sZzjhyPrTQGTuLrre2rp+BFoZW6n1ZJ2hmLVFPTtSTUf0kHBQ5FMinFts19kmaR/yZ/
eA1Oe3BzCqiaOqGgcFXyw43c6qlK24iSus1J90dTYLd3q3srEoanb5Y4ZQhRKpv8T27JEPJrivb3
/iAxobTpXkMKzngkQn0iGbtGXW8+5/0EjRmf/P3ZHtwCA5w7/vFjS2RtBMC0jPcPYfMoO44srI/C
YAmIMDVT+/JmBFWP9oTbmCKW7skHs4Yl28mJmJam6c5wNfFKMX9flbGE+54kthw59u412aEnaZ6p
BFdPFm1oD8Ikrnh/Wb0IvhOdxNq3dzZRlXIvN7TWUn8vyEvadoH+W0gPwoWrHjR23TA3NQgG50T/
mo98FTI/BLIESQ3yzPkCVDM/fZsb+5+KLULaE+NVqiQ0IUhEOJVD0axY50r4niUsezGeNybOqFas
LN/wzpXEWf+eYZWiJc/bdP0GJx8uYIGFvzssiRVa/AySKtih8TWoRwHrhhgXPoT3acUDuL02eHO/
vdUjM03LpFUaFUZBcon2TSNXqrpU7YCpb0BgcEsiOQwtzyaOvTeYhlKrMB/iwHWi9rgiJ/W2Geip
GvBo/NqT7Qc+vBy6Z+pqREAmM/BxMEp8FAXHwMoxEvaKF4d8Xz1lwTz5qBKmisRVX+77cvi0TC0k
OIxlBX8UNsbkxAAmvyjd6UGE4eHA1eitp07r+ZpXmwrpt55D75pgD5dsIYZ2/x+c7XacD7Ef4vO5
gmIUqQnHc+ueDtE5wmhehrAAxd8LmOZ8t+sSEwf/rbXMnSCYgDa8Hjpe/x69VS/JA54ORPk0HlLB
yRFHcLpIoSHBHETWqockTuoh2pWVnnjF2P3W/ueFQEAjon6Jz+v5/6uv/Z0UUcilZPH+yGXYleAK
6/Su4lKl0maqTd2ZYmCO8ORl1OHxnXeTpYUQcDaq3jynqI1GFXlqOhZbs0REIIYb1UsQ/d3+DtH1
+X0eiTPL5U+IE8XCzmzW3ME8ekZ9/uS3ZtcKkojpLi+9aK0Odx81wgJzZZTBCEP5IWabeKWSl3VR
m5JSyQbVk6fWyyPNnie46oUtAcby7CK88AeS25YYUPjRRu9TeI1JVMrZgXEIxanDh6WWKjxXfkB/
ruXhBj34L+VP/M31xAIAyKNCa2vKM6JBbf+LPtxCAhPuv+ngcRKDuIHYZilSv9UHc5jpugsXfg9C
ejBKR42FfQQZOE0PHYucgKmDrR90IwM2xMgIMf0AC5Hn2sXRT0YX2jGAgUVNNVxYA/drcRxLMPDJ
Vtcj3gb21q752P3ElnxaPT3Bliw2K/xaEflqydknG8ZNsNBTfggU9YBH8t/qygBJbCaukK7IM1pa
DsNajXQ5f7yxzwUU/SokckJaeyPuu6cC4rfXX8L6/ld3SYxALcaOnAWJ2xVomoD6MNoAD3tM96Y/
PQsoRlQrpGDsw6TSqs1/jCnjCG/Ja1Bxti62rlMz6jktnlJ423Zo21UzfSpzw/GBHZxzDOhgRf94
Az9u2lK54bUAI1njEjZ5ROIBZ4pmeDI6obBpeh4Gd+nsVlvKOLq4yDd4/U2CjE1kokO5vSQDQCR4
s/8i59NDoG3B3p6b40QXkqK8TwhBtw7wdruW081VotzRzb7OIJRkoc87jNEn5G1/4NRSG7gFYrkV
zx9NkpfFtV1LuKiSrbtgttrUBeI8HzhMUlyQRfA+JvEmjqbbREXTaET+1IjvHfM1aCYMMJuEySAn
qTMyOYMA9+wxPP6mAF+ZXID556eJgqg15ZH7vQrQjG6wM1ZVcwF6qio/ZptkLHEN4EISB4LR/8/Q
XyVWwch9M2ynSYyt7xkIZIpqHFOfHi0zKu8MqO7oojE2PsmlckmKDe4B3M6HH8ouejAeT5rhrKy3
CpSIZDT8fLZYjhxv5vjMAiR0EVTT0KFt2kzu/X9papuZ631Y5gfgzfqJRtYSocIG/iuXneeXYOxP
8ibIAl1cJgUK/dopArcKv7OzrexfJ8Zdp8itgZrYLKK6m2pi3F2Ccp1NdzV4A+FuegqN+ejEURr6
4cgH7xeCXw477UyGovd3z98XDdhEU8tEm5CJzJdMxnK9FFI93ZvQGrr0PoQzFV+2A8ewttxftITS
+LEwwFOo9dlcm3q26otrcKndGee51XYB4Pb/ZxexK+9cdwp1PET0bDWcokybV+eRD4vwFwQUfZb1
k0RTcWhSc+vIFqAN2cHoYRC3wdPkwWYCTimKA+c8xYUgc36JS3U46DMBr1ParODor/2UzGU9qGoo
YNbLguFZhB/4pE7nzdvAdSdGy0E1VIowX5OZDMf5tcYnMp0WNzCo/x6IemfPx4qsEQtU3o8kiWmk
HxFrD3vAiiK3su5Yuhr1pHFOzd7azO46n0m4ud6uajGmjXPjoZQssGo1p+UkXRZ2YN+NWA1IPCPM
sGU80Xco6yxEVgxOm0q/uu/CnHGHmrJZud8V1oBwsD0z4mTBhqUapNntEtuMiRHznsAx7peYnAPo
Fqshf5SolCjqmbrFX6XgVmtvy5Surf9Rb+/ZoaG32tIrlIAYmV5dUWW3IaO3ajfn4jiLMcX2wGuu
pYLPBD2d3cRahe1c5R7dWB8HF2PbATtuL6V/pivFkPMLjZ5LtlyvX0v4zApFkUp6G0GrshyPMp7F
x/jZhp+CQzlI6dCRgMS0izD5/hL4+UShdfFUyBkLYOihDBqa9K6yBWowBroRHvDpSYUG9mDR/9Y5
rKQf3ApG3btKVg8LnayJUgScb0lrp0iOIKs78A2a2oCMvOZmJI2BK5dXW+CaOzhoPMME39WgMOGE
vmwuSU6qRrTSP/KUND6Pqd/cdA2NLhCQ6Z1uBUsWixqe6N2r1u/BdZr0xcBCoycGTKI0ROzidEUg
r2wdIfp+xMJStqQKs+zSETxCEk7wjuI8YWGi6RriWq0+Na9yWEwS6raIjQSIw0Apm7REN8alb8BY
qtEfkG6ER5To6QkaItKtNCXWHM3ByR+7SRYKOqn6AprR+NnH8LyXzpkQa0vgodHG7JvmvtELcl3+
Zn2/DZqoWy9SRDKqZvMiWX6m8rw7FiCs8QYpxlBzPlTXoaolyHtFTRSthGKhZM/Aev9eS51h1WiF
tDEcAvsxAlM0oFfKa1lhCYB9DIHSKN2LpkQtkG9+PbUtanbda9l/CQGqeROg2HMRoCZy1G31dUt0
VEHJFYnaId2+cfveYd7w2RDykOFr7TbvYs/CiOtK30GcdnwCAzYvaLX7FfwS3AVtL2KblJZ8dCDi
UplL6e+lu9G2azI9LW8v7RTYf+9e9zkBBHdD/pwyOSL+K7LpNaH6eMkt0MG2Eq8RCBP9DsTncZJs
T07claUuxHaviit4HJe95W9+PXXnmMJAdrCvJ0NmmtsaTPoMpdY3XCWATZFs8XtWiN4bQB48VJEE
wRrQOUm+O4Iq5DwkQXLjy+6aSlVWWg7LRQtV8P6NAxpYeecoocGId9QN0ol/dC9rP/c1BeWuW6YH
HAi92xiu8C4ygQRb7qP/njWcko4im+qidL0JGCLsHxHpLKEO2+IJTUOCH6P53u2+TyO33ueSd7Ng
hM+8vBnL6Fo4oh/j6/dJ8svNRFylmpmMYBi4vZ03tRcP8cK/YAh26ymJ/szRlpBK44/T53jwtLqp
zI+Rahyy3Z8YEKAMxW4zTcWlhZg1QUByXIC8V0hl5lpOnq+3uS1zyR6N/FOYVGphhlsHVWLS7br4
yvkqL1b7fiNoXE19D2CcosIOrEqL7v/eoeqYLmp9D0jubj3hqAofmXkJLIdx1YEimCK7HDw1rdpQ
iBdTz8u3BBAukkhLpbirOZr+oyr20xvOqiVvkvPI1sF0KnMcMHWfUXD8z9PHhCucqVkTGjwXAk8l
Q98XntfI4cIIDu5gRP3GD8c6uHB043CPP+pqerHDyOa8N+z2+51gpqvCvuyBZdk7xLFxDauXdfgp
GRt8BI1fUMUsJwgeCzzFX72JN1Cxhu15dE3wAYnfXFdwClOHalSqznaj3qjhfN4GwQ8T9dpegdnZ
KJPocYbBV6Anr6LsRzNAgEBTXbIA8C2AG5KA0Lyr9A82POnynHPWcSYHyqlXrLW6V6cGT/701rtD
9L5pknO89ydrWB7QQc1K6Mr27gQcZiT2kjIY4MC7EH82eo3aNto3NYH3aT54qlOWuoe05yCDtK1p
8e4c8OBn8WBQCfpNmPHbiANt44r2x6NqBxLDhxWhXUiuusFPdChVdSFMOJKKWWIvZOQHZFO0XcQ1
JqIqqhD/PKc7AMKGzq5a0fInKXyPutzsw4Nt+AzQfWPUy5itdngWToNQT5yLm0SuuUKJDFMYOiy5
Xn7Z0urnOqapsd0OR+IUPqzNl2xKLx8c/znDcBwUqYCRd/PANI2WFpxkAJuY4u/h0/+Ss7Tu0PPZ
W+UkJJ1qUWfnh3xO6gAUOroILveiSrmChQApmfxNrSFxOyPUYSi6cZgllGBs4RIZ5+0S2IwE5T1j
ReSHCpqpwI7iVQknpkuGPcP+MADxyCf5qK84Mi05Y10Je/QUZi8E7qeoqRVPgK9wYenzV798BSrr
3AzlUAUfNuTJIYkIrziXjVFn26TeFo+6LFJw3OEQiyTAJsubu9NAmmo8fi7IGfwEo0vgrMNCwwwL
OHSe6AOMzpz7QzDd0FtCHtTfCskPCDO2SG/GVdQzJ3mA4VnKr3caALxvgYrtqfDL3rosnVDeX4rP
Wn+uDNgYzRb2FINMlLCXbX986r71Jdufo4IpCpwCER9PMdiEgfdvprsEj63OLsym5ETTa9V8OuLp
WbDcU8OoIbYYZ2B2R1lfyA1RwxgvOo1o7UNQR3KmnJ6J2bRMW7RvDwOhAlTpuuaXhY8EpoExrnzQ
qAYC9GYu1ntcIgCI42XnzJ+lchjLggszvun41ZkISnsCMToz0jqZfFppgPnjtXsTYOHX/50Co5ix
p67H+Resj23ieecDTAGhEKMeQRMWGl6dqs56lJZ4PTL0GTY+JvkLe+iDrXLdfsY2iKbwx5SJkNiE
6CWSR27V2rS/RL7h96rv3UcvmH511s/5SReKmxRPR+QTpL/OXf2Tz4NpIQldAhwkGeFqfsQaQsPu
cqaiwF13MW/pbqs2uZfqU6nAYZTtVT0MTolJLdTQmv8lux9kzVYnpCRs44FdOx4GKKKq48xwvhgg
cLyGdLTDP9gowJwyQqurgVkfqozT9P4/XSKp0iFREg864nFOtQp7QsGadpSSbFo9S2GSN9mTm7AW
C3Gud3GF53wV1/SXeOnRiCiPPhBjxTB19fuOLol9VfnAnWL/J75YkqHnvwXYcvLWkUsPqO6mlCco
XyH1gBVYvnpJJDIJMq8LFO2xTBvNUkcM/h7XgbQ8D9TH8SuHYpAb29qTbeALFpeAkKpLVzSEtEXJ
NWbUYfruDx/b/3yApV+nPDTELPPrqOYMCNrDZTfDiWNbDa6az8O1jJ0uHhJAbU1Z+tD8zbL6f9/h
hC1Jj2luCysmvnFrk+LX4Opcs/OB8k7F+mJtvsj4xMPdM6DFZF6gkLILEeMSZlq7FAaV69qvyhYG
g7y/winMtapAQDzv8d4CM4PtOFYHPPpM8aP27Etm1ZzkCa17s9GNlgLXxz/O39ir3dhw9fPnhrRn
h01m2AzY5kBQW+nv1+3jo8eNEEASuZlSfp7yQtuhhBwp6uU+K9OiJGuibZWP5wtR2N/HmJvweJyO
UjPMeBXL3hD8clq9Y5RZK+UtM3c6wJiP6BC26LhWH+xWhLcjSR6Twnvp2APv8Le5qc+mqrZlRRVt
uzpsam9mN6k0qPpUlLAsls9r++d8ww3c0Uor9vMD37IVgD5/UdeJJPG6C5TCZOW7Gpr+5QQeYiYQ
4IU15nAr7ZAO3ltrmBSSCijNaDM60Fy7wYUk0hO0GudcdwsG0PjRiDdcVamJTEso5EfN3xoMPTFd
ykxr08zLgqM3bm6bGVBXnZHok72oo0YQiLEq/3jYsozh2qCoUp1ZZfz3z2ox+cmoGFrNzplaFjvi
g8TxwWiSi9lgn6eTLfmMw30B+PRdcJd+0UtbpKUZ6Ma0RET6yDg2COLimg15JkBhtx/Um8yf7AaV
xiVGSOvrWh9kHCJRWkcEJOPvo9tmqpIK4Js2W7JLgqaoq8uNOQHNAyh9ffVtZSj6ivP81vq5v7Mj
p0js/bqnrFpSAdotOv4N2ASdCqFYLxhPDHqc2mYY5abXRBXfFiBQe44A8aYm7ijOIsSmeOOsXOC0
sKIvUD2szBMdASoaqyfjJXujSKEor9GZkHo/7ORR0GHpiBlpxECndVovoqQay6TYNIpkc0+3JSwm
NlY5eoZoaWaqObOF5gLfDo0Fm5JEDEnqTXCHOA0WUd9EdS1oP9ViDghYDStJG7QZdD/UKMcZd7hK
o5fkaUi4JL6MtqdQZr35qZeP24OY4uWoxvHJDCFGMh9GSqgBcZVw58e0tJzUhCcvvwPZ8xeKuMLX
ABOocEjmeVCV7PqbHF2BrPmf5bZuvbmpSZhA0YdpPz9GnHegLtERGYmI/LCAwGis7peUr/ztN4+T
Z7I4dYPg5XqxUoKaT3Itmc9BuamYH5oIBl6/8UHTcVEHemD1CfBHcFDFMH9CYtQern6+YV0VVQ1L
RF/uPGHerxZ1C1UewBzIS7ag5kJ0EFLXVO2EYanqodrPNZNGCIveHow1WmJflXnnK+9l5co38Hql
efsU0jRJltNlimPv1iIEwMzzluoUnstnrf8RDvKikubMLG6AWCHz7RqechfoVpYPhPuApDQFua+y
2QWIpVEL1uvlhF1BhIOzkcERfiPZqZR8hycv6NPOS3yBRPHHeRivxEyJn4txk7Oupc+j9uJ3mI//
T6TBgON1cX0xsf+TZV9YFTm2IDbolW++lprfd2MNUAV+LoZ1EeB/UlKQAPKoSdu9zsHl5+fhcPTv
KFASF30vZyP94UbVROGBSWvUJz6lIpxz++aJDKwspYQyh7hdlOOq8nigsZYmCfFvawwlytmOZzOU
jRt6AWndT4TZKHyoTMndHfWZXFSLsHTKJWsaPHagNCfdgfj94U3XQr9W29yLwUhz84JGgkti7F5E
+t9pSVzRDGnSHg2wPITJJU6TWh/7Co731Ps24r4Jq2A3EJVa6F1G/WcurJOWHZ1cMrzSeZo68h4+
3p8A4CeSL5LwCN97AKPYDDBTLbmt8hNUGxDLGpfxk6fZtCXd+mDvxvCFqZ5NcoC5weCEhoxHBK2g
FzIxuTSQl035I3NdiX/2YNuHJ7Ct6BahtQk/egIPeJKdPStH9XBzApqrUYBCjJUw3CYzXAr+kZEF
GXhqxcTfhdgxXjk27U0IKNeBRuMogaefgt/Z247msUbCzgokjP8kxmO0zOar77I1UoCXxnf0eTR/
+h80emVXi+8n0l/lLYnMhDcM3AbWgVUOPtiqCkyI4F+2oFEn8CvpiwWwEs7E0HeU2WKJMWNeQhOP
VVdDH8Kse4iYVqSJLAiUy4Gx90R9WI/IOtCaCeutlUxmvtkHhiqo/5FvQ0KUp+ZYMIcE3KD1nUgM
IK7ZdylS4IKFeikv0w9Q1V/sMYbDUZ8r/lNyBAeij9sq1TG4sMWcy4bY/j88fR6kg6/9rIZMML98
gknpVPaRNikCY/ZIr2gvr7XvQVFxzy/aQ1bZ419R4GZPg609BneXv+izTWvA4sWcscRsuLrkP+Nf
IhpTDuE3sEXfIzVwrxDbr3zxFkaZ4NzgkxCS5qHMjV3PIXuj/9dAazgUSSKdPCCdhmRyFPeqYICo
k/9GPy7F8SH6+cAaeTnaaB7QnClTFmbIyHwLQMo6Pxzn3YgTrPXX+w39S88uGmKsKsESRzDQ53PA
1AhvBwzIUA//Zv8zg09XDsjeivdsy/tzKEFpjX88Ng6qZGKsv49sQ/m5C2OZmKQcqCZi6rE6xSaP
U4Mq9phLP0XgU2CWGIrjn3bbkXb8I4cB0+BLHkkIvjNaCHNXYeAenPiLv2XgMfQDjoIilJX5cPdr
Q7GJBbwMfHszCWVF7osnYi/k8iihEXnqYu5frv7bQsA23gCKDcIndxbElo2pa0HmmhZ1UZAkcdsj
BZ0O5A7cvH/EmAY9uHyibBwU27F1uyDqI/Tx5SC/kzGXiwN/3/IT3Idd6ua4HdaL3jSnQnHCKHbx
G75CdnBnBlrSuUTzra4QrFT3CMmpk3IReoj9vXtf4UVa4QgG5HcHPBWdPV0e7AbUp7oy5PPxuL5U
mMNEYe+nH4ZvS6Q2+SWEMBg6azIbOgQok+6WTh39r2JUZn+UObcTF+mvJ9/9TrJVAns5RT3OcgMH
IW+oOyxmr6NV/iQaFPhYv+rofkTZwcQa5bbATQl6WQfCEQ1xu1zKw3lX2WVwuwSQfSYuNYMjQzQX
VjcmfBugwXfFckJqtG4PXgSotlMyVba9Ap2cN5HkqgF8hBY8kAQJVkZ9Oz8Pu+hy4oUCvxhY1GwY
Vufb5uMR1ui38ELjl4bTbKm9ihx8hPMnrEFZCoefz/svC5YWxVgIsMXm5fexYk5S5zlpfxO0XZnC
DAf8WbYyP3Cuo52Fx4kHHfiUj3EqBT5dt0iZKFjoqZlqyx0raJZpxRXuqJ2K3bAIMUIehQO2UiZN
PTOcmqARSQb3kUB0nhrpANPlw8jXjmvncSfMw6Hvq9Ajxrf7DrKjaQHWlVd93N4AtXyxCzpwejKe
9QWjnuIj+RCZ8dRpSFcbvwFfqzQNb3Wdltyh/A2AAaI0ZkQGQfy8uOTMpW47/XSuMvIatuYvgRM9
vTtHLmf2ngnebEOZ4OPEhrZPSVmba3llawbrIpXH5wHuHYgL/Sml2QABnzvJKvY021r0n3r0Sma1
DdEk5US2MW0Geyg5pCzhQaa3S5cFeqTQnDzIG/Ianb95Siy1wJZakMYiu0g6ZJg5BXLULO60Uzoi
TvTZ5j64I9Oc+A5xuZOpNK70FSSuFf4fZSm4k8dL8cZR6iQK1lFbcoOeDh987QgYUEZGy9N030e+
hUhSO/iKYNfhwmlWauS9yYv4b4gI6CPrRlXXDYGGrGD5ahuhm4EkJq7o+l83xAY/RnOIkpamQS/W
wS5Ak01bhPWdVx2nS941o0Y0I4ZfauEHXmRDgFGccbMZ8Yfj3h8s52z4woqHwEYCsXTzZy7F9Fkl
OkpQpD8zSHooznrK5Rf35sR2JCHEkliml7HB0HBNCi0KXkjXBCTx/13NGCJgAVxc19kEP42Rkf+u
J71JOcrHFztUFjsESBrtTJCo92/ITyJz4Db/3lYUCr6IyIvxOI4eHG1s4k2+YEcQTxBJgQsGBLQM
GyDJ8DXmiSnCOKZw71h7m1aATUnHguwPBEyER3Z5yR7/Sv+UhEgz1YtlkE78UeehR9kQ/Mclo8om
ntqUZ2D/gPzk1ucY9qmBxdshiqt0u+Jum/9aoJY0Zsxf80kmNtcUWGqr7COXD0HBcwBsW60aB3ep
gLpnvNb2BOUFCjdwAkK5DQmMietkjn+Bk2XlOM9ISvqjOYmgCup4rKP0pkhQ+WJEOLI+gvCDvYVk
VGTBdKXl6L08GjubQLZdXRKNDWjMcq0FlSXo0H0xkvdzX6+NW2tz//FZgGjDvNnES+7TWOO4HFl3
GVJ3IAPDztXIo9SiCKTqSJ232smYEo3/UZsaEyaqhXoZx+HbbVFoI/uYmxvGzjoZSVgXh1tLME31
zXYlS1hYBxEsdzXD6M8dFqyEauPaRq3ljC51nteMhEY/7KXi9ieKy1Xz/pR228D1dG/OBmIJc7cU
7lUG5ixKpjQyG5apc6488vMpxMbtSQ5D/GVvJNO8IO++vyCe7xRvmXuIsBfgMJSbscW24aXypsSU
V061fgI1SuCh7QXz0w44rvOfHBtpdzr7yjRhhW75dCaXBb3piSSKkRXOJt/YT1L6tE/d9DJLLcmg
tcytnWK1KKQ40VYamBMnZ8CHOM/7IunSvik7rLjUZgz21j91A97otjf8Lx4n+aN0S6mNBcjks22b
9wyWcRAAa4INTUkN9xNRNP5mM5OoKVX3S5fP3WX0UG/7Ze+ZbSQBfmM9Kr2jH5HJUPpFJyH81HnB
4IO9KM5TAWBJJh1a3pQx1qnZ5iTYN637t8IU1AT/9/CZnaqYL8EG2In70xza7Hsp6zdegcNWzqVS
n+0fHpXqgqgF3FqSVbQaLjo39XUhm5Bv+TKbYC128IEn/msMnYr8kWyfG00VNevLhHzVZ146tUMt
HtgkLQUEBBB4mQOVFTW3y+jv+lYPTgM1zssMwDFp2k1lBD2L6/CdMW72T3V+0mGTcVyaEManns2t
ReWDsNLWDyuqUOR0unQ7zDbwAc3qf/+iUe9MxMdmdeudjbL0/n2mdGAs9GEwR8hOff5+k7HBL3ar
hhZWrKbtEp+UMBAyH/oItPXVK3p+r9v4NGz+DuZgvWoNw6PTVmCmTRAVABSKsK/+Z4ABuEYeSQoc
/r+m4T1qriFowSiylWfXeTmTyysowDvNKvfsGpk0ZYXVKyfM/4n0YqYlJFJPWCfwZiiBOquyhaPd
+DBsoiJ1Gnz0p0Kw7iAwqQXCz15NA++G8YSPACQiviYgF0wGvLP/q+FmGLTS/RwXEgaAYmIMUevK
LTRQ+YfJlLj7ixktwAPGhWQFJ5Rt0BCY4oiLjGtEt4RgdYERkbkzsW45e0wf2scSSbrUoY2fiy0z
Ofc3JowoHOinqdvRCyvNRlO6TJ7KW3BnYZMMUdUgJ9gtI5C6zBS8qCAco3fZXYdka/A8ipJo8tgs
VYZSZv2wtWTeHQsYgG21sg2w8grFpPBZAvSuWzNK7cgyjPLMubaP6L2IYhpHsEQPxwn4vGZOk5TI
IeFioaruPq7W7BHn7kFWSPO+VC0HC+xPcLW2DyWQ+7GrrrHdWz5knJ4eKaW3BMA44vrp73r28Hbc
eMxjhoibwSXlifDN2vWgsfY9RK5C3Y+/FoSaumkdVkeO6ZXrfJveCLwhAmTghEzTx0o4k6UnbQtt
TkLIivxY5HZjLhbrTr7N2bBexdGQqsFwb4dJL70iuWNcb/BIadLC0ZHDS5HY2k+WPHMPURlixEjX
o+jv/p78KY3i7JK9WvXj9cMB4WyVK51aUI5DePuoon4tX11GpgvRRg+6RXEd38e8wkJoZyZ4p/R1
UpyqfiV6IwA5/Tn999YBYHuWhGD2k0DOab0eb4hWLe8vBmY80eU87v5QanedRlRTGLo3ZARFOZBx
5TnSC04hAnbJBl9dt+nodiZFnyMfSdMDAGimhQWm6WKsSnJiAG61RJyupRvOsOZKe0P05ec+G9Kl
UP6Soa3xTlqeC3pNZe0+yzjz5eITT4/wmZKeOmj3VmXOA/EKyQ4Q6FJUF7ML1jmIvOdB5znX5Itj
RM/67q4EEz/1S5yfna0KMtfizgcifFB9CXTWLpGLnAwbh4rLtSqMylXLiT411UEd+d6njmRdOGR0
G7ZxP/IkxEZ2VDC/PEnUioLHgOhqPVY8N1FPrlRe+IFtsDJnCBC0rOC3ubvfCImJkgppajCguE+L
uQ/5SKM5BFcRdfnKnOGHLSoJoXF0xUpthaJGye5WZfJA3HiAywa10OcrzSwbdb6GFk7FCnCencoy
qpHWqMfa4UYEi3ERhzSrEac4A8KEXZwyaQUV+zbgV1oyMTiSeE04jgNMWlQCkje3HuU2+HrOSCNp
6ze2yacRojOj4m8YcFIOkoY0NyvxCivWoJq8lTSHnlto/G3hzPl53CWBzHdntvrKO0vV0O28Ur6K
45Qumoz6knVmH/+cxYb6ffDP+VtuO6kcyXqpTLm6BU+RjS1yCOiGVnTTErKI6SiLiO6Q1tywf68p
mp8ZboeIS2ZWS48zmSJbmdtkhnMMuvvL11pQrtN787rvOid0UmLRkxEd2ElkTYlwP58Ldmaem1va
LNH8SKA3GxZVj7LUi4yR+7eIy7oZvY7/0m2v66NgjfpbbJ42GNChAqLTRFjm2/ElW6jGleDuPrwp
I1fFU7/vxaXSq/8wIcvszX7tnFU1UPTvln8xO7jztxCeL+94/aHxAPz2zsla0RGiuKT0En4gAsO1
jn7IblfT3avB4Ihn+yoQGxqjynT+nkQIWU1selAl2Ci0L0veVoMUt6qtfyOCWiAXo72aXC/0UNKD
prPTjVDCoONSYbzeCuOlgSWYfcH7CIKhLtJFKfjsGvvdyGqgByxcaXQVkUmk81+BmGsq26rnzWuV
tHyT/1PJTEt7G5W9Og9OGudKjJXO2igMC0GnGeGJjJjkZBcCZPp56I+66JBfbsPWyh9eih2SJzpy
9xiJ/nPOY4qinGclT3kN2oE7pBWw0W7Z3LYx2r9EyiuPo0xV+d9gqPowrPwQSnN+3m5YUhBRwklH
7BqfzGjZ7cxXhUpEoeRbj3H1nEnXEeqrUM52VBcUXg6zNKddEYzenD19ycjdTFPbNzg8xKKTH5EB
nBD2MSBfptyKX0gSRvZlGvv79ASsJ+2xbzNYgJGM+gn4BbnSodS5X2Zh+TPeuEVqgqZybCyBQ8Ha
voSZ03uj2pvHACFXwwaHtTZyKE/tnHB8INiBpWw9Gei6SyHtayGg4jAzWhHsHyv0QP+S5pRYxqaI
bOnsKgn4UqLg/Cb5kKPr1Mv7gztpaioyMBwrSSF7FE1EYCBbgFOc2yM3AbJ+/gc8zEyQmPqnUVeV
jFA7f731rnpQ7CpocDOHtbatQRm7a0NarRbIRKvLOqESBU6bAuJtk0Ff4VGlJd86ENw59K70yVLY
CJK+BbgsCESbVXAA44OUngTQdZW8dVqMm23AXxFrPc3hDNUsFZXRKM16ohJhJGDGhfy62WXLcXXG
SDDcwkZYcBWYl04AB1amHV9yjp/CsGRRKIb4kU/nDTg05LTnRob/86iDlK5NFAlPGTmYRAQUAjXG
gMEgsLHNcqtkWvyTvY21PMr25mKiqtWZO2OWeo9RI7jCcR1a6AnuQp9d5YUBFgb/WsL3izZICOwW
46bf7n+nOQZ139bqlubJQnbF3upDQRFGU3uCiviiG/Y3t3i8AMwB6QJy61FRDnFYWiyP2iU7XxPt
Qti/59oTNu0kiA94X4mwOecw0WsFLpakHn8tlBBnEPE11wa2OqXLSnsW0v1pZ6ezPZsUd9sb/XAu
sMdmtdLkNIZyS8xLOVaE+mlWQGHaD7ro67Fkb1cGJDMvxj6zoE86c3LDf1qcWqU5ACvJKYPCuirf
0Rng53HluooyVvoGzrwANnKF7ndxyHXUv+bCBUPjjnUBrp6exfe3ZZsivHqIFGxZ9FD2ItKrBDXR
RuUGZ1YNbXOJgvUpFb/YdslTDLDsj6PHZndkVEPZVthNTSRbCxA1CrGoU4uqMiDSXstj9VdRG1xN
m3z9PUlteggr6+CDUk+A7D+xi3QO7KdE5+Z97BnVqv2WzJSg4SlFUWVVXBZgXKF/zo3ohV4Lt9i/
lQIRV6RsSA2JlXf/qyvj6azU7Uwl3GhC/fC6bxYkzwawRdcN11/WPjS9UP/sp/C/IRScL67BvE4a
HFo4zynueJPflnu4680K5Ia0eBm74xW/c0Eb0oKY+wBn4medzoVa6QBkajmpB7pEnAwNV/7s61K5
Ib8S6x4lhZFrPnmCp3kfZSQj+2ZQsaG4f1TKYyyaBfLnAexxP1wsucSoaWT53l7P3qMdDpyxeH4o
H+ZzhSyX5Iz2ln/ShRlCcDcSRjIicNuc914ctMtuX7aMC+hukzF3TIRSZ2UXcFGDlAw3Sz12ueeV
yM91w/jHxogqC1iN7vg3Ujk0yQYEITRYrMm5VFnCYP5XI3zg5q+NQbE0m04HIvG+Kz4O57YH4NBF
r7VASqbIe2fuHhYBz4v+GksID08AuLvnNXEp/EO2chKDHo9j0CBTwEO5zW9i9xcN1VBF0rh/fNpA
s+tsZ8wqQdquU7+n7FAmD3UkLLPsdU0faU0DouZYaYei7m/vcV5JE2xts8SWjcnFhmCVkYC0qaa2
lxjHnx2gZuDg6kVKbd8xUUXyAHFBR9VrayDlPvvTfZ/CwjRsKmx+9BKkznkWluLsdsW7mADJPL9x
UmN/++d6pKpGCvKLHHYNERkugjVNoa95MasyjbaR0Q9XWWoJEIHZF9Yl7aY7yr3kqvt+P5KJ4663
gmdxln+IMCVwLfaUee5Zo1khXzd0Z/YaPntveeoZRswnIoxkedVFsnEeD8HRNROZ5coykcxMumaD
DcjN7klw9p0UUehiaXN5mvwn3G3VM4Ng34FVWTGvH2i9roiD5cKXO5RXRApBMTGan9VAfKiGFGWp
KjKNIVSEL9zomHRbOKhnrWv3QOlLFDk7izGc67laJe4pXaP3xC/2x4VEdw13h+pdoLc38Z8xupKg
SIQ6N4tP+igUe/GUCYdmAfw7eOU1VGpbw/j4PNu391gB147xRZWU8j9l4iWKaFICBfHqoup8yxB3
c1+K7Pqejdwmpzq3Ap8G7Vd7XrKt6f6RSyzSXMqsEmCAnM9Ss4fSjcTy3KTZcde2gHfKZI9/rwAf
BSUAhtYaJL3lOCYL4omBQ/ng1sfkZHNuGh64WqOByrakzOAPW3bx0nhICstWGigVbrzorZh0dYgp
2RA8DzHIkP1oJtSNU/Hr+KF3pCXq49WSKVgfeT+8IJ1qOnUq9GTLnQQ39ZtVpJFmbPYe36R5AqAP
i/tIcAfS7YKL8FVXStfIp2UI147UkAHqB3YtWl8huLosIrVCRlKiHyyykPtPECKJAggvo9hoe1BS
D6AB2pGgt7n8JgrJCbVMB66lJIlVA1w142E0XyV8nYrIdSUegXEXeBQB/zF4TCwhaQwvzFpRa2Cb
wn97GjDTDjIKeSrAAQI3YZx2TcuOffiDGYDNluzP5yv8Mf89/hhNXVr/hK3j2A/yzT2ytZUi8OhP
CtajVBmA4I6gLlhaio24Gs+HrfZSMnPP10bgBeRHjYnv56fSRGJc8xR/SYXPtLhiK5UbFc/GPGE8
GZcZe6k2b93F9oQcGDNCK/vP9QpW3VfeV/5pmEe0IfQ0HU/IvM/LRn3xBHTidT1hZcgd/FGQskZZ
OO0pF6q301q7GnqMj+HRtkfiDfcp4FHgdPJKQlGhn1vu9RGwS+RQ0B76jm/Pvw5NC+oNt8a0+EUn
XfkI8/Xk4BiFlBTVgJL15YK4x4tt2zNCodQj68rKCqvH8QusRgWqnFYa8lOplrL5ak9OD2gLUvYO
HnBACKt4UBi6KaXP1xtWVlqw/yMXrYnxmllu4/kGPjvZ0unuzugsToJMiZdlKHnOIpgs+m3EURGB
Zreo90FW/ry4aelBTcXYLhrBD2vbHYZs+mKx4YVfY6NXfhI8TOr95opZV8yz+faQjCjFHtde3Ygo
rEf8Cqc+OEYD5OJrh1T3kNLi6xd6B3V1bgUz92jLkQ/fKKkQi0dhd0e9S/Lj00Am70cZXs/jlMaV
/ovUCOzHfkRFmwdR8NfSg2WYcsCTgcTgI/bB5MUK2js0c4v6ZrOztgn5Q3DW6vzGt+p70u/iWpVM
d3EGsz/LN79OEChpeZcOFxfz+7nVOMMiPR6IaOoHCPFXpECiJr4geAsLCRgXrOQ5NonKV6RHZmLP
qfySmkFw/6ttwmi+W2zcAeR75J8XgJUwJ81DX1+RfjST1daE7eKFL8bCrbn6jy43coEsAi0uWxdt
NymiiwccADPXNnxFfUHOPZ34Eak7Foxkqidp+EULOXcb3YaYw0sB1eL1Z9wZmsJHFvxf0jytwJE7
ow8MwBsp+kDH14+xgzp6NNWx7ol+wl46SfGk7G6Vfwkrfe1+7lQZkMXOs6zJTSI2S3/jCJ+Dy45a
0G0C9JSkHMHwk4bPlrpmW/Dgs9xzDXGelnmjyAGTm55Pzt5l9TABsE+1fRNTBJXN4hphmvmA8A1P
BGDd7LCIPiQdL9jxLhfkBxMm3wOYFUKuu+rUCHMoEPYvnct4WC+cKBu/Ezq1vEQzlYxhQUz6Iq/q
vhFeJ8ferIa6dOguexxjdO+MMqzwmMapz45/+ZBPCcPlgaVtFhK0wxHHJ7o9KQApPyvAePUed3so
LZo/eo5RN4RqhdLFlp/0+QjS9ssosPQW/KnNtn3m1wqEX1bHuuNTpuq98qhuLzpuMQmAYK4GrPMc
QzBut0lc9q1jDW4rzxZ44Kq7FmKC94WfQbBQrHiQH/J8og5MVPdvXUJe7NHXvFF5nnaQ4oxHddYf
io7JeInZ0LvqQ6uAL1cMpv3CAfxPirordeZnMRk47ABSzMktsKhZvMC5vbRiHR8NlhZjepyVi2p/
tEwtmHnjBFPqZPMAnzgx34aiD+5UvrrDlEdutYm87ZQFXNv9OHozcAiPDQw9YFTwmxcbzdboqqUS
xqIG/MJs5PerDOLvt3pEs75uJxxqyGtcsMB9Jdhfn/L535BnXbLJkutRqRRpC74KXW2f0LAhmkPU
oFRzwdWO/RK1WsmTM1LJklh+5j0KPhovs/yN3nDLQewWQ1kVzQ8xe+hEMoQusiARSDeh9Qb/M4lR
TuCivsbas57VjDpNv9Xvi6Xa2jlw5BH9cmzEwmVdZY7PcjWJq8Wbe9WNklEdLWT6DeBqT+ozKFuz
ETgQG70YAPC5PX0+0uO1hm82Y9EhV5V3RmHtYp/fndPMWIAuvSd+Yu0k0J3E691mpNXcfc+SSslD
uj46jCJjJ/PCDgyw0obtcavC8RUmyhRpKkHpDdhAuZ7Efiv2xe1dO3rS8tdi29cXcQJA59cvWCLy
T7n1Ccbxrs34IXCfM5nyGqd85X5jTIXdhZVD0cdZ9e8TFWkwtTQJhbYOpOKS5qLH08FG81EqtP6u
DupOW4VVsXqclcsKGn7sSujgzUpok+4sHKa27HAgNNOY5z72eMbt06FHvtmdsVL3dI82Ue0PxnYe
7jjxyA+r+SUNvjiGXHv6cS+iGWoAYvwdTVDs05F49YGVhfdP88QGn3QVDkNNIVzKIcGq5ndq7BGO
hC2mp3xeMD7NqfobtwT5+LR9mF9NzJOuxUegY00sGSHDL9jDcSqaRDXPoI+72inGG9TW4sdzxhbl
1G2d8MnlV2kOmZFZRl3IVfVaK3Eh66T3uROd1CWVR1fCAMBMUozcUcoUOZ2YtlW10JsaF58u345T
Jl0b2uPW8ed55pnAvVOnfzY+oylqC/VFDMqaf5Oxl7h9VAWkfh39MkI7Gkfx4KLedkhoquoNETZn
8+fbTKXJvLN0YO8uw1NrCT8PoCO/e8V8PjM0MO+yfXrVuU9CFfNyjxO2KD2GnVO+cGMWiFxcT4M7
azJl4w/cGKzakzOoamPtbJY/qXoxl1rJkLb8IINy3xIEMW0HsLqE7Ep1cKSlEWvRBxg92fbj3FBK
bBFX0EgEkNlj3iDT0XKxn60tkrSpMAPX+hHkjLJFEjDIrdP5W3f0GR7pycLkYprwEcoNIvgI/H0I
yB3x0LbQ7V6EyOWKgjo4fes2OivZeHNEJ3bYjRgn2zqyix5b0lqnQ2djZZmJSSbZdhH0dauLiqEf
jCB2y6qiZBgDE8tCTHnAEWyyXCTFWjlzH+ubaYblIblP5PcHqwJqjl0vEchT5axaRMe+hAId40vE
FLbu0w1JTCz31Yu0foHYxvXnkfNoAL1+M/w1pW2xA/bAjP/pfK6rM6TgswkIqKGrqKDwPdi9DxKt
5OjFlndKtIDz8sxNT6el2W42CoMiwSmubGnM6A75g+xRH9vMJ/l9s2SjfCUCjTjhVCcrdfzhF83A
/lH7L/CsH16eljcrp10aiBMfWuuPr/wQ8yjO5ni8Lvz9rAr6Pv2quJQWlwk7C99k9qdSJKu4coDD
GFZUhtSFwnnXosuLijP4uE7rw6LhX7HIQGX1KCitXBwVw9sMT4RdTWkgGTeceYrspt0cLReEoNxR
5fVCZJXnaV4dyJ/soW4dqFzjeDq0ZhytI8BZUPlDT52vl5ObUipnLaqp8KH1hxobhHoTTC01sCSd
HcL+26h7nD0sdYoK6M2oBuPDgq376M+QbbxKYvHqjaWjqhXt6HNHvh4OsXS/IureJrAmndo9qKEk
XztkI75iEZbac7ZH9CISrgs74LJZqV/V8CYceUl/pb2kvQbt39nBWfhMgZhHLKy1QqOel4awcAlu
aSLJpea52coB52rW+G8cwjuPVLsnOcD4i8Y3wPjbTSy0rGCPk20VWpwFVkMErMjw2rg6t/O3AKln
VQObJnI2s0H0J2bW1etQrYTpKW1tJjIFQ5r8BV4yHKu8rFItZEqSoFztE/8+N79DasRbcc3GF6ao
7uUU0TzF3DWUTdjWeMzRuwgkfJ334IqbWX6c0E+LKInzyGv3AkhW5Dg7a8N45GplhoiOoLr3F1Or
0Mby5MQ8SyC1QQLfH1a5mC8byUl/FHQ2Cj4fH/3XrSUYjAHoEHMpBAz7xTKnsjn5TVsAE6ylTqZE
pAK0wwGUVVx/JamNNQxAcmUUg+wPKcL8u9N7IdZNCuN5c16zjRPRawyJz86CXA+sS390wXXTIN52
niSdMmK45+77D/tyz7ahAd3g9BkFJhCtmyIWPItosmgFxlmHs4vDaHCiNw5XEId5/p0DTMLU5DH0
mZKC5labTT5EiXl9TYztJ9I2qAEF0JKhwDHhn413m7hZLyTXUqVWakINJ5SdfOW7OyXL8VEAf3zj
z3RBZBiA3gsOLxQJO1JTYEzO3+GneqWzUc7ugEZj6VN5f1ln0pweb2SVJg7rkHpBtlLWKG+JQE5e
ITuQJu8Ig3U6wYgqJgN2c3yhl+1uusr1wDMtjxb9lWIZNa1zK/3Aqh33v0+IqWTsp9elYwd1ZFJL
Hng5i3fs2zM9YiI48zHP7gzCMQDLyTplNNd9VIH/qgnIL31sHcJDbuWt/hO7vVzkCBC3umgWbQqr
Zkxfym4RQCR98Y0R2TpF1pFcwHqR3qimeYkxgX8WyR7ahByyePtIxpgSihaq6CxtwkwZacoZuqTx
KRdeX0oET6Fz5sLcVAybMCi0pM1HG9Dq9rlQSn8uGyvTdKn93ZY7VDJRK3z2JVddZb8n9MIXGqXq
JKbmXtgP3+FFKm5PVBC1oaoSKZcSqzJ/T/CFTOYh66RGIXkd1uc8vN0Vbvju3c4n+u9PCF2as653
HiLVDZ1VeWluloXBBdPq5RRJBevIotHh3mmQD+FioyFKDqKQqfzAB5FlYsCIAWrqmzz80YhS3+tb
n0eWv6r83FL1a9Akd6voWiZPuUEkStsDILsCprIBZKLCN1TcuQmmaDTGrpulISVpdNKhr5x1wJka
7Sg6WFvYhT4cvxgxXfVLc0X+iam+oZGIPxryFQmIfTRcXpkTwOkucJ3t5I/dz9ZmDGgf3yRverjD
cyiAOKrD2w1tMXPZ7Vhi2LdzA2LigO5ggOcIOglTBe4w/i0zteHSUVMm6Z5UFvcMCzzx5J1+fvXn
cSJTv3ioO4ldj8uCzgiRa54e3Wsg+gzgUm88583OUbE+OmjVjpKoPoL6J7flIsZ7PrySw6wS/1R/
6IbT9KIoDvTFVoXS6qF6reLrr3Bz+SUpzskH4m3q8sd7Fb4pA4RMSF6Baxtm1sl3lMdZni/jmhmJ
0OM7jGxA+KfwzPMULYdV12FwSlu+aHgVJ8voTq1XFjDrFW2ijwmXcPGBuZkzl/whiOgPR26dUfWl
7V58e+JMNbkXV8kClooS9x1ZoRhMuPpinpKa6Ez0WawiN6IdlrQa3iGSoyM9muRJ6SBVZTW0fBn+
d1ntjpo3/+aMfYr/4n4+OAsvb1bhc3XTHaKVqM0avkZcDNb/bTj0IngQINh9EnGSn3aH0i4r37gr
qaxMu5bHri6yolXOqCwCxCUvENJ2d3ucfpoAYbe3uHES82ws6ruFq6qHICl5zH6bT0NTZhrwjC2R
Dl0gfPfZ25SZgDlm6QrzqbGDoRX2nz+rHfXryIYkB+S+jEKVLtiTYlSpMnA5R0MyJeyZyX7ldiTz
ErUNbX7tAtuxVbyjPYEUESTlBcYzEiN5jF66DcwSqBp/QKaXqGyQ4QNYR/izAmeONZsM3qYw07XA
yVgQuNdDJfepx+IIu+WD1hSglytScuYn8LzHxqcjGbZHwyMcSohnvNZL60yswznqWEe9l4r+2nKd
4oHToVSoNqNx/qxtsi0+4tVaz7ByKp13vEh+LR3rlbCPFk2+yfpK7CxY0mmU1sqgZOSf+grwzQol
iBAwbLvmZ1utg23+Sop6XCFYMgCOFQrBprNIK/eiZF4MFBMFNvfnwQQwYrVg5DxHQotjuwKusxlT
MDKieUR9PUsYIa9KPepXScxZReGiPITtv56HlTIWfKByWbtMtttjIcc7AnztRXbsXR7/f4yryMIs
8YB7Ob7Sh4Sx3jDz6lRg7GFkx2qo9esMYzKYgNf9e9XFd/Cu1Uu6qFmu4UBI0hAZEZ07mH4ydlAE
LdUfa2V+g+tlXTXH64pL+YfhU3LmDQ1ZxaJAVFqs9IICXTCz2RkCWf4kV71f7Y40WcXVfMgpyvnw
+Jnu53MKCNYdNBH3Jp9TfutXcD5XmlUHvSXz3N4CvbzcWdzVW367QOE+3FsIBnZ7u1zbncvTDgpn
1uK3Cm08FW/Jl+JM7GMx4Zyg4UbbyoR5+4R72YKF8Gs25syd9Yna+Phl4ZIq83TCRiFgzk6FHfBU
7pgKNn1f1amb2wv0bO5Io2IZNYSa4Eb2b42GZFEaWuWnBX0G0pFi+PymsiUXZluLmyHgcM0CtIIQ
mK6q8ftIfhTP6T7uopY8AiS1pi9oiPcYq/rAyB6XeKbcE3nzVXXXS9Q6koLQruBn7+n4XxZJfzXe
R9pFgeP9tMPBvpnlEAynaFke7ymSoINYwtN7voA8haqA42Vwzl5Q+6YI3w6K0WNUb9WkwW1bksPr
j96pNQGpz4qQzO/sRSPMikkAqnDAn480/o/m5Zw5yWSGkLwd7VRTVbKKgRWjp4yQ92OkYgyfO1V4
lH2V02Q4NvyvszVgIav6OonILSzh9ipjHMkXF0ojiSuJjOvLH+qgSHB2F2jX+Dozi6OqQl4Fv1lz
HMKVE7LpVfXzr0scvnIGeW0p+hrr2Oibp2WbC0qoQFTcDS27/GLh/Gnglcy5UlOus+YXPTOUJwnM
f3vBdg6khEHTwuoFmD0E6dey/jBJ9pPQPKcpvrDvp/cKRF9A9Jvw3e/GiolgC99d5t4NYxucxhLW
feFbqeV//kxWXXOG1Z6Y1sBuKobpI/MZLXwDkfi5zouKD5rssZDs4323ixziOK2AYhKV0nUZgYy2
lJi2Rog931wQNFDnhJPkaxjia8jt7ABIXyevKDbBy6/BQrIgKTemVnWd7okSdFQPsHoKIuQl9xC3
t+6v6BcKgoIUd66jSKn/uWiVWaaFpBG+dHX8pNHPP+2pf9mooZTq8zD1dJ8POpaUc7QibThUW7pJ
sRLWKBDfCN4auw5HEPiXxfVaXRBAAye2MzEZDn4pTSAvE2QfXUWX+vonIj9oOT483jqld2gY8o1E
5yFR7lJJMQDjn4/LxTAXKEZ7t3fEoe3Yv+KX4AxFBDT6f6Cg1EM1BMQLmN1cc7voPX1u+eojQniv
Gu+OoLpBYejcU0rjtz+BUwj/eU1bLpqYspaOdp1CJjd0b5UgV3UnjQkqDWpKfZhhkuSqbRS1+Z7T
xrZbjx7iIHnATmxCxEJs1lPuyh+BN6NygYplVrKHzUD/nxmvCg0S1qg1DfBk1ERcCUBUlY+P9/E1
0Tm8Hz7VZczCX/W+OFvnahGMSls6b0pujJJkWTZogOBLsBgxOJj/VdMiEHBEB1Mq7xfu/l/+nyVF
juhyhScMYYQXwRaIvkZMb86Ya41H7p6YLdF+q41Wv256E95jhi1cLQNoP/nVfALph7LqiAYQp+Ik
nd4XnBTo8iY9NEq+99y3ALhYxtEILZ0Gpq1IGKQb95zov50HM9AyE6KpTjDOtKmT0CzhX7A0woeu
okKD4pokhBt9vhvI6nH/r+W1blDp6mePCtzyR9PxiykhGFxuEVVcQF/K+ISwVnSkK8ZMEyfbeIPC
SlXg+bXvVIhsDez1XtqbUlphrISc+Ydn1cvoN37wNYHUZgVqls7owhOGa0ThJLbkQ+0w5ZQ9T32y
KMilYCxhOak2ypRPuqG0GbzQJsEvyzJUY6/KgWs1Cn+gSOnbWSTOjyG8YhdS+dtK9KN2WxCeeXMI
3cZgsQQNjMd9AH+fBwqZSR7P64HhpvWCeT1J7ZpHIe3jPryDOh4Y9ZGIPpCw2DdF34o04DobobS4
JeL/C3HN5LPNvhfi+RzwNgl8UHdJb8rDzna79wA6aYIY/1MvBVKqmQUZwhedISbjGhydi3cz0d02
JF+shIa7dsxxnbZ9IYOvaepngolSWYP18o4qrrn0Z1f1DvDfmpiwl4+MVtm3JB8nmsrByxsl//kT
T5mLgQmd6z9hVvlP/bWs4xuIc+QuBbEhOXmCrXUE2BVvXFoofMLSn8q/h+qoU3l2qGefbTLSHPPQ
p1qvWYp9AONjE2YR0p+GFGJqIpw8FcKYW/EMIifPADnCLzhf+s/gIP2VdHB8WGWwvwM3KQ6nJSu3
+UrSo27l4u42OEO/8hk5MSH/kSGH+Kpn2XbIltui67rqlOBJTQsFVO3GGlRwHdLNTFC5gr0QwxRN
Pph5fG5fWZmFVIzGHqaopptwGX76rcq6ACGWO/mAAfJWi8RsS330vntC9hJSP45qptBsSx/EYHn4
+XT8hrpjs2eAJB+f3rAgPCjLUEnGB2bS6K32lkCyqYB71tDiY/Nxi6uMf6qt9QqgdpM9gdhrVIJk
COl4qsk3yjfiJoda1E1LLgnhnBUbn47KsS5aTEcrVF462KQ3PYuCkmstzE5D+wY17YnWhCadRu5z
+Yw3JypXJS7Io56t5re+K2tNunon4LbtYYiLmRz6VQUHbIUCdO2tdq5RLl1Bl+sEUS9NiFLM8Ui+
SOStKMQBS7+PXmMpS1pht+3UjvQ/ATrlzzEH8nRNlkc2h2giAiEGNzGGU06t6w7YnK0y8Lia5dKe
+92zvdje9ih15Mck/U6xfG5Mauv78SHs2wE3aCrjrhgJ8Fro3NGhMGKpiNJu7GGP+72a8QZaB0SN
SLYjpZADUdb/2hCZMvH9h7/+Vit+yw9ETQglrQRPhicByITDTzYeYgzb+1Zb3jZfrfHb88nGRufg
HS9XKeAYC5JVTEq3D5B5I9ryUjdikN1PS4Kl8OrXi5TAHMiPYt7H9OwOveWWsFW55MaZqy9fqJKH
PaUitYs6gU6xPzF7VxMSLR6MRIACseJpFdfD8WVaaqV91KAf2z35RfrkrfZQ9fbzjzEuo+jgPqXJ
cUxI4omwtp7VD+To82YFir5zVkUI9W6hKsnBBXipvy35PmKQuoKRO7LLw07X90vwjKoDcbvTokLB
A4s1jLSKmAUqPDPnRE5k67+6xz4q8uedc08KfgQ+smpuha15hy38jlucsxyVh1WYjkve20uKWYKB
ka3lR0yMypLPRqpDkv5NlvrX/MpXKl6E2hzjjbBwougLNUqdghbTwRON5ibxk/tQjev1ydpDqGKG
TBJEWWMWPxe0r0qO1pfaXWC+OSME0nHZFoE3Ogih3tGRJW4l0uiLtRz0OyaViKEfoi8bmyCFsbzp
1+L1Iz+tbrwX4BNT4FisQ3vbR51KVOwYOO0s5xbgzll8w/8EBjGS05jA2Wc6lITFWJdKPo9yZuqu
oXY1zoWSaOAejndZP2EkXA6utows2TmtiV1aXD0SHBxw7x01usz3mkICn+tYM/1VFaG4bUN/MPhJ
BGuyhbZ3/FYsuE5MboMHgHy1+nsSGLTV3N/zi642dnqxLDQHt6JEb0jV26PuK3lhKzab5uDI4eGy
qcDmKIY+Sajyc6P3a99rMwby/Sf1vgS2cyO/dQPsc5SBmAYnHdxBxq+BqKijP/4rwV1uMA654Q0b
VjxXrmE5XZ8zp9YvtGBGkqAD8XPA5tr/aAo2PDY0JQNL7UUdhXMAhd9lSnF7Aly2aq/lLXO41yzc
z61Vw9PwWILO0MMCy/adi7hSQRwH+0ii8vMWfqTbP90spN8BTKSsd4DLt+zaaKKNJilJAedWP06v
4qj0wEpPW+vy80/qoL+PGD8DZOhzxMYi2jlCCF/QnxY3PuPRD4BUw1eAe/+ov8qxCLKTMD2A5QD2
v/JIEoPlEv3S0+m1DeMcJNWlJBI+GprDj5sn3kwW42u0+oCufAB5Fc12MvofGOmqsR7oGYUNbDHm
d0GWmKZlpYd64Yw75QMVuS+5xtMIzipiAvrSAO62JGJGgd9ETuHKdEKSiZwXW3Ezo14WyOKZ5SKY
DO2PL+sW/OmUL7GfKi2Sv6zFG+iPCsn9LuCdUGRhIiweuDIR3p8ZLn2n4lQkd/su9b2GkrFfcAqS
v2jpfjkGGXa6wpNySkro8Qy/GcmBjnKF5t4waXFRNaY7jlq06MvekqUHmJoaS4DWiYeZKezwhBxv
C6+SyEeY4rcs6yKXErkDNzzkFOnZAMhmnFZ3kqPJRK/xMwOBV5Wy4JHRi2X61hLXKwZsokHK+vUL
HWqOdd0KRsL5PsVUbc9eYtpFGo8utuaE+K8HdgQ5kNasfMqEx/cEraab45mnYt/ZG6/wziF33woR
LNoOEJc9KTaA3dFEpZDIwgDKgUODxm8HGr/VK7y5/rngDLHQHpvukBVehLixvp6Cw1Qa072f0bWB
6s4ZLMUbowyJKKHidgd181Fv96eQ+I+kmT0DBO9uIGB1FYx7PIxv8Rep7ykRwyRUog0FRoi5FARL
Udl5JaGcirEMoeXxrfS+ZsUVkDZUllqfdqb6Dj8CTl8kDHGGmqqL5N5ECeA9FX55gK6fFhOSPcaZ
26tLxQZ93AtQbDeQfpcAkSclXYrK8EJh0a3y3+dNM8xrwaskB7HyhSD5XxiJ+bTHKcb50pGvw3P8
S7wmf2qYnmhpjhJMAD/DnAF0tBsdTZPqq7u0RoAvksG4Gn5RrQyZkooGvAc9dZUJ95Afa7aFGAzH
G2+z499PK5rnqDnsajrko8jmY0kSDqDGsoXIRr1X0FRQSsMmylVd2qwTx/Q04uVrgIKSvj5LPyt+
wlmkDZPnRgYZiUhLONvUng1WDNNpiJXP/mrrhGSKMuBApKSOj1U/wgPkKlgg5157MnJUx3RQYwx5
0Waqr2uwDhRoCunC5jgq7D4omcqII3cccD6D/0fq9iwZ2Hk8X4PPUXG1dQxfcZmwVMpXEcKUlhJw
+QlIbSHIFfEhy7m2Qn3N7BaoXhDTzC1qcHCOC1ZExgvFPA9VTkN3Eg89qFUoxxK5LkQ1jK+U8ZFJ
joA6PhjTCXYOdRg5BmB/axC/j7cNlbSvolGPFY4TqVkMjEvlZEDUEgscx9uzelNAzrAG+cosCnW+
atUUTHgJn3dF4tfK+NbetCNc7+YPmqqiDjGBb3TPGGITmr0YCDTcq/IXNefBDGVHdGcO8S4ywVtl
/l/c//x2bablpgEljO83JYIIdXMi5iHxOuUb+rBQhtPc2dgzXAzsh6//DHsUn8AjTgevNy8b4whK
1qhRK4syU6zQq6WKSXdOz72avykvdnj/v/1Oz7b+J1pcJ2GZWkf+u7ZG2/xxuo7lOa4wcJ2Wu7h2
93u8LeBHvzhY2g2fT9Cul1dmoN7eBcql5dq56k+cxG2Yu+9DoUC1617JhO1G3RPljUKRNABnDLJ2
8YKPMhTs09tdve/SF5GpUiP5qM68S/l6+sKPLSQr/xSkSyt7V4bNSyoIJc6J+zQuMXKYKF5KyXyv
DGIXSYkj7KxK4kHncIcNclpQ1x7iZy+rQAEkKDpYhSmMuBUIg5+79/h3X2zGti6F4kdo5Qzc/c93
eqvF+r9kEgNwQ8Mfp+jdEY9ITzjSqIcr7NxPKadvTyYLaSQOMCV7VTlwJXnF9M+JDmfJZivxNvjc
U/lsWpPpQoq503zXi1MY1nCMIGhoY/4wgrbce4gCMZzJhZM4CWyFP6mbZrHmBw7QWHBvTMXm7VGW
e+9qBKWAvke2qriqz0uj2fTqgLI3bWqByoGcc2YiA8DWLdabob63JlBmcj4Gsdgn4BvwFH+IJdWP
ELq1FIGTVCNXLEXmXs8gb2jWPAvR6YC0LZdTV+peyaZ2dIBCSF3XHaemXfVCTBJE6a1NeyZAyszq
9j6dAgWLXfcSHi7nDoN4inE9yHJRY8IwGpjVVUjAmQ0OXIAA6DA/4eWCOhCb+4hhCYFuAgTYuhT5
ozItDaoRrKwn6fa93Gmyxn4Tt0kxegnq/obfA+YfiP1VU4JL5xkKeleLAIkJWKgTlxAwlgZAP5Rr
erN3jDy7cGwDLs5TUoHsk0VqvI6OOZ7Ee4yv8agXmoFQoLrkRAw9cGkcEyG0u2e1cKjENd9jbChA
cUPFe3t1iHXZ9Ge1+iTydg6n48mpN0amUT2Tl2zUQEzi9ye2swCW6j4lcmioCr8uf/h+9+5hGQyb
Ke++uYqLXZ/g41IDFJuFwpbhM2xTs/6fFBr7ipoSgsSjmPu8uO8mpsYYM2bc38m7kzL6p8RyLQw+
bt7zf9RZS08lqjrRaTAuxZdXQOUKNc/cm+RwBbDvAi6r2DR3uwX/2RiFyNTe67azaOrFyHmuF36A
LUh7U3xtH1+KVzjfXtKiFCEOsKdA3lmussXXcodaSyhcSjnuQp3thQ9WGnQ22af5M1+HvnnZYO2V
gNEVXH3wnLmZAKCs34YBg3G4YRkUvv4fAVeKqnGqh7huOsZ4pt3ttwxAFiRy3UgyRdrKmFZYabCv
W6QkAArA1PGZ2oQ07aliukwdin/QMdr+YbiZLW/nA19g0gvQ9umzUyYrsx1MzdXhrE3rqm6AhU8a
xptHoBkZ7IuE237nhT/ooq6yl5BLMzHINVHtiqiuP/jOgpb3XpiKikV9qwVwvwq1TVFeCI2DxiJ5
20b582hv1OfHS1FP4K6G76CFpBVtCziLHV3ssNq4yosTQjNwh7y22d7ZCwPn+kZZpnQz3CRRjvtr
LjQihnfPVdMCAJU+/CElkjqSxMLpoSh7O6vP+OXZRI8YSR8+tTE3oeZarG+gQTNMLvYtvb72tyVT
/iD6+yzKtkXf7ela+CZQ5TTw5fhiRPZQZbzKUJbV+JjiKJ/hvSWE4hc5dc2EnpkvAOfWqannz1N+
+nkyM1NNthPLpYKPDPOapo45Mg+g7/ihd3HY6BjibZOe6P7gi+afF3pzPYUaLFxZ7joV1gD2C1FS
XfpsKTM2nrjAM6xaX7bQFCdGSPxSuDpARRDB1OPdDxomnqfoTAMZIsddTwzKiA19214Zdw5qF6BI
1q4spbo22DdUH9KS8kKSd/qlkkPRijjh42AMxo0CxY3rVXbZUky/L9clj7zaoo/QAD5y7OK3n8mj
4nPfF19eUUyjbhtK1GVDwGDeVBpeqStkxtIfL9RRfXWLvke9w7xbva0Hx3IOTbIQyeeQ6TbWHL6D
TsfGfuCgaGb/mAwm4qugJwB5tnLEKlPzSvGXIU6HfQaSYw9Y1zXzj6CiA6ZwMAs/1EBSZPnR3N7G
CfpHfabtGNMnRdLnZij1WMrzLidoyP25681YqsB2mo5Yr9UqwBjZRVdfOMKM9VOTyTCRVTks261x
Klqrm5QCC7Dj/FJelCdXELeSSZt6YnD5+vVidiKkAfI9/etsuZqgteezGC5it9VNjYsihe2XcNDv
SaPa88o+DLzbmYw+hor11RXXOG6SP0VIMOnQ+cNYuymWOqjXfQ3kl01VYGX/fUwQXd1mgBN4Fh53
jD8Y9jLxZcRMSAVDbwSARgCMuCNmI4lLUmHF34GaFCV5+XFRqm+FyaA/eK/7+CTs8dgfcNC5Yg4o
3ECTUDekbluVw7Sd6I2aqkYb0yErtvH4gnjKPZkD4SyiDSqgzgSjVYh2MoMXkaStrtM0xlcsEH66
iugeXvyloiOk3TvNlAIo4mblw94UO8H+gPx6kie1ynUtmCJp1AMiitwvZ6Itp0Nm3DNxbVR1jJ9N
+M/yGWlBZM9+Wi1wvyKCo7XcC2pBHWgorUW46m3PwWuXXfP52rYIR/mKu/g1FqWxWKcphBeHRfWO
6dY7TlIDJVAjIChErn7hsTlzM/LPt8vxJ0l1pHANct7NAxAT+ryWgtrpz/7KS9px11yae73v0DhT
mMaQTs0ZAGR8qpj0S6a1bn4r3Pk5Vb3vGAL2dA1JG4bdcPplHIoZ5Hx4sYUjTCceyMb9B4G80oBd
rwnYr1BkPHNVidh/vAcif2+TzYy0z9K+uClK17j4Ss1qAeY32TKB9Za6z65FenyyCPtFqvoM/bKk
pmToOhgQ1DvAjfW7hAodakK0AabI+J7gbnFccuyg/goPKZ6PakGvRmnJSK1TNAIuS96c5KseAZMv
xHUoy956le/MAqg2Oc6nBCaTjbvohRvZsuSHDXRAKkLoavQUsU2LeeBwdLaiMeLfZ4EPN05Hivc2
oXUBPLQrSgFEiBxz9au08Z3x2swSQuzetPagHbdATBGaXzqkQ2rmkhVNH70AxQPrYZkxM0s6vYK4
WYPKLVdlYP6KhmzibqDvSal26drvfZyCb9GM0jkTUc70UfzEFj2qG94xfsldMONt+7l3wLVTy1a6
PtoyVzQIcEcR/zo6/e+4wAVstIEVgYIlf8b0tqiuTwp1bivRelYNkCOKaftw6KfeYhTa45MPpnek
tW+v4UMoIoDxKU9K9NNCJ9859Fk0ZabBUvoFqmG3e7d9FA80ArSmn3ZH1mE2XwGNnlJx/R6r0Vlv
TOVG5Jym7UBOBU/aUf5xLpIbSnGMrnfat2y0h7CqKZ2p8JCEak55if8uGTWTLtdkAMTV+J/mKZrz
IgdHqRbN34k3I5mjwGxdobvG9jCGC6ZQR29NuA+oBe/GYjCh0/tVaymbmnEFF2oiPTddNB6SGeGA
4CcdoOOFOjJ5G+k13WpndSmBLPZL0IefcBnc9O+j9TzYZ3CiGUt7ENFVsDFtoK0LtzhXpC4mNU3x
flT5Ml/YmfQ4iOvlcLlL08XEt0BdXkZZGiV2J0BV73i5AKgNNgcudjYxrsIZr6kgrFreOfnropwt
e9UvHwrY9DbhAnU2QBBjVdjuuhcMZALPq51PBEHjN1Tf6NZDiSqUM9vIkzd9064lwA3w6TXRckQm
nzp8NmQ3/pWSea/7BpAfM+nNwuhdSZKtJueK3FF4Sf7iI81j+ky7Edtp/9pO9lmYmSTuTXxCQQJh
AjOknxNjUtdNOLTJdCWbx8c6BHP/GhmR/R53syGNHkYh4vBnaWioJ4cM9zYJkC04DbNioAR9GHyG
9z28dOoLwhT89ojYYLxpIjPPAp0SeYyoZhK5Bohtu8nuwqXE4lxyUQL6SgG29YJ1oa2cKmn9sA5M
dk9wXTbRXuK3Grhf40bdrQaODPEuGbdj4pXKUK78+CD4Yf+7HJkMmze+bJFNDVMPHIIKdDsw0GKa
GeodS0NApil0k41pNfYp7AKhLcz/jcczOtSqKmnKCu8b0QtgUBmG7M1EfU+2YjbHVRMX7E9ez1/d
4gQ+UcPxJS3Z5JjCWHFWGzuRRk6XAi0N2+90EvoTyosA/ZtUuIJ/qeAWCIQ3lDsDTMKIUhcVDcDC
JBjwulJ5U+Eyjc9qtEW2hJq773QfF9n2HxnSN5CHrZ3/vO4sn9DnUyoqIFVx6W60OkcJMF22m2rp
kmLHgkcdH4qPHtKmU8m0/OWepcQ60VVoFfVabSrZzoZO/dTQzepMikMVBPlq964t2RJow3/NeHfD
uivDXbzo6oFc+lFCpwddreu4wW3hHkxXSST3d4ziRMHQFLNXPnc61zXf+PS5/iWzwNXd5RgguDdx
M+EWnZppCeqEkpSTWXn/1S/4KXhvk7909Wrc9UqmBfcSDHXcogp1YotmN109s4mCNWUjQts+uHoF
qXMS1sMuIhxFIrrni9OyDroRs04RzgtrWrLZnXi0rRsxNp54tU9Nlvzram6XCur5Z0/9TaHA50cj
AMW1jzKB1YAV2wBidpmc422yHUR3hDe8YwdBIOX8Ka6D6VoLU5HpXVlKI+VEshI+EklNlh4uav95
yLeOE4HyvOLISnK4/HnK09CNHNdAL4tlpQ0sTfA9arJ1c6Nr48Kg9iOpWn1nwTPRftiKOM3XtWdn
nTSVcVP8DxhbuS0DJ7YjylvAvveXkly44bVnxDuOjmFXPGE9rDIp5VFWa8D2Sqly0puyP3CQS1dE
MPCmXyCSgrWiR7CVybGz1wUoVLgSJDEQ2Rwn7gXb9evnnrPP3IdjJtvsKdygZ65a7Kj/X1xubxWR
opWJEAVeSXLrJSXb80JK7gExhMmJy9zOoAf7iOLxHO3yueE78d6w/GY6cdh/RQfQgdyuEhk3oWGl
mfx5sjyGebqcvF1tYn0YVXHvqwi/nSuXj7nGNTaRYvA148hltR9aBZRWuCZBWJhh3cCUeS47kMjl
qOy3I/8W37jBPbjMvXFNjHpwse1x67EbnVPaVImo/tSzuYjzSCZJ0EEF7Y74XOineRm3gE8rLHo5
Fj1y4htIoNb6Cf68S58cpi9dyF7CvOkzkNgY7MxQBjUaSyMA827cik/DbfX2W4f/sWVt9r/M/Un1
6GtYNQZ+bYqrV7x64WhqwQM4uzDqgL/HcNvcjtt5jY6qqaUsDWbjN6RMKmGGBYG/koTi8Q7VHHRa
eLBBZbP349Z4xFu4OJunisyzHCLDxo3muK6x+BaXHi6Qhoi6kvJN9GCzfGsnTNIsM6G9QEInoTbq
dNHgnuh8HEEdKfBR91qkpkqzX5Uvhw/drmVCY19+WO2rIIP4cmo2mpWb5lKGIFOHYqwpUdueEuC3
pnUbjhbOKuZXhve0QzKBEURBvlmMU9yrFtAQsVNeA8WyWkitLeo3VIpl33AbB9cz5vtkX3W7OSNg
GEdb5qbZ6E8CXKfooXLoIoJ7h09VnI2EY302WAjyy1WnCfNkNsoEhZv/7dDfZZFR1LnMLgRCW5ww
rk1bvuFc5D8/aEXz8v887pHxFdpERfceleZoLOUAfDVB2A3lifYPJJKMKm98RMEX9abwjQPpukxA
eLxHor+FyvxqjlEthHfvhiRmh4SZ2syG+OpgUWMZRoV03pWx0rzdNbAowvewXeJFmWc1IIPR1nag
9pYhJ1BjhQCICjcM1vbzCy+9BswtKGrVi8S5d3LFndh/efDP/AP7xN5tWZ5FnYLdIs5bmixk3G98
CV6OFmmCZP9KHmcEnIuh+QZPKX+7wqEdjNiUU3xiQjBBHu2MF4glncItpQ9JhYzdtTqeVWsSLVcw
abAsodAAA06tBTAvlJg6yUr7ckPDLmfSQXPLbC2+79MOrxZ3UjTACzipUYl/AMp4IXmgKvGBV5aa
WOHgsGSDZU9U5/TZ3r8GdE41dr7asv4XAgA8fWiSzyo13m/PmbXoG/jLwXIA9iy/gapiOIcsSuXU
is3xlFqFy8MB99iu0DY6YOJcN4GEcyhJGbfRHTjTFsq4Jztjo25cE4byutmvL+JuK2HIULQ26TTe
5qOG+7SgMtHUmCGlEeOsUI6Nti4W4V8PUY4mQvdG1SLWgALOGw2ETcTFhBjMKwGILLh0eJ9RrnjU
6X0RV11JJhONiN8SwIimfgsU88mfFm5XInh+JniUxz1ZcOs+L91eJ8140IUw7UZ7mXSCFVrSXHY/
6aCUsSuBVbPsJaSksn6vRqZpOBUpn78ASp7bV8DJ2OlAFxTRe1T+75P1xdS6LD/uZaLMk/HawzPw
URapDCyg0bvHgewKUkzOr1coyQvXEE3gx7fnHREHPy+4ygnHgemerUlj2QxATQuiXLrg3C28nQFs
DapRzIyZov5YTzLkAgSwynNErtq9ySMvvWGaoNHh4rtoB5E1HScuzfVQjHt0HiRGV2LeRxwPLi8r
/U/Q//48hOOTvyRlUtnLRSck1DCOIxJndhr9JFGoOIOuknW4x+LvNWTqNDA8IO5W1MlVbweIrpMv
Oxuw8vorptK95K+uskgx9Tf3pibixC/HujZRzeoIRzVP5M2lT1G2ByBgOVI5OjGprClEbqJ6qDyv
fAzEYOsrdXLj8f+4jGzatl7SUqb51AAhBhIwvFj0MEdhmSCuKsIZZ8JYzuQlgGil5z6kg4wlLa5H
9Ao4DSXFfIVx2U9bixNVltrMRoKKZscXidtvi/fji26Ab3dy5frDhuOD/NxVOVR7qF79Mq3fJA+/
DglkYcoowLAVvFmcG2ix4JDocCzlTp9GIPVu/Uahea4bUqYY4YR2yMayMm0OKjZN1dA00Y4poXJZ
bYNYi7VSLd2Gv7ZR0qTcDFOQ2nvPJkWhdykFlQo06tRCdmq1NwUKWhLVgWrJwVW8gHNVo1qKUtrv
eDouHdBD4VwwOBvacrVz2T7dBp8QbZfYOZlGdiZBZUWkxk5U6v9ZoqJPAFT34UglFzO1azvNU8OM
h+mf26pCrjjooUD1aElYuGTQeayyyf7swh9qsRm4u4j//+1YmM2UB7kR2GOAX41f76m7sl8Lyqf4
eOdY+3OtX4j2tIFKeNt9WbJ3ddpToDM6YVV9IOtIZD1WBoyoPzxIjMPubaHZnCJ0DXo+KKpyInKm
HIKqSHFezLbnfDDy+I31Rxa+Gd+s7ITlO1L9zSB2MvIq3m0nZ50q6m2TC6HYSoAKAowXY+pj/Tg5
jlNigOabQu1ZtiC+oRUKZXLQeDAvW2c2CDB2ltO6flx1mwUP7Eaek5QceVlzKK3Z02i26xLB2xNP
+foQp5k6GWDuj0sG/B+Yl2n/gWv0xpZ+5tn/ehoKLfzZSSD/fkIxRIaxqs7xxEqythu2RUyWB2Kx
OhArUFdcsTsCxtdkIEcUo9V3JVeOAA+89B8ItrQV+q/XpNdkBeBDuiP9mAa7jS8MsUC6qG7fGZvg
bXvEts8a7gTTjvfxIpZehOPD7bUiwbwjwo6YWo77rxsTv0YYaXCFw3nCITULOA6n1824x/40sACV
GjfVrERLm8lNGugOjy9dFkpihXAGd1vnvXSIzvqXadG/lcmH+IKoKiwdtpDyJV0M2RgeR2qh7INn
DMRH3ildHcdAKvmkTlVXxm4SzYECZxgfPjFOPDoFlb0FHqw2TrTBQ580rq4VFIHWoHgY2Mj7peFb
OMr3Ee+E0lmT24H6XkrQoUuYOini8mwigmHVf20onUlnb4PJaRlpkd0h8jYE3dbx2/FDCfdpk1pp
WAtBsfrtY36BPeZ9FyLy3cxmWFltILWsCn9Ihw5AcWUyAVYMao4kw95MgU3Ap+ZUbk6vHpWDCGmu
BzBHLKqp8i9mzRwjrDmRJI4iLn81XVz+TLC6ZVJFWHcBTlImM2EANlnlkBtdQDmURtsFlAMxX4gQ
7rJ29tt/QTwC6b59e4aDYZQesano3LZxGsA3pj6ByDIFqO4gsdlDceH54ZWZnaif7X1/kCJM7pWA
0xU8loNocTICCJJ+BPMUYGrvTrwlsxlswUNtaQ60MqPjDmlatb57/h8XTsSvQiITDEfP/CiPFPI1
L93rDZCAOfq6r3zjmo2kER7xKl8MjX2OjNuWWK4aIfL4GYATHVjo2Cyed3efgVIMgU76YU92+KRz
1JQdQ+Ky9f7KmRSzCXKFeyx6rQqjY85rjFtTkSnHfkFKYgkSyyThUsjIE1at7TDpUjyiLTEoXVjz
SBGlYd/3uD/ShjKiKfBw5X8zm0fn1yac8LbJMOZP/PWc8NeOWS/CUI2ZTbn9y4nY8AWdZNukL9KG
SMBiE6H4V/bCjb8o4I2N3G7X0irMPVyFpn67K5L5adjmJCnvwBtzW7KKUD/96uiFGp77cZnqBjOy
sE9/3xEtvryjv92TiIKgp00SmrLxJqKj9xAZ7fLpoeNGNWnOvUsDLkUWJoPwB3DZnt3HEbg6UfKU
vqJ1Ffz9DX0bH3YGLtlBx+vo3PNB1aiRW+mwRD49P16a+AbOhvxmbBumH9fsA68zT7HJdN8Ba0Tp
B50dg8kGNpU5tluFmj40D535fWOf02JsHww5c93bEAitYE4I6TdahnnOqhWljIj9DGE74hCbjxLL
KHQjEseY71RyAC6kkD9Dc6BbYnVhIWNr6cfNXwEGRdPEerXoUG12WoTq4sA2D1HfbGMSf7Hmpydo
Jm1NZ0ddF2MYBioVgOqKfb79a/QNl2jbme9Xi6DCsvFBoOFUkAmIxCVJ40oXea1EcIqOEyrhT/5L
G+8GOtuFARhivogG7iiFwiCQPcphBEnxceh7WDv2aCbaxQ/WMad7vlkosFkEqigO63hC9CuDSp0m
9m7JWwI6Hf0T4XwU8D1t+OjkOnaPc5/++P/wrXkQcvJElDOkuF5RN9qXDgNU5h/mBKhew681Pcro
cS1yiCrRw2uSEo4MjQDwvcLM5w2HuGeYfNMmcsy8zRW4SvdG58zaByEqUxftyoonubpijgJDyyjz
n7Z9n2alOD2ucQ448alqwBtDk+jKNdaA7aQhZsSHkt8W0AxHvBAQKxRIAZnI1+SmFiCkTcMdxAco
yVjftgjSFklkkw3k3YJqDZPBoKgyGaXwqVhr9/BVO7N/gp+PVk8rubTmlFUOmalr3w641mAvx4IV
I1cYaaOZYhVBA/KJX3i9/bVu/GfwYPM17yg2gp82B4EB/XFBy/J/0pkRhUJGtdMYmpWugaxjeLWx
rgQ7PsnD9rgbEcIKj3JhuTe23Wz1rAvBX4uRJgJuPPKFoQr6bMngjW8X5whVG03gNOMBPyLmF/L0
9aCwSyyQM1f3sfOrzZTCeGRAoqETYca0fBKd/zefhsC7COOtA9ITYa5RyqjvPExy3+4mXje6bufV
yI7KK447l3wqZUJTGMxEO4meADkMKc/zUVQ/1o1mfSfvkPw6HgCi5B4Wuqhz+7cQ4b12klcawU8R
8BipHHuUE+eAnpMMz50dXeIwxPsrA1/LqLTaOHYr8gY0NRBVn7WfuP/VwuzHoXQOts1JYYElEW48
XJ4Pyz7bOUOsK6Hw9qRW6LL+CwV1T6ZbFwEiSaDXEmFl2RlnwPtMduxPg34/9jpoAIGuBc5ayGwU
mSCKHmmHIv/4bbs9vcZmrC0HBqsnKS6FXLsZdZ0C6wEQ36F+ZkxDdV/lVOHMWEiwhd21vmeKq1ko
UUE4/xPFRecNqYyXZS8CgUZWwJJXp0n96AeFeX037dC5hGcm4Hs9YwXf/1O1wBo0eb1hS7+EixGs
V3jChYtbiyzh+LGn/9ayf1Tn0BfzgK4u6uxQDtT7CYwbZ4jSNT/JuIIWLDEskYLQNGmaycsxeKmA
sfhkcPDwGCmo2fG+la/rpxJq3TYsH/e64vbcK5KL07I3xAFTnhUEnO213wHTl/FbLBNr8mkGH3RO
yOiobOIEwWQkONFpzr5J3HgQyiTlta1nGdwboGAwXtIoThz1+aDi1L6nLE50ve7FEk85yjDCkeHz
SSm5oVdKiOHsDdIdDURYKQMXl52HBABFdToxnKuLNwHUWizW01kbvGbtkBtUo+9Q6QK0/Bjo7VmR
vHgM7e6Sv1OWrCqziVGao6HNGLV+mHWjRicJcOp5UIUDyjVmRlzEAeLQGrHcK3Ubw6dpRv3pl8bp
2BMQjr15Nscgaf7vryFZgH9kQvLyIt2jUon9Ljs2mNxo0FdjM2qNQXok53dw5b3jBfOGN7JFsHUq
XbA1CDfvd8mKEkLxTU32zbjTrTao1FfbF62JVvlf4Q5tqnE6gy8tKq7eYXEWqgGFbs1yQ2ne+a08
MEu14irDwB06T8fliYmoAdX0X0qTKTWDTNf2HQjLapjMhCqOCYELPkdFRO/FvcBV+UZkQ5fadMV5
wW2KYouQ1PgEAwJHBqcv7wlTc1pdHtVGCe5TfttY1AQjx0AvHiUBrDRNWTBRqlIZ3ZFJuS3eOK7r
5uUK1bnV87s1vVOmIJ38+ZkPqjAX6smx7Am8+r79oJZJvbryuhe+9h9HKuX3SGlvAbMcIH1aT0Vm
eKuyop0OD5dLbPug7uChpjMjKEc5dWzIyjos4VGiP59wPO7ZwtgaaR8IdW273g7sNIIkQJ3IFQOT
ihKQiuwsU0c+dwCfACBIZWbSZVQSr2l57Qtz+2pMy181epRVazh96EiKYqW96+yiO1Xupm16EPaH
ANFaEHOK1bJ1iStoEtcQbfkcALhstbQmKbajGJudkRih7aoo15V1YJJVlk9X9mmXqOse8AMq6mib
O7jjFEWIxtEYWKgIvuyPmOfOF2ybASaDw+5YujByQJCJgizbb9Tfcj0Bq09OqOuodc6nUmbTTRwr
oJXFEJi1fwkCiEQLHGXLDMosn8GDZM0C9eaIpuMNKZ+aF5q2om5i7pbtEmEEHWzXX/wpjqGqiBnS
WgFHpbFgEk4vitblkkiORs8yf7n+e/40n9nVxxBMydOI35/L8+CKfHaEqCJhGBshxyIvc2rXfDg4
zkuTy0p8calDFpk9wkAeWNDKImnSZQa/2UKF+A6PU+9hauoEm0kdY5xU+v0PO+8vhsjf732aCT8A
bZOs8vuGSTMMrwWPBu7sDqnABnsMNdNtpw4duiwXD8kMRI5UJHZ3n/m+RqvyxRIiSqvBQ4n1s2PU
sTdBu5EV/1JXcfyn8OXU7vLGMhhqrGXlYjeKbpYjEur+b1TnXCtg4c4lC0rVpmEy+izlnDMx2wQs
jEidiXkbOfb3PsNSc0o4f0buIV8jLzVObllgLWFBK9CaTd6CQdDBHdC6qap9xeRLNHPVlZZsi3es
NAc4aJHvaeNVZwu6sbqkeHSLA7QQbl2dpNNnKGq7BoFz6XiYsNker1zAAjM5CyRS5oM27ZDb+waR
DBCqjV+VaJb1zo1t8P0k9fRufe6VZXTrTq/vd2oCQES1yoCSi/DI6uJ7hQwSONYYAA9UxcLX/mJy
KuwBo2xqfz3Xd4uzddAiMwhlI2DlvJqgHiIGL64fJ8WEuKuyR7GSOTqP3k0bE3i0appY6iXXVmWN
qzemztUogqnbANuUQCRnFoqurvV3X3inGYgirHR4d29CtNJxm19lp58tTA3fCwmwab01MNy8GHPw
pu1KLgu4KwLvRObwxJ+zy1+zt8gjs4afMSHNN90/592Zo1RL49QwSOMFfeyr58+bpKqUJlEVfllK
Dc0TPsHHzWWpflyGmWfIV3j4tShOn9EN45zTDPFWGEdULCs1af/+80PFIM864gJsWkws1DNuYxV4
IK6iCiAbTUWEheB6sE5kWwGOGiLWYQ3wuJ2AjSI555ujVLI4lE73AyJR4DJfEefKbjTbOXvGlRg2
fybZyexYRISceAa8bD+8YkBtqiG03FMC0K8rrYL5ZetXvYBJVjR8zyvgWQF1cynoEY5c0L8OypdX
P6MNmLziQmxLbM1aaCUfUzmdMiJQm2N3qgkhl6Wx9YXqLWx9f7Vn5ccpDLgxhyP1kXBW9iLX7+hg
4k8HtiU4DYLcBEX6WS5XkjyjcOEqEtJFJxWokFmOE541wrk0bHouA8ENsC1yX2Tk6x5dalXafNak
RMQ69fTLv2qxPMTq9S7T46cgGBWWeUGSY9thjg8U5TRxuSa0C7cQyp0nfDy7/njTDvDNGxXrx1Kl
TJUaMA8qu5aCRGZHSJAnRUvk2XPNR0lzIMscQS2OaF9DrX5bDDdWL4syE9fw7aWiI5ZEIMuVR0+j
rgook1zvDlO6dgiadQS2vWK2qy6RLCm7X7c+J0cN9logpas9s//43BAci+xPyxwTEyO2K9/rpiee
DvHq9En+Nn3bRz173lb5pAbOdiog/jPwXLbmC0YAoKqq5C50xXeiX2yDbBCYkYXXb6Yz0uTUISh8
vvfCFYPe6PWfbaReBheFY920NpPqw4mcbxGS9CaY8obnRrkE7VxIezDesSYwqgxdXleQeeDIeprS
Fxa/cf4QWTUxVIwEBjSathBp24bjGgUxgUMoYi1HT9ILKvvvVFveNzqfz/kK0qVdnCW6tNXIh1rz
Y6E2tbK5INIZeZfWLQenuZVM8J0sAUarjMrFOa8jrVuAGdnhFccxLSrAe2aDUT8GXFSdhUgT/aCk
7l6jpIjA9D0NnQERNDenl2rBaPpUArKlkr8zeDksWbiPqSxYhS0J1RSSf7SDf+rRnqaSSU+xg7Kz
J24+JsaPjs9v1gODofwrxrkDSiob5zi9TylbMjiEiMJeOQUBSgnyuduZAUWmuud0k4wUp6NzhWO9
OMsk/t4cjwVrKHrluwK0HIKxnv24BhNlSOHxjmhXAFpvtdIeE5V4nzvC4PbcHd4ImA+guVujJanS
ZaxJvwX0P02mlvTl6EqcgWkjozqVnrU3sCzdukFmowXckgnsYTzbPj6HiZnreSHdqJpsTFwyPI1d
BVkiQaoPRk5Wxh3mHpcGEzppAk0RE0rNI6H2MR3wleqewhXinOdwAyQCCBSveet2W5st/R/zvVtL
ISbsVZDNRIB6ltQdwTwImKzprnudWezx367QEuAXqVFjzLw/InMFzb3cx72PK/jOxleEzRAl59de
eoo8i9oldi8gZ0mlHMe8ptkS1gwipsLgETUd4livlVCkazm9IZznc2H91pvr+ECB0flRr/pAADmx
pRGScgsAGBXUDZJRE+YNH0Xenm3RudKDdUzAMYbDDAbQTXPJ5B9MnFD2SpDgZFtePYrqJ0a7gV+M
9uRM4mfqpDn9TDBCK3QhwcQfvZN1HTJfR+DLRzVf1Klqp1294BHZGnraL3lI2WLnsFt6E4leB6e6
tedLLb16BLHZ8E7Mh6cnV3QmexHWfL69Bsc3QepttDS4cZvB75S0/hgQwtHWS75zuXW+DJMiONqL
ubbr06vHSitwDc6BOsZIm9dBNA6S/dtfWw2qEPdepeKKwH9fgAF/i6HFly/k3jF2VKdcXkWrXP05
ChoquyXWQEPuKmm3gyytwd4/h0CKoy8uf4Gb0Y2ZfRhKdkoLPEixdceOBHwMNxJ2UsvgQvltx1TZ
wtDN1WLnBC62FZhE5BwISqRTfQrpXhDBFouzZYoF1cbfD4+PvukbGBwHSbeTcvo3vKBlCNFuj1qI
bhEri1cK0kTMRqOc/hDOa1whdkuR0yyhMjsRu8Ox28GmdBx9bSyI+qjmo0sTXh1hIhd0pcgDSI3p
hyE/E2atOKlmxaYAbZQIDUmauiAu2nG5JcrdamRQbG/q4MVMz/YTTylwz5n+X00nj5OmJU7LbcQJ
hjQntr6CtXjrfyMGE/dZHWvskY9rHsuwnLTLVpLYx/2zS5QwsHlh1799MRNI5ZRMUJfXtwaOnzGE
i8VB5A5tZa7u5Vv4PDS9SjxT2DEf1DIhXY36KsmsAF0EiGNnGxX1HOS8sfg6ElmmmHo7NzoYskTV
a8QHoFB93IkYU2hSJ/oBNQ5KgKJ++Ms3WpsZYLPLsmYUcp47svtD+47Mvt6XvB5NcuNFUAw9KVlQ
a9wCdOHVzudEJ+yUodxcXzqSGHRD0/0l6bA9QkxpzJAvKn9oStFbx3OE85uOQBoV0nMd7cw+yTLw
FNz8mJKoB0xZwONMN6Kjw+AunM9xxDOcP3kXutVHwDy+nCpn94Zpab+8WyhThnk+lOzqo+stZlFw
8nWXKZnfSzm9BFtZeu1VXa05G9TQyL6u37nErUw7v7rQudNBqi0hFmW5Rs3vGiobAtKJjxxVPt7K
W2rkRYckIgbn1WszL6w8hwSIbKjiqT2EAESSUo9iUjePLKy7kbxothq6LgyhZMLj/yo6bzXy1VOD
5j8cf+CQun9vEdnj/T70zYo7guvGsd1yrHnm2yu66NBw+ahcqFsnkaUGEhKqrvDXRQKvnhldzTRF
pnl+3hHcvZ+VfvYD3tjFglm6vXkR8er6SQ/5iEM+Lpif1P20z8gmyy4BnWTjoLJDx1DIDI4684oq
CfzOOxbOdYXRquSLZhZ7VHVBhJML09GItdWzD0VdXhGdmGEWClTlsGZni+lDvKJj5x/EcX5I7cT9
uLkJYmJg9JOmhLyPekx5OqHLs6J+qQjuk4WTemHOknoByyy8dam8a5IB38fBjv9yQtxMspcLLZPJ
+MNgiGqR/JeWeJz98gTaffFyfNoxijdPXwyu+Zv720/L6kxV5rgJbCbtNHSvffgNEkHXYkJpurEU
FsXm2kuR95v71qPXUDmfkWxl0DldmMXfNZDaeZKq/LzljvXtkhyy+sr9BsF5dBLGFnQiGMxj2mjE
5BrqvcaWqS56Os61UZoGKqOA6a92JBfEpDO/QEVkS1sRHQG6CJ39lkkHtap/l3s5ueC23qMV5iLX
clTri98FJcDcD/KVKsKMOyfxqXqJicPOwYuuD3gmfVdsxeRI/RKeH9SsSpYydqg9fNOz3l/TlltR
F+KElUcQXVVhILH3/QDlG+s5BTin6RSsfTCrfsWliiASDpoFUKCkCG5NIlMGdSTpur9l5YzIsoGj
rG8gnymykitgUUqvFJWkrR5Kf46e4wJF4rNFOvozLVCAiDG1UP1qAkWcWgnlRtdTXGJoUhDItrYg
yBup5r+EpBxXZ28/McrWqSS/FJg0cXBluDFInEpaXb4d6EOhzKqhZdCe2kT1Sh5RB0oAtouRDImR
YiWJzJbGooXfBueq6R/ZYQIo9BaZJ2JLyItE/4N5kXgf5Lm5YvUqTC3BBw0mLOz7jd9+x/2aMd2T
8+XSqY2gDAPr8sL0N+4d7W53d0g4SYvJ9j3S/IEMLONVf8wDDc/dKZv/k9BSKZ1kmrouAUHOUXAM
dBekf7tUsyi6kivK8yY7jiTpjRmBZp1ObftPkR0zEgxyYfxEBv2tj6Purg5K5yQaTp2wXVv9hN2D
YlisXOHEqvNQab89GaGXXtcqwmlpQM9xiMuf57c74HkI0UFNonALLBgMYHNEBBwhU5Yye5fEXIkf
ol8sIiFYWjvg68n8IZVw/PBxutfSBYPJWqWW4OKaYi5xaznl4OEGx+Y26JWEtlnlyRdQgrixE9E0
u6iK2RYvhatpBL3EtFhGeioTavnLqzlnGqBij3Ai0BgMl7BAxQWm6evs69JXSwm/O4ep0inJy4fp
jzs2eJtMcFeoBBCqZ0BRlSTCkGrZrLZezH1yoC77NeGX1MPABGkNSTzHudDqwB05zUIasmpNHKFc
GoSKyelLBveul+ca6Qwnk4s7FSQalbTeLDq3HX8Kt+9aYLMIoQgpq8zAkM9HYPkkklyesyx2lB5H
RVsKbfoNGj46pZY/6eHymgiJ/irrqlnbN+Q2Wl9jBmyltGnOa26OcYx/tzD+QPAcdOuxlGbEZy1Y
CMWbS6X48d5bMBdLgUi71cucOyW0tY38yoEB7K+xnpBaTycjwHxk6Y7eth9l5BlX8JuH9lcrI+FE
X5j1/7YFqvYy2Qjj06m2/dGnxCCZZDqur3bFdLiqNuJQ6YCFs+yRqvJ79a5GUAmWmoz1VocO+CI6
saad2AWf7N4chbQKips1uQff7YJMem3x1XRT/7v0FkrGcG5g9CJRNMJ54UtLPhBz5dG+yN6yXWF8
ayS0O4fT3qs6eZgCyCnql2nj+H7UBu3PQAV6lzhNCXm6pAIfvTzDmtmMUrzlfp7GC/raRNczc5DA
/iH37CxHlsoO0rRrfpBUbC0KO7fc5iFan5RtqMI5X6MkzqTiJrpgRkq4BkrgwQwSsmQJYVdvI4m0
X4j2ikh2WD8TGETRhLLvc5cxuriVQdlihyRObl9ZZ8P8p9UlsmRH2YMebV36/MvnzI0HlcOMpHPr
2pGhlSNrYcIUaGo8+V9GuI809PgXfUG9nFNCbG74sFKsxUQSB1KvA4XwhDYIZ91ii9Piy8nrA3NH
UculvwFfcPxxwGFUTmNvKRJdzvBz/wp4U2Xew8EOdYPl8irK7gaZJ0IdK5ZPkTLBolS8jzIt131N
jD7LtU38VLdoxv8fy65njp0ZJFGS9TrLjZMXtqjoqFRFcfCyuVB/xnHeFm8x3Joo3B/0HHGZSrkn
kLPJshjy5Vwr22+g1lN3eQ/PlrS8jeTpCwk1tdddOpqvLlcEyMQvt3pxMSGRcxTlM+tA6Qsh+EUd
uK8HYIJEoDfmJByUxA/fD0hbh8cBeakNREwS5la6mm5tKi1dMAR1ZlMf7MuS0JcYcC+GRPyUW16e
5IQkazWE0fMmgNvcfVBMXZlQoQY7/h6ttQw87nnB2Vs+mGRSky9eu4oXw9YHE+6bQ8ulnTa/mYMv
Bcn+J4xLMnCEAEzzhr7JVqn9FF+79A6TMDQQtD6NtmBlt/+kVXofP5oDVTMhRWn+4BOKBF/AvBiS
qKg/qyU5iQ5jOt62CwhXK/Mi83JRhMCpI/cCj995OdA4J1eH61UZ3TfeSIzEc5enXrEtv+Kj39Yi
Ep+ZYso6FHqM6Qy1YJoPUld0vF5jbHMNSHtKahwIBDdXsAHkM7oEktZiHvUGYR+t0PVSQ8ORl3+y
KURTBrsgV6/aAuJCk+b9m7JHD7JlAcB9pbGkZgtWfs+h9U/HhhzOepWKldH1FBAolfKsJoTyoYGj
V+wLttBX6FNiBhIGWGw48sY13R73zsG+gbHanFnKY3ZCvcLibVzEW9TBTGfEv2O7QInTeMLx3440
qiXyENrlU3rCdR4PNRNHsdvJ8QTB1p64zVHmmLiwRUbtRQ+YZ1FWZGhMwQmP37DD8IJKrzve4bdD
49f1bc8pDh04StnXvt+V7tRJ46DvSEfftdNDUv2mT15BYy+MiC2xRavErvA+vrTXQJiLfHZkOpoH
0O1/8S+hZtXju0dCayqqzC2kL5pdFjxQKVKwUH3DZNCSWC7515q9lvlI+6cje+dvTHkFgeaC/lNG
JAJ04tNMeVaCePMMzGxzvvq0O0Wq/S5UPG9MgxouVvd9rtR5Lmx5dFqsZupSTA0EUfCeHztp+um5
JNj10DiyKOOFvAMYc/cO7wf0Si2BJsGPic2kanmni8E9wfgNueS4dgP876JaF9wPmXvT3Bk2Wh6C
C0cO5c76CHvPAuok4LVXY7rKiT09EhK8GXnAznkE0DsMkYqqXbnIVinepW0EU6pq4yEYyjYqHOX0
GxALD0smyQrVY5yHHPWOcLLoW7eFBlBBZqruIHGrlrZUOohXMYrMkjzwwidS+gXY4I3ySZ6OJPwb
fmuv4hb9q6Sm/TKSY4zL15vd2qaqYD/ZSqEHFu0dnb64qImqlvo0FXbuLfcCWG9BJfkNFiuC1ISV
FA4jSxQbAZD9+XpWjdtQ8YBDg9MI4VyTf8aQUFCn4pBMH8HoHffi1nDZTqlgSs+EWXgRtUh5IGty
lTXWrCvMnCQHbB/zo7GFG87HhSvLgntdBssm44dQRMrI6+T8/87N1j4kzHoZOQD2izjmhB9yFa8W
jYMQkOjs9sFCxGaLirrBcf/K6ZAbUGfaCPmtBPI56jjBYmxXgzVzQyrigvBaAqrT+1RTFmn8n0P0
te902OGV7rDgl1W7m+G/1pTe2QxPIY5a6odIMTV3R32aubfDBHT09ni8uTqoMOOvmty+1tfTXvZW
/uIbHlki4JplxxI6wo0b1fCYYpJtepo0Z2vyFi0f8JnglxbARHpazPlE2WJ2bQmJpDoXen6N8324
x3OhLbBuewJ7n/hIdQbp10+LtAFUbEta1vXr+K8ud1qZnp7sAo1Evmj8C1QHDeD5iczDG8GMhxLe
O8uEzildifdXCW6MZcNjCcJjPvNCkynfHErzFfCNOzlg/e+XgKVh1Zwc+ALxb5EWmWN8pDxDYIdV
O0tLSRI6MwGZAdCxlD/rrDrAuiokA6BWEMOuDXzKclSKY4qWuuIpp1mJ1GSxOYF/JMO74Do7qhWz
/MjOGF+6G3vIfpvRn8vxU9LkZayQ0mGVPIj9j4gfknN6NgDtrw735M3YgWQyxYzzNPLmd73/Dehw
yXgMqh3ocVuEUDcSSZ8WU5VYOOZKxBcLjLiBOW1KGXqnvO1LN8cTiPPdL0BslPcYWnvspg1pqI+A
jkftoMv+zcOjoySQjW5AjZDi/2QdiAzNOfCBVeQuiZCwoxMCrxI6y12uTKFJ/Q6z9fyIVBA6lPrY
eH29FLFh7V0/rB7IUiYUl+WfhN4EJow2+98VbkC7319BQPUdQ9tvEu1MHgtoGerk4KPO6IhkveqG
YAMmmC4Bj9rPGTj6F7/IlkR1OooElpjLOZjiDaCfRgil2Thcbly1rlxT0CmL5Jj6BiMh0obbV/bR
SjmGo9ZCqd+SQk0OEdhPfOgZ1Jzc8nnp+71K9FQss+/kDM1rG+YhsvnWbMnmQn5IMD/isTG56TSd
8aOrSaa3ql38OBbrx0MOPPH2ZtJgJo1OL96D/aIV5lP9H4rNLBx7ozqpxtOGMb1L9h0AORKFSsqT
qvYuULV2DhCVClFMVJjmxkCHzLXe00ak36HIohlUjiufzvKfpV0S4XdcCZjCxgaHmWHhRzI8RjRL
jIgVlaIGrrcFMeJmimJ1g8pXPgfjWLjNcG05w12dvNkSDB4KSjOjzOd3P0cRemWQfHVngzNWMNGI
DEnjluYv/QIKUeOHnpLRZh6kvF1tH5SOj4fzc7VXLk8dNMR3XodfMAWWXbo1Z9wDsMhVRX3ldHmB
N2Gv9sCaqLOjvuMW1B2OrPqIcHvuKASVclXgTIZtWu/V6n/JnS2R0gG98oDO/5LfzV9w8QmTBLGo
gzqedz1QnxvF7RZGaGAqdP4e8Ws977tZXSvor2Jj2ThZQHr9NHNu+kt73QsS1tNIjyQO7lZUPUEE
1YTpHPbjvA3dJWc7HHGojkCazDgpQmnmddxNByhhxwjTVIZ0faXT+Ure+X+HwIpI2IhxCZ/UmFJL
HJMQ+onZMaabJD6qR0rkRlUY4h858RETaN7SFYFWG8nUadypgHYeI59kskg96ZxfrGFSbOY/exc5
ZPdswMj7A7ynSc3ziVpFs5HZsf++CB+SP//izHspQ7fLv/laqJFRZ0pONgQRjv+l60GZ6tviea2e
ZuqxqGVMYiV21kKYZS8sz5cwN3Xriklwhk/Yo4cr0CKHbA+b5ivGZylMIOsbgp9O1Xdpmmr1cDZ7
j3KhY/K+zcBkkvCYj46ZZYT29zS88cbF6L8/SlWdPs/vaVvvq01M1bMTb8Rcct7ZB77GAj+QdAO6
JpB4mDdK3dRxuEQWKw5Mg2EUB1LG80u0YENEPrr7vWe6Tb8BaXNQ5rRlfGBWE+J/Oox6n2MS3Nx9
CL+y+CiTnCAHNAD+t5RnvB3y3lhIx1gBpXeQOnQo44OvM4g/fY9/0/DTX6MOjZFFVt+x7BNDD0N2
/3WkWvhacAKwamOHHsWmb32BB6zsaQtU9plXBC+cYbwSE0p4inuXwxVT6LNcoBK5Dzyue+Hpupd9
2NWn/cse36sTunWiB3WaZpVH9HzTFIzbzTSNFhcnJIKCI2S24fyKphtDIdX3OatWdS/0dKESQWt2
P9fowC/XN0QHbP4twoQJyPlXAxRTaUNR31e51i758vD058b5Nh9KNJzozCbgpe8n3gha9IhQOAAU
RZtNjci5Sbzijkwk5sFm6g7oJw0OClRY0Vv+vQFzp65T+JtlEyRxgKvy+w1DJx8IOP73KtgaBtLy
gVtNWz+A5dt3fFeZoMYXfRXkwaRn1jYA5gyWTp+3bWQDoQ+8fpDvfZ6GZMfUtNrGoBZbtHueNXsX
1UO/MZR9hvGP1EOoS1/kKOf5etudp1CBlQ2S/YC9AT0i+EazyRffcECJwKgMFfFHfXHUC15nxsIf
2pK8KwIhF010dLzY9rot4o76vSboitfDivi1u9AbQTOPsPc3a6iVTOvu7DmC1+up+MSGzA91l1bO
GcCdTHlk+S/Ao9SJRZ8oQ3J5Lk6iQLHIe48DV4fc9vpVF5qqZ3++V+bF80GAsUs3GOj7fgucUZ3a
wcIIZtJvYUW4bfN8bpuC18Rsk7ejez2QTO+KcP6bBw+uR7RoOuuXwlJc/f9K7OQ+2YG+coZ6wCYp
80QvWvYj8hy4iPmOVH385LpdTw4mDL1gv8eWKI7pfA36yz6B6+sh6TyMrRoEMIvwzvuzKx35Zrvs
AhYE+GpTp7Io8c9/yRSTU+KvyJUIuiEjoGwyuw12QHEh3cRr1/WUmtwCdV8c4HtD0O86lU0Dko1v
WvnIrbtjO8CUxxEmnQL4owPY04E9avss+RDNgnwh7H5UF3g5ffJE4MEuFhV+XvIJcB3uW7XL8xhm
eP0Fw0IBkv3/UXAi/FXvJrE1Uzw5Alcw72/9NqCaXIVhGEVMn1TuR6tbtfPE5lLhN+Rxc/uCvdz4
waRVtdRWdOQ24C+RwtCZMPlh4lKtRNxA9WZ9PXZZOgIu1AvCTwmPLoDnjBrFqJGKLTKDg5px6Fcd
fbjeLln5q32LI4PGqZ2HJeiL9Sp+lzSSJMllzjLxzHse4nYkEZMDM1eNlX1uCJpCngU7xUAQgmjH
u95VeuW5iEi14CDao1ngJHwlzjx4RD51e7Fs5bLgfLMHcMRKnVzSOZMQ15YhT/MbkGNPLizVkETf
Z9VIZmzyjyQVrxeQKdYHHR+8dIFWBQNjK6ijYmeDt9VLU7zDxVJV6KMf+9s65+vT93vlVTEbU3mP
7x54ZzZhlu6bxXsIV4v8JOaln1y0DOtkUtv503K5sRhMUv7Iz1xONPotpgZ4Cq1/n8Vxv+rFjHM/
J7MWu/1H35E4CMtb5Ku4qkPsRrAFp113LeUQUVyC0kQ+N9GD5GAKJqpQDif78i6a05eryeR5FJNs
Kyof+VJuwAasO1bZbHruL7aWqCCLqg0ABKNvKzPRrZLT6USXzGTvvQECVfPfenT+ul2mJRd4Nxib
tmEIRamMUI49zSxQd6WWWyNiA43bTNz9DPZcwy8a04w0QujRjVdcDZmi+ykbGLgKPzrokDWfGwgx
MxL8JttGhLFmL6orUhfHE4KOuUfuI8TCHDd/nGM3Pdp30yXiIqnXdQ38ZK0gPOW47SKAORioPsqr
pOVWluuaNufes73fWfGfYf65Pc4iq03RV+Az91k48vUO5ee9v4PgDDtNXh548v5sL7RGGQun4j/U
djfceTqcpbzHb9hBop4epELyE4lOF9CpfI5cLJ53MNHkGlIg4+nqTFlvvVqIJvUIEZM1em3FAxZf
J93ntiyVvAXMR5EO/ieYX2rZYkDuwBviYYCKJF3RoDqosITb71SCSSvvkSfsBVFhQB4z7wSpggC7
TpURIYp9w1g/z017l3ktFB0abhoURcsLv7MiOyZz+G3BwiPHgJLOdmOObcrYXt44SjTBR6B+iy/6
DjHmTp3OUbHXIP2uzVpjkFcmc7YUODlcn7SrC34to5iMJ82JLM2J8Z6Rqjv24gc4/jiQaNPYw+eg
okCUbBvJ8YHcien5pfF7uT49/NZpMhFKJvWyrFwbXRNnKFbL+HX6SIUvR2DLM2Nsa+aGEpnw6rL9
klR8UxqaAuiHd5POB5wERciFYYos6xwtgfi1x5aeUfcX3djVPDTp06ZgPZY7yLzwjTmtT9XWrc6J
9ThB1gd2nBXkncZIDI7ypxlA+XmxK9ejKJuBfeP4oh3jv7brLNivxtsC6wfK7qEfdeaUtYzGh2Y1
SE+4AnSq6KCdyasK8ksUXS12I4Y35VAEk3PK3kBIFscQpDEcatn4CqqJTlx+RUCP1TZVCn9XCAQM
MxaeF1qqMGkMvyNDas1t+VgaJjTzdcmh2KM7ZJLazrmTM6ZH1dm+ojlkrj4IGMuFCm6Fchi6gGbx
XIquWznsw4l7xP3craxzQIC+4mPGhgZcLfx+6tWmDXQ6BvcMYSqp/BiN0UZhixxrnlP13NPF3uMQ
SdkTc8yDi3tFoTeZKHcgnYv1XgCrEcOwiLdk6vHsfR7a92X4C65wBDHf5lEKAyeHpFUia2rBve5l
ysHYxDJwg1flRwSIba3D2cNKRs20vk/1cWz9C6l3HVr3w2cJvXfPnZaQ+rwDQt1wrbtMaCXOKaGV
xb9jhWp84M99s31ZMFiMi/f+jNleT8CLhI8idWF2OklUARPA66Kv+Muj/H2cHP8FNx+B8M1H8HzN
xp3HGUKtAJaZb6LxM7Xl5PeWrcC4kHP134aUCTvC27dzZpWQPYpYwQ2F1AcL9tvAjMj7ebAGRaKY
TAZ7gw5QCj+mpzEAxXtByIrQQZglJCZY6bP8AxkEoe3FinrhvOABoW/VEAQGg1cy8cS17do9dSyj
emcm2LF10J/V6WxO1Soxy/AbcwqyTegvkuATZKRyBdIjfW1AuIeHEGNl4tnS8kzWu7G9jgoJCkS4
MJc4F9g147UoVK1aUKIjxTTCCbGVysprI3grKuw7nxhCHh5TjYO7haRGKm0e6b/Vge75nZuh4aYL
I63uSl2Na4SOXi0E+vjEybAs1Jz8Dfkl9bdjshoeDqKSp4Mq/FGRNtgQn4TGinaI2OmLg81QuyXA
5WjLyX6DwB2F0jb4aVE4/fZhHT0Oluv/H9HA8bY+XKvN11HMKXDncUbTQ4zKRXBDGBPsDZ3KCGOJ
KWgD14Ftq1HIqLReKc+qjc4WbmzBdY6MZU+NrHS4gep/dacJZFDYp6f3iG+rGEACVWbkYzZtNap7
W8tIePIbeApYHU1//eKSycagoTXIaceS6bJ8BbRY6xIvjIS/tL1/Pbdx18+wCe22Dl8p0t/I74Au
oFMhyNdh6QWlRTR79X2hqdHuiUZxUFpyBEsBSgGpWJEFGKdIGEeGmK5C+bORsrJvYaxZHL4JzHNj
Ukbx7vf3Rc+ay9YN/107TAG9970d8TdNYj4noOGwGL88q4ol0VVXP/DGL6GQFxcD603fWT4bxaVD
COZQPSazN8Q4kB4aZKxPeijvWK2mwqRVyAHbQyHh1YVfbi8n+DNi7F/0/RT4ZAOvSwobMSNiv2FL
ehQz4QWODaTBZL3b62GMK+JUxshegw+B+OiVH44IoDCZ2/av2aryIwtfsY7RZikTb31/mgsl9EK1
0Y4nNgj0lPOkQ4o8GtowLm5M5NXlOA292yGgocTeNGxyeUVQnasSHpZ2jHJ/Yh6Zbl/Vgt3ppkvm
u8pnKN9mQUzHmCkHUi/UEb49B7t7h+zKF278ZahJ3RxiECuA8vBaulL3iwghnlGWSoLAjezO+6Si
kqFaznhNwYuwQGbC1xa7Weg4RPs2ZKS/v3Lao9L6MLP44eL34uO4WmxB0EGIumUunrVXQUyB6sLF
Um4wgmo7gfBBvGE/8muRI6r6VbPMdEYr8I2EVWoDmlJTaVOrpOy4y5ZGzxdNla6/LlwpEAv78vk0
jHalgzt/T9odfy9EoaRBaCK9vCrYZV8ZbCxYh4LElzSZrfguIgv9DpiRuUu54n19qXfxnq2FyMqL
tjDHmmIGPAEHW1Wtsa3GrXVGip0RWn6JEKAJx+++dpWNCUryjpeKdZsb4vacEA46EBfOeOTlywwL
QeyWiPyHCuZyhubhggyHmvY9lEGOZChmyw/j2AU8SdR9SeGZbip8e37OMrHjU3DBL8tt54vJ1Qm/
n+ahWgTuA7MloMRGkNSqW3OB1gkSD8Hora0eErIIphg2UX9+ee/LbzU4wuTe+HkwyYs7KRTNK2++
SV32I01S1BGvvP/DReE25WaRWGdzIBiC9yKuO/CvkrjwnZBnoUFOB/2mJR7EEgAefoLacIwh5BHG
fNeqSMqddOcDF7T1MkmHGJs4Fy4k5KSQ7/A1NOCZ6z/epfe8of8BarfBLtGrvc+RkOSfM0FQ91sX
Kr0yolGBxZYu1XsmggHHWJURvjOzELZz1uNdgFZQbP+CRgTaGD73/l3nOtvKuEx3phNWlz8itYvo
bDaUovbb292drxB72NuUFG75A6NV7B+uRlLZ6ImQOtvuNQDt5Bd2/J6COTvnGocDPFXSL5yyj/JL
/QB4NPrfGxwjyj/bobD3WulZL/HLJSQDSCtca+f17gjh7UxkDkzs4fV1PFfixOl/Tq0/S8abiM+w
f3FhSNHvFOeQ44kwQMqibe+cS44dxs05Hrwc/83UCFfnHvOLH+0ueNUQJzETv3YczBDNsGK/wBEB
FLLzVHfrg/yPw1O4CkuZlLfQBjZO4amK4i5LU8wxrnOCHS6K0/E90DjfYuDUMRqDFBIWK/I8FcRA
ZdbdIh8iGUD6Yjh6f8oUFlou/27MJplFMbe+M7i37WpEpVuQl+fQ+bK73Jhi8Nqa1/Rq2Ssuzxy9
PML+kEBSbEIlml5RPyM9KejiinC7G6asZ4lEIjRGZJ36hP4rTr1YPWEvU+mgbhLuwZp9lFH5bODx
7nyG9PvYbV27p/jGGfn0RELRix7LZD8jiM42MfXTqG+ihb8ARCu9rT5BsQbm0aKQiAISdT1z1fa6
fDmn/Qbgnyex0T48hsnxFXCcx/wZaMQ9RJrZXuQqgm6c3CWL6B1EhjKmXHssSmSFY6quC7Bp+lVP
JDZL2em7b5W7C/L+Z02hvu3zCUZuBjNno9FWnpBAWqAN/StyfE1gQEHf8xBuPq7GIwAS7g9aWCpe
paNiW3aZ5RbO85ryvmAj/XeQP65i8CAxjfEGMIGov0xAGB6X6WV5M106MAz9aZy6CPfXiPZDoJ8M
FWKcUjJw76M9BsoJpdkLZM7AFhNJRj7BLF8CaMmx5/yAV42URkrVV7/oecc0uhChkexRBamMjyvk
NjFlhP1JIBNCeGooNgPV76dUpxW9NCWoJbLwYD5vQqEzYEPgBNiVmNVl/FAXrTGUKbx7wXPkKCdd
TFXDrUAW8i6bFos2ZhnYHUNHxOv4W4BNQOK5pZmVLDE3vGTepXsiC8HH5+AMshluDZp3mlEqDpeQ
3nXsYQPKPOTmZa6WIDQLT7QUjANN+OxDdNFSuxPRwf4kUBhDtiNr5gjaTkbezg9p1q2+O4Hl8VT7
OGksMiWZawd7FZexVK4+Rx7ofJUcahAMVE7E0B3eoOxxKc6ffS3dTT4ZxmAece+/yx4a+a8iPWG7
gFFV/Uq7fAsg9WWGrjuffOPBqb9nC2JE7bdMGCcPrLafmUUpkbAKt/ijihb0YK3Z6lfK8KkCcb7Y
gP0i2msFNZbsE2v7qKxM83JBsD+eAqpRl3ssWY2KtKEmBvSoIj29B4lVkqUjtuie/UlXCqRRPD9q
IIEjEyOdMMA4JztxBP+XoAt+d8x4+DiGm6+HcdGAu6NNSz/ttB/ZzoRB8uCYx+Zu+2U+DIlXh8Wh
Zm6rR7CDIT2+EAlhONNSzyOp8fahmKZ680E/+LJxv4A4YmH9VlA4DiATztt9FijK+JaKOXEg792w
w2RwuALgmAUkGImHV9ug1RG0Q5jLy0OgKz62mkGtf+if97hOZZz8ZThj6Ub1vNxO66eEhBF5qQII
Pl/eHE2h2n/EHIU3JOjAJFd5ox3XPBzW5z/mDZS1/i+ekIDSSqUZbxaXZ08AFdO2MI49zW3whGdK
6c2BkcC9hUBM7T5NOAKDpsn4pPca/aDeIw9H1Z/dFBNb+z+5kZRwO5IbxXAMz+v03D9KGUVu4mQS
t9KTOxaSbg7rvu89nV/DEempmP2WzqdQUK9In4iAsAoCg5fsXPB/1Ff/qp6raP2Eo6KaCr001bbI
ncaI+tXgWT/RwuJ9q2+wKEOg7JPUGOUNF8EL+KUgqlsIUMSqeGOQTUqD3QgDRXnteqENum8l8+kN
EfBjWuv633qUBH68t/Eo/WWphOW9EdGgIME1WPscRNDwnCVgXBTZ3RZPPMb3V0PkKGUTiThAKle9
2gNCE8dcDlV+UMkL+ejxRgpLIZVcEyFNIjoYRuzmTRqX3OGnyaUlwnb+RR0NoyCqlCyxakJLpB1d
fyPc5vCuzXmLKDEZeJXfBcoTSeM4XGRmIMxxU9LSmB378MsxeS/lJvjL7kQZA+ifbbq7wTvfZVio
qHiNKpzSDi6NZTvpj/YE68m5wN/wdxEMqlrrPTYPaCJMNdGULCVDBvkN1BlZFqdbAJxKzpscyZyE
22sW0lmVYOqdu5+VRRAx1qw6s8wQYBPEqQAh8Yyy2xO2U+chTcGgfi7WRipULOnUR7bIoTt62qK4
U1xZnaNBCsxW7r+3kpSENcTet1O52prm/TSoOyxdZhkxH5xfTFuI0LYCmDmhpoDsDhpL/9Weed7Y
Dwk3qB9Tk5pG6dPWX8MtdTkQw6sF5VxXecU5KBlvWTNbdIbcylr/R0dZZtwXf+3OuPtMH0jVGBup
XgJ+RSEDWQHUl+WA6KsgjtI9YgyUgG0h/ebJZDwIz9PyeucoUmOoJ0obBdDMNtGokvWdlFk3hs6v
83gD0semL/aFxTFbJ3EEiX6p28YXiswp0jcCaUxnyxmStQWxsVycSw05ImDKEz73L65oQWiQuchW
WsYfzEZ49L2gXNR6OotjHjPoJn1U/z5UYzHo4GFngrqbH0JU0uT+zRyX9672A3VIN5R0ThM+/KrB
BiT2H6BGUzUJKBqHi5ZdTngYnbAcDGTmwYk1EmTvMq37OgF2dG31h+5A8hLG4f4rviKKUHOcA7Bs
pvjn0BAirprnUvhtBUlTzZdvGO1H8AaHcDSMV2tLn01Opc2aFVdlX62mjXRSd/CMGV4PvaQrvZDo
aCHUvVMYtKPhD1WokNCihgyfWad3knzV+qdO7ZfKPRdAbGvtAEv3JSRCo5HxfSsS1N5xqX8TtNvA
XBiyx1xYzZgkebRG+06hcYNsvq0z89OvX96Rx3oxuFPsEbGh++3BerkLhCvnaAqnaE73nMuq09Px
axlKdxHER1ycLXWyu0psSt6Rd+UrWa/Bp76qqp80rqaZl3g9bEByP46lTK9LKsP2ulimbBmPeqfm
o6QZACmszi2sTgP8QPrzyWTLIYXoOhKDw41reDnzgYgC0uPpDQDJWC3m9QE2RzRds2JIfonZk3KF
XjC9hf9YZ+a72HKLtEYwsx5Je6SQo5aP1c3bYpnXrDS/c+58he8mXKp5ZldMhJtEo+MthQKJNI8U
auq5yk/gz3zOQs3YnNTB3hxukKse1y7YFEa+mjOt9mKJFHw1KB+3Gr3GcJtIGH3An6/zqOCE9BdK
uikeGGLXD0b+V0MSWqZw4iR8HGyA+WAicTH5LoREGMBNUhlasEDrXjHwaVzS7l4/wivI4MyKBhvW
OBulj0GejqWoyje4Zx8jDSsFcIQVm9sc+15oJzZt09owaX8ToNiT9FTlJ2FQbyBSjfol0UWjoyEX
5YV3Evfa9lhDoC4lq215UcjxpmL5F3z3xtq728CsUzus/4awwa3ahL3rpcmCJwVdbL9y/wCMliFu
nLFPy6/0L8oN+Zn7uXXh5G7uWANmRvuBlpYmbFxJK4fa3CMpxFgzzAj1+5C5AjGqlvKFIusQweDV
V6NWIPaRSiosvjzHBvoZTvZRjnxBpjETogP5B8gigeDuxQKOgR+Uv8LnunZyPNW3hGSp0trsBQs2
NGS+vPFEpbvOB991APmh9x/KcbE/QVsEekwo1ukH5qI8nYaHNdqhllzD/saOmRnt55YVgx5AAvDD
bYQFIikesfxYsL2odWcXGjVezNdaXVzyJX7Su0gFupIzRBG020n6D8VQ2DbOBBpq1bA0WoIEfFXI
QXivrzPdctF5RR35HQqXntVwLHnz1c7uvyhiyJ1veVpEnCpJPNb/iRHERqwa1CMXalfGBlOdY9mc
Sw0BThIIluaGOWcNhko0oiUH6Dcy7pwO6ov9+PgaZCLFIlES7eaC0jVkHLO/lVmOHD68r00A0DZU
b3j3j+BRgyJtjL/YdXtbvoc2aY6uB8nn9DUtsdudbzkFGUT3vgssahIwkrvGJ+hBQbISr9KMKIf5
HBn+c84aTa6WPl9YInzYOf+cEMridnDAQ2QcozIdpdrCKgrncUzxvrpbroRqdW5zp9jy/tMV3a7Z
BfKtaLvpihA3NUthiPe9uzmN3ZnlmFvkKPVGD9TFurkBGeE8RrXkcY0icAhtSe+wAemZhcYHuRjP
kRS/0vWRq/qfFFuBr0grjER8MnKXx3fLEpUpoh+JQnwu80OE9hGfYac38h9WmHqisZ+g7izvl8Np
JHBtcsMESQnfCswsvhrjIetzf13Kk5w7W7iBgf1M9DqkUcwKYYZaB+nCxVdoma04gYLHM3qjw81W
kFGv9/JkMBr6jM4aDEu/2PxfHYbogBcYvaV/IhEZ6kORlSeJ2dPPQYQIZfAit8NCby165V1vDPEr
TIz9j9s9Otzqj9J1fFMYPflzuk0Krwp0aBuu25AojviCdJ/d9seTiqJ4W72Yo5e5r6XyTzt+q/BC
Im7lTXsKBAlJjymOOpikdNa1pTH9OMM4jbMNiXWrPRb0+CM8/c38hshcYyw0FyDy2SBTPpJXPuo1
HdXVxsM0pT+i2cMpgnaoVRbK9yEiG0Uk/iFu7dCQziZ1RqNw7skIoauwzoigKf2J+BMqOvPdt+Sj
GYH0fmOam3wMnsInIVWMx/+0XFN+a+qUc5KOUNbtq2fTi+S9huWbkMB86x+qKJJrzs0zdeN1L3iV
FTPsIantoDVNhEg4V+X7XrsuWfU31sGHbig+JAYiSb/dkvticbM08b4RDsIVgI2UXvr/7Kzg/xNZ
nAeKQOxMAtViG1AIAkw6OeiSjY21Q51ZtFThaaQR9A6Q0gQGZ0deo+ZXFkYslAvW0SRMmd9TB/W/
4fXs4bBBxXF5+VDr+ArHzd2mdagwItbf/CW/kP4AF+SDLZ6B0xrTA/gWfGGCYJ8P0HGvneUpYZSs
JZwmxubpvz6fisr1oFilpuKggNxmQbP7YFV2k3clQnehcC8Wz9xTNr/dvSliethrAKD8/V2OU5Z8
jLq7NYvOX2dw8BDSvGnO9/ZPtUE074Ry3p3yZVCttoulFf29XlViBnIzMoXc9WWu/UmxBn1LDIC1
D4Ki1NhYWR62FYkg3GDRkS22cfRJX9yqianFpeDZzlHI0wNj4/Hj/iVpp2y/HI2gscLdU1xJt5Ft
tncBreGRALUPA29OOo1drpxZune4kutRCmtkUFz++MtxZzWL2xzUqMLt4oHTfMzmVkaSFffoyVB7
7YLu5tERoBXWKACymVCG4D5sUBC63aTUYpSpLXeK2KDu/4bsGZFqdQ9fVrAQ3j2lHafP9Rbps6IO
hvu2fs8WH06rq0z0xhObptnAdw18yd3ikxhM0N0b/36vv+PT9CzVercF9rWaOsH0Jo/KTK4lcJXQ
SR3KeRxPOLoEhzEg0q1k30G19LJn4DSz9nEoAXJgq28i3wmdeDpnzxCLkPVs4b23ZeB8shm/ro7S
+mxNokc0PaJTyQekhVkkulwaZLVuaxw8NDsZDVS3aBue24i4Q094Nx5naLKaAL5xZ8ojihhB3Z6E
V2JzDGsBp/FqGnzs8CiF8vaHiR7O6bPULeZ7b/+SOoZ9DeFimpq5x2+LOnwvwN4UfjtG6UEkLQHe
+UI/zlGRvcE44LR72FRn130jGcy0kdIJ+rMwo7jk5a6JZfaUa5xobaFTzoGOhp9PJiqmcETUxli0
PSL4QCWWLergzRjepDhDitC4tL0aX56qR/NjdPILgwtsVF71UKeaM46AAiXcb6z68RGnaR7CubEA
dtxWYilgwtOWqRyumGbnOeBIsvrr0RiMBUiZJxKM9jvXiBfZLovWOkG0QqM9hfjOhCf7a3otfUmX
gFNOpsGJjdPBCJrwp9qdvVorFA7raIw/3afICaB1xHDL6ftm7jouE0PwBFt/bAjHqOPnhk86G62Q
dm6kOBsbvWgJYwvf5SkbrfzjsPbS2O9YOPtj7D0zZMeAV0MJNL9we+tinGa6o+R9cSpB5pEixXgc
xTWSJCKnmfKo693sxMfPRo+GxIJNqH5G+h7wjv0ARs82BzW3BECRnq38Oi8SBHBrTfR9tHpi2sSz
MyaS2W5UaDL1bt3rbNsIHlu2z5yFXfkFP3cQmHyS73BQFCIhgvkqMacI4AvfxxcClPLnAyi9jckX
r2pcU6hf6EOb73PfVIHmVA8M7/Rwr+W3kxcz9WeJW3QnKEJoa3GrV7G/l70En3uGz8XAbL57BCDm
GMisnHHM1CUCEDkd8Lbd7twM8tRR5q7xnhvgayfYQorjnHLielgtes/XBnlNmI2KOCuA1Ja+6c0W
O55Mo240g/whY8omt+Ksfn2UgU/wV22lcNlm1cWOMxCGnRV/F/FAVvFgbWj4R4CzNNwCN2pTxxjs
AvtmWGjnkJ1EKhJQ7AB0SmMjw2+iGVSmfNaLOhaja9QEsF8uTk/kuPayU16ihpHR7OAUQ3ktQ8iq
kt14WIU9pB/UZcP6DYjM0SThBq397wpdSqxRhSSfJcLQGzyCy2R6mAI6W1R9egPwuTSWADoIOGRp
31dbC2lbyvfJwBmrRAUd+RoNv0pSkBuVOcMoP1/skKookxT5w7nYb3enxxLIMzGXVotvSNgpBekH
EDJ++rLfZRJTr2Ev09XV+uEtJ+QMyUbTVTJb93YA92xW4noLOUbxsqv2gdWHZ80LJGgwoqASfAQI
LydEQlOMnrmEEOMx+UvuWrb4uyg6kzrckvcrjf1melVeNk/K/hcA/AqdHr2nYqVFZ/zhgALSuQXN
vWYVNrBnaTrSkZRbfRPRme+Vd8ebrbNXPtm2bcuOo/50RvDnvVFXwg7g8ztDwlCRWNkOQFVCv7Kn
Rj7Un8tnDWY8KTspt2Zi6BrL7VSdFeu9zSVwWF1B5sMgkI8yMS+JIER0pK3t+vzoZfnMHNydev/n
yuBY4mOn+FRQUfXiNsn4V6mBqYb1oP16QYQNj3wVmC9W9XhSuIXgvAWE0W5tT98W2jEpM2Jvgt1E
UdFjfOqfiA0ePS3UoGlSlDi0dQVJ+9rWzpz0eQB5MhqI2l+8a/IYyIdAgNUYYh1A9S6m/3ToJr5C
ZqDYgPFnLcU+Fs3iW6/iNw3Lr5ZKQrl/YGW57xK6sCX80JLSqZeWVqXEZhkS6K4sTGPllgfqf7vU
WW5ZJ6gpUOG7KVHfxteEeYvwmbEpZ4xIQIpjFbPmmS3ubSpPBKR8DMJV0CbYzF6kYmRZoUP80YTQ
bjjpTYrwjs0C9JoWeGRCfT1K0fkhKz2WjWVwtm+gOHrsJB+31ZpQGZinkJHtqziac5UP7jMIESAO
sedWSlCDaHE0PXRypMZOGWWbL3DLA+M1Kcpxjdqp3JDx+wlnY3/bbzFHMdmD9K8LOZxuFjouhU+W
oSRZu7zMnkBCSsx9SJRp4dzlYHdHOGxI3sOxWgoiqUOiI4tHw8hgYYwVfvohwZ8jesKdkRNeEn6j
QVwRc5sC2jWuj5xfbIMjYlzCOQvRr42lLJf3a298j9mRSBZPKwdZ7ATkBItVNkUBAlb9x8dzX1gK
xYbVANAsykJs2+zzbULoGTYwWgLy9Y+wupuVApC7BRgn/wiW09RmQn6mzQwobPIEt56SSnQMF7mR
ePugoiLcTx9sJfepMdSsFqpdB43dI1iNUXephweQ1Fw3nzoVOFoPqrlxgZ7UcqNWqzsKi08oX7Mr
JYb7tn6qwlrxJ96O1lcQB5J+TJQMa+lye/ekL2aSJ44LxxKikxGtEelBx6P8TN4dTraZ/juJAYQK
fUlx/9HPLKuE/hR1JCCF21q6ReMAvTvx+T1HbovMkFpE2z7cQ1A3S62RcIAtuU8i+Oel22NQNhHL
UFPwajtN//GJiYOSWbgWYS9z0FuhtRgAO5jA5fij5+1XiRy+DYpAfORazxKd7Dg3M782u53YZ6S+
sV4oxE+MO69JXOTNRO3t9D93D9NHfPfhgt0GqmZ9ziqNXY1s/l0Ij7vOSt0jeJo2i2GssI8eCwVL
pE4NXAVu1zhCHzZWN3ZEFJnp9pMCGZhxk8iNlR7c7kHMuvbfGQxaygdfGXtsRRGJqQaeR3Yq5GGp
ZEsV+z1GpozcbnCIcUCjBA5PBPBVK5s1+/P5glg0Mq8qp3ooAf2Au5FCFM6GPSbuqiPZVgWeE08C
QssL7/3zTmpernponOj2lHRI0yGNk4BQQLNpQAdD+ZdmaCMwFsyklMWR+elG+jFuhotVrkCmjpSS
8VTubPCKW9OsZrrymHRVy+Yla4kyqn20fRdaRTdgNW2HIkvnGyk9tvgHrSUczDChJXSDKPG7R2Qn
0o7FT2eelsFhM6tCLkH/koPTx/kD7UbS41C5fCPY9SJmgvj1DL+ZzjXWIDnpcKogsGXKVqRcsbRs
tZYSOWCp+oIbA8A7Zc14aEuw1ZRpc7wbJ3MI5UGbkTqzA2C9jCOeb5QpoFWvFdaIDQBmHXYlXHzS
dcZf6/JrrjSMCiYeHgU4bOm6l2zPl21hRWr7hC6ZDOaugdaXDnzCYWsfVyLAd6rFUfMaqOhGShla
AcxXgKqk2fFJ4Gibqiewgsq1MH8saXwpEg00wh6m1gudnOykkzTlFc1Kw0o9/EmyV+q+alhc5fTR
Xb+5qJc2f0Hga6rQvg3KL2MEvNGiJ+9hrlIysXqPu83C59dU4mC8dsE6RC8X7MyHwCVkc/vWL38T
0PAKBr30IZmy8JG+mmkNBLIAG4NtvAA3bsuAbRR/zNqX11TQO5Te0+P2AwHSgBTqshTCaJV50Eh5
NB/apx+Zh9/j5XOKeX9Kp7g7qpz7cwjMQm3orfKkTvMl+hCdXaA4b6KqDfMbZvyWGEf0Nc4jkd/j
rCFbx4RkcYP9tBp9GHmDUJcCNsC5E0LeaiV8rk0fL1mNvCDqfVV5z+COtTaOPAUyzHbD3ivKi/xt
75OkQxyd69zX5zBx2wVmpjTe65i/4GKt7VUu6Wu1BYagzKgqgUmSqMSEFKN6QaAed6RVVEnDm4A1
F1aNmJiGmJMZd8mdU8nMhQnuXd7YAWnhORkF/KTnxk4OSSVd3vcLpTd85Y6xL751b6EF3T1MToqF
CSNtf5lED1q1qelDw1Baspkr3xPkJ4344tjp7m6YE2ujQRdiYqUg2P1FcDYgfTjD+KZO69ybc4Sj
25x0rY7frT7rQeL2hycb7F3P2u66v5SW8FwfV4g3N11HWgmGkwsnZ/QiKPA7YTz5MjK6cy81yHOs
9uUwllJ6oIwEkfqfhd5ujD7OmA6MHSJeVTJu5sK8CPoyOYZUa9TLb86DdJ6ji+Zv7i5L8W7x2RAp
ZzXESb9yJl1qQw/tGWSxSq3jsuT5u16VmvWVca2UOzDALFwr266dTxwr5t/HPlUGlC/5PeNtn+uT
SSSc8FFtpD0l/WZbPrhZ4xXxYZn95R2JUd+IwArAxOXLiAZRY6dvua1UFxHNXUI0sFPpTZyFS4Bw
RBg/Scj5kKaO8CQFvSLmznuwUeS0gyJElf1Nc6EqlEj5Rl61Lr/NC0rlU4Rl4bT9cQES2BdyGeQ3
bxJeLIpFoTFlOF7ks6h9ulKaMNpxWrMyFBZG5uHrDoAXp4LjG7WAJQsfe3fL8c2urSKmWZV6TH7f
+eybAQw1yEpduNp8HUPQVN1adjxmFlgNMSprlk/0vRPv37nqe3SyOnXTL+fOV30I+vrA0lo/A1H3
X0eB1OWQV6ccVvTqqJO7KBM4cuvmu2ieqqekEOTVjWNpU3pWLUM+iGCgi9EzlcX7WWJWEvONfRvU
VnF+3USIzvB4sE8pQ5wx02ExiDIIY4KDahw3pJ9R4yQ5ggacfHE+tCQF38nkbk+qJmayEd0+r9zr
xBVZtitscI6PyFsmdsQtszrrKCx0wjIHnEG6CT7vngSYBj69qgrhpj5FDlicCaGW6mbefvIuY9rG
Nuvo/e3pp5Sq/qp5GH/lQD1hacWtYU2TWmnENJv0zaqTIBQEnTebUKJrBjPau4BdArhx3F/QiBQj
NSuhcHy280Sdt7pa4AcxYj0tVLoWT5cg52RC5pvYXtToFtffoRVEO/xXBVXDUyLMIAV19k9/SVYo
9wmv+WqF1Oj4K7+uQ3Wo+2BuMAlyooFGIBgoyBmTgtKbiYK88JHUrDVsDtyzSyKxoHfhz8SuNNlU
7LfeSCtWoRcxgFOHOkcNn1b8eE+gPF2bzzgp3ks3HvtsfE8rVodjj1/Nnbcyv+hHJiS3SPG8Tme5
D+FbP78oW0/Wx/RnJv8JHyS0rYjSotY0V1XfoaXnd5k3jbqdSwHBe7rFeiGAMykiW55RIuK5tJE5
XxUzzs4MUTJQ1wT7qF6aXU3xukVKSNiRzAWLZnb4GCVv6BDTMFM9vg4xxLmkn/KUsYCXNHMzXta7
v39EW8eb8FHa0aKGFxDoT3Onu93AhiXHwnS8DAY0HJWBHe8Phj119hWyIDoUmN9k+d0CM+2pgZsk
kC5VUXUxyKojM83YlWh/+DTc1poMIlWexFRr8PSnJDya7xt3MkIGitC6YNHxJjwfD0Hk5IpOB1Zq
jJdsplCe/Z7//D3kyFj6lsPkA9M4mB5ZIrRl+NQxScED4q+QnL+gG2pL9XYtMhU9fYs42SeIFG+O
fr0g8aT/2MRzop9id1qv30s2PgJL7M74Z1xrXzQAzmkaopq6rMOzt/1Q+BLI9yPV51gMvQ2szYrU
AizbgEztpOzy+Pa3pJxcyMqPy5AXD4dFEUUhZBg50LV1GCgd6Io4OsjGdUviNtWcrKxuyBOkS5Vs
KNOXUQlDrFknEgMYZ0/HR85w9StkLn0WX21JXceaDfxG4L8fE1PvGgiTXaXHtgtOURiJni6UqDUx
HjiI6iI+X3r0jdkEy1RvLU+33Cc+6aK6kMtJMtoy1ZOzZSGxiO2mrvQtiSxeZrSxPsz8aJpC6ljx
z2VjzELiSbwE3uIQqzL0ow9MjRodGuncEHcKl9z6ZcqdMBv+DxXYpv8YUJOEEBS21L/X6C7TER1B
glsNypOsubrfdkfrfjZIBekzqPBjQqfP/5M260v/yvFBOaFdRYStqDIyKnGGinmSEkIuRZfGc7IB
FqKJEjoMDSZe/ES4x2DfvlznFYPlioG6xf06czf3YDUEz4+tvfco1w1wKfEDMkAsjEL2DovqWDrY
dmhl1CLytaOERI+RxK/ZFGPNMNG0PL9PIXLuTo84C37/7a2gPLATwmcKwFOjuUOuQFNDhCuMEB7q
sWiO9Ho3ftWB0HcMpN3nyWFIwCMIBYHyZWnt9dL/CLFZFPajSegRHW6D34UBZ55DPKzpE32LxycT
So91AfdwLAnZQdH477aVlLlEIT/h21IERuiMX/N92sWCSmjjgEkkGlq9SrOBkGjDUnmrT+NFN39s
7Tjc2duEUXNqhotCN24raC50ozQhkzQ+mt2x7pwuj6Q+3KGh84juNEcykx3nwRRBFC1RgyRbuKjO
Ypzd2w2rZtbmwdt/uXoDzFBSzYU9nMSETgSL8xjQZqlwigdaHzODIhGtMzaqgLkuCDhoCW5aG7eg
l5IxPYs8w4RCYtIJpFPxJ08meKq19iMOKgiw/WuTFJFT20Hy810oRc9P9Zf12Fq9POAwCpsRIhug
IV8Wy+F7QrkjctS9JbEnTSw64L0pLbwmcT2kTK+sFLAWDLPv7pBkV8L3VFHeilyhAcjM1ZHcPrim
Mvxjm0iPjUbWDk8dyblKj5jPoaepNEjy6pagsa2VoNpfehZwN88vtzwyaCOxJfeYZzUPSPSA3yLQ
BMYRaiWfCBjnZs6u4cp37P0adGQljqSQdKFNBqm8ypOGG4KpSV/S2qWiU0xjugamQmjxA7NcAX4v
CgrJ6CMvvP20gzhe+ko3Nycim6zp5NqkoVtSMEsXGwB9dKAw1Pr4p6yDsQSBXAfyGxmQPGLkfUy0
5JMvJos+0FW5cwKtDGCWGQnrchlPsCnrkNCUGGp4+vKbpRPfIFcQ7/kMwC7BHe+bzgpqR4k+vade
kriVCQ6nNqgTnlf2hMfvT1AqEz06pCYArDtdIkfmP2an7pa8jbCjFVDM0MN48yS0Cu4zkcXqt4k6
6hCRU4DyyrbpO8GvHu9WKxFv3z9TEcY380v1Nxnp6btaH0XuOaBprVmgYyXRvvM7nq0R0YzOR/xf
+w8KBfOXhrQHxPdI+Wt+5s0bK/QDiMooO4XMLA2CdKtYcx9bX9MGeqhb9CBdfDk5ZvM6iQCEjReR
DDZUx8A5f64usv0R9admcfvkjtR3dY2fOYPQ5fTvvqAXHjQk9XIXKlFxzIunPj2SCTGyw4HQEkyb
yAINYfI9Z4KmuIVnlmPP9RFJR96rlqZXBwbKpGZ1P+6aZUO52PTOqBo9tciSxSR/BeBMgp5OU5fY
tsejOoIkLJI85eCvOeurPyzqjnrzC2ujCbbqRKoVJzLgfqKVV1ssOPeDWpH+rCsC+Wxx+zcAZXUp
Z4TwgzDKs6IuAexUTyi12iB8qUXd5D5Uit/xDHxAx2zDbAI8E3HRAGqA04vqMixyKU5lIDrL+IFo
8i7A1u3juP2aoqdM4bj6bSYyZ95Q8wrzKrhTaKINmMbdNnrXPXq4DsI6Cpnh7OD/IPZh8yGE4iYD
9hCcBeEzwgI5qe0U6/6de6eplWpiKaWXmMQZMuqnj5nCjadOUFxFvshXvqjdHA/qbWZKNZwxcjUG
uhgA2z7xWMn44zuKZoUNZKtb2kE3rVnTih3dAw7ssyqDqxdW1qLXquxDMET2hChTBvWVgpAhOCfT
MV8w6xN3FWAbcZrfyRdST9yOPgAE9zjx+GZLVySFM3lTDmCTRL0eGOe7fCuuITDAnhwuoD//mCZd
xlArEGG+BD07xUOD0Wbh9S/q/2lDfeGSoFHQ/ttcDr5OGFaHf3r1EYdC1gORANIhoUqWSDNF774q
OTimvqv/FOilPxPgDw4rMa0vwtZmepC18Zo5ai+3muFKBeY5CUZpEo5Oef7+pp7HnszCeOGLjKFi
i2Y3W7pNZrYk4rktYLAYjlfXkVxeRXZo0RsQXwEspwwxe9EIOzLsyLiW8OwJu5GLHNrD0/0vxc3J
Tfif4jhjGXDn1X7daOmXfBk3TE0dQi/aCtFq+F0JESQjmt9rMXmQfC2cQ5vRFzoq2mpjZWF7/nsk
wvmHP2XZWLL8Rn3mlSY1v06uIif39HWe0ONBxH59CeZx044gtFJNx61tyb1tIByYP9hcEN1NW4ft
zATcZ/ThhrwohZuVblWFMW+dJhdRV0mgzwBtAmy9VYLkmsB91gavniYqFwmBzwBZfGj1aFbsxFaj
9MysFeuHECGz/+sliIOklPDmAIbsNDEZHJQobf5YiofMLPATJYGJ8Q8aDc9xLKN5lHy6hsLfe651
CjIhobPUPLJZ42a9QKrkWAERQ/eucTFn040M0Q9AKfZCk4Ri0LxqYE6kZbE5/vGiPCNlWa+vP8G8
4ilq4DINKe4bR3+KGv6QA7xB/u57c6aGwbQnKSeEfXfeLWU9dOAiTuIxGq1deeFrYIMqKh38TEfs
hA/fPEggxN4fjShOxmBANGwVclEvbtA3ZnpntWjRq4j//wcuV+Zyc4qdbGRJudNK6030rKfkG7pM
8zU/KGSUMqJWM5CRfM+l3l+W4kJLnR/+ppc/w3ypvCynd6b34nQCVc31z8NrH28Q7otcHKuOoFgu
Al8Pa4yh6jPGRZQDsOcuYgGURmMVzreFfySyZZd9Ga+wtrHNfKQYfS0ducWV2UlM6J+IgPqw/67m
BdhsSvT1tim7n7aHJ1xu799sxgHljtij0Q53By7SF0HWdG7mAqapgPAGUlIr+lHaWeovsMDwcJl6
UotuEEbogRhuJJmxK6+MVd2CYW5upHrOivAnlxlO8teyAf4d1QPma+1KasOpM/br6NKeZbPt/paH
cfksdQBUYYMuNCtIj5Atj5UY5XWnjIOBNabCYCKzV8oJeXomJWOZ9gyM23pd97YGDJrGr5VEBw2l
GXER1HH/D1+lemSL8g6meMuNLxbytkgAnrM25IXmaes683Lcv1UYJp4c3Bie2NpZDm87qht7Mqu/
AQLBs1rNfajOanzWBW327I/7YRnM5Cl5oPiyDAvQW8ZFs/ETpG8KH8/XYCQTCT4AMzIDs1kvxZum
SmFj0y+GsY4NLVPOFjz+0G3Qo3z1eJBbkCB5tu3AUpozegJUqcVVczoPOlAiYOp3lym+4j2eC7gk
HsQjsG9vXsINN41ruxTEjtj9znlQRRy8SU6EbsJcS3VMqemQvmYjcS42KfPypRIxDoy6Pf5k3nfD
awmc+IMLL4KPF0a3zPEInp+3rM4aFPZ5o1R5mFSrRw6JMuSgk5Wu+UhhqazuxUK0nJkwYtBaAM8E
DgQfJSxg4dqg0E6cHBovuXETQPmqvQyFlzgUT0qA93Hh4VjVIuQjX/5ltUMJjld1+DzrkfZe/w8E
SY1sW37pPviVjD62t3S30qoUOdngB7sgJodgQ/TMyncfKLCX2jt/vam2+cIBx9tVEH414E0lwNR2
Y12eRrOOMzOWORP2r2II02ERtz30PtkRx+Uvo1F8/R6vhpp/YDrTjerqfOg2mCrXgCYyNeD7DTY1
HpJgz+ofmRAcL8V79K3vBlC0c5+puPrEiz6nZ6xHL/dR5HyuZhnmWKI6yPHSWuTw5+yRscIVWlg8
s8RhNV7xeOPbDrmUy7ZWyttpRXW8U6bcUokwpmdHsY2K8HQVxgVZNd5EYFp2FKJWZZACqdQVV1mq
zwAf5gJfTPNWzIEaMVMhBfY+wR/X1ZxNNFWaaDtrmt6KwBsBZ9W50CyvX4iQylkeNoHrJK8c0ADV
uocEtLkKmjjjKSNSonwBLHyQmWDzINwx/an0P3dw/bcYmxrmWIPL/O8tGbl753PgDeVsFp1VpL20
lPlvUdPOj7GXeZwtR5ifvwaikBKEO3+EcGvPJc7ecOY77ODPySgrW1qzyGw4nTKqFVoMSlhPdkj9
GQnsFrYmjZ4/RFCJzQ8fqfn62lL+fQX6fQnuFwybzzaWzI1gZKjsAk2tHzwPhxo5BaLgQ7+60A6w
+GXXOW186pB+KVndequv9u81l/4b3OZosM3QlECFkowpLP3B45OHWekXrfI9brwGf3hmm6+YF1h4
nO7zqxn82wBcp671SNkgyz27/Ovx8itw7QkFhGs+sTBWpRI+iM4y0CmjRe9pHihXdDT6XPs1wyew
NuDXbKjVxMveVgw6ekbZ5lI2/1K0DS2Y8ReGQfeSpUyeot6bm/MJhAiewzlzcRyePxvZYNnS/lu1
qxT9MUMA92B43oxNlhKEAilrN7fw0IL9FlPJe/zfS90MO9dwcIauaBeR6oh3ufPGe2LIRUXq9nVA
X0MXoPcK+TqygtCbASbL3ZC/7lGw9v6oYeJlnXM7tMvQ/lBSazclOqPP5gsuYGw7YhQ8qVpF2vHy
mXH2680CuhCZd9xdnjGBs6waNIsUWCiQdwHp+zVIPIWGSBNEMNHrX87OqgBajmzbRCzOrOBJP2ZI
C5tolkuqEgRdEiM4065yfS1e7tJ5KsCnYgIhieRbyFapuwN0qweo9Ar0Rgf+T3dkts++99dIFuvz
bOKjtk3Qu0UTHyWQJYKkHDZrg8W285hkz/zFWyyYjHjWEsxOPU8BFlU55YfqsoBJDZNvKF3ZbTW6
dLkhFJ4XoogGeH+yIUTUQGKvyhlP9UbGQUbnY+yoa7dYhtENAS6KmMG1bY5bb5o6ueHGPFurj2Xp
7UwbjLr3kNK94VxWRYKkLo/ctlvN2YpK+C8S8EAzsCZYRTgSTJR+8Fhka5coFDgb6xwwouCKHLFT
mOGybcSX0ZXd7wDE/Pcys3uWJ74lSa8Qo7Nvj09s4/RMAHtecNrdfzFeYd8PT3+i9c+HwAi1VrPr
gvhqJcxQIv3ue4cFzeB4mdQULXx9kp9toA2o1fSCEJPCJe6XglT6Wkx5wBLtUHykx+Am3SHMJR3H
jQKZ2SR3W8mqfwIFyX4RkpfRzZIyMf0CjMHFEK/SY1k7iipQcFwK8i/2JpHZwGixhl31X110RgkD
rxXrt1kS4GtaaptsjZtYUhwejceJrx2rNi60aoaepTna+DpRwSHh0wULpob/21S8BVd2vNTN2rul
tKSoc/XiG0veZkgTgoCNlekCR4yesaQhREAYd7av7BPbt8oizDcTjZ1cLTNlm3FdAbTwV2g/TuWY
G1dkGGh/xjaYhkHYmP1aIWbA9MPpOkc7RISv/jRgZ1Wpghv8aFzB11K4NwMRqZtrkmbUn7Wc0WuT
ktmO1hpqMSFku1Tz4uS0WjKENFOlAC54JlTzSaiJVENBCBHzZoSgXXTqEZdlBb+n++Soawp9U5Rl
l5piemC+MKhuUMmgmscSFnEVKOLIWJR7Z3H7aulsxSNum3RTJkfGjsMDuSiRIXIePBK3Vr+C9hnq
VBVALZkWcYFCSK8QR5boQanwRIMeFiIJ0v474H3yfx224HY1wWrKR4jaZMqOsgvblFR373Risgyg
uenpnd1OBjKCw7DCrlv78jRRDTqfSB4eWy0hXKcSTFeMEqEU98jcHzUDjFDzGLi2LMD0puSWZi72
SCaniaq1DlrRiAYlQGVkcO+qSFYvfZiz7FjPGUe1nHSNQXATiN7jAu+pckNyr2++1WgnGyrkHyGm
AaUmT0XhS1W9lH4vSH2wV4C3ksvu21dn58Ns1dKSXAAd2bkUPuEdJZFaeNpU3KRoDj8tQdawLze/
XFejcBxEpCv7Eb4I5ar0nnX2AVTCGmV1Cp0b+PufGiL2W9SWQ9qwINmkBxd79dXlfikMbIW4+ZfI
LIy7R8EbcLxa01GuR/yedkjleJVpL5SVPberfP1tTrocsX90wBK0U4UIoTtkROvMzGXKTwoRFxqu
PUiY84nj0xK0qMpigox+gXUH/hap25tZQV4W2LE3+7s6sfzHuVjFFEEr5UA2o+1BUCbUNrELlX6H
Lv4SzvHJih4T9EbbqslXxIZeivO96ZzdmyqPcU2zVEs2LVoAccWB2R55kLn8kNLF27WM4azDU16Z
WflW1lbZmvfIdNi/RGC0Ug7U6r0epEK18+yDC+9+s2R549gjWe5Dv1128N9V21T//YnxzYyK4/2h
1AZrxlvEKSp1slTeRO2sMAjlaEY2qmVBQ1Me0VGpilfbGBOTcN9173eAh8Ff1FXXjS2xMLBawWsr
o9jrfHsHKYeV6/eZrNjznSMqKZ2cHF4l7YMjPeqqp2n6lyDJkl4Um/a/XIFw+tPJJR9z+0cDMh/A
AJ+5UhQb/gJyLqivBcnXiN6bNNQM0Vl5HyPq9EaOwrhgVCAl/QGvg6tffTFO2/QaEym79co/vCKr
HCETLlL21IiuN3n9mxBGiyWx+NfkCxOiItmGrV047RltD+4EyOxhkng/Evtc6nni89rLonUVWCFa
5WGcOCImpJsLDFRzEaPLXEdGnD7Qr/VNplD+rd0xUETso4ZJjKYTck4qIjUhSbY1MtQ6HAWiUAkC
2m5UPJ3Gc3MIcWd8br4flucUwHzd2010DbE6sZlQijqvGUJxs1CLq01kzuqJzMGZbrXtHYW1BX81
XwleQ/FsDJaHXmsQm0TZxEKorpHd4xHGZs7nRQg+IIrfWE6hQCL/7OJ11QeBbWzmz7v2ZzBaEM6O
mIUqznyKvq9vkRGUU1UTvyqEn1NLMjPb0W3vM1M3v1IKW1aWCm/gngfl0Wc87Io/7Avsa/yG+0RT
5Kl/2GdJ+IlvBsJYcOM8xL3KR4WrmAsKdD/5Ao2Hd8Pq6cjCjjVxJrO5A5HOmZZUzVflYdRgHUQr
5s3s/zNZDNZq7SRubzcWcXyl1so371LT61mJLV2KvpFLp5pJa1y2yXgouWm4pDLizJb4uvu14Yd3
QtEHOCxDu9yzRAFgGsw+MZuQ4pBwzVlVA7iZot1HT7cvxpWwiqXN0YtRfnd0iAltJX5SftDSDUQt
hMOoP3Lvnlur4pnGWvZkvE8H+N2ayk+3Q+/hUyfp9CqNHejoE7V1rtx6sXtFC3jx/x5Tv1aAQ420
/VBR+QSlYWZWjwe0nr17bEEFeA+fiWRJe2k70RrYzqGMIjrrrAXjVNzhe4HM3ewsQ68qsDKfRleh
dwE5QqvyrScKhWd+HHNcUpXjKUfdVaiKSbhS5PFGT2rY5yY/YJKZjZTm/8D1mTKotwRLr9d9urtJ
kAGimIwbLuxSQJn2QiuvOUXt4pqxmJF/ZTIWMQKDVDLT6dDyzjcbUxXXKyIbhS1mfZj6QSvWw3vy
2tRrP8h16c/5JI1PQawqPJyLmRTPakyVLB2InM6vPojHT9YUOAtD65kWMAolfghbwjR140HmvIpq
4oxEMRiSXzlpaNvsYEVPJpiGO2GDgvAE/3TBoUu3OnOFW68CDVSwns8FYsZdT2ZuSnEiZhnVOn9X
e5+5SwefgSZhv+QFFfx77U3saBk8q4/eGfumyMak0dQUc5E3d4/UVhBRI0rfWVpUAtkou2Bti5rk
LGTxSkP3QuOlloET3AQf7xIhqDslmL839m9WHoJp/GtLvFu/nrPwCmKLklv2uK8Zp6yIqdQWtLr9
MMfwzXvMxgSwZ3PLcw6Bs/6LX23JUUwYqIM2q3VCJTlAgMuPApRFG7pPoA1mOrc91X/B5T+94ZRs
LlOWFKsuFqBk6Gqh+N30gv62OTOVh3M7otOED94/58wAkacYZLc7Q7i0iY8wkZczHNuB+8H6IyP2
XGGZKIPvtRBx+ANdZquyf4BL+RV82pvkTmgWprUvbM6Odixqs3g0PxYCtnf0bpK2x+bpYKqK8r3o
6GWObOmg7yurrLqWx1NkhCRioxAL1dSnat5221ks3Aw/j0LBuokeOEakiCgcimehSkuIodVAGoGV
JmoxoZ9sYFTM2XDmS64gW1EwNMrhWxJCOz7wWqASpOarhcf7dXCYvCSh87V5zkBIdaDvirLanLBH
K0XkJs6wf5QOKUGa62Jyau6CaQWnO3RccvQE8Re/0d3JomlOc/SB3tG8gj+gK7zlG9prazmD2yu8
7x/yn3kMkxrcJias1afHGyFG41mws7vqX309nyJXx8+tIlDZqXgTpsk3xfM6QX/vXd7mCqtZRm9s
WfmKe+Z/1I0QCqCE78hNz979b40V+hkv3Ga25hA7/0MHFiuFjgduIUjXsGEPvgQwFh0rsnu/75Lz
fmEPT72U2DHxMNlZB8OHsRb3pzFZ1QpqGhE0/JHwh51IgCo1QE3zIgYXG8RpcThaxImuZyEag54W
nFyYMe+VGNIJoWIHSSWqRCh4mHNvgI3bsbBIviOsfZt4U1RlxEjr0LF2wMTZ+B+0HvAmxLFsmWQD
vzUVlhfHzB///KztfTPHPYsdBsfFAKPlLu1ZYTP2bU/gLd+V5NXCGuJjPnwRdv+m9Kn5m5cHr6zK
3aGLZR1wOPHhK+KH6JogbKrETnXafAXih2L7ZEOtOGE+vCSNscHKpbLu+DT3HNxE+rZDjx0LM5io
S7UxQZkJN6ph36uO91glWWI9LK1CIUMVNoNwKt+Zn92OUtHOsw9ETMp+Z03rcwmO66lPk1DCSy67
hQFDKFxp3u07JrNxMgoEkZiq2fZuQM7PFgi9wdnD/TUOk07Lgi5OTYO+o0yWdsp8KM8Hff8vPsCd
tCjOAC9bYffOp+W4kMb5q+dn5GEFMovwlzdtdlfRMqV0ggKdUnPbfRtqbHY81n49mEM72Gz0ovIi
f+FzKtqO4dYS9A5eCxxthKRn31DXmjT6Kk5JG19waakrZt0llUyUWDKmor78hZod8JukMlDgZw4D
O/m+HTbEAv0pVOCMT9Y4FDr9zS8DVwrOqaX0EkBP1rxI3Sxy9LfxujhWnXYS5Ga3iPeL+GWl5OG7
DDqy8Qw/XaszfZQ28XREkMNZ1MBzm/ACt4E8CShXV/Ic3e2TWTv3sfIppcfRVGEcLxFdVynngmG8
4x7bleEfiYgh3gA9ZEPz8zrEWOoEby56gUE0RGqN32yw+WtvmOEq3zwqMS3sRj+f5UkcxKMhONpM
suujvcFOzU+ha0oWsd+rzr2y0xosHbZlL5Qt8aqY0Y4ptXombRwpRdCZZ6XAktXtrOoj5IGUPGZ4
3Cw3puehCClio77eZ9DONk0PW6V18Tx8+3pcYfGAxR55dl8l71qaMbpb34gaugAYwaSlb5xlA2Di
TI4frApOWmYf5aT0JhlBUA3sEriCdEPP6I+Nc2zF1lGP7u/GlN6/+67j6hEWxvZvKqQh8GnD3oG7
hajQbXauBZWVvL+oKKbzO6piMSyh0g0ERJFBeooDNc6uE41TsG11w5HqWd2ugiRmLOXjdsG3E4zc
icaw15C5QwphSzi/1Rm47kV96kpwoMPeqhTmB5YWoNRT95qv7TmRawSESStTm45M/mdoMXQ21EEE
otOVqJq8yazl+rrsGkNAZrfT5w1y34HDHx0tAPdn2SSbkI44heeKfXCY5fZOYTF8Oqy7pvyvJ/oM
R8rMAdqkmK4QUr5zB384UX+qy0OGc89TpOAOAdhj1NfJRSPGHtxnS2ILO5WfntKfa9lULVk9G6NC
3nzbEZsiF615jOnYwrU+VLk9DLpMVvAvbjNaRWn5uvyNKDrYw4LcDp7wi6TFyLb7uA9DyvRobI9Z
NQ1w94cKVVZGcBzOVvmkUtEMeJ15r6UPOhoqnCZsfItbQdQxFC3pCWMqz01O9z0eW++JnP2N8uXA
NVm7uvSGyE1P2KdMfxiCZuruHpHQVjpAKAtfzqHYGpmT1Q4Fe+A/XPSYUgLCznBnSepJFVIQTGmT
Qq8EIyhFcrgYt+65hEQLdOxvY6rAoOhBqQ9lTk5PRPBiPbbm68hms29V5AxWL0U8ykIzRjMxmCIb
OoXVrnDwilVI6J6a1fjHh3YNYIG9p3hgoluST+h/WvsrDYhVFAMqSJi9d7I6PW4hJKDUk03mcpnB
r/+EkrzPRH5nenk03HzMnTnj4NL3twpC1h+qg3vSM8bINoDUVx+LnwXTiuuOIc35VJ6/GRR4A/20
N2LX7yAwyW1aDogGwwM7Tbo/F8sBLCdTjqqNqrHYxGGcRBStj3iWr0+EesJjm8jVm20bHBVQwRE6
y87PYQsAyICgRJFMHloZygshuws5JWKRz+Pd5eQXEZ7w423afjEfG1dCZL/v+EwrFmrl3jQKPhc5
3seoCSWx4sPu5H6jNyo9pHhyrtMLfOp8VsUEK9R0qzeW8ffqLVRliVaiPvM8YeN1pEho2gH+9xHZ
PtyPbi3f/OmRW5zYeFkvGgV2amNxXk+a42r26dKEJe7rj3CCeb+qdgWGrVyId/aF+B0VpRV9xVci
q7Bhek+lxIBTtZFjA50fiOPD5Tv/1JHn35MOslQMt5wqsH/4aRiiYMCeHXA9viRsyVIfP37YoXNz
FmoEXBIluwClP626c2NLa1eNTQuiCXoW0LhBkfH/2/bQ0qjKpL6yXt+vK5+EkEeP5gNlX3csxz1j
rFJW7jA9yJodYT/+WU2cN3AZyuINIuQeHdfBbPN1iYQTvgXUn1cOTkt3hMANRS3M7njGgPFoMSKY
MUCwVohSYzV3RDwPLPM4ulJkqZEvLcs8/9073BbErhJWu+UbXEk0afZcUh2/2C6N7RB6P0QUx7Ns
O7zoScQUX5MB8O5XA+6UWGvppowPRPjou/YQiA2I197EapfmN3f3cpXfINjzv2ymdE4u537vDLR4
CjJCyNerIG+euRAQVLnEEtJ+8+uj5yPAGrhsYGNJEYKcomAu1gWO4Srx7wXq/+5oNXOasZAFpnT3
366sHobqM1/hra1NJ1NH8ZayoCB4vBcBkt967BqeF5wqArRcmsk2cTwvMnzLJ3eH5+DjogR5QfAO
5+qlw97K4lGjLQx9uOIL0dQeusZ8V2wkYEThN5xuwEjCV163JKEsvtw41DtPcafif1JCiYAM1kuQ
th7pQkY00AmWDdUK18wYozIBjRM87ijQR9mHaJjG15G6dt69E7w0PaMy6/DuZgHBYkApjgroa9LS
/a2SXdjllQW038dVmmUJecyvMgBcO12KVxF0hWjB4uecGeXxdexoOEaWsrQ9o6LVI3KoIndxWEJZ
Nns40GPD+CQE+ZlxcG1IcuDZI6le+owRFRHTuU7FeDjFz+ijfYI16m4zCS/j9Ym6y9ihRNESQvdw
DX2fEX35g078U3G01B+w5d3ugQJQ+n8yjD02FsXGgJcfF1ELPtTDPLmSwmGLfnHcIRBYf/QWGyQl
1Ub4DPjN9VV2PB8pfX8SuZJCx0BRy2HmHrYHdZA+HrwwfFxXCbOSfV/KiYklQ3nKyDfKDrnbCZVC
TTFgt/hib9CuUJUIWjx8rrbmPOxThowE/s0N2+wXdhFiHxOkE57nF3UPCNj/I1R+lVaFbxl+bTGz
4fsYtb1OQ00ABw8NnKs7DFM9sEeRkgL8q9G8JSTuhYF4lbFs06/RZnhx5uZ8TtiMcoqFjvy8g273
4cDAxARcFBg5E0Uw4OpSVnGRB1M9BhTcW2laF2nPuYv8FN2g3wkcWyAtL2El9KSn1y2WVuwukmra
KGbWkWG++KgO2ZQ+Aw+wuOMsT1cP3J+/jrjL8oaFf8Qnr3VriAzxCgALZX5TxFwGreMW3Qj2emj/
VHBazcxGnp3s6IO3FQk3VpKwwlPcCQc997v5Kjzry9dvBp42iMGyUdcoLoGwwm9qo210SExKoxcx
CEDMXGV+T8x1SAoAzaBzpf6Vaj6t9KtloXRMOZ6vFwx4cFdaplct/PVFlDe1OLv3znpHSToyccv3
l73KnWCAAM+ps2c4IGXZ8t7tkp4VgVIi5xoCwJOAVpmXJ2Uaxv5VS1GEbv4Run0t001L2TW7igy5
iOU6qlpirmEAMYbe+OTTONt5JRtKb8SRBXY+E+e1l0zqkrDDl4Tt6J8qU4CA9f8qLfnt56aNodU/
xWwrwIvuouPfrd18BAsaIV0P+b4Xgk4Q9Y3VOrFt1fTuNCBG8FI+aXjCq7p9+9C0MBVtZCnNslHH
csIKqJvawVYOrgUB4lH1uL9/DQsyZSovKq6CMId+rSK22gd4H+Xnwo39Nt3jQUkVCV362fidqbdu
kpOyo9ezG3hNbREWY+UzQnHv6hH6VcARoc0U73//r1RYVJOCHs4018c5WT/XXKJnCYg47pUhn6CG
g2SdcVyNiHQLoCxEQiCJLvmp99xo8hv/65gz+Pv6i+ybcQwlrNpfTu0JQbX3F/doD8VlAWh1bVPZ
OkXINHRTNluxhzxjUEDB5cGZsUFOdX98GryGWD5xDaeugwXheaVPr1Nb6+M+SBQyq89kz0PA/9i/
jIMjlJ4z7AmE43LXJyvKU/k4Nr+ZfgYN5fuT6bJnyFVytcNXKc4IRAPlTa8/zfh5kY/tfXnLqS6O
RGqXkdNdS+Y6R+IjvWq9gzL7SSiiR81wUy0LMTZgetVikESo//lhs3OUs58DeE7G6/eL9yOILc3t
1j+OE6RvaSM3JfxuqERZJX4Qt9k+Q0bZmLijOUlM29PhwX33DVmzGcqMAdWbKcJGzTE+E63+pLIg
3XY2Kgd2XswXaJznfVndZhlH/Di74AFcgxw7AxGwDmBsqesiE1cwyqEAIwuJebVYVMSuyhCCkdOu
S3J+9hCROpM7ILNHMjd7HLtG3YiGjdkLJijh0bzAbW9NuZpBHiwaAvhZJFYofTx6vaFNwnwsJg0B
JIvSZJe3HwH3nbDHI5jymDREaM6b5IiDNVQff1oOQRZBrcZjsA2ogsij0eFksONZoAYkjXtYi3+N
hu0IIbkoKfNdIlMSJs2vTx8f8AhsFIAI3t7CylkYPxbyf64Yj1eurdCPJm66bdaYRVX49uArV7g3
YzeusD8iDoqlfmiWdwR1mMgK3f9xTyAm5xaYFrRMWcB7j1SLVVNNRHH0STV5ndh8iGmF9xDncw1W
CA3ipfwXLl2OfdhknnmRtgFuwVMACfmaIfADego8oGCjzL0DEgc3U6HIOaTZbuy4gM9EdIZ2fICS
tX3gAFsto9KicXiqus8aAmf0ICfVcvyF6y5Kbazx2iZYfPbQ6e6QPQD/xbnXCUYzetJbcO9BFFK4
D0V/s17oumlS06Ho9N8aW2sS4L8bPx1yyQ1y4oxZk1rQu0yRIiaJRPclmn2IsHwY7QGX7NRHKeeD
w7CV+gVMCFdaL0HOpYlsZz+Tlodut7RENm5/YJLxR29c86fAW3BKQCT6VY5r8oJiCUDiiRcN6ZRa
KAd8L4g0Z+pLsIpcCZZWuSc+CwD1ysIpfxCi4Ks/2aigE9MyhodZ+UmiB1d/C1p5uHHqcjMl8Of0
/LKS2v4hMK7LWeUjYMdtybpSAfKxDgjRBWpMAWAxNDfLJrLDC1YPk19L1kcdoK3tWDqWUL+602P+
3RhLLqrZm3+mBwS/4TZF2x89Sai0bJ8kePWimfewWUuaPsxrac9Z9CdB25MrnDcPEGWTuTeaSntM
LsizPdZ4bWkJ/mYbbzqs8JUKSE0/LdXLpz1G26WCrEdFRaffMay0W/XxfU8NtuqmjcnEZuGCX1Ed
Kc17nsGt8M+p4ldlW/dgmXhQltEwOrdn5fiXvO+M2htSLPdMhYK0Sa7PW+vUN1Lf/3LFyLgTd+HJ
0gvYDxIcJBAsEg7h+uXenN9IJ4i0UgKvj/BFsBzRCwko5R9PWyD7a5Ky53fKUuRzOhQx/vFqBEni
dxdPlnTWkCZbHYeOF/3JbdMb973pq8ZQpcHhqxPhXpMYqVNrs5JCqrE8PGsTkEfUzJ5dZMEXJbMH
fcSKpIaPHta8oJRtQz1OGrUoRmBf/4TKTPH0c5erARiyFverNys0jw35yohjZuGgSy1Sfd40g34N
Cb3yiCfKhxMP5y0HqMMfXtO0DInIUOh/4VFl82l7IHyY7yME1aaWHpqqzTuw5nY4d0Mh4er2Rme6
WUazxXkuHk3LMWpJnAOsXYXosXPQuu7Og31Ns5JPxIAuW10OedeFO94/xjUDHQrkjdaNFWYndAGQ
RvTT+ORBiZzAmo3HfmBEmT56+Dqe0OXQlnqHqmSe0kc6L900Mi7oXP7Ttnp0vmFtKVXOd9cNvLCh
eJg6jkAGiRjzsJBFQKSW0pjaRHCW38mM+IH94rGOqyhWnm/YIyL3W9QgegB6yWXdGYXIBbZvIkZz
0VbZk0uydkf4myBssvbZyboMc2QTfEpt/oiracoXz34wvWAn21r131H5wBelxlLvFQQZEjrRmpCs
DuSEBX4dBYbguhIkxQJy1JuOLZ2rEXHFnGcl/gLLqbde9NFVxUfQBI7M7+GKih6n/3oI1Sk1OyAu
BhTi0YAGQNhKSFg/ZWEW7lJ/9VATTVodew4pUImHoXUClPG55eQsegJyalLwWODFZT/n2ae4a20R
1C3HGkd3TEspKyA+fFLxhi23SmRK8mQzv0povkvqZh/uDZcwH/6c0kVywUr0yLfjZ8j6VVmwNCrF
FKcfdhNczAamp7h2J8SZ6+cpCkCFaNjJQ7Re9SGyBXwv7mtyVCg0x1Inux+TGanawaZxaxvX1saN
RXCjYq5H8rQpsqpAsSpn4QF0R1AK/YhMgy2wlvBQ8nrM9rsLu88CVzK/FQ4mkDyeoKUoWVH4MwLL
+oYhq030CXTfBNd3JaNM0djiF5AevoHlBL03hVNHHEcMmrtudjOLVeHU1hpI35YQOypvl9h4kySu
QkRMh/HbVw6ABgK5X45AVlUfKS4KAhLhMxwJY/HRvxYFX4fnCSYFGU1PSOrHSWyxCjFNcGc2ZfG5
bhhL2NwlsnNkqKCpJRUWanF77nFTh30Jwen0wf+B5hDOpWleQKNBJNhaOObaftAQrVQdBbmBZgVt
dyqXXB8yfDC6AHBKOQjDpzuWqtetwJMoWzPVYX2UiwUYPU6lA4K7wEvmK9AVAHK/04MAh5V2EkFA
FssIeXASKeBvJ3wt67HnhhSj79kUM5fm6iwV8HwEEJo7kJ85Jz4iwnOrd5wa6PtookS5WpPODfGN
aa3TBSL9+5bxxBzlgDfoFt5QvGgem2wo26JdNPxK+KnxGvyXmhv0qMe+eoeaQjZ2nXyQSL3AHZFF
6FKCaVJMtt2nFayh7xavEFWJyuPtnwI3vr649Zedp+/KzuP9aRFcI8kImmVfyVmGpkECZ9aiTBcK
1DESYXTbSk6iIjcnvXCEuHjgwJeKGPnl7Epp7bYHPajObcrLP7rqqRk4AtdbRjmQOvRW2f8wKxkT
Ugo05FndgxaiH99/UcZRaQrDwI5ZMJw6yzlpt/k+yv69Hi6wpZvFk9idoFM2qmO+yRStTZ2q98ti
6D8MsxzeCvNF9UvrVIYdur8cK2BI/8cgNkAeZfT00Ve9n/pY2WDwUwmLIXsaJfspa0SHXm7YzMks
qj5EoupT/f+apA4thXjCku/60T9421L+CsKryVyKE4+SD9IXfzaNk0YEQ4HRA3mID5X342O40Q5G
ChFgdA3sAyPn9FFO5dZ5fwP2/iC88YlzCQANBpd4fC3FvPml8DUuWzy5gmyaXQlfPAz7uC90wbJK
3GvDxeSRsdjAMrFGwQUXiOX2pxySu5cAT7+fbswJd1sIqWm+jrdoKsqDpNLMtqDzO1+71KPGTqRE
OfZexbZiPoCfQvPIlWRK8MIuU6vXJrpKZjLJnM+RhFacH1UMnhs4ljoT0bfK8gwzXeNZNrMsQYKk
djBedUQW2KRqzv9s8RSWGJM89HT6QDLWlo9b/zeUtgyQbKlZ2uI0PKNs0D/D0oQaXxCoufe4C3aX
vSu6O1dllRdueI4HWgtzOxRjDDMS832eIOodM3qEjAVbzyHnHrmSiq3iQUaM2IONNuKxyZsHiQqz
9lLh43G0DOdY+bh9oBtE2RNDyq3lPKzEo8bxkC0uKTEi9uAbR5aEIdNo0UbKhh+vEUoQNvPIBDJB
4qBhwT/vKiLk9n/Wfv+jr7/GpxXfADeWr+Miwz5YT2y2PzUKyu4EgCkdg7o3MwFyl6rCgTB4DCX1
rKDvIdLiZxazYRqbLuYN7CxzJcRFvN6b4L8vDQpG9ss7Vu/4TGr0Jajg8oBau7KhQzKLmgiPLqDV
bK/gEXyV0DI0Qtzni2CFIf+KfWc0AshmerTBwQ+IJSN/3MeLJcVWUs28ceRDGBIeqHe0aRE+Y/S6
2OWxBHdvZTByxRwExmSSSwgcE9NSsJTLphkk/93x8SFJhmDmspLSmD3sx2341opA5jK+8T9DurpQ
/GC9ycSkVxRNgDugO7NW4WUKeJAsIssdaaNQLAU/O/ZSEpmSfUJMKIG0HQmDjLE4DYqruBJaJUec
WZUV3ZCYsZcTzpO9M8LwRBHR/WuSAwG1uSgm/XabOg8PBxRsUH9BbvEe/ZkAWDecumnO+AKzxTp5
xoSiTOqHTxzkRA0Ul7Sb+JFTLUZUmqOUNgtm8KylxkqbgX1pLyDfIRiYhcClFfYr9Rwkua3zzY7N
ioQqBzy/9XEeL3rsFjXi9utivM0IYrsVDHUwlqNt17+p5EnN6DFAVygvHHAwYOErFZdfLVyTebTC
fhyssoG8r0Yv9xLQIb8n/9Rp24104SSE7PR7fZZF2u/6JLPtG+bnvbehWJ9Lzit5yivweclL/G42
94K5NQjD1p1oy7y9pqCE/nQjrp9eDxLDk8xE+zMEjgMmLpPCO+VdCyeOv4xNC7yX1g9gey4aftkF
HNJx8+5L9v9ZmUpeCYyFWdbCWEDo/encQw91FBVQqqghqNoHZT73kCLX+PE31aTXVCPvdEvA3tlZ
M3e8JXC0ikgMTPNTaUai4HRxLzAlxkPA/+kQ2+AWZ4PCKto5ho+ZUj7atmvAi23PgH7s4yPeYk3f
qFRSDSlFvvnzTMW5XWt80zX5zGs7rvIIca1XbcJfrkZNO93/vUNMFDospQS+7uOUhA5yfPQSLF8j
YnaNJmdGx3BV10q7jvHNL28wD0zomLR+CAXo8yLBPkoiux2Y57w1OhC81huoe2HUGXmfYSd+yp9J
mNburbt4NhzSJ9kg6zUcBcolprqExFpSNDnf4ZXKIgPbjfQ9id3u+MaHmOYfYNLMniGpobH3tht3
35DGdvheT4hsS/tydrePOIE/fyMuYm5fKIQukkpOrud2HhH+fXmV4kYkmDgER7DaqceqJv3THUYi
KQ6poT+uMhKz1TqME/LT3V0LTuf2whdRmWXYyQ6NDs323zwxaDPA+MBR1u5hyEyu8PFWjbyCwWev
Jm7X8I4oIf7aUXb9YzNcB5VX7ABptgpoqIy3rkSDLL/u/Sdw9hEKtzo5FaVcnT/xeLOBf+KhYYmC
pbeCfWtAO7OCfggGKXi++Q2eyDt5TPmJYelyolcHxiCKN0QEVM8SLvIR/O5Q8E+DSCp0e+VcY2qE
j31gvK/nMqxQ530rEjTRh6Aq3CA75e1nvEQthjXxJR0Pwf2FsY1d1xReBo+Lk76GxaCYTFNAcmKU
7HGqPMRqIoo2vcLTka+ZhcdM5/KRxowragCKzzh5R9qBmpRlMewswNy1EHjQ2r8UnVYUbIJ+Ty+i
9DFeXy837gCJFTRgZ3Zb/15Bue/xh0JrraQ6oTDZ6GIYUtXxxD21xx+faVUAxePN/euSY/57zaSA
kses58YleiPqUujcKRBCAnkK2dqEeIu1og2W3RrSH+hJoR9ubdUu4BrGJgEM9OUCaBD6sObPSs1Q
rFJFDSUGPP/a99/tAweXtwcBo//1Msm5ejkwLRmVjwxy8APUm62/Q9l3VHGefaObQYUxtvJxiJR+
80yTQfm2lwOjG0QQB7YoSKRTwRxBw/Fiape4448Y37WoEkJCKTSopyZ/BYSd1pvV29pzPSlN/u74
hX7tAG8TOm1jMUK8e1Cli4sVTguGiEkdoXzg/CmV34TJEJMdb4IERx93aNY21J1AKS8Dexrdhi1D
1uz1rdmcG+fjyPRjYvvyE2yadu+W2w9LZAToh7Xjy6A1Gf0zUaBlnj1Px27khrIwSp99bk/+ty+B
Fd7z2nXKaLbaDbryUPVIqjOWqPfIWYc9zwxr+05+OBWRR30QR337ewf8py93veMFBBhKfxKgcZE3
ey6SUU8aWz4e3GZDOOFjHxKMCcrXuV87B1veN9CXQ1JbzR7OPM4/6LYVuEMGOx27WJc6aSw4Asz6
nG5DZ3he9GWNaS9VTwJTzs1t9K5AlyKEppcBZ66Oz+Mtc//1DVxiVw6uLWD/88/4XoUH1S93fyXG
fNfdHJy1DfqEuQ4dOgX74ECSnChdYdbZI78/2ma6yWSoB87hk0bDRtMgyk5lSHd2/96wnpaUZpze
8Wzzh1bb1vf0qs9iq1v5nrX1ViSjT3p39g3slcaMt3f0fDzNfIoUaln8c9xasB9/voFiL+Tj05HU
cdc/nvbdJv6ZOoxGli3+4fZQl9zb9f/xRvND8I4ozAQPOX1ZaMzFuKbzNaeVwjtR65Aup5/I2ubQ
IjAxhfj+zQXGlEpeAzB9Gv8KNfWJzXIu5atTc02dgEuUlPNlqnW9IG7qLLMoFBBJmVJrW1TV2iXI
5zaNxiENFimufi3ALOl3JggaFuPveuJs1ETvfnuIRiFKjDzc2PCFQ9GFcCdZ2/J6W3UFbU2xCvZZ
x4nkp0Ike01HCkaHEGUQ5wdNNxriCnDF4mJkTZWgunFiVT6XY4cc0bPpOCAvUF6+IIyU5S+VJv8j
wVPGVZkIO+/TEGGubzeCIYB2WjcX0LfLDhtFfvdE5DWQuWRUpPIzk5vFfn4A3TsiGwii/NZkP+6R
jNddpydFpXwg0MMmNROCLoyn7Bm/eqCZtvSJOOL7FAPx3SKejSoBi201ArjF9C+AIOZb2eoaeZss
0Zs87PE/e2rUgGfvRF3zuh85Nrjjg2TZ7h0tgjBa/8qp28fYNo8sYZVNHUazSHt6RNkkEjsojtQ0
j7EwPXlpCkXoeltvrwAme12SenbBczElyW2+OJcsEQjk4/cScu8Z/w2n6DTlaebmSuwCyxZ0xkUz
IFAqYfiKTGndcbl6avYfvZyJRiE+GWlRzskQWdsT2Nx+0gmNfB+cQFw0BOY9OVEDb9O92ACsUZR0
rLLdnvOHECwa2CxLvVtmtAV80Zx8EWfaIUEHInICmvju1RAV6KeAYQnO3li/pI/KzEZIRysjx2ul
OTSRaaa1/fw0MILLAi+Onsiiv7eRvIARGwPS3MIyjR8SGgSqqcNIottaiLkTm5DyCIMsw4vdAb+B
5NWXMOyobCdkzGkR1dQJsIPR3IeQkw6UUjEbm7yFpx91lE0Dn3OzG+WCvrK/EZTDmtUQyyJNVtu6
Ppzi/Ohe5SusSxUmL8j6wfZNSupdXjKualMUFwkdtRSy78mDaLfRFxuliMio4nw0HtoCftMUIFMp
W4trr1cnp0IfXonL5OfsaWmDhtJgo4wJ7CVW/Pp2rEKptKfArlztiTye6LxKep9LLYZrHaUFTOVt
Nu/b+o/cScPmItAAGmTgdzc5kPDHO+5O7616OI7uP7rezf2fl5y9PQWDZRTnVOLy7pB20j/fnE2e
zGf5cmyv0hNjI1aLTKCpjSAm7jVt8PVRqqcaLWGjzu+iol4PELbdfX6HJP887Q+TSlN6/zscPq0W
kBTLwvl9zUsXrfpSbhnelFQIW7I3EjX9R5VNzYcfke3HCQ02kszgfptMF9gsRMwJggwRKWqzHOFl
veFAkXwBDChHLiJOD9T2/ehQwtUC7jRvmngXF9W2HrOz/cVLivc1TbAdOw0JhS+nUw2HXyG8JUFy
2wDLjKqZnUoXvUh8JIe5wF+Xf0GIbyGSrGthvay+2Fsn03kkpQtct87nhdS770U9TGWSlS/CbHfP
07dHrmR8mSMwmHAFcQ4egBgMHABQuvN+2N5ct+Yud81IdYg/D2530emJZtwF8eQgKBw6sBaoaVRv
pMDP6NrDNrLz3qpkp4tmXssvb9lkSJkZMCpNL8q80uHKgT6/pB1x5WcoOWi5EWPr0HEnJR3NAcMy
4RrUFgiHSbHDEfrse95MhbUlw5k1GNH8b3NupH02gtFKGR/ZYP8IWpwWbZb8hXNuaEPe6Gj6NUhS
qk5eAyhb6YDrbipTSgeUX98nYFxx8jeerd+Vt+aUxqPRHGrEGLFRUbkv1NtJfCPLSQt+a3NHQCnS
SL5jvHmDYVhvZ+RCSWAAVerw+ItFZRw/r3FzYvN7kjR+/7m/uaTgDKWTgBeRV/AVK0k9vOv7IOhU
z59RSW2HOf6c0attOOygBR/L9KlmASpCSAAVw7oMklkCzh6xHyH4X6ElQ/HsjdN+uZGHsNx6rW0e
QayvQ3fvxPiNcM+HMJkPCZ99p/q6oT3GppehC2iIbz3zZpThSDOWdBL0LpAevsymbledz8BGTqi9
NZkLQkpbtQqvFs6McrKWSJ2CYzWWTLLRl9xCCtFwgIyZJeqRJCfvWQj4g+IKoBxaG7WhjcWD2QKX
Y14obGzbLjW84j+DiI0qpiOLtrY9vT8L0be3mX+YChi0oNZ2y6Rh92jsFsy0l0OVXZCONdoD0ex+
NLW2cA+ZNFO8x1CfilstnOBwtNv3zzKpIfKfjlvyj2XmqTvEd2pHwJfkUj4wwOtHnp/JPoWQzfry
7fKvvFRf42ofXQ3K5MnzH3uB4T20eB7QrJtrRzVL153zk2bX/gDfJluh3DelebLok1hdY1xRy6dy
thNUexR1HptuMHTeBKvL2ZjjApPyVM9CSQEsTW64q+n34kmhBZOuUHcJTYhsy5TnXh54X0KDaNQN
iLi6n5ySE0xN9GZPTPpYArwso/KGFqaJoZZMzVkf/h1mbwKHtxhZT5zT2/TPshuy9fWynI1hixbG
+/4mh/WiwFdpUIsrXRDaPW9KBCPukkfDBFFouqg8tfRFs/FizHIE3WG1uJKNzJqjhXCLhDBIwGlM
xziZ0J2Q42bq1eqMsi8261K1ty9i4G05piKy3QqZvCpR2PxADy2IoJlWCuxqvK5yAGFasDipuDCE
uaLmWiiq5MWmFcBjp2F87Uf+dwKqRcdifaggf3YfR1FBkPKReD0/PbTS8Y8jOY4qnvxFeLWcUKu0
T0sidEBdJ01Yp+7lJq2kGI7sM6R2sTve8pT+DM1mxEDTIr4MQIDIY2AI5x+yMkiTRj86x+Ob/Ju+
/XXH/MoFl1byd5BmozpzZO2nyBN41+jB9MNvdwAfMnZl9vt3AJUSQYJvJFiUELT/hpZlgA0faDyj
0amgkD8zeRTKGHpy80eV/bcoXBymcv700MLfxQS9lzcgth/PITZVFEVFbNWAASZUsOGK3f806xPp
f9kVaLFJqtKh/1GBgrsa4FvFuTk59YFRps8mCAs3xgGJrJEOG2NwviJ5Ef8BXh6K3tzDv+099xzp
TyeWcGuKAzpu+kPJ3VTgKicKXqYf4pL4TyDU/K164hY/irb5FCghCYkChGfai2B35bGb/hfA3bVl
3PGfctzgoHV9A3zyFaNguejDXTjAJXLMWrXlWTCQZlmT2vyfDktvWaa2cAkzIB9oKVLcbIbZWwFf
W8cKXZ7R0KiHQEdNgH+7AoEqI8xhWlJZbPkkDRyklhdIh4G/FHoAY1Otp4Tnu3/ckp962H2WCxLH
HB0X75zrGM9eHWizBxcRTVcpUR5gfG3gljJUXn5HmL4RqLzjK90mzt4w/2LQfuaP3IqWc9Pugvja
U2lGZxI5HiJDLk4kVWxQMsVmBlIqjIO8yBAUEYAfuV3QZYfgAkzXZLeLTMvMbPjd5cCm5K769clD
iGlNbRTWWrTEExmWinOPaQLlc/WCPDWnciwxZnIH7BTT3xkKDJbR18EDFqYoCFtX7TIqCCft1k0O
dOhtj7gOYZKB4dJHHGYc9V+eLWjmWI7s9cJxD1zRrMApwrABI6KjDXewjxdgLLhquILiFBJku1Nx
rdI/GmsQ9CIriKutj/wjWsoq7NCk5Y0V02Sdn4dkdR6oYaqy1dSjKwGNQ7EbNnj8b6uYAWjAWYB6
4qDwY+O1gLvnitqM0dAeEFt+vghfloK0QDj+JXVIRM+to8W7JPKnO+Of2E0QbMLa76DmZnaJudOM
dpBK93T8RbdUttH8gzg0yiaVPWMKXI+NlV8MPIC7uUyiEBRE9xYp8dAkk/My14wAgw4uf8SDXl7P
WzILciSm7t/zTMXdHJGCTPiymuaRauW/+N8KEmZelmv/dNUi6fNYgvsybPg/b1o//suUl9yoxijY
DJ1uhQD+h6bhgjBG7j05R27Y9mIVS5sQeSzvREfmk2UDHn9KsB2RsSLxAOumvm5xyDXAPR2Gf6Mv
RWAC60NJy8KUAWKJ7SdlNocWoXAjIFNNCFdjkTZj41tZu/p6ZS3AmnilcaNoXhLX0HiA2rciOrKV
wxmelc+Tgmvq4JywMHmHINjoffGRF4U9uLNRpwp2/hWPgo+SSyYdAdWjcicPJohr+GjK0rBbkJWs
rm6Xyz9uvBuhvbwrhAJmra6YPphSOGVnMAFWBV8h7Wf1tm87nL9BLl7Z+wyVeTahkEjbpLnVbCnk
pe3trv1wdwj/nFxSprc3Ydd0AgHkJcU+HFTDqoaCPTwo9bljymQq1MOgUuU19tHqoPXE+vaygHrd
yTbTF7uUsZwHs7BStY7aCXSZqPEDBpsYRnwP1fd5Q3bj4zjpM0o5WB5otren+81qGcXdbORwzUKt
5rjPbkLABwekLF505k4z/jsMXsutXUUfG3MEppZ5q+5XR3c9Ei6cLepAeeFMDTNnJO5r7CH9Csbz
YrwCrm1Ca6fW98JERXv7sgFmg8kVhYHCfCd9SRgThAj9uipRgfElTEaBDoSATxyc79NUYiBEkRb4
JcO2rKeibUJ94sOn9WDp0kG911uYlRMkZMJHXZXKg8yGWFsP56s02z3SxBwTKsvWFwhDGQ84KCRo
rVoHeYRcA/0rwtTxtso2aF+cZlI15Dl9m/dNpg1iyEj+f0AK+CIt4RCmUMZ07n2Rsq5lQ5Gq/5nK
ofdAObwXohtj42bXN4p9DBp8srBl2e/0XxYp/+vFW+E09KkeMp31D35S2cILXzcDt0tvZEa/WMJk
w744d7pVpwRKxgzNzm7JgHFJOuhQSOdSlPwwAjilLWb984x0QXn+YrJv1xhjIWPoGKMOQSpbEaGL
memhKb2ZQ8PQYjU5FpIWGZXaigr5PO9ozBk0gRNXCNCF7z0zYYgeNAYy/ZBnesqOqGVs6vMumFpq
aUjZ8g+1raO3lKXLcMUFrkihIK29Ll8wJDH+D3k0SJdNQ/wj16e8n9GPoz0ZTust64zmkgJAtaGJ
5nCgnLD9eoG5UthiRI/sko6ex6tBWG/pev6tWgLU6BrDV3lukmS544i6ISTekpqgd/icbSQI6Qg+
gY79F2zqRmqEPqFarqTb3otusqX2Du/mKBp9wT8xK/soP1Gej71Mhi7W47jNANVOV24OyC4a8uYB
YAsMeQlJ0INle83GGzkX60K/IeqQBcPZKRlcl+g5xZ+pRzBvn9VWwXQAs313zomUtPQTdO+lCKfH
NVMPpQBpTGHzPaBWDtRDR8Kbxucm5V4Mrzk1cPHxVCHl7OKkejLLqUWH1mcai/g4nzb9AYAzzlUI
xgDdSMGp8eFnERa+XH/l48h89vsJ5IJh+GQzzQNBDl8+VJ/F4JJpk/4Cooqxs2QbWnWWeoG+3iNf
kIvEZzfCPxqV5tnKbxOKln6l1otTslvGc04EfWAgjKdgTuDoh4MtyckFBQ+3TnQbPaIlt6HWrLlU
qlNWlvzaSG6hXF5aVkobjMKxnLhFZaqD8Uei/oXN4aB3M4f+KUcaYykBjbQNqVTMpGhppWbVajHS
yGGyP1xQRDAqax4WwbA9XpEC+H5nCGrA65obUchZyo0H66Au98/D1iHfqiQZE91HqhibBbZ83R0b
FyfjXvn2aUSYaub//a/QNHdPSnSaTmuXoXhXIl53LEgMRenKhpZfNPpUiq9QepTvv3PYNCI1nBPW
BkEuoGYpv6hijrb8oKTGIeygh0CCEr3RbvjN1HZrnr/Fn9z6i5FDm+BEOhI6/ilMP8cM6hNteb3v
yKmaWyQUjnM5Or1QnrsasbhTxk6XMNhCDrryBnfGgZeOJD+uGp09wlIwUeP2Dr1s4FkiXp8fEbjq
0hNfECZi2YOjNa/bhA+fWOfcs5KgQrgI8hXtXa54EnJLSlua8GW9Js6NDQ6xLXpnK5tFiSUReEGi
/qujrBVKo9C8hdSbOmSTHYhziQ1p9SbyY2Gtr4fqpW6akrYFLJhuO0jsXO85KVxwQAPdSBdJ/NgN
jq6cGlpzL1WE37U2VcUR5gE52eb1e1aOvGxPWVu1tzNx4sqEkhnJ1cbfW1qFwrsGp0pMc8+UclyT
H/vKpS4wBayvaWYwyvocSidYb/0ToNZc4pzCKePEZ+ugdMO3Lr/BU/9BrhAQ2TbeOSa2oJZDkbQ3
KUFAbOilbSZMuQaNrnhvdzSrv4HwQXHbJwZ7FSAhGpcgEPeR/zDU4TFOKpB2FRFLwUd1mlNdJMR+
flKwJhy+rEnqBkLAkNjpOJYkPCQ0GAwr+oyWiPsBf7o8l7MarLQtNn9f2Q436U415iQNGJoW/Nor
DVRjrrD4+PLVdYfiDKfoBlYR93M+RVr0OCst2aGbkvKM6WumjnhauCLzvpVKEXVx+fyp9dQFZP+a
4YnrlSjMKMTocqP3N4SbWciE3t1SBKKEAASFfChTWG5a3vzOfMkwu7x5xzSIiKAgQ0u47dmI0/Z+
oLzHbulssy5gVmMHqZy6hxKtQYiy2Js0j3XrjmIO7AhlzJGjzkCQbhJ0X4iVKjaT1V9xvzVxJaBD
YFLXwxqM3Vug2bClcGC6inZ2zpmhQJ+HYPTrb9DSDQmRuqEE6lcd//BdP1A2/vTEg7BNJUj2oMzI
U5zYBt0d0L2jonQyZ2Xn2oXH7bHGuRAsHWfGeP1eAygGnjlAEdosGFWfit7MY4AEWLqnelZDjRdy
O9iKr++/DywVmWfp31tx7wB+fcel1CedBe+LY0JcHEBPGxQRg3ICQUmivAvPAjWzkyurbBJGgPfJ
x4okikIOPO9SJgHGOXGNxk1vUda+ckVcobGtxzDnhLcISngXpBPAzlyIap3xNnON5y7EusS/MXSl
GYvMVek/sw1996Xr0W0ODLgaSMDX7DNtjC+HTEzrLnzsqicd1PLt6ENJGU0G8LLNLBfhBcIxhkiO
Yxn5f5AcCQ5n2E2FRv5CoKxcrmSOLPw+gBUjAgoyFX/1P2IbbM0E6TppgPcYg6YwRBXK2g6gTSXS
gwcZzoE4ZWOl3QC8G2mBzZOopWaYgy978EwxnBkaf5Ypo1oUwSiG4zIkK7MRyFiZM+sI61m2AMi0
rolMF6XBHQj3XWYLWdlU5qpNcH2LvHnkkRcuCmPTrpWITzYSBVN0ObL/wB4ult0CUeU239N1eHQT
qEFMUgPKeDzcMkmbiPEVdxbhPn96I42lJXgjGqIEi+c/5nIjaZnsjKNHFqhsR7vOEO738GxiFihG
wtfCLqf5VRo72l+fCFNZGwlTqgZ7v1Lr1p7uACoI2McJY9egMWrN0QkEjhVg0oPMN2RtBS7lgLqx
ytTIy04chyk4OZUR4BLwOncJDfk9xlxZ5pj5ooF/VQdaM6aCEpZA6wcVoCkHXltY0/bcfjQU94gw
F2tk6Pnc9M0lmkAbFbVx+5zETWsAskd2qJh3OUmhckiKovL7WLqBBfq55OUxmT4S+OCyjqb6GSz7
sz33v9ApevvaBlhaxq6K2jFwECkTCvNsW9lh8G0DCRG7VqyayIGpHdb+hkChkW5NP6wRkOZBj42b
wccijDU5pYNBqTt/Drq0EM9MgAlktAOAMU0xvsnV0FcnJY5YE/xVRtSf9ic/5picH1A4DlFgOwZw
O1OrrDdTNxVvPuxS+DRbtJdu9tI7x2KBnrbW2bwSq8BfteQdUjSlqzVKkj24kYR12xw5WuR1ULAA
oJZuX6KY/crVLJFZqgayI60GJIc9CpqoT6UAft+NGSdMXNXkRXdpscZ3268x6o/Hy9Lmu01r+v9a
5jR7kyeEYCo+jc1ApgZo9WD+Hp5qfHACAgNGBZqZA7kzWW61lqyW73FzNArz5HynnJicqTmbf7bO
rYxZqbtsBE9McyqD8Er6Vf+IQgE5Ejulc/5N74tPr5govDPnYphJTRRYXhz+PNj2msdsks8EmA+z
zg3C++LVaaW24XeWTKeNwbHKlyw6yRVRwQn1rHDG2QvVYysULzz5bq1ZoTSN+pSw84Rs+7mK9+vn
Rq9r79sF0lZS96mr4bhUFySVmzOL9Mz5VYjHA8BnSVjuU7qJRhnq7Pf637faDXP1HBkK8c2GYDqP
H0FOb52Hl/xSf4O2Ve/xg491NLXCCXpsp4o8qBzbBfGZJWDGLIB8vNHX/s8wyWHrdrsWSs77bmuQ
EM6wq7zkWuCIUPrqM4+eM05RkvPyL/s0D65aPb7MUC3h5pn5e9CR+sQk4AGwS203sNcDU1kfvMVP
LPP28SmzvaXmGsUm4kKvDxNhi7b29eNG/ifJp7NOcNBwQnbMgHzXy2bau/vsuLBKhVy0nS/hxqBz
daKVOXUc9ww/932FiTadEwvixltvLurNlBpkWx8Q+oFtx7UiKINsm00q5rePjKLQLhZy1DVcZgdh
YM947DzWuMHAsO2+qzTB510VveKvPkwxEUeXwjJFeL1KG+seMkP1iCBTyEaWsFbGi2p2GBmnmYXE
2IRA096YZ6NR1Zqp7peNe3ouclkPEtkr97Xn0n8BdC6jcI9H5PlG/gGo41PFzlrciXHtHI09rlGO
qlrCl2+rt7/WT/s5TYhLwyPx3kvuvm03DsW3I+//gMuosLY8p1jIe9N4XIp4vqyiC4iH5eFWWm1q
1D74pgg2PFp1ikBnhE762cdIjCKpSg8oF4ELmO8MJvfSkfK98TL1JL96VgucD7PknbAPcyrjaRnn
mv61KqALUw5utyHjTg+YQibL3VvjB8qRtptw21yKWwrt/bhwIHraPc6SGkPEv7pXT/v7RXdEnVLa
gTA+ysdr91jaOtPmo3FYAx2cN5chbm/wqfuI2JTPP1Whm/cyXIN3dBggLvyvWRNF0EsXtNH9jEle
zRY5dULx/ViuqfypK5Xv8wCs2SdH4/MWGdcTr1T+UtigK2mMKcGSzv08tlu4/hVouWsNK2ZaDdHi
MSSNgvObRJowWOiafO+E8Qi2uXRewVEoqIViBhLT4tC4iQcOVdNy+O2VFEh61raxyX5QQw6apRYY
clXW6ces2/vZtRU993riG9qf9k/T71/bqI8cyg2Yp0pykad5GMfjyoW0Kw/YWouZf9Yeh8wp6ZWW
VjjifVnKfW+BEPTcFhb/fkJM/HLzyznqNXcjgvYjcwSqzJJwCsZMMvkIxLQ8O6fvu4vuPH0P29qe
afgmw696I2EHE5+WWIIL5Sq/fVV2th7rbEGeBrh5hzf1R7V6zXCO511/efMFSRUfDjpJcw05uVag
8LSs3AdSfCaLg3himRt1cz3YM/M7dPTI1+VsFWxUC7Ys4dhMf2Sbn5tSyRSYEpKQRKMMKUX0L4iw
UxO2u3gGy06Asoih50ESKaEhf8S/21Nmx0Wom6B9E6WpBTIXzmKItOrlGiQmatih084ERGNpB1Iz
GMkkoUJ2RJMXwkPiBEE2gUaVxB/mDIOd+mZ6zSrlh+IjVnOZRAOx3nILiCaiw1LLu0foIALOtWCo
PdD7EvEQwDxLDeA1UPi1b0pk1JuPPvoanjGV8+pv0xfStfiIKS/37cTrj/BPn1WEXwNd7VGwUj2g
eNtBWGFTRs/atzAr6b7ajWhE/ld004zs7uljHPaF2J74PNEKaF0w6ITPB/HWr0LJS9sq85wC1+p3
vsA9t7qLQHREXb3A4N/SAovjNBTeaVcexKo1+4I7nbXUWgEFH8/GfBeBmIiutXXYR3ISDiDd55pK
ykK1zBoAFS5uFfavW5Cu4H8qTlF9O1JvshaHibDd7Usvu+1J/MefXmlKVHdt+p7nqKmvZ0gVbgSZ
gEEu8Rs977543iGfAC3dNfoVzZ5w2Hpp9HKMfFXEXEJjesu+Hz30Q0t3PAs4g1T4s58XlRzck/ab
aBx/NFEdyHPSQu/1MMaiTEqqlUocURd+h2PZsT8zjM8Hlcp5bcbfPEsb1mn3HCDDW4L3BTB2L5TF
jDuPzhI1PnIXpTizOFr2uu0g+OAIY5pWgJC66cp2K8GyMM9WPMsNGf9CFenRsip1hCnYY8s9AIdT
7XLT8wzaowifbOG3DfQf0yUsIJStnGt9rYrUhtzQytQ87UyNDGq8yy/+OtaM6ZjTLF0sSpSB1W51
LLAYSKo2bOdCieA+UFURq5whLUlUbnJcADy2/uTL0kCdPVEdveXgvr4R7MLnp9tNfAnaIRs3DJm3
TBTwdMZIixLrQIdvric3M8Ph/uq1Zveb2tqwbFzjDu20xRV+0YXxGE0QQjl8hPgsbUrdhcovAV0N
KkpGNMirqQXbOleNaiaoJpAZgYiJdczC47F8TQ6ndasetcUCLM80gqvBeoUFQpm/wtp7hjntuqSX
kOR/rDHm9I/y8rS8+e1FeoKhGJhDhd3CDGOYeqcmS63HaXfYlvA2OnSslO6+LMmHLnNwJdWACUiU
Ctawma6jXceTueyhBJkKt3zxONTuikNt0cZ1NpWc6SKGwen2p2Rs0CdWFWqMwpzjcij17cQw+J3x
t1WWF62Dp0tkd0ZVSjI3VT7TrSm/2Rd3gk1MKMsOKVu66W8/nYHIvGAwtQay1gYeLKazhVxq3ZfI
JaIa5x3VQXZWqEe8pRLluQNU8KP1oxAnxkufiNzn7Na7jGQrpxSazgKcP0WvJNs7N0yW2AFfhdKR
1wj4aRxXOM99dfofSKFxWTC6R3puKWfanWfwHJ4+HTas4O9o1inemJCVUE+MfRmA1Fr2M6onOJKp
CcOp71IsoBZFNGSbzuY/g8X1YZWvdcqhTF/ylnWd6vDzYCnyabYRwAYkPxzeJtWDdHbS2xyQS1pT
NZzSVpCuH1FztyqdsUXUBXQQ03RCbaoLRkLWFbj/hxKjMAQZq2Tu53oapKwnH4+9BrN+D6sX3KpA
VEn6AtauOT/tqWdeYhuXLp/ECVdFiZL/2sjTVRDH7GnSl0F630OzaNpVAvIWxN2A+WN5bTutTvvw
ZLyGcPy//bD3z5JTeAL7+2ZdwidG0L46SgeL56zpRlyYye8ceDKYjBrdL0P/7E5mGb9Al2+49qVj
DraO8FlxobAI9UMT4BEnt0bCJwhSJLj1bKOxAwbyNxZO11KoMfBHVDWfH7RnO/kKCnRk220RAUkT
zDsxaQTC73iD9s0JRXFj/f7siir6XQ/WEwJKjYcSQejEkee66S7V66eRV3uaI7fhqEmSBdnJzJUB
I/JVesn+fNGQ5u3c66MigAhRo+vbwOrN+D4hLhGCvyUknek2wk/qWHauXNjHvkY1mLxxyf4rZhXz
dtMRLSN4+zCJC4SrSyoO8q8xGE1++IxuukMJvD7YkYpuS96VjOSNtqToLkHPvrGddVUe9HJVNYqS
kAG23AOo29rhScZOl4p9lOLyfsxoETe9x/FIu+Qy2Wb+HV2YBDZU1FSAJjNN75SWLer6TmDHRhYt
BWIVlWCe/WAimRxVZpI727mJeyaNpZXyydYnoWP75RQCGqTh+6yrbB6XCl8zXabsClq1n0K2AvTS
ZK55iLU4yHaSUc/mHOtf+DU31xEpOeSJltWzQacEUfy9NOO8wZosOteWCyyK9rWPcCax8NEeAmCF
nyExGTybdbAhBVK9PpIP6K0HlYRjtqOH4MdfoaH5QzgcONlNjAsTa6ov3fqIigNmBWPLHoKb71bG
VwsQvtEdhwbx4qNBaMV7bDTrgZXJlJfuajGUhgjGR9fy+zLNxJ1IZa3lrg3+v5j9llHPTNUO9NyN
QFSnFQUuq291mtkmmzAm7Q45FPzX/ymq7snG6PLvOJySVkXTD89ZMewBQxpWNZHaxEr6zIS0FW0M
7T9XR8kRb5a/Uk4aRBv/ehOitD+/hnBi15HxkadYXNr/hU3Lj/jf9tn5H3RCl/zC7b81c1DP3m2c
6cW+hjBjgrXfuGRG3VzusEk6D0hjJUaLFAHFcwhb84OkFWVN1nMEcsGH7mTGo5BPO7bFhW+iQAnZ
6r5sppoxHIns4auyR97MbBv51ZG/bmMrK3+IH6QPrO9OgtKGuXZJeSmLBEzLLerSU19qz/nlhNNB
YSBRWiQU3StZlcgYwOb0U/26oUCNITYYS0RdiTJwC9yBB0MFS1dVajhr5wL/mGbzmvFb+EaKwQdJ
8pTVGv6X4dIuScVSfbmNcFw7XHYjWXN05afuaT8YWNwElj+ysJCNl0iVkzgFHsJVRzdIvQrBlycG
3fdlaWJnmF/ubKOdIRWkxKhtM4xmomNZ913DhKSIK6eKKc6XECpnavo2w8SBnNPLTFuWZzJwpwJg
4ky8r0buGCzF2Hxs5jYKWGLgSptqRumB65mYp3gZhx7Ec9GQ6zBNb6rFQ9QxxUTjLj2tBmDYQVxU
rIBlg5prl8Y0UlzfMPGccaOJxoTgqoPb++CzCr52r26mBSyxVLbf1HXs6T+MHmFgVMIrCFaZVz9F
FCN1ITdTH6AIWoxDbYCUdjszAYMLW4tDRhUjiOMRB7TqBT093CXmCuCAdKKWtcl884aGEDcjqgiD
kjqL37j7aZpIAKZy7Aa88s5XEuudkxpkwg686Uu7b/+7I2TLR/x14oYv43m+h/8G3ZgiuJTHlLhm
BdLLZ0SbUytW+6c2FsnJYp8QmceFmXLM/vg0Q1NiWgEyNoN+cF1A9XTwa4caE106m2b8T3qP0nhN
yFmyNJbOR9Qt8VWetG6VN0f9/WfOpsQQcf/cWmCcsc/2aRab9taMbtl8HJ8Z94NzNSzHbA1SV7vP
VFjb/Nl7swnt6Sv6pe4Vw4OadUKUj9GGGFTPSYvPGghnRSOatJ7dhlCxywgq0hLWGGujO0TkEVqj
BIknIZIdTPnJpP5LrB2sSEoMI1kjeTGOaNYATqZkiJRNPCPJ2SNwAgu13ouHqBTlF4Zi3S7eHTlE
Q00Q9TMzoX80sLtyczA5V+wocN8x3hu+MVR7LtibwQIkPr738yOqfVkPmBiyn38QDCZ4SodliSWo
W+OipHXkFRJNbtT8nndKrThLGmvO/Y7Yv4eMxfdyffubnDiPdNoLrLQYke32A+e9Zps7OXHNloUj
bsME+Y8LrT6iZMGC7WGdepilIwVWGVxwYbn2GmnUy/NBOW2SrDAA6Zkth71kE5DFpRHVDwLbuLE7
kNCFAlk4G10Q4jkD6wSEzSi/sbnRnf1S/L0RcmI+TIhDPaCoB+vs4UTQAbhQx/JBBr4F6bTGaQHK
ncjyAZN7xwuk1Z10j8AkbCSukm75WLiS61uJjuQweMmjWqgTyipbxDyWJhtlVfzunDtO6eOUTUIW
qOy7qz+UimFwQO027H2+KBehwfhqu7L5CnJDcs6RMXBNmUz4CkEhTOOsS4lv15QbwSF2K3Z8wBzy
0oWlK/gfBtbwfbWxzd1KVJsXzHxYghoSWHsC3GE+qjFilWMNh7OjxBMlUtaZxdi9Gu+d+0+q3Lef
2zzVv7QIQKCqiX/YValZifGZCeTFqSoZvKZ1JGuNwn0+et4HQBmYKZqy2eEWiy/vF2LEAWMablc7
fqxY8fZ6sv+oOkYgMNu4m0zYxz0aEnkeCmMc29DLltKJ4KrHiWwSe91I1Q9r1PDtkGNON9Wv9ref
Nn2VALWzlbpqTwdrmxTkg78eG2tpTLu7ulKOvQIspnuO1Ws5eqgthevwTV5jc056xcOXkDO2MnIS
Mo395uIwJWJ+pVc2gilepcIQ2ssYy1dLE/KF7S0UDNyIgmBtBSfgRFsLohTcRomiukvqGreyJRWb
NuuPTDqIY0m4Eh8KxGRvA0mh/AYSNSvIpBUkfcteOEarkWN8ICoZPoQ8sLoLaT11h63c36AVLfNd
/RArpCkTVOmZRZlMxEVFBebuRNndJzq3qjEN5dGUWkpX9N6c6C++ydOm3RtUX8+FtcGdhU+TeXWK
Q1N5TkveDgdKkD/Do3ltR8GnufojpI4q1QiXplyo2QOsiG9ZdbOn2xglBFeO9N6FvzmovJ408boq
jHDig6bOA+envoRxiCMlSV4z+37D6TGHwHTp+BluYnDmBVJ1f7ctMUVxTxXEA1STxAm0bQSo9vjc
+pQM0IjjSCZhIt95cgfqZcYsA/ggQdiBMeKNbcQHKaI7kY8GZgZe3l69BNxMI8n3jvAi9rQwl6vY
CO9NNsyoMsn3g3RCV3R2mm0dkXk0tchaO40+k3L1HigjSJSRw2cRp/4WPfxHU/TL+F1fNONre8GM
Xmg0S3wFkP+z8zxli/zOBFWmp6po5BygQ6+W9Zpzfpm9k0KOYil6rwKmId7VlnhFJ13ZreAOOkDK
+e51ryzRIpH4crS96qK2lARsFyubp4knzulvXr9ueNliTWTFYWl+vTUJSNZ8KlTV5jyYnzd6iFVd
W8URr0rZvdWifNLTyJ/H63vyNAc+4NAnZlYst51a/0CZeCoXO7gPgVbFO/mEE7uOo4Jk6bn13hSV
ZXiq3Pl82OVsg6elitrKX1V7oL6y40G8CT0/zCYl1DM6ko6IRS1YEu0Wk7n6yYdjY72HvxVjRrc9
QQ9pSZfaVBN2Vh363S+KST/bL2Wte1LytEKJC2ut5dh6A50AmFvu/hyFUzcx3dOAkSmVLR5+ILMc
6MiZoZt8xht2CZzI8AAajkDZNWCOm+p4C3H8q0wLfjcbhd84RKE4QkY+btJbJlfcbSHx88WwGTHy
HvvR8SZMbLMzWiQHkxqtgmQiWxwywk5qTUaknZlx6X6ZmPte9YbdAszfny+F1ampDzdZ5ul2dU7t
7AgrV4RSG9tTlkFpKtgRUh/p0HcNzmrH4qf9tPQbZTK8ivmumFp7Ieaa8LSWpXJByLVGI7gdU0Ub
ZONEqpzt5a0SAMuoquw1nP5uDkRIclocdi++MhaMUcXX/vuouNPtck1JbTKoJ5zbzzU3y7AmQ5O8
TDYIRZwX3mZex4bcvlNnJ4kEQCQPUOqMuDZ7DuYywZmy2eHIZsmYoQR5gE2a+gPc3akh/Jb6M5Jw
Pr+5I+BpnnXXHI+WDqZmy6XxbGFbNcHe2dBr2TycdPscbjw9vqPo/SMuFWMc961VTOxKMOeB0pbV
0TwPnYmDUU7qOhhd050UEy+kgKZ+6c0hP4gvPvvHkhOtmshFWmR5+n9LgZoCeeru+rp9nvTtLz7U
5PSVShIuBfPtbG7FrhVoMaRVJ2/EDOFQmlYO3tfTLdkqcKQEFSmF98cWhnvDLZL09stnCqt/s0ZV
3KY7wH7kAcEN7rSdyNpkDSmENwFTLHJAI1m/bqAitjOEVGhb1c7T9ie9OU8wMuZlXeXCSxtTLowP
X+pXpZeqTfAWl4eM5YcjqlBCGWHVH8biNMdLwyr4DC5TY7M5usoVokzMKsHRhQ2NqXXcefxygDAf
PVPjqwbif+EdD3dWhuz4aknnmhqlZBXPODs3kp6xr2M/QfwnZpTbJ4NSH1UeuGfYaQSNtAoUhCO4
kK+mhir9M3N0WH5CXHmS4I34/8urp7R2lxJUAVVKjb01dJIgQQuRnYsWWPHbNbIjPgtkuXy1L92y
bUWmXGs6IyXafND65BOlvQLD08RY45rGjstntnGyiY3GmrtMLGmXf4UUJYF62YQ0kaxH6oXlu3fu
0zXwe9Om7u4SPiYy+k9DJnMSLCc/lwHOOabRkQIEDj7uDAeQfKgqtMw/4AkiXAzDHfDdBC6BH37t
tAcXhaAGCUWmSAeuRBAbm1x2R/L6x7wCxzzqZMxQaRpaXwslL5QWWYu6D5aUPUgzinXL6aTNup7l
OOwPbSK4Qlb+zpFU0IMqMuvsLjbH9MfvJmmVgMTTMIn7El9RLgwPceNzOnevOyYXBFFBpbIKpv6F
PkhbklznrHHOUl1QnjoqnfoiwBzC0s842E9Gmp1HJ6KoYSYk/2i+0r0pcaFYxQA0yYdnnVX/HnWh
ZLvpd7lAFQqgf8/KzgT6K3xfX7F15+JZVt86wwxjG9O06AUlPXhTk4QsnYIsPB7hsOJKrIRzZoGw
JY2dqtsdXlDWeM8XeToQkTj6epB/hoAr1HtqQTn1Im1md9pBU33q8tlUp397Rh4npQSZ/foScjiO
KQa8VWfsALl5rWFyU8DWG1whLS/CT2qhOJEo1Bjzq8gxfrp7DlpvMTsUMW6PwKtUzq1AY/JGZB10
4YV+eTiro8k4Uy2easyXAit3LSrjUQsguRmA2GemUYouibVlDHp3LOwbxx8MdSbeBv62+R4OFVTE
rePjWssSpKF6VZMxC52kwHPnBSwiKlRFj3Gk/1XXrbyI8ZJZTgWtMY/6Mst6LoDQNsYrSi56EKr+
UG7yasPoEh4lJSwU2JFwNHBMYVUDr4aSsIkOUJkupZ8u9g+OPgC++ml49rP+NEtDXoLfjmXngvDZ
nAtN7WAO1Hqt2cJ0OBySD0zrah2vYtMfcNebnj769o6SLSx0zFCWiHAOUqAcDD3aKtdtcl2pE1pL
50Xe+mrho25vqZJoluu1uqKrwdlk74Gg1G4NbMXIN1S5M8oNginkU19C5yjDUAcvggBF7YEPgfbd
rHXie3ZG0iW3Tfv3mKYk+wVkg3vSsN0sroCpQKUwHrEsDSvkUceidIlw6AYHk0PrKSsuJqB8cWdJ
yBRBz8nR1n1iAw5C1p0dfw1XuAyp23ZaxfaApoHsTpL6NlJDde00D14hk0D5UgbyyKm87frkkWEg
xwxJmTHipeZBq/PgdQkOwf7rUFJYqajGsG4NrGE8K29eFSRGnWoN8QCR62cXrJm47JbbWxIaByED
GhLgGq+A0UFj51od6DRdKje6jsI2PZ1iyxjjTFp4GO7anXH9w8bKmxp15W/DCEwBUwzF4GqxkWRk
vT1dwD5BfvzkgpPGMBjKXzB3GT5MsslqRBSv0EQYLDnbiTiXN0BghXQMfcVBudpuFNQoIEvngXFG
uWokF+hX4eHgSy/N+1NdD/N0+EXh5lx/nLmkMSyU4DR/KvOZN6+3vfXg3Yjqc2nc8/hOOljpWX+e
Z0V/3BikLTvWoxW++wpR4PGm9G9DCBygfip0snA/cqXA/9ssDgdZB0NfqBHrKGndfp04Kr10UDkA
u/HzB14KR7j/r27ngUQCnQWieHz1k78wDyIZx6oos0O18sSOnGMqEu0XhKiYhfBq6WmpTx7liYx0
fwWomks0xndIAJBVcSXr4ic7nwYBga5y3k4/4tX9iFI6r/nZ7DNS9d7bbtwS8zFXS5ADIu7PZco5
9vVXW+85mtN2+SKfZlfNL7oTwpREj8pafMbN6WUXP7KuTuBUfCTiCyFNkFKXa3Y49JjnO0g0CpAA
BJP0vvcn0sIpxPQ+UcxPLPEZgRLjx8MY9EienLi+ofsjGVUwx1HgceI3I551/zn5qmIgEewhWR/i
bRz0V3b28Ukcfgo4tJvAlE2Q3zsAIAfXhi2Kv8IzR2jxPFFRmJNPc0ZK0hSaQ7kIlQqL/ySG6DJR
ci5SPZrRY2NOe5P9dXFRBDj3kOroQ+TGQeF33H5Nadq30fXkLhFy79G8V6EIkMhhahET5PXNnSv3
e8EBvopXL/XlLCdRV+WnrQJwaaJZ+8HAH1aSf4ONtgHHqRgt18nWLqYBHr8NxtJz/qkdfXCjFGih
OtEitq8Jit/2zKumPikC09zSDdJgkHU/y1jyK2EUOQN62P0oPnmFnOBC3ZfAPptauHN7Jc2TvTMr
yCqeZbnePNea0XKrWaXcb4vRJ7H3/8gwQtvztrk/gP4m7ye7QhDbqaK6vr1va2ErxPX7IqiYW7pj
RP66sZAILgSImFwY/+zoOsyFokxGEIKgMiygaKsp28+h2eXjYbR4/NEyGgxdi4528/IPqA1+oZsb
M5/S+Isq2dcO6BJBfJqJ4+ntmtkSHKja7kQCQGMC3YlDmmV9J6FV7BvGlm38Plk3RfExRyhmrFTe
piAzo8vgxoQUz++9Bihc4+hjgsHROZxLKiEssmNBAq8XZFzksf3b3yfOcleE6l70Nx92H6b5/ccs
Co+6/BmH11NVVa8HekB9xQAk3iPv08qcfgbGIxgG8SfUFvOAtUlWzE0N4ge8c869Ic4Aaldrs4GO
Z5zDtPHreCdDcLunJd7Nr7NS95yLbtm5N5C282akoAYv3TzVoyeRmZfzRjHwpJ/iQNDSpbsw51Jx
UW/7i4o5CK8RplDZTPF4ozKW/dppOnjQ2SIQ5H/Jzu06XVFCP/gJXZUAue1EZBwgJRQwFrv/eAJt
SJNCnJ+SkZYtIxV4u5fbRpt0+/NWWXF+zqzL+3ziJJY5/Q3Vs1PX4ORinZ3lEKZCDRW7kRrmugnX
AiU/SF/scI9XgnU717EFaQgdezOSpLkYUMvjFlST/tZPWQpNqTvLF6vTYXeoSQ97gENTLhSkkuwx
F042gC2A/uxfVZ+H35U4eVR6lGEY2CNGiYFGsXfZhhI2sRTpoC0j8EyQkGWp1dHL4LzfGDWeXfao
9aIU/69xpYW8z3lk0acMKu7Y4APhLobuvSDmsjHBzxEOPMTOO2O39afuO5ILB3sXK6jVZeRBV1dH
kldGikBp1Cot3pgb2phstAtt91KzIoIUqftAs5MpxdCJFeF1MYbgrL7omqUCB6HsbB3NydDmcCxs
KcCKjuktDIerHHwguVh06wFwARCrxlpyQYM1z4WIB/ZwvNHKdFT58vYjDElvpkdc1d1dKTH9IfWp
XN7HMcw+/99VCJWEPIVBPPsKg0zCDXV2ccNDVAffZHzur9ICuGt467Z+mu07t2cpZQzQPFELXGBH
GYL6w6deRFWDJdhQMbpequChZ0sEORHzwQfU6HJ0asLlGZK6+s0T84zBqjhZiA6CnsRPq81T0jeB
Z1Neo/tGupxTIUHzas5LCzPRMgm4qFqzLS/9tANX/90h0QIZu2m95YLx2mKoOxXGMNFNb/1PZutS
g9jp0s5uAJiN9aobNGS8TcKm0DjpqXR7HZV1qvbExJq0SkMKU3hFruobf7eSEz0cfPEZl2tJ0h1L
AP1cm5ZbI2nOi+0rY+I3MlBfIDrsV5jdMCwX19U/KZoIj6kvh/TViURPa8ZQzjv4cMWgrZ6Vf5b5
2wc/B11Jq2TC1p+J0aJVENVUwjBQDieZbhsR+/UHAv186tZ9H0Lp4qSzUb/vjv3GzM4YfepEzWy0
WVHyoYYxGhUj0UHTjkSBPAAINUAJC1TyiqFRLDls917LXN2c6iFhaYEuta65UaAxz+qTXJMtkZD3
Uouim53qAj2OJeOey7o899UFPefw3unKI+DFTdSJr0vR46vmh8Rc6nkfTfEFByTSaOm6Eo0CYAT+
Aqa6VIL26wO5P7MKzxiL9NgKN0L6IAWyk64zi44x+wnLzMOErdTwhtOsHYz3/oTs0V4gYL7wUWMw
LREEFUSdpv7zQwums3cVhIpl0hyUgNdDl72glOzfUkP/vN7BrewH6SLcQu+PgFObQtCqT2zwY4SM
HiULNXzVEeVmr2L+l0mh1OfXyuLa1gPPKdfE8QE5PT+qhsj+FSzgnY8BXs1X0NDyXFhOQ3fsuWbq
d1dPCJyBr1GzcA5tsn7rC+iAzy/jDIIVerSY1WYyOCJ7JZY6WT29Ud5anWL2i5wcgflVweISs7KJ
xMjZG08Yd8tl2RXBEpNBbmIFLdz0gxrl5ps7q4M4Sixsc0KJniAam8GjMgTi4AwWTkI5Zg/sfPBA
L7LjdmYk/7FzsJJfbDvZ/qr9/xFMGBDECJZLGp2VqicCiDbVgcoMU84WFFhHV79wcR4ieETZav5X
kbcnDyk0WRFUevOh3kGYSgRYEe+a81+2woPlHDzVrsphcQJNAwr4BCh2FW98u0gKVQc3i9x3cuht
BlSoa+HwzOvzx4lmoAHMpiMhTDHOcC+xobGWg1NTQiJEAw4XW4/bgSXq2FFdLDEohTm90kGzkGaR
s8JgEZGbp6ocUKSs1Lee3CIEBewm541EOatvY5JJrJ5R//VHPFw24lx7kePFE8baV8RX/dOtOk0t
eDMgEti4f8PVniYrMz1L6VHChGQUtrup6t6+7JYhXLyObPMzFyHPVmM4wgkb8YMDkMM2PNwuAnPI
FvWBZnILaKE82kW31FkYKWYXlJtBQXsWj3Ut7MIPtAi8Loar6Z4yzR+mb8i/yQwUYIoYCNf4UFUy
1vTQ7pviqMaYKjDewcGtq15pWp30YL49jpnoZscupJeZh9xT3IWyYjO/9RYlRLJWkNQ+2FZEpokP
EYwDP92Hdkq1kvVLEo7Eu0/KFHs+3BZ5pAgVWJPQtguahS11X35fTKqRzHxCzQA9bPyzfnnjjhXQ
GEmkxXd565JjTbDO+vC8LV0CJGt3Pf6Cy+uMs7FRB0sj3RZh4e7Zi6qK2H74K2+Z6NCWL/RoH8gh
SRlWluFeGrpV44V5qT1pG0zBFF3WbIg3HVOoS2YwLjsKMCZ2VfbUeAnMKtxTsuTh5JnF6re21b/f
QOAdSY/pONnuSyLiPLMlv6X2X/IFOcvrX0DIpJ1DIEHYXCD3f/8MLvbce6artNXFmaXRNWrajLc9
63jD00YQv/uwOC3QOsgzqoAzw3paWeddy+EKxFS785hOoMKBuSCk7YMfp+LjHv83zqJQLqfQwYVd
M1o3IrXQWr9wUBPV2EJEg079RFiwmYaukBtymg/qD3mmieMPKMBX9G5myz33OWhGaAbWC6CESAyM
dCm7ea5IknxkRjbWFZY5LOHqTgbP/Z3h08TaNDAtqClLVOIXcL2CWgZRXRSP4tuBPbR7g1PH9jM1
cK0tFQUZ6GG2i4zKUJ1dyF9cXWM/h8aFabkG2IWxIiDWXmsJf0KChJHz0Te9HFoQkIfsjQT9nH2R
4caKwbbnFXPVincybyv5yK0wrEfS8K20DbXxz1wbQB2DJRlABILNz8ncAFqfcsPeUobcLL9B2tKR
b0GCFuCI7cjIDCDORgb5Ma/hE3QQkZZvYfmZUeH2ncQIVR+O7N63ero7W9d0obYZFwrzDlrZqrIV
L4DBFhaZnSICJD30jsxr7KVW8OA5/Djx+KPnpijoosi9uYPRHLcgJpdVcS47RYhqciEsnz/ANnWb
1s8WEyTomh2GKhbUiQQaYzwgsxMu3LV0/i2WFZDosaqEKNMmcNi3mQ4U5vwGGGcT04BPo6ZilndR
1OBBYH6Ve5TkyKw5cRUcWoLk/ocv01HjNCZSzNoL8upzoQi6ZV0G8hhS8ozG7L69U/N88DL4aK3X
3oUoXQXWOmDU+jTdE89d20NNHVkus6LPojNK+jT2X/JE/PKd9FhMYj/H4cvrKc62rtwOuX7mDirC
nCcvjdeWpsQn9UCaxSD6P59XiHKr+37U3S0duXwkEbAr3BaS8WxtFJwdTzcZlcMq2B6v7JdxxMID
8jFAz3iZ8xnwB13W5VzJq9R+QpdlD1CGPZBisgMicnyj7NZhdotxyD+7So8zCrgYfb1M4ZSZr3TV
BUTprRaEt+RSBMgG6YOXdwNXEfypCqq6/aAPYzEzpB4udV4wMb4bxWuw6Nf6t0OZfNSdPke25Fok
DVR6dVE76pUlveWgXbZYli4apMLPmpU2aElfAygfr5oSMmdYS+nIce0CR1oLOOAR/exaTvD+YfGV
Fg1vKPDoF75X5vEvWg3CZqX8hfAxUJ7gcHA56k6bU+HZM/ZIMVobNF3ztVq+s31RIvsjWqdhwYtk
rlZyH8gZbPRUKBPuts6v+n00UbJwF6tbg1f6IXYxDrYZd1TRvmcxuOoHWXgks8duHOh5k48BnYjx
pLRu7hMAkifLUlTf5zFQ6TN3wIptT1ZfDXsW68V1RHbXzHEnvW0Z/l6qXy/17zKAHrHNN9j2nliJ
+apYHeEsB2Bq8mMz+8+KzOSC2VvvKz6Ro1EyYAqcGNsu+6P8Pwm3tN0m7uXt6KVcMO4Vpal8mITW
oV9Gl65sZfwO4kqX6fK3wk+Pm7CqUK/ARaSP2iSLW12+A2nHE26oVh3T6CXTj4P9jtR+G4vIV2bl
LHG/n/cDC2hgYV+IDQa1ZT3uvJdX2PoBTm3sBh1FvzFY49GNakGdFx5pD+hFnPzVoqtSF+pfsDjl
QBcxMHhd+A/cOlmC7INU2aghV5piTe9/Bck8/x8EyOMGysxpCX+81b0JX44rpYT57K+T5xz5jyyl
o6MDIBww45YwzVHgw/0qyI7ha2PTludd9cX36lg70Nf1a/lQi1h3HStAQTthxkA+L0UO9p3o76wl
bVyLOUCe4JcoVaaZUdBgKEW+KvKrLfM3kxYLB3ec9w9RhvIrsPJ8XpQOg8Fr2DoQ1WSEOXlFfdzz
0dB/56FHfHZ3qGWLgRn1BAkuahTv/VemcllxbR6oxP0A0GNVw+zCh5C4zayfC79NfbXv52sQC36s
dbC4g+q/ONZ0p4u9Lev7kBCGslYpF4KCc8nMf6AodOzUn6d6KFR7WyCVQ6REqycgjNodLVb+/Wo9
D6xAeJ+Ewx3W5j5xSoCdREaLZvZkAO1/l8CtT7j4YB6t1Bd9FA5m1jJkPjqnOueIGEgPQs6dfiAR
Mt/zhckJxJEhaPPt/jb/iOVbOagPQOk2VrPQn0bQSCVRMmZiUUQraCIBcJLaK5mprS+NZ/XME2Hd
7X7AOeRR8UDevtL2dM1vCDWqTlXRrfIn8cRa49oQ8j6FTU9ngTM7maE6OhWTc1eMwS/AyKt8MlPY
Swqqu/0UGSroX2astokPBpDth5nw1rpbxqBCyBTBvUNDE9S0hi2LYCWXbHksSOH8nqAHkHTHrvEU
mqIzbF/j621HseEnEQsqrEadJdsxz5n/LW5N5r/hMmNC/1CnLDdSmTaHWvLQ5KGfQSC1mslMCM8k
GEbY0aqj5PIvOMAujoPHOpmkMKBUne4kpP0+mRrkIjDAKZjC7Fz/19fckoEyCUD/SG86/EgnBPEi
75pDsRl2C22VYZCpYFoN9a8Ic7988cmSxCPs35dKCTOK/LbmfDU9M6ssNJtzIM2f9bOjY7RBU934
QX8sHlhCO052uJTl9k0ZNzd7KAm/E/VaTkkppMthy6Z6vmjEJh1DauU4BOef3PeiGQTsJF+HBGB1
FrSHkwh8dY/rYGk0bPqTx0UKbd6NgUIX9ARKKCeszvvmnCiWWawma0UdaHLeaWrIbpuZjO/nsyob
SHn78DIxZLgHJaz+7xi3pzZGwoADMjlOtD1/ocPF2KT2fQ+HlGdGYIl2E9D73JKgKJrwDawPxXvC
7pHGjQhZ4vZMQA57Q0wSUwC4ukG2Fjzq0P2vm1NeIKWxTaJEk6qNvFZNf3wfwkIAfAH5+84Y0ivD
Ui61yi0f6R0tag9ekxqk+t+7exoGbPSi4x56TZWsl5gIdyoVXcAaJW6JuzJLcA1+N2CDsuw/Cqxc
Qhc2pGz/Px06rkjsdtAjuDqHPE1EPjrDAeWIFcsd2C4xEKdX3PccDeoY6bQsfurWGNVMVcX5uD/P
zs6BMo1SXmJ2TpxlN9Z46dTNR7VBpyj7MqLg2HI8rQW43/VYqKczXi3RXcNA4vEAIdsvEtNDr67R
dlgIP/HRcltnH6sZj0S/bzni8wcGFnOpm7qLgxDY2MDgOG3OOqFs4ruD93jVYojUVptwuK+nhGEs
OuF1E7c5cyuefljv0Md5lAeZ1f6/B9ISTofpcVpmThTuYvFnV7AsG67wJjhLbXoGp8+MZmqJhWGG
QWkcggRBs334dCwwST4kAiYviCxbUNyW0B9wNipTmoKYzyiEQERiTvO1WzVZr0hMKeacLsxBi74O
EoATLexo31trzfyBFTJ74fId56u3AJzhJyzFqQuxtz8MyR5shtfwRLlFHi+4ExbwKgRf/sed4Yep
cLNVADkpulmp3XhlBAjmVl4PdJmrPfO6dEOjFWmlmh04ajBZKbcRpzA92anz7GiUJupQZs3vjx3j
FK2ebrMMYFvXyp3WpZc2yGKtls23IZeXTwI7dPGOVMEtNOE24xFOPbSYF8ccbiFctd6twuqEWofG
Qzl5mzLa3wtQAMliVqOzqycQCQTc056nDMpFK9JG/0RVovIQNttm25buNOPqF7XDVR52cPInAKJb
j4SDaypX4HFqCpbbSkfKSIJpEb7OfnCfZp9GLrI3UsIzLEUDgbecFuyZS/nuuniidBwQGkhw8/wY
Z1X8g2iTAZ9+H3aHms+YDY/DhvaR8tQgTO+8pQijsWb0nKaqRMnthpQLiS3Ut/oRV/vwCtuQgJCO
6RofCFbApTEGwIDS/qOFuZrInR+zCwuwnX91IqZOOS5ocOaJa/aeGthUg7dRumKB/FJesK1Eui4X
dTJTPBV38ckWldTfDonnR+3k0HN7/mEcXnxePoaY30p0CTnykAR2PcjerKNOrOGS9svLzPsGU+iK
8414KKPeFPBkOjLmEKcgDTXZzBHez6kSKuV8vFDMBwms0ceFS+ALJULRWJPr80IgPUo8S2p7WFjq
d+GlXk/klIRQRXQ5wCJP5KqfvnOHPl8wyMfB87Aaiy5z2+eydhME7kaI6bu0TgqTXlJQSeCEUemm
IcONUaU0f9W2FQi87662YgpiPmx50AfTD9GjqdGV/TC1StwVDM4jcO9Y4la3Gq88h8LXQjVog8Nv
VB8sJRHHZiYWf2RUGJojb0qtg0Ssp+ylp4aWVVzXjuNb+8ZApIZJLz7T/PC/6/LDO3H4rf4MxkxK
nWrIlo5uM+eYVMCjb4y+ykXguUqF59C4g7JOOWKcaVhe9JaBqVCf4FeBq5YRprTUi8GWf/XA/xXa
6EG5f7iIZnnomfOyjVCGymqXKW7m4A5H8z9tNTzQf61R5O28Zt1GTWpm/q7FwjTDJZRnZx6ABmaN
fyx9Mvt1bURk+IKIQiTe7mQPw6SNXi9jJREF0iGozUt868dGq6yWelw/79eLPvcy378ViBAt5G1l
6/hsdcYWDsx4G9UYdDiJjrWoA7kH2DP0L41IK86VVKOtVxQ01hQsNIuawlig2ffdULMhLiGD0fdz
M70Bn5LB/wpH8eId/+1r+zootEQRY0+15uUTv6Nby3ChddJQamkcjIbO9WjN2aQXmqFsq122dT+F
hDQCjVWrbpY/TdaMVVqaN7sU+pVUWrYKlyOyU6qL4qpn8lCqy48UKkKMJxjw5MqJXFV8yoJ29jnn
36/ms/YQiw9Q1LTOIgzdcjZ+G0fEAqdUiIWqcqmujAnBduZWYphKZK1xoUXHN6Hzs4eoLChtSHql
UpVTSGNEa6nqE8wYU+oY0pPLv/yOZvVeIfg7qXiT01p/B0ONlN26XKLBtgQV2nWFJFITOtciBf3Z
HaJ+glFQvCp+h3uycHau7GG+h8mgifM7Q9v/GejPRrM5TQSIO8EG+UvH/DhzpCY6JwZyex8+N7z9
FBbRyERg+cCQ/yMQ3XvZTqIACsckThf/eJXfg/b7Doq74uC9LPJvgNPQKRH9C74Y/JK+d95UBepX
K3+hW0U3fhznLotOfDVHDcgn4j81B3e5BNpxs1RurxJFsdnAXRzD+ghQc99vZntlA1jScph64duf
jkj9QpWHchhF7qO8X+CT5E3vfQjZffX6OV5lxDYgjUFtqPpl+rIy5NlNWT6ryIRBbtLwuM6sfIeL
a2tt1P9e4J9+KU18qDyDB12kdcVS8LkWQW8F2RxjmRQDxPnCKkl+UpR3nqguwR7hhk5BO+KJeeHi
jLOJUQuv1TLZ1xiz7nPiEBs7OoOu07M9bY0KQClqvC9N8sLFZLFZok7LzHMfRKZB+ea87fit12PC
n5wFMGHQNtuG1L+4iiXSnjJm/6urybqru1ShVGgJY4cIzZfY1nond+A6cdc85KETZTjd+s6S/IJZ
JlWxRDYoiHtJpv2SAopObL2p9CnEJHjET27/hqlfOvGaE5eQD7ZXYZ8oYxGGi0yJeABR/jJOdDL4
6eSpKdvbUGziKAsdwGPk0woE6MDjUU5M2Q0SiGCYdvQ0D4y0OAzp2Z9YSAQ82tqJoGhLeGivF/wk
piGMMbTelOIcjyhKaO1t6ybAe79X/EUlPobvugDd3+6bW8QTcE79wYHBGe+Md3ZDastZQysD4sAz
5i3eq0uGod9pVGOmWJOwCXKdfyEPDPRThYRt2QCjK9mz2CpQEjjTTQDqd53aH2dXOs/EhdQ2HZBb
8pskY2/ePtTO6psF0SX4GzIJ9M878OpsUftngiAn+MyRRYmkphXMg4ldMCaIoMT7gEsFkzlEOXj0
EQrP8XxmTaDN0aCKrJI9FJWO1YFeBunxU7VX1QrYab07Fv6TuyqANe9B7hYX/UHGHkadl0QfpeqF
89jwk5cq/nArpDgr5ovDqJZjjyS9zbK3+67mDh27vgHgKsuRC0TE/Kj9ADS32Q6XXt9aY+65X7Gx
wgpxYioYRL/4ZoNmpf0PppRTl/OLeu+wCS6821s5NYbhkv81W/vX8nxHEoAGLdeCq3tsEfT/hfch
s3lvHKuwEjTIt30Dx/kSU9uiWqW9tH47Az2+dh+Mtux8VsT2OwXcvAM11uilEqjkpw5ZWsqbIN+w
A9lvpcyVrL4bj4u0/kZxX3YKOc//jPgGgGjAvwUHLyuDK97n3gXjfpfgACxIBU5Ep6tNVcz0wlRI
EvU0aarKuiTOnkoARAnErqTkMiDo4UKd8L9yURug9r9TTuSyXBngWAp3A4o98XqnKkoJPCU0T6dh
SzG+ijpZP4FalXQ9ecPu16e1vj35A51EYc6RQ9J5qt3AKqDkNoLqsXEBE6ryCjOJzb2u1XROFPiD
cbZhqBV5Tea2GAtXouPROMPV1/IbenVxez0zF49U3PTqNp1P+McVONhWL3U/Cv1l+m8UzIX+FVHy
XxzqWL5pPNYVwg10Xi/RdAVZgu3kOwt/ZH6FTfPEuTFeCrhrXd1qIRvlEOCpAYeCe1IJbJinVRMR
oZuNQCZGHZcf4dx6mCIA03wl8npTvWiSBr7vyVRO/iuAHfDgoNC9y7dq1iykRsYzfs+gGhf1wzqM
88JcfuFlQ3coumooHESIJ6pRgXaAndZjUwff1H3IhIRANtSENQe41r6YLcMf7zeIDNyYcR1yXh5U
Uk22LoZ+ixA58LASB+1MH6FwcwKY2q9BnJOFUEzlluU9KifmzIewvAVGoTOdr2hNMh7k0Bbwk0kA
bRy/KdM2WFtJYBz2Gxx6ZBl/Z54dT5z2IDDzSBt+KB9Z/QbfrUfTz4Df/u/nXx8No0DthswM5hra
6mAF0E+jL01apmpDs9DLPEEKG/zIAihnjPklm9IuCmU2Cq4Qb0HcvI0JHJetU/iEg0soNF5CR2H4
TST92/9qZ2jBpaIyRTlte5dYSkh2cbbtTKGU4VFp5KKtqDhMFOmTfaUr9+eL/CUsLJMm31NL1YDA
Ua/6LJQf9w85aZD9VT1emncZ6E6OIwrNcbQD9c2GiZ2rTDVeAjSI8fNy/Hi8hdRtAR9t6vjg2EZc
KkIrKqFhL2GzycIYnlvm119x9CjvHqVi/X0yG9+E8lkent/bwGKla2jNbNcL/Bm5QrjoyYQ5mLE0
BPnYGqWvmun4QblHQrLS5b9miDTF1Uy3Y+WK6BHQWBrFnuIxKAlbodO+PKM64dvrH+xwdJbWWsWE
ybdzAKMpPGgEC2Rrzfdi1hVPZeRE9B+uG8qfjsRQGsea28OqLoeWF15EGnJkUFaA1C45qo9hkrW7
FFAqNi83PzkUnnR9Ej76v5NJtCfw9seyvc8tB66TH9wwBUu1OC9vVgytKkLdjyTbENw1RawhMjug
IHCk9KWBuR67m+zDo1kiDgYS03E1JC8uzkLEP4g2GRu0roVedX3ga8KVVZJaAqA16OeJUpCIjaA1
IGJdAbnY6Hfek3mxZ2JLyYHXNst9IKkzn8Est8RHZr5t1E2uP5smLOzCnWYFEK/GHXhHkfX8WPKU
9fYcsBB5zdxjGbaYdYbHpxxZCzenZFk6TcuXIy+Dqyp+DzFcQtChPZPmh8AlyS061goa8ndN4lSV
6fmiElwSKBx6eTenwJk0Gop9VKkHUy01oMgOF4anxyqqz2nQQ6bVyN9RtK2m554qLM2dDDqqmRfk
XHV3BrsydzKVLqV5mQiQdSGH0IDB572cCNLCFZDdbpPYThQVFLQ1+J+x5VL4qrMBchr9nMxxyN1B
uSRQYDoVTT6XW9B5jD1M54SMs2akLSiDUMMIZdJXi1XQUfDrm1iYB6E4vzmPzpg9L3qgVKIc8YBh
ub+cXWnRfidXcIgBt5lgNbj/8xXFIGs3XZNyll5jzcbaU/v9S6pyacqP/qzZY/mV3TovhxXODTlI
LfBS+l/ibLE2OsigYkpH65Z++cPD0XcWbXvRIamzq1t3WIL5MynajbR4DB0O02xVmcKpF2F8zGL1
+PfPl4qe8KVKbapBat22DFQEb6QXV4muHMKFLuI+Dr9lPo9InsT8Ydufpv0/W8uSKh5VhE/zue29
AicGYvp2q2Y7l+Y6EsuyAJhCrWR4oz4bfhXjqVIjvT2rWLsQZFpvsBzBPczFDSYzi5rQMugouMIN
tEYlruCMZaSIVziKE/6yhxQvCxtzw2acGwcbJfvn+kFM8de307VMynCIJNFDOksOET3Ng645wGeE
I4+PCyfdLIygaW4pvvObz/cL0xZ4ly6Fn1sbyvrEV6s+K3Yx63ERk+cpwG38sNLohz1m0iZumTmC
0HbauTZ7ET3Szkt+u6muGu8DOviqWr2it1ds0Q0N8Ra7a9VfnT7FeRqqEZskd5+7gIySNW5GrJ94
mHGdL/xWjojBXijsOaPeuRzqGRmng61eu+IdlBh1cXvyIFUXx90wP65336j5/N91u/M2wDFKL6mo
4uCF9rcczyrYXpjVnKyfC8lcKy6HgLE9U83p8WLjcnlIHMa2J4riEsMltsx6auHHY9O4TAeCMOSq
WugN6kqBAR4Zn78AGGw2SdC1/77sAxvI+q+6Ec4EfCMUU6hT/iBmNReZ6Zpd6ddoUURloqaDT5W1
BDA5FhLAzIJAaA599fNwW+4BEwll78WGtWBm4/sbRq4koHI3pjnqF5u8vdcIy7ZPHL+w5MmNXElt
5PTECVJBU7aGwlAqEwapWGNQB0ne8CsbcwIjA9MOkdUusph2p/Kry1HuoKXTZoKo0MT1kOL8UZX5
Yyv0t67VCrV8NtWm4tN85BzA4QjjPNCWRbok+/o+R/552RfkX6mttJbUNgKHZ5PfpuOP+Lu9wn2j
nvE1sJniV2yjdkxJCJgoUEFkqEaRPgTSR+RIok3msMZHrJb7HlEqXCtA8oPuUwtQhwHsNX/P5ZW6
5/4FI7PmpT5dVRZBuG48vX3yzKblZfOKIBoFWR+oJ9GaLw929wVefqzQfIkrZ4gX+GcqojQtEGzq
AaL5+/kHTKGrtx2ykmBBW6CeOprXtSRW07sXxOyVjwNlxsKLuEtjO6dzJF9YF0nY0o4sMSVV7odC
suiELJhxCYhf3Wx0YMQzHAGTg8Gwrp7Rzx2/e623EUnSZU878qf6wsDDUAm+C6PaILyOH7QMiXaU
JR31QJUCRASxx5hZ91OcN+QartSQx7skSMMgV2TNULMvzqliEmd5eF7CBuBT/6EOIXTkAy4INnwc
C/VJeB4gba9sIosl/rrmgdbTk3U5FBXGj9Y5jLDGR8ZzVxLpw57P4TfwYcRMU/vYiRLK17e8bqxR
I/xNjVPYFnpcIi97Jpme/VgoIWK/H/ZgnqcOqPYxd3qNbFYnKN+qt/Gn8MqMjU/JK6gDBrt9K0Ky
Hm8piSL4+/bsiNxDl3Zph83pkmCTLHPtW/I+/Xkjm2yptlSUYUDgD/t8H6EIiVYVpD1gqip1VWjg
OKjukJHNvzjX1h5a2GNs7TiUPulPS3o6yW59KUVK086itTRFPodO68MLMZvo4s0UpH+EyoKa2FoZ
eKWLSrHAwbuk4HJBh3LLaiBYyuiSTF15384mREg6HviF5ePxOdnNMtqtA3nAHq2lrKpgBQWge2H7
r3rGZ73bEnAXaZVXlpXPOHM9btUUt6ypdyrHZGesWLleh4/2O/SYNT2VVz6jqEtfUqZ+8SEuahKK
U6ML4D3fZ8qJRo658ehuKnIyE//pX8UJ4h0QWlUtvxQDjJU4YjeZVs/K55p7PNNrppFaMNdm/ORQ
CzBgvt4D9NAjeRyFApFXNNlfAVIsgGAPgKXkX3aQy5qsQfna6ehLwn4NdiNv24V2cHk3X8rdEXM7
ZlULufBqKF42gNHszRSsandFCik7coObD+iCBNCzTyt6lPW0ZcQS+NgwrbEKHi3qf9KMg5yh8PXJ
a48wZ4z8xeNHaGAYZtwxxeu0art11b4QWjfm91HhMhpOcZEDYGvOmkbk1Kh5Tob56bxtT7CExQow
RJkzAy6sARDNyp2RXjX5xHeBQYRYhlG1aO3JlKuL7/vkps9YY3ZNvMdJUEn6ym41WQV0rerVk/40
EyuFYIFI49ttgZbmhhkB0ZWbVpuSSzmEIwEEaCM1tETe9l+513elg3p3QvgHWEnFDKBC+qWFiFzJ
k07V1qL1ZhsuTWyal5wfX8+Fo2taYMlIAMRY0LNXEmIup95S+er+cGRoMVgpdJuoOl4s3C9AA8XX
/MA3Ak+BSAAw2xHm0BRP9YJyGcqaQdZzuH+oVZJveQ/STusqgAxoS5dAr68SQsJa1TWqOFRs4Ei2
ndVLHltIaO81o1YiTs1DhoKSaHS1Fpe9fdYSJhwWaAGt+6n4v7Fixd6KzzgufvlrQ8bi3Avy8vzL
HrXkaeCP27J8AZNLo9RFfdc9yV7ai9zSVdgOrL9BfTcXBEG5DK5iVPRjHrOmJgp4DNpLEIiVpBts
aoCvNyo87aNfi6RK0uarAvvWqh6Tx5f9JqNfUT2bqkEiY4iWvdgkpLBEEWKyoAy9uNLXAsQMuBL6
TnzlmctvlzG5/+9yhKTm2Olew1B8GbLCGSBU8fhv8E7QLiQoeor4KmkasACO9APqp9esnq3yPURB
s2kpnms47g3fxpLhWCQOjQRpK9j+NnGaLkokrJRSiZbSDWswf9Vu5zeQr0mnw8vpbpUg+q3NGo8w
YSc6aWLBRkWdWV8xGjQQIl7qXsBf/zjX2mJLf+kir7XF5AH3x3aUOTVDQpJg2JWdh+JNDiCCczSJ
9o/YGiwuh4b5+Ck/O2uYG/sb4zt88y3Ru/u/YSgezwRel8iicaK5TecdQUONLZ07XrF1hBhvPYQ5
ltS2VfnPrp7Z//vqdeDhyIsgaYrOJzJkjE10Q9xx+BcTCpqc8nbznlq2cCK/ORlwFts/U0U/EBGl
k50O465iLzg1s5ixuEVdb14aY2NYv7BR5fkv8HiSQSd/VRsGnJYniRoDH7vX77gci0BziDc41uZa
XZ6+4VvgM4RXOVtSICEuNbwlM02NiA/nY85xuz2xzzKafMpzb3sld9y4vJWsaigD37zJZmi7+7Wj
POTNMPpXHU0I7z68RAKjmdidBwwt4bi8CpcM0/bTAAitbLqhW5GdX0/bU4KwBrujMkpZaCcVPM7c
7kyCplg3dmg5AkbiiWKxuh//anLqPw7eaABBerlKDrv/vxAjAodBFUGKFkKF6l0UWnBziQ1rfebm
C8WiIjp8ArevgKIBQWAToTBwJFeLqKWtKq4g1WT6YUnaxBxNXTo9eyiem2WegqivSCsiL9aPfYAM
k5UZ0C4ZpVVFAMXKE3ezdev9X6oGvIDVNPs2cX4jwizk2MqEGQWXWP88h5NejuHAiVUWW9i8pr+f
6v6SmIDeVelhJ9C71YTVa5JX0fXQCDOfRTr9ljXwxmuGgaJOp2y1D4Xe/d6m5UcFWQ/1EFUVnO6W
cASLJf5UEiW3izFcGfWEG7XA6RwPUUAEcBqTrUQeTozf3hNG8wKYG/uHdXr1tnd6C6n5aGDy5xbM
hz7Lw668v8dr/TImhjmfiNGnULK6f+nufBnrA7B9lqqcLywUooUWC1QQhLLuUIrs+rZvCB57eKI6
5imMdsXxLrrxulsx1l93JnLsbA2AacB/Sb5jw8GMtGKn/pkhoGmHV1CJTUoX1ahW5iNbqM4ausfI
X3HimrlaXzUYZAavwHZSXWggpMUMYRx0Nf55/J9aCK7XylG5E+sQotuUA2Xj0Htzss/OVvkmbkHM
wWz8LZ4wjBvLiK+4TwNga2YPRGVKzzqlrS8fCrHitlPTdAK35aLMOwLY0DoR8nLzkcvQjmbqOQQN
ieH/D64JlTJhkX25hLk/xmamKnd/qp5tWMFfMCwk5fKrgOGzN79XX15mqkJ55l/Gu/EcCeeNzUh4
fhQQs1d0uHMq5BtcB2lWRbBKZAW+gMcFByuMdc1AfPvyPMqAei6FV/0Va8UW86QAS4XbiwfbFPh0
ZwDnWhT23F0gxen7cH4+VksxmIonc4Xp3k6Drp6b/ByWlMWPA7yFZXwk6dqBKCbYZZUowP6iOHEB
MY/Hy8Ez5VrPj0K0hEjZ5QaeFDc0/YTlIZUeXgGE8ISsQNB/WbZxfEP1NOH7chm4L8WF/jnqsbUr
ksML34aL7BEvl0h8dJJBvYKQ8Jco4e16ur5nriifWQKe//V0f09ElR5LnzpQZ3dc9qA/PZXnbZDU
8lqt8n+aIcu7bYPxAigd+KUrPNMKraZSQfNl0otIsdxIxroXt4MsluPboTplxVl2pwEujPugZdYV
guM+yhqucrNbOGetD9qhbJeaDbFZUtRMtzTRrHlOEl8+uTvwYKFTHBERnAMpNJzADbn6AoLmT8mn
Cc3QoIB1VeSkWjLArtAbxmth9C4Rnw4/MSANBtrLvfgqjaSYgvKB7krj78sqsLmWR/DnAlQn0MvH
WG2IIR2h/Bue5DiMIiuxXjjesh7LelZiP/VM92+cskDIG7O2CmgfPX2udlvt0Qs5WlCm6Qj+fjms
ybGvYgF3S9KoyhSv8kg2T0Te4Jin4NkDmq5SJjWkurna95XKGVrpiquDMoRU+Ee75doOIO9gjULH
TwflNi+uAg/zaSzbg+4P5WM41+XQE70dvVGxI1vn52PnhbNOVML4t8FgRALU1ec3O/xpeuDxqU+q
zicLa1PzbQrAtAm/JinSwqvtfatq2jyIX0iOZViVEHMg9oORDLYKRUdXON62HtpFgY+2cyQEwUd5
9m77D96semAI0B7zhbJa4GSacLFuaxSpgWJaj7v+rhFf/eKCfciBpx/9pAgHY0t7dUkmwtT3TsQs
A/MI8CQS5gdRz2DosJFvK0ZDFLeK50gGbXKlAKQWZRSy7JQNuvsHcIRjwYvAGY0nHS6PKMp3mJl5
fk1H9pAHXDYUPZLoJL8SyuTwr1FK3+up27tnHdO9XQBV+zyh2negRupD16alyRZjvp/gaGa+wh/M
GJ5mXoku6kDPrIsRaBcDnfkVfgtwCw5wkz2zTIScvjeV7VjQz07yOEyC2Dlnn0/TLaHnJNhZe589
merpXkQtCdHxgYbpfvRV0vJ9XtJbWz9bfR3ftI9aA6A4L3g3+t2xjcKTI4N9auLU1hfXKu6WIBpZ
9QIkPhQSE3klNJ5FeJZRw1R+2JDWUMfdSgtfBeL0tojJAROBaDblh2BoKb6aWp2ZxDez8h5Opdjz
E6umqLgw1fKoN8Q3HaxQXZCBX/yT09DrKYejJn6DIDGSzQQ08kX92yXPkBXFSKQUTAsht3UZtSyy
ulFApEqFrKENjAR6sdb/AP1B5eD5yQ59769WMnn8pSBrtG0/8hTo1fYkUSG35eBcFuFjALGqQUak
9AsCOv0wcjMyPmEmrgXDrjVPMUXbOXPYYCt2AfhL7dM76WwNIDVwlT/Ql7MN1udCKmfPtRKYM75U
/PnlWRYyDaGn95VRVgBZWrYSwSd4a3iCsQ8WE7t91afv9xl21VuspWZu6yq3m+/M3sVggR2w6YYY
o1oUIEoyDLk8080iHiB7x9k0pUEC57jgcB8Coz/ZEFwok3JzF5O08D/BVd4Ej3VNmRuNMPmS0STB
VA4HOv8jkkHbYXzvNJYx7ywOTsgUpNOOGJ/XlaonguU3f7/aRaju66SqL+k5gqJ4+1em2boN4vs+
YbvUkplDfhxEggUDptg2t0jyBzaCnh+V5n4ofaoo8b4j6Fc5IOgO7UqUBP7nLqG7Vj8dh5XCvP0O
Z99R/Y5BTePNAtkdBkI1If7Fcu1RRbepMPkri+d9cTn3aCOXvJIq0DSmFlE4L4XdcLBDBU2S+fJ0
L89hnYOTZ4NNvmq1DshP4IGjphFaT4pDTgI4L5cs6+nt6T4gfJgdufxpDGaUr2tD4MqLK2Skman5
BOsLWO0bcBIU9UUds7vNq5py7UctYOvE6kZd64uJjJZ+YQiz8K0GWEtCCoVFo1nBx1uQoNlv5L0p
PUwlLxkYpiU4VKs2TEfuSGVaZK55n5Baz4FFFXlu8z7HWCLiu1tDv0emTtsbQgC7KlMbDXAzQPap
H0XUZVWt1RjKzm6B/fu9vExpQIR0ErvFyANtprHuBO/B8dSDTIDYHord+C2VZm5ylqtzBgensq5O
87FuHyaADG3uYDCp2YiK5PcmbrdYx/+AXIuU1b3Fr1CNG+38gJ7bHoy5fuko8oeC7/m5EDT8R6sa
YW/GDzV140vB/eM9naqKrhWL1FEZ41gCrwCKgiPYR4SkdptXoH/3esherW2HlcjERvq4ICsD0uzb
7sITGta8ISmuQLMDCRGOD3VjW8Ti+bHvFlRKrfG8bCVnUjJunWXUEwihU4qsh4GwfM3b1ewdZUmb
mBIAPrmRx/GmgBc2A4l8Wa+gmtL+zGT80qErkXO1waYPXLBFkgkn6+BUKIeXwFaRou3SoQSAWed4
oWAcnJQsDhMBhffG2B1kPreHVCLOKOgco6jYaOLrvRZO+YRjCdkT9yBwiVqV0CYWa9syLKpjqBaC
wmxjZdaTf0s7kIbrJnp8+L30n4Kgjz26viR1V/A3TeSg1ynNuuIDrtbfyLfGKAXNLQdJAvO+v9uz
A/qclF0USvXbv2VnWg2w9RTEHW1TMwnw9W77dV/5TysK3qQNlBOONKVA+mKWRzTubCq/xrGaQsOg
jF47YwLYQNdtJebIZO78BXelxB5fdagRdSep1lsCgACHo8GSbvrlp5FvLUzIxfmh4izS3uOPg2Gm
FQdPgh1oUMHYJ4M6Gz0uR3lryRM2jAV0WjWvvibwCv97UPinngM8IFZL9N+likvjEC0EQbIo0Qtv
uPGangFA6TgFLW3ByM0M06zyjzSKepiEu603Tkz1w1HMizpZKJoeZL+95J5JY7EgJocdQYx7E9Ss
40oDcfUa9IfYuUQL8ZZKxa1dXjrWrLnsz9ExLDEc2ujRdSsWe2p4HqOBJ3C6bpign0Tv/oKoPAXd
b9oT4TJ/Ns2d/RB1tUadm3WWg7FSw25SFJxnxdLVSuKAvXlh3wWk7DX1/swqObWOB0IqhaUrPsmM
CHz/pPYurcX4ZePBuU9Bo1zPA4tM0oSpHM6nKpGnzJRsQ1aMZjrl2WGfM/XDT29ieTRZETac+w2N
i6Hixnv+uDog7CUUBYl/xwf1Au70Tdi4bQpP9B/sLRZLhE3uH0sYHqlgV6cXwVWyPOWbKjlNAiDT
HCCuNwjxepYU8+NggF7WBVol0g+SqDu2NkZK0spKGrLfitcpCUy6Xa4vegkWcabYqh3fL9rX9uxy
+mfrwsELtZeLhn+ou9kYAKsds43AuvgQYDyTWHQexgUngf/zfhMHlXv1OWVhq7WlQqBnOgkFUViH
P9R7htjnvnEEii9VDrQSFrNTsmmOp60sk73Wm5rmenMoER4n9xeBS2wK/nMJGBYg4BP63MbwwsAT
6cm6ks5vIefyWpu0y95QZJOnUzctqjoP8ddY6bnlinsuqHNaVzHFry/IiA4w+kf5jWvfwZmh9feO
4rvI8SmNRqG+1lqRa/rhBkWkOUz4YDEW/SYFwp+aZHc6/ikNxCLMxcOmmuVyaLT8Iq5nARibM4YR
uB3yTKNJlUeq3q2vJsF7eBEQJ/Y6zHqgdEJJUtA4oR2lfy7HBsVpcQO5ab0SXLDl2oovo1hxkMnd
j/XT0jw9t//LPv1lk1T1KHoDcoKsvhvGa3SOpVFUHlwI/ADx2Dt7iE0bt9L64u0tE0W3+pawXOM8
b6JBdAhxqY00VHb1g8U+6rCLy6FQ05M71amqgyhwX6gQZl8EspmDqtlcegj7PRWXmRSD5aDSmqTb
89b/rAHi0T/ISVKYAsas7TkrH0Poi/GUxx61It5t/TMc/ArXCo70pR5f8LoM4JFgqNpyYwcugZuW
M2O9j29RrQ/ru5npEG6OsAoU3/LcVqxBt7azDwDymu9T3RcPM4HxuUlonYUxJTaTQOGHzKI63vjM
Mv6xM/s2Aj6nMAzM+29ko4sJLZ3KeCwHE/2JzDxZCsSynRmNEkC4jEoIWzVkmmjjAVmjdVWyBLnx
HWjtFxSeCWkcG6fK/wNmncywCEfqsyYivbncWearj9smqcGTt3tcmV0H/g/DLViTEFFyHhVKWAfk
9PtHBhpRD8ai4O3p2xsoqEisyDd2F/N43RTC28DUMk9WtMuWgw5COKFzJFU7EgpqfDiF4Zwn99uS
8tGc8Y7hXE1WLlj3EPEam2uPAQDbPloC1XCc8fjtuUbC8O87zk2eK5bt+FRmemBTXqNbKnw40OL9
dLuWWeXVtJ03h7K08m6JGzMRxIqCanKPaL9IUT6mpCxS5GrIl+LmpiWVOZsp0+VJNzpjh+dvfMI1
5HYnTvcJ73hJfnQHHgVyvsqTNA7LnlHrtjcQyVXkdOaWE6txgQtX57uBoUaklpEhB+rEVPBBaBSx
p/d+aUMl6Ce1BK3P6zZd14i6Ki0UEv2+q0TjUzg09tzdE7jJUNsWm0uxYKerTpC5GnYrB71FdyxL
M1pa3XFaa4Img9yO/iD/gWkBswWI/eRmMiZYsnU13rD011je5KdSlpnmYyQEm7kYhzg0JchrheCe
yFu03v2dVc/SXR11EHA5e5pTImGNlMC1QX8zQCt2NSYZwqHQMcAu6EAhpXv97jcQ2liH3pzzuuG/
F8jDF28Ca1ZiHvVlIBfzv6ayCXm5N+ZrAP8gmt9j9GOlc1mx41eb4+078tfWmwoin0EjYlMI+fbQ
1/+T3Znwc+2TdCZ4Iq8gBRdQIJYbKTEVvi1DzksrHY0SouAkU9dy9eUApNpyiP4MKNo0l4Lk2gAx
K/qpeRcUEhq31zq/G7WBkQeHswUo2tsVZcM3tfMK8ZC03WPuTbTfRr2WCDA4A8um8wJUCvuImmBl
Y9DUdiejhnb19u+gFGKN1oVOD5RvsLrpLjGeMC6TB1c2bcqftNjPka6MGf0J1OWF09nZcyKPwyNr
06jsypKwQz9cQ+8Ljhiy6nqGC/oktFjc2ZEeFBkfCqsC4LksGpT0bevOVzyBdSiMQa3Oj0MEWTLX
BFUYecBPBGNABHNY3NDjZpqsA3VPTYo3tpg8dFau4HYBuAd+gZIsL9+TPuS8d824wCZd/39/z2N/
6BoxgZShyyxEmifqrmZsu+t8GULG34194XVyJmpLEAb2ztMJ83oToW2jQinKANrRFcz0PiZMcMKd
xaV+W9MJzVJrr/ytdTMH1RhYDJNGXqwbO3UyUtmR7UQmnevWiHxkJNb9RhVvRlO7FkpavRLleuBP
3xyFSVBTIqZ1zFYgBnswObDSP+cjrdsFDwJyjLp6NjwPGymMjiVTkugyD+UsEHCyRqe+kFNAcIk9
b2Wb11w8Av6T/2n+6PxVb/Pe1IICCaNGDDDE3qplpNoeyzJTI/pCSxV6N5DbPWGkPe+E1/gFIs6q
Zcry6Avvi4bG3l4kbubEUj+/wbm5bXmIfc7TdtSnY0Y+pUztxeXKh3KnEXSNI1xpWJ2dgOF/Y1UE
4GOOqmHPOtsGZV0fv+Hwx4Yv7OCPtSKMuev7lViHi9QC27IvLaHjeuzX7WTcYpT7OCVPM04wcfMi
fGWXAuJZ+m5T/+ucCPF60tqlIKlb9/ktUiD7z/1ZxMFVrjXTdXESvzreXhkp7AM2BNggxT4qQ9Cb
u05N+UwWXDOSB+pE7GHIVd+gSH7Xc9BVMddoO+ezY/IaaNOR5mneRqFZlrQhQE/r8uoMw60ybdkf
MlWlUbNdptvPrZ+MLCnmbhtic50cSBs18ZhvQLr1DI2WpAcYFFZy/SFG4Zo3r62+MHqpibZrGElp
NpPF/PIKKGLQAVEVRZU2JTjhRHxDZGU3bfmZjiwecKDQHSMt3kvZCW9yT5DPtr5xPYhJKV3t8fDw
1hWN5s5bT4uCHJrf5+b8qWJjfzxYOg0PdjJB4dB/NzBCqLJg4D5uZ6sr/WOm+vn08PnUYYSYE/jK
At2gIa7jGN4JMRvXveEe/X1Llx4L+HcWNZcENGS/qUm/7FgIa0SA0TYL8P9JCG21j4zLaBKKTbmw
VaBtNemz6KkO02REe/5ZAhf3I6MSGkuA3gC5TgTQybDaIUv7sHJy/+WXZaH7dJojZ5ffxVzxM5Dz
AvRAB7qtVDLjvDUYrIjBvGE+QnwjNewuIPkQzfyaNiIFT7U/mWzksI+ECt74TLnSkbt+uBjD3JOu
QWr9GT1SkKuz/4Ofyt5m7vQkUGyykMcmj37VOinNLBBrIfO9N0GHIWQMegiTyCxNvbR54oM7AGqF
9EpFUIWJKIG8a4l7SfStQwoTWj1VMropY9EGWRtibPNlaRVE3TxOdrOTni3Os1EBbWl1pGOgdSrK
XP0xJY+vCoxqPwxct/7dI43/nKNyAK9RD0ZexbvkFcdFcA0fk5L9I5pptEToJ7vQLh8Vd5swj4g/
Ghmv7m3SYF5Hpqv7WBU2tplbCAvJ4iAelbonHbkXeUIX8hIBRE9cjmMKTCPSu0jTL6CikvnV1rrV
1k5Jl9q2nd15RGdA+uNgdPeeY/dhioaQFk39E6khOLW2657gtz8Q9WACGm83KWFpPrH2ldQaTidI
qc+d+pj8GYEf/E0E/wMCod2Lj7RPyqBsbwldCrDZYvsswx/qdnLhxGkN7UgZqPbbFntSckEz9D6p
n2ONX0ksAYEwxb/BlnJ9R4EvXHZxVKL5QfX0TKMCzofT6j/tcP0Aud/IC0PXXfqgEDIdzgD0zn7k
OTm6+dmrjHIZUYbWfNI18AjxwsAa5c0LhnoCeXGg/xrc8mBzQXPIfgtFXZCPFmMUUBn9UlW3Uxm4
lK7BlbGUI/xunD79fqeY6iEQ8MwIcVDuiAgu8rR5cD21ro8HRNbNRIHVAi44MHG0vbpg92uF8Lid
C/LmcelKxoOkvSj9w+a4xgm6lklRqGeacjHmx6gA+KjvOdXKTK5HHwnVxJCP2JRB0WV04oFrNK3G
aICa6eScbB9ANywOGn9QrW4VGK392UVMnEJXkBzVzr2rQaVDeuXpb1KJFVGBhl/T9oqM5TTeTtK8
5j0ytPK02XqxDcjnToUrr8uKxGp6cmCdrCU75jJ/zG3DCIxEWE7FGaGbNOujjXHSwNBPKtY7te4N
XDUyOIZ40L3CanXGkshpIR9quE5IANxgmCN1UBFMJb6ndgWKjt/mSrGihB/MvRGhVw+m0XaFrbUP
A2YSHCuErsHTr4GTccQlkCvEE7AEUJqXoumvcY0YBfqQHGKkjl7+q3E1jXH1Px9LQUB6WkRN8HAt
lel6509OPvdN1mN/xBjzwSH0jwTNM54WWjg3MYbKCiGakkOSC7KmQfe+kP7NW0rLefxDz7OcbUGo
+JSPWsYR5ZUyrgOkrkPM4ethTSG0SAkXSBS+m/oB4ccZ7nbz5AZiZ56402GcmoIa4O/cZJzuwiiD
S9MvFcAj5TPhsJT0ZIOyCphb0Pzni5iZO+2sSKvqq4GS5K/gLROxob8V0aRKLtFNe6wuZrbsbReL
NAXazOOid0fRZ8hTl6s4Koh9u41y8GeLOT7forhje0uAqqHqGYyicvIb1c6HeGa4TdEwLfmrsFpA
fuivqY3q0aDnUCZr/uzb9kL4EW0FS8+zMTd9nZIqyxkBckpCvglRZsRda7Y+E3iBIiIZmYl4Rv0c
h93emHvHz+WHJ2LBaergMGyq8IT376B+YkRK2+OMGGYowHVZ+Hp2X/UrdiJfL1L1BTRYt5j87U5B
xZQNYjgJ543wikR2JCm2BhO+vur1f4RCWwGnqjuoBf7m1uRsn8fpokMhPuap1JPXGoL+MSC/exFf
hRIbb386z567lt/OQDbCbobCUfbSb98VVqm8BEsFtuhQXCvIDKSatSFeLV2OEwo3BBAwuBIBVs7K
uZIfzxdCZO8FN9u3TrR2xGUJiF2kUsL49XMAeKk7trfIerR3azlok2Nycic3LyiY5KYFYXBV+ZW7
WDSN+PvXvPbGCpFUbYYCzgvBlwKodloCuc+PjRhzPuHcSuGQz/3Ilu9QWWRPLfHwNyrQyC4luwvi
4E5E3l0XxxWjQDNIxHIoFn6S/I6V7Y3hpjOFm9qO5P0gK2jisJpxbCI5Cv3IHe8gJs37qtL8M/gZ
OMZN5rNHt4c5rAG9yqzd0TvfuuCmuKJfc4oR+giN5lgnsA/6NM5z6cbzeivpz9lTcDc4Ljz5dP3A
d9oGYe4U0Fhdl39BX65Z1VmcreU3fHZByveqVgRnREDueV4/B8qaAlPdbXiVz4ju4aPTnRjD1aMa
30qmcvxZNgI8BmtC11t4AH/C3um2Efpp//w8Zg4OtFQAcOfnYyLDsoMeNClBIM05t+5Unx8oJCpW
c65TYUsBaxekBWAxUbCe6Evfaj23SESlcUV9d+lQl4/oryUUz59Mp+OofluwwkbckFIXB7q2OIXa
Bzfba4nmcjBMd73L1JSj0wAUocIqSSVIsFCm8Ne41l2c5WqgHylFZPTB7/l6Sn7M0QLTodW/BC8b
9WbCp093W2jIJDwKGCNZsXiUJA5tUlrSvSgO291YjjfXe46kf2gIAjimqS/H5KLrgVtuKZQlW4v9
8jd/4sxDHc/cuSKRokjTcKWwfjmyEEXonYiNnp4Rsf7RImB6riTiuz0vD18aMi3nrHCfSUVrFCJ/
lgKnEjm+Wdp5viklcwNhJ001jGfTRF6qgcZPrc4qBXbUoxQbUGHEoIim/1nKQab7diZCZEkRoRLa
hcmzyNG7P44MKY7sJGJoX8ZSynihDALQX0dlEe1lnT8R8aBILWPW4bKMZpHxoZtw8uYG8PLD4+l5
ce/B7tTqXfKh5TbxxPNx1bRuycLAdIwGlDjU0GCNHt5T/hXhmFGc7+16HP0hjg2Mf4/9MptiiDJp
fwbvRu886ZOHG+NgjfFOUBG0WJf4FtaBzMk7/COdznzcB1AyWDdP4MWVk0hy8oc4OqSKbCFG79r0
qKvvUHDAP5AUEvQdqlm8kcQoVHmcoLqPR+sUow2qv1HQ23UWY+3O+JmkbBy5YxbkPLNx1m2Sc/Dm
Xzm/hcbNUWGLazHIFQSnSkpGkHw0g0ODzlhuXfTexxmGy18eDPtMEc5J4qXImXkNBJmNMNjkeGed
aZXC2aVnPVCsANRslWG0GX/SAo+Xxu1wo1d4Vn1xHLwR5arnuFu7TwauQPzmb/Vxvb7UjDKigXo9
Ma/owPI2he40nICYr9AItTaCCkK7LHb2eF7UkF30SQQWxVV8ZlK8yfsYtQOxJe9hiOcrRREFYSDw
/kt2RQ5z/LHMPmzB1T19Zdlj0SVKUPfufLHhbA+MKv4xo86XgtD69O7Pu+6lNJ4iqn6tj4UoSFjU
H1/XZwbVZCKUoQJGLsFZBSEFq79gRWuR48AF2xSpX6REdPnzeReLYAsJWAfAgY18yvSBfr19TeCS
DOZ3ZNgDvef2a68HNtTJR3LaKdSiH16sN6nhB3Fc94RPr9jLTEpCR+2xsGQIJnnwDrS+zbS+B8ML
VR7yyqXaOEzmIvYssQle7ncfXt32CoPUIbdaxjhJRJMJ3bkyiHplg/4z4e2HkNDuQQr1zXe8WT5C
w67D4bVYaX4I8R7FPllTG0LsENuFKkg2F00PlJbOTa+iRH2QoNaJjmh8EDqF5SxOwsi6ONpQXaJC
l1LLot8u101OMXPRZhsbApF5cuV9dNbYxlM29aSxrlLZE5E1eCxHkkXKh8hN+U8cWN1GcPrgyTYK
Mhx21tgsST35aqjiwnfrrb7CDR1PDYXZmy7RDTs1ouKxxUX/3SOGKlNvWzJJ3l+ewhpQJQpjGatk
6eTP2qFyNU3bPxxLAHofB1V5HScIs6GwtkGdVu9SDPfHl7VjMXkPg291HSmxpi/+SbaPLeDUcgFY
2x/OPHrKDWevg1ucn8DpxdCH2WGd+rj4xez7+4CbNrqBBAfUmlzCPR1aK2Q4lENfkWxNTcaHV+kU
NPEm+CBSh+um5ZiW2L85uELAQ6Ujfb2yzQZ2FdXYULxZrpZPv3XN0C2z2bi4JPrCeCTDamr6JOkx
TuJkfciT2XpBIMZZc6VkfOzXAp7r/3bdOxPIN/3Iq0GEJCBqjyuPAGC8gFnJqhOjdCIS10lubsxc
nuV7aZPRJBojsd9gVManFIUdjCrXr02/HrrQjFpO4Yx4BEBZSL5Ac0t0oU8wZ58HoLMdyDd42nZ4
iWvH3oF+5BefXhn8BDk6NThZRVKPiUewadZ85eknwwQ8SIWBzKsQS/H4oR6f8KVWKRkjpxCRAOZb
qDlqK1147XZDsG5gwOZQUJ55mZKFfoRv2nkYf+5+FA5EDfszWyzRzvPOHUN6IN6r2BOpA/DUcHD+
Hr8iQNH530nQnYo8P0wx+aLUNBDR0unHZVnsqBtK8jHSWuqWnYKQGYjibf9bC7bBJYVJJddgOQch
D/bmHup//mCsF3iwhPUIr6q0b9Y93ODmogvzVMq2HAWy7T+0yX1vfxIO3abAv7Wij3ulKFXzMNsU
0pV17uzyxLKAl8OE7gWK/hQ0lFDdxpR5ppKtIzjkLa0QJvGqaJ6oCvnjh+KAbMyA5LjDc8gZi8I4
RY0krcTBq3DmsZfiEqlvkiLom+Hrcq7GFSGVWEDh3bWh1F9eatUqNzf9QxQPY6zwMWj33hF9xacm
sEpFzEY6frwdst7wk6/zqdSLlSlljWkevdzH8WEXLWGEm0X9qQ7I03AXEpwz+AcLy2Qd2IsZJFy2
pxFBGrYS5R3t6Ds9rtkZjC+SkL5ijW88ifcvvm2NM9FFPFB0+Gcvf/qL4SzyPUd0/EYonlgcZOCW
DFW8fI5OXhMkDjnjroewJcfebw10zhN3kNcxVYPzixYdI/y7oiHAZWCgCglIUGN5UPPKfMWcIvOd
lk5l2EC0ttDhhmlVbDKDiXDuYw4Mpum16nPqfhzH17/6X4nf+4S52Dk/cYEMzfXxYzQvuhvVmJqY
tLsW8iawcQj/wyZ9zOyaNKlAYKQPPkFqPZOPb/3h+lHF3+CeQvuqeCN5N0ZJkOAyvY335IBtC23z
5JpIvrGTUwUsHcWjbUy0DlyPYfWP6uw++h7KEbFp2O1M/n/+bCKSU8+r8JAY6KjWlm6C7Cq3MKfM
UwE/b/BvNt0qCM1IwMC3jSFjXoaY1Tv3EEBk4eL24oGHMDntO9DQ30/H3/8Oe+Ems/PXCjMSL6kR
oKBgWauns5HiM9x4/kmsMqZpbW074JL9dErkgsw4OCNeztC32XgJhReI8tVNueZtwvQMEuoJkfNk
ZOFjbuIbnd5aKrsV0rScOfX6bvBlA58JZFdhi0K9UOMecrOW1mmLqgwtmIGQ9GkHz+BFszyR3Vzq
nINbVoX+p+HigspgAlAomse9zyafR0wJrzijVw9HrL1hAQvQ9WZHKUazb+BKN2afrmKE1fEopwpZ
EBZw/ffZKLQbjHEzC1upOturBCsiBJQ2Czawa72IyIkYC11OMKidKBH7Ub1DoX10b1HrJtE6LHA3
+ATGGt4wgx2QNau0OtSymMkBMhQ9ZhxyB0cvc4CAHwgpWda73jTdMiAfE+XXSc8zwAc6G86ZpHwi
C4cnECZYP/nAwzi1ClDvhKV0oMxzXb/oJyOJk5fQip/dda938B5jLgDQcWKI7aR8EPgzKnmo2RUp
xohVg9keV0v83lOOKT8vTME2vHCQZJNvxnl+2hu973cKrsJM3j+DalgpAmgXXDT274Q4GOZHhH32
CpEZn795d0ggRBeyTXRqQ/IUPSFkNBk2wyewhJR0hYmTkTYYU44MgfJrJyClpGEvdeOutohl7NWR
f+cpgZpht9VZ4xD6HXFBeMjKSMlZR3bl3K4iDVyNtYUtHtG1ojNTaHJQ5e9LnhmB1US9yksmElXv
rlSlk2A9/gOXonVgmqyTCLXkkUbQ170IdYWKYDzpcGS35MbpkUrdRTlnQnpDmUdJY20kF9xsDs/P
3aHlYYp37BPbJp1rn866CXapwgKJZe4Lo8ko0r29Wjke+ZyS2WSlU1h87rDc+hS2wyeMinYIZZJ0
OZ8k+TEM9BOWy9qu7ydW561ePuPbGUGuTlGsJB8nVD25OD4nsBBb//oK7nI/IXJEDMHCjCFVjsnK
YWpQlderkiWIYtOqjwmp4LDUSit8ZWevK/7bBnu2+2g05DBvZqFjzhqoCrl/gYUGDXwjuE/cvgTZ
rR3zhUY33Hzz/NNKM+IPri2lMvn3lS7Gk3u0sNMFiPGlsvkjvJDBwNhODNzd/goO+Wzv1oNmZ/AO
THV6YsLTtXbJJZxH+To0ZsXhKUIyMEE5dF+E04xABBchLPylR+ZQAjw2AnDGBQrQDSYfap7INUOK
1b957p/NxBNHDf1N00vG/B2bK9TOQB8/VD5b6cTpMpQ8YBtmIf2KATNyeTCOXQsc310Y6kKv8agC
YRH8e8UdRST/yE5SHwu/BRI6NrO21A2CxRDWhVuF0dwxP4GMErrUoCBCUghzeeNzDsyhn4FzXjMN
NqCO4TEje8Xpz0CQb1lEF4apl7khDte+EzWySn/zC/k/FVrnon3pHbsaHpT/mbEeg7ld1Fhi2Xa8
UxSb6TD/VsQT0uVTyiY0p3DMuAIr7FW+O59wzGW2K+TTBHHPBgbtDiIA+OSa/647UWoAGtiOSfQM
arGIRyIQ1264AGBdTMGtCL40Cx0k75Y+xpvsW3iOYKhp3ZJd050sTPoMQmeRpksm6Sar66ene2i3
qCmzX0bkgev6yzuXREoBc5G2GuO4O9c0yK5VJ5D3EKHiOOwlf0ZSrUNEjUDKNdCHYxXv7F3rMhQV
NEhRUx+D6Zabsd1I0pdwM4uygOamXEy8NLKHA0xAn93cXOXQ2jzxfLJEgmfhSpQhjL0VBPl/lTkl
ZCt+LffosBMCqxYtrGQvNGPZ8+EAYxGzFWhuIRBWfI8DlbcQ/ddIVKrj6HGP52JyyYQMQVx8qJGR
QOwy3h6HMrRHpRFIVpOgdE0vZbbYBkOCiR0mkQvSKsy9/rMSk6W4UWci98viELUr5mk5qmxq7LEY
glWDUU1HzwRblC4oY4+HdTr5xt1qW6G+i8EsmCTbxG2IL/jORSLhAPTwPSVNjdHAdys1RjgA9++E
YHl7fJvNgdeC5hjWM3y4hPIgHC49nnmtmQK+Cmp6WUo1DV3iLY0glucOROgsz9xJ8vtJ3Onj1Qi4
FhLoA+FMbcAAvQUbfABbfwTcJpladKz7m0wbzdYV7jgJyOBgpxv/+Rg1DjFd2vfcT/B/iwpSE52u
5bPeUPIG1FvSxGf0Q6EazU4mUNINR/4bghBn4ckpgS/0Xm9fZzFpQu8u39m+AUSaHFSV0sqFLF9J
UByPtCXkSUsPUzGZhNpH7AtemltEKRA8m6oyJrMQTdjIQ3etmiPJtGLZ1C97cOqAVukLi5p0j7hg
ANiilHuVze2ioSTzjbdCP6g465vyz4Xcs94eqmBC29aS1Nkq+VJlREagWyKR0S18i3Imm4wj3Ev6
jDLKSHaWZ01JYVgK5xQleQE5nEtCP2QHZgoyhjMzBrgDa/c244OjVT+r9tB0xw4Qx+85NaJbs17j
9uKkttH0ZE3EK0iMXnyr2if+Q/ipysBKRQ9KVYr07F22PNrAFxm1HwSavKZMmN04qdbe+OIuDsGH
mVDRvzqRGvFwiEHKLNTKm/0UO6GEPHi3WNLckNZYlpxPdHkHJhtwUoBeNN/Jc0l/pM9RmPAKfwIa
sEEmZWOGA6/s9+lpoHtuLIlkseIDX3vjS1cCUY0ypPGaGE9VKCAp4vy/v8xUzbb2qYrBHN7VYAOE
oAQXMOAX8ACB3fs23K+PJwZH3B6rzOzHzS3wATx+1hSL5futuOjx7d8GD3X/FpsZklpMyi+3hmaW
5YpGNCPCj87udig/ctwNHuKj7t02zKP62YUDUWmWCwaMGXD+Gf3jPKHNTmP5sx7zhI+QvQK38G0S
pGJrA+NnYGu2T2jMxzpkutyvSCtFSeUj+R/TwpRk1ZUtr9fHyFdRWCY7R5Md98oWMBlkV7hAVzwJ
jdXHDjHYl5u10xbXJTXjOHIxVG5xi8fpioiLlYPvYNUNm7v4h79XBzzR5ivAOBImk67w8Ze/JImm
kmmvjHDJnF5jQKY2ztGtS9VQvMl3EIDtuBraT+lmlznZoiDlLfGWpuT3LIWVs5MdPmIP1hITZXai
GTwR9GEfYxlfkNeZqcFCzIaYrm/9hADc4GCPuH5YMw9p4G653yCpRUSJkiSrwbjWNXEXwG+bk3n/
pMiWNxngfvDD2+lD6h8LNAKeIrTNZFXMxNchKmvcrOY413zbwjca6Wlbioh2sAnN1NAwKhSykp1L
Y9rZFE/Ghy+1H8MTnRfLjz8L3UyhDQ2mdnseTov8BZDLLvGH/c5BLoj8yLbXGK7AtNFIdQv6i8XO
MzzUMC98ohlvf/G7LZm7WL92iDv0a466EPqRaesfHdtLA4f7mLwwirBaWYLfl7OhDWOYdc9G7D7w
OrnnQjGMZCPEp7KiK4ua3Iz2d1rt+G/oYVbADf4I1Sghb/W/qe9DXE7kBF2MTQTxo4zxJEi5/g0+
QA26ktISvgZsNWnx0vxQnj/89KBS6jsAh8kMtpIWEzaHm4Sl/lmMJk6B0j7A/euOUXlRFdXatDf4
ojM276MCrgV5LpvwMGe0LutpBsUjBHn0jr7Q/JxTbJdFb2FjVxIlLvaiU5P8flGlEGn3GohW8icb
vLWaKKlus2sWJWzlM5q4Jo9/4AHS56JgDIai4MbP62gt8/sppeKuJCJ8JxbphmvJoshb5CaFhfnV
efIUkjnu2KDxRGhgJ56ZhC5DgegzrFtMorfBcsXWfNXSYkhZdYmcya3jJw1SHMval10wrOob8w4V
o0gie6KVoul7z+Jd7FHjgCghsNCOE9TAZgxox2YsvMiVASd0U96mtESNH1pZJUKdYW/Gav7k7L5X
cQG9QHqwdi7KpvD1aNbjVpgeRB0eeNjl2kXc6WnHqM44F+Lw0S3rfCowcIj9SqMiOCO5BQKp11LZ
WXwVt9yWGpfgfpK4omd1kdTRbk/E90EIcfiToT7S19rrIHOGvzB/F5emGKzYm897+Un6VYp3hdhv
DzbqUDnLd+BBOykL1imSrp7xoRDpa1mqmIXu5YmFSlO6lGULTh4Btw/9GW8jcgDhvKt1ZkwY/Log
STSE1uZ+iblmMN0YlHQAn+v5zSY8sADrWJwrCK4dc182prm88vzxf+M4FQroejnf/7Q9b6MjVWZe
OMWCsbYIKZZnp5gA7Qcn/yatkbBymAOsHEX9pwqiHBazvMGaZWHlIOIwyc1zKUy8QOIWvolanUNJ
OHhZrqimJeRvOwClCIBH3qVgKreRMsMFpg2jTgqfNWry1Suw5QSvvdYXg7VvRKktmThayb8bJA9e
9AvBZ9MUA7F4RO95FrKv4THlCgKch26p37Qc8T/brWSerVN4RvHB12fHdtkRPxZk3Do3ySIlScXG
a892PXp2CXSDsLdopk5c7eR81SQosd6tUbqQ+bY6/AuKOPrLThpZUC8b7ORT7kXq7K6poDaUCfDg
+SQq+qy2D2iJ1tPVs0upLc+RdQGM4kw/xeIKqXZno2spvN5ZdVSsN5Jb2GVGFgvDH2bA3BdM6xm5
XoG3FyFWe4yhaM+n9m+1yfljVpDh8VNyQ6p8OVTbULQ/yhBeBPJclP5NUjnu0NY/9EoFCIQgwiFt
Zd/NbjkeGVpzPT0O8TwOp+zrss0DiPz6UpnlrxqQCwEz/6fOEaIJMpGQr4F2Prv3W6XuXhoB5Tnl
EozYbsehaOjl4dDPMq0WuU8isVOOMAQzbqS5UR3lIcj4UeQAJtx8gjhvHplwEjypzum385VqM3cW
7HLG5oq5qlLZG44gcVGDXCBmr7NeY2tzvn7LpV9bU+tBq1Y5l53/h7GjHy2l4A1nexY95yHqu3ON
u47O+jnFr7ZA4LaE56SFMp5nas4PXV/52uvAyXsZR7IRpvUiDWZur3Y4mfNhaBmTQHv3zAZi2q5h
r0e+77mjCJfC8so6nG5Xcdd9p2fr6RvGunC69gS1cy3C1dMQiMiitPt9R4XEtnUiY9GSbWO1NsGE
KKrWtJoSQ7zz/f1nmMNd7lLNzSzp0SzpeC7BXR8WdRoneLKPgX2dOFb40jUTJnlsya2R27FwXp7v
ASlwPgyQJJY72+KiGaUCay1Tyu4Hszf8FK/0TGFWUhnRkpivRfbJbP/cGSc0aJBKtOzEikp+rZHz
MHpkZ8EXetlBsvblUJXkG/XYjIZTj/QkJSBbfh6RaAQdtTtfZu+2ljctkwzu/IjqnCwlOlxEyE5r
0wTegr/mldTMSqOVzLhnXHOXhrfLhbXc2RZj1lIZquVN03xi0TvfDqvw2TnV0mtI2Y8ASCbbtDsr
KijPBSmwtilrJnA3PjWNiYjFtP5sQOYWRqjFlhLYlo4jINdouY9iLd2nseDz8ULjC/wTrpWXkGPJ
4THtmvyM5GyEMcZ00AbqL+p5NQEIzCH+NvQKnbfG2S8+NTz8meW9tx8dJB/GMTDaGsJauwz0zoFg
wVoR7i3YOYbPkRQ31aiAVEQhqyhQaWBjD6XxddWFCBRmQbqZoQoL25Y7uWqy73flwEBwJpnFyChI
ZHQSffSG4vyxYGoEa6w5bibAALPh4q1DOKTBC7timchQF08rKvtHS9ne3WYua4IeInkPk9eG992W
cc8XBGbQYbX2Dd0VQ7JRJLvk29rL2W1+zgN7GyD+MJw5MKN9pSmkO8efvjye+ugrmocHGRR2JjZS
0rX4MdSRoOBlgZrR+5qNzcDyj9cX81CNBcg80KhOimkVqetacK8Ufx7QKU1cXUsqx24JGe17Uj8J
GkCzuLOdMsLvyyQ+M9C2im1YaiikO/tNHCnGqX32xIBxsjKktUnGpqQmHWz1sLDK3aM3Tqt2gocJ
A+mjPteKtcMd2oJDyICx23JQs73fcSZuBlk3x49yKSVSWAgQbUjvF6pKEHpo8IcBbDPndUnwJjng
Zkh420pnz/Y2gsM+avyhONJtiOIVcpJCjh0ohqG91+4d4s/g0VPlzT/irO8yQCrfFTYV/9JaGRQM
JdI8o2U0R0hAIqlAEIc2YMszLcM0m6VNNbFQ0veLDEvAv276bE3mVCL6CQDFCGS6TBT1k3vbQHe9
Lse5zpnRpCYqxvKrmOJlWo7CxOYHdhR8JvEhche0pSIqOJYj41s01ADYkFUlw01ju4eEYtLXCqKJ
UB+9bTPanSUBBbJDKx+pACcE6zis4nQJKvH0mbJPrXucPfdw7WeToXdmdZfbWvp5CtsTaS2JIMno
ELsOPa884N+g9J/5okPbj8pKXYqRWpMHPpIjUdZpRNT3tSAxpAiNjhzd7qquEcCi/FZNqnHjzuVS
iQPUUgOUzU7JTYc8JF0Y0YFpNp/3ejelX6iyk6dtAKTe3eE4ADl6TK45AyCJQoifkeJdxRqLI1V/
XyJ/V4whp6UbI8AshxFUuoTf+F/Do97Hsrh7UvoBbP7X4M5NWsq56Ch3AtDkm9SOjLHIJkQh66SH
hhIOt9C5wKGccusMnUFjE5tkenvW6IWX9wIPh+URIS7ipAjRgBkN/En4bQODVQbGXogqWooFXESJ
bfU3VOa2R+8TVgOmkAyMI/611BWOeHQBoscpDwKPzlZgTSDHZ1VWj+Ta3pIkmPHfSnieD5C2SpYA
SE3p/Z+m7g2qUuPc8VUz13rNdE7zqEPwSIH2CLvJU6B1oldQ12O67w5fCgMr4BbLJwGcaPX+B/Ma
BOL+M9BzWG2J0eP+z2SFMmRICBOIfAiULtSOCmjNGJ7dwcT4CsX/0SWDcl5DQyVsVcLkCQlnLqFt
VQIg5Y0LP08azWEJ1qMkAi0/9dlEgYIVJUotOixMi6zLeQ1rjgOQF0ZF3Zjca8PH6ZfbmeDhdlEU
Y0WXnTdD7OjN7DrD4vltiYCtyqzleld4q4IcVTDdudJU3Zu/HXGilQDgTAOcBf4sK4UHlMaul/Mh
kNm/VI18+OiJWcyOuDKYwzlQDAvEl9W0kcwNXrMGlVpOhVWk8aasTvFJUMSd6rJ2+SbcW4Jc1RTz
E1nsLqvde2nrrl92/Q5r3Yf4TRGB6ryHfqQE8SszOsmJvheYEhymI3ZHVbm9QD3upLWFICUg+CT7
ppqQD8vsExxQy0kcRLTQM2vg4Syze2a7JCMFp7pVJ3b76TBzAsRzb8DFWcvqkEtc3XsobTngrM3A
gR9CnaSrGjAFDTuV7P3tLp1aK3JmN4E1xNyBZD1hlT8lW9uolu9kIIPEEi5A4SFf9o1eZRfSQeqQ
9HKchIWMebtx62Dmxj6QgZ/BekTZmiN5n6iiNIoO0YTXzy4wMuEGkpgUfo/M6tWlpdLrhK2KIhAp
jn9Mug67NG1eQIrN86kujYcv2YX/JBfi7DpKkevtSRRy4et9a7ZFPfSshYUH7NXIFiRO0470QaR1
NKaijd6nAsmZq6FD4k++cR6OGT82w/HcfythrmjZxY4h10zw9ZcLmBGjcWm8aqVonteIasPuDkkY
SAdoULdXnKLKI6Bbkptwr85Agxw8c2+aFjHaipW8EIe4wfLYCvUugKNthjEA5JKUhjvFDWca0Pzv
p+Yd8RwGfOiV2hGZHxuEfr8q4vnnvfXASDu/tituClch1H15MIEh5R4XTU+4+SzRFle94LO8zYNH
9oO06Rn7Rt3uG9ZYWtUSmyDve0u1Hpj4ETwOky+qyr0uVS1lpwVSfro+nZ9D7B3qySycslHDj3/i
XkihbuBQD5ApQKAWdPEn4M9QHah3XilJljFNTJoz2DTSlv7hmbDCpWaoVTUvhvlnYh5gC6WjQx8K
qrCAUq2kMoUuAD6sZa4++b3cytvKkEa1B80drw+QcCP50WG3N3ikWwRyK3Zq3lq/nwF0H7DBZog6
NIlqHs7tpMsYLv+9mpb8O8CqGS2OWokSZfjq9VPnj51lYVeLvpgQ6lZy1hQ+2BhEp15pTOqQg2WY
x64NlI+TZEvJ5HN7jhzH5a+cVH4yloXcSeyIZhaOu7RHGildT2bssnQfmhRY4roSWh72oQLJDJy8
I7m3zkEBO3WN9A6k+t2InjtC8pyAF4KTf9NT5LTGpFQ3+VPEJmyf/kzUq3igp7t86uiQGN4zwF8V
4yQ46eOdioS8j9/Dps2Cm4EDIkAAp56NtIkWv0DBz2DNeWWh7sfnt+a/3ysdJLkd+G/51/H+fXTS
lyAX7ApAmMEv8/D3pHT7YB/zUvRFKMz6Eo0RAmZHr7aoXhdz8N8ZilYa5fND50thn11VzFnFzy0B
lanK6WyQCD9txlgLT8xHx+Lee7zyxKHrLvAxJOxrQriI8kTg5iERIhfesnOv+HQg5f2TtpETNobh
r41ghtqpD0YrVG9evNcJNayzRIktYANHHQEmt2T15G9XYmU65vXbsQStx4E1cKHED0QV9GvCVHhJ
Gvx7rQipzfpxOKBN2nsJ1Vs5TKl68cT/2LHqSVUR5UHw2WozWolDAFFe7t+Dd4hz7LP2a74KtQAN
MsTxFBZdpD/z03xY74Y6BOaCxo5p6pU8phdHTbSCkE9HiAgnHQHiV7lUJyiNekO9Ra0wf2R2hKZe
i4tVAIhzMcc1Yb+kN/4cccEOOb1P5Z3DqWinJ8EO/qgWulAnSIN1F6WLsR8IthQI0vkH0vNIRlKQ
9W3zZh/TMHwXWdQboVvcxV4U4gPjNGr80ty767H/Jtn8te7ADxxmSUcOGC4VT3pnLRw2eWm1rfBX
nbCe9vDELqzTlVRGDaUqjSUTvIzr8wPU6pG+mXd7nXNiEkBjh9VMQIwcf+IHNnImxmvzzu3c7kwC
7aOSJ8HA6BpRpjrF2zh+Xnns8QPfNZiMNrbBpepCH6KKj1VkNqTOwDV/ZsdeHgmh6uVqsBeWUFr0
ryyrHAwf4oYpFYIBKxFLYFrX7LKN96qOowi0uGUQVRNwgN3iMPqYWdH6HtFRrOWq9hldQR9uRwcC
4anXOxBfo7oL7n4NmDuiD/bRQdoc9hNeT/LKZjvLG+8Qs/MhAn7Oaaq37P/UpTNtEbvMUXIIC00R
fzQST9uwsOT9c0ikN9OoUMVdnXNkrpGVR35aijthYjHMTPZkgOzP7IReWpzkQBsK/pOKeu/3Zo+K
LHFeg81lTzFnXwrJy9aKxRvyf3Pt6tN856NjqB4E8BZv2Kj+23FJb2U3q4pd//9HLFwiUuOqTRXp
ekThRtJggIGYm8AshO8fBDNIaM6UpD/oE7wWHbCxpKN33OMeT059CqtZoHmycwA6bLxMST4+d0Ti
+6khm6CmBxdRdlXeU8VtLApLfvedRvTXQasDvSJWsw4DmBIeL4BwFW/FHzFoE+2sdWFdCN8Io057
+2+lf/Ps3GEqWnmitkS9o80QDOtybfe2Xj0AchS8UFBsxb/ntZOTzmhj35vjMxRNNaU/bOJQ4iz1
h1SuxVFoUrQnZlMZcnXoU7G0Sqb58hOS+jfyCxvnIIKw4ytG+I5uWZQb6ZVuIVRzTFW0ACHf1ftp
lXtg7UHOSDW021VEQTM6qUS3pJa/xdJuft8vVCc51V9YKwZBC2F/FBEoEZ/f+AwjMUg8Gr4fgQpE
MB7HxwdZzw0D0GxQSiRJb9jtLpJJ7B8r/2q5yGvgSGvQjsa6ND05WsJuzpKEL2lO+axFmt09M1J4
vsJHHRkoJvNxhAMXTjVF8oTqMnZ5NScbGdGNTkB29vPG0A9/EXgX2uwBgQQVlKTvsddgkTGl1htX
m2ee2o2T8pX9eaI8FuIj5bWOUy/O32IYVeKUocEqHrt4LIdDMAz+9raqbTEFZk8zKa7B1FnAIQ/K
+N5xk0wV+oJbG9b7CN1wRyvIK+wRIGK4D5fydR18i5KITu32qymNrTOyCgu1j8QFGq6ErTu6CC0m
Z56y3lsBCFmZrWzb5+OJtIP3q2vb6HtL2O1qndVOgXc6Oo0YVZM3HcoC4mqzFwghpvDUaGfP5v7d
L/wC4j6tPP4iNYxPlHqI1+RHy0q43M+jSFBqOcI8xIBPcg5kR4vP0zpi+qbleQTBCYRX9SAqSoq/
7nfkDZb7C1xk5pLTi1kMV/J0jDNGQKaLUsI4bv+Q8AWVGpHwUq6swHrOGvjCe2JgCNDVEBYF73UN
CPiX67pGr6B33nEhrcwEgneiQjPmNOWYyQvqprV7qQn3BO4opT+trPWLfbnPZr6D8oTelxzH8Y6c
VN8Yff4uk3FMyIk9kDdqFGlUV9M77cTkwRC0bgS19cJzFYYamTfJkeWKkzFkxwOVmb0+cxIrPfN/
+4+HRieBBJmXV9+aNvoQ7BnS8zzYN7oePGojF6BqD7NuXNKa35ErWxmNDwplIY4653S7p6cvdidz
ZGe1kY7KBhvUr4bJFD0T/Ocf1usl8AdcoKhTP3BrE8zE7rbtR1MIUarvWN/yYLrrV8mDQ3ANM+Ax
YAQidLSYwsO/sKxPfEgX0YbGenIeeWsu+kXaH0iLjWRW/rZUjE/bLuv8ZzbCflVxFdHrq89dMTR/
bcck2LN+DJ1k9+6CYz0ZgL4Y+TkxBzVL5g2PJpMQRhxmIR63nucY9zSdkzXVsMCZRvVNXWPtJTBZ
YmrZwl/uXUjKW6NnA+09HANswZYzgVCluUhWu/10hMdkAWHpxUZ+AhVjUx6ij4sWIXPk98xWKC2z
9V+bkFtJBvbbHV/dWmDyKLBy8sX+VXPsLA70QXDqjXeIUByrRGdlH+FiE1fbQf0qOkDpjrj6nQKk
hFHOh+T9PVEwQs0dgWtq2ZUK5eYGjrZrxn3wmAPdMxuNtdhrGbyu1z2gKp2iMActqGn+0+5MrWEp
scNPaunPXSAOxr/TDhZBCJcsjGnkYSCxhw1L/flIheZUv2WvTtLVtRklLEPrO8QqBNEkT/Ep74Re
C5oE4suVEio3QYO9t7yP3iksZ+gYGpvrwDOPLoY+Sjf76Dz924uihBn4eZi2v8OZ0jj42NxMPJh5
zQEWv67xqHh/cpytB1Ki9Q2VCnhZjPJBaYiPkt2LZWUc6Xk//UarsYy1fkQvPn2BghQVFMax33+q
pdwJdBzcqQG67TRcczUmhpFfjQROou32O0ObqyIkt+97lsQgXZvF+FlH8Lbn+gdvMVB/KjHS47jt
lhlWD0XGtbSLwiKjVfkgujQwUiKKIKNnBhkj7zOyaDA95P7soHTZotvcQEEEF1OkuDRRugZDQV21
UoH9wPf7KI8B5XEoExl0I0z1hUQDa9aiSAIlUyanUegVQRqnSCsbn1tgTMwgTjJn+Uvyh7DoI+Cz
2i8K5hjsml4jjKJf+P0/EdOQ0A8FUZNLkY9ST++m/JkeLgmPnKCwArey94DE4hvuqibFrQdV5clb
2Sa1i1vsUhmIUYaSrKnIIvflI9QxLzhv0NOXaiNJjOmLbgWnBZIHCoQpAarySBLjjqmjXpwbGsTJ
nqrBIEMyLUVKjbdRlz60OUHXf1H+XAirwEee8ZnSJbVzFbIBM3T2Ch5wwjXGYS1D77+93zPC8xXt
ZZBzhdnS71B8Pxhvl1C/WZxAsdmUr1egWNqrWAuYt+DVO2/ecU6P3Ox9Wz2DjdcDR2g3LWELnX/9
xNW8rD/gT/iG6VzBwXwzVvL5IL6ptUM0pOAa5LoKqjC5aI959/cjOepqSETMaJ//She4U+8lbyyv
8iT6V41ZzmM3fcpDE0g+xCMgLPdIulIaGyS1q/g+H+D6lqayLR1/zmbDS5NJSkTabZiem0fp/Swr
A9qI4LbSyqcS0FQHjKGdcusFA7SXMiuOqU+/pE4Ya5FYihI8W163kgotcKubVf46Zt9y+z6CxJrd
VnAK2GpIi5+8QdcLV1gQxxlFgH6Q2RiIwMcPhd7XvhPa+mhS5MehlrKWaKkqu9DBJolJeNu3YCRH
hu2kjebabY69PY7tNTbS1bodf6GDEH+n6jtzb54Ib47MPqycRD8Mtyxvs0CkIdVauPrNd/8rz9LB
ZMXX+XDR+a+XbqM+ZX7adCWjbl69vfEhmcfuIGJUuxiM/OBuHktdJdSSKjT1zEOKKyTH5dZzuazr
ZIQShHWPu4g97EoZtAADu9Jrx+j4d5b7DOoZJj7xuOHD8bsLA1eez6ctz2GvqV4Lnoc6wNlSLlO3
HfasRMTQK+XM1DWeM13VHw1m7EwO/wZWwyusMvfq+tEhraZSC2cQ28UXBOcr5mPS8tGLYRU9wPQO
rHGpnBvVZ1JQ4kpyORtOc0AK5o9wKEkxqVLdyudkXvGnzoZHQgB7aBs+pmb7om+UVmy93PNqV97P
bQygTcVSjJX5KrTt5t42HclXGXzbKBqbL76leFI7Mjs+JkIAN/kJAxIxES9UrjRf87uRlENSbnn6
U/XB7lcXnYM7tZSA007OZuCD9oGdc8NX50KXElWzaJqaLfi2zJkTBb7oh+XLJ3ZibWdZdkwsZ9hT
cDctlB+pCrNFUvxf2CZsUZSmTwmiDi+jmvERukGCvQ1eYcebALdWiUIFrUH899sDBbyE6j2LkkPO
EWDokHNCsp5K7wMYZFaOCpEW68RybM4n+PWEjy3l3AcUQjesnVllYJaJuACrOLWw+hfGSs71uHUN
5aP6n2eqmKFC5IOwiCFuI26mHLRezqfdvKr3ckCBVvhDZnaMWM/XqovmWeRt39NUvE6d9b33VhjO
0nqXJp+m4dEg0gHl1QZtxKv6PI44PVtwuCaF/+1oQA4dWGtELOxeChwXaDGdaa06QzOb99zpa2yQ
1XnmQqLNuDArfsZ0L8+oE3H6fK3RizVVEFJx7SxyE4XKpuTCwk18UH1k83tjw2GlqhJvfmHIkMaC
jrIbtU+2u60pUys7eKOOQgRf4/7DSgbr5X/iLecaOsN5nt6kjiAkRIDNfLmNsdpcQBz1AlBqyluL
YxXo5Xeov+mvfaiIqXNI2tMbxxLlIWphNvYGEuv6vH3p6wAyNAW5YHQoAbiVRYlk5Ly4xblcJ79K
yxO1eVBk9lcpx9OezU8CBqmK7bmKJBjK5g9QQElsztsqe5/+IwV1ITp8fsaomHQoFSBlqrebE+VC
gbqnYL1LRRkUww18a0v6wT0QjqBy+axctnJ31MAvhAt9qoYVQdpmNJmw7FgJ756GVDKXJT1IykA/
Yj9A612GuZzQehoyrLHf+lP54bwYhDLTQMwzpqSzJsgwlGTZuBTwXug7UrNrhxbNn8KttesFc5Ne
VltfhyKl71XZWQi4II5pvPgEPssDuqJSenZ1X97WoUNd/lngblikHt6fH2NE1Irk/VqrlJfDy21L
PwqCcSoogGhLJW8y5BuC4N9IL8Kmx+uopPOStumSuYEo82CiA4V8+eamXSYteSgHfm6qZ42+ixC7
fWir0BoSOTQkrv43vVczL+isRFcoQFWWxSdJ5Du/UVnp/N0YlgWS7m4FYOBrHdwABrUw1BTghs75
zr1WmQ+pJJ9TC5W55rux0+Ru8devaNzKrBUglhUUiaYkGUTLSpJ0M79bOX0taz14N01zjxwA0rwZ
bqWUdju1yFBrT9VJy2dhAyQk038338kD388gB4TM9GxUASguxjPbNOBbsusdyO69Q3d2hH6/USJf
8bFe6By1fIZ1yuUQ1DXu+siUry+7Xy+LxZ82YNGBxontACoX/k1nTfeO2YK1NsZ1VxqffCAlbCcd
EuNVgUKz19wsNkmAta8/0jcbHV3nX6JJ3TTj8PRxV+UjRWWWEEDZR8PreOeNGlyDF0Se87QpzFoB
hvSWmh/CEprXjTxsB5NkF3VptQ8JyrU9SIKi8fvz9TDkf6NZK8uuzeiJU/SHagbKvr5QoibBLXUZ
hz5EMOnTwZA+sse5JGCGfkxCEqpQoyWRsCID7gUXAJHfEpUv5q92hnYAw2xcXWopZhCq5HTE1d2a
4P6etxoLM4GWvDe4W53QRusoVcpoAm7/4MKIPAwnxqAl67zarJF6uuOh5y4DMY7PE/kJQBM1R/s+
g/htMTUCAYlQp6hSyuTZWSzPgUBt/FwGH3KZDoOsM4ohGUKjaWTHEwQ6lV2k/p984MpppAT7n9LT
iaCUSmbJxvG7k8NUFjc3F993M7feom2gslEZjfRTEgtx4wm+sn5J/7CwM6xVXf6SfyPHUcVGQmM+
HmvhEvYGm9dhdaTYHsuCNTDXpJtDwezCUD6C44ZyZnODLdyvG7ME9QaG3osf3HmCDJfO08T9pNOh
w0ujMPPEjNXZQAULjN/bRzK+k5iJFTIq5HmWwTYx5CMXoaUcROCMyDIFay9jlATJ8Ieu7iG/XbX7
G8hW3fMQQEEcO2Jk1WkQO7MKrby4uKL1YDXE9Hs6+NA/Mk3nZnPWHoDyQy1mzLV1VtVtwg8b18uH
RI81MNW4RaoPFgdgEMIIb3QYssMbSgrVCpUplicUiNaLfK1aqcTCqDuOWU1/4/1WuZdF1L/SD1p+
LgIlFzoV9r1bmMGtn4Nq5AofmXFmmqADdZwGWgEoTxCY7l6+42F47/3DHi+/1blvJp93Rarp82LY
FRSH71JeUNtEWEs/mqjUeRNudjfuU0mEHJf+Dv0kIjSqn6KjcyTVnjF7QL3x286ufjVLz2hpM+TO
xydzQu8Vc4oup9ZyRlN8eHdkhULzW1eqaaXfCQ9eYnOfrUWQf0BjlNqeFhAa9atnTeV61c+tOhgf
RPJGXABbEcswDikYOQ5pqnZoowiTGOahaCMnVk+z4OwSr6e2XIjRnqn9OYrK+g6llXo0h1tyMg0g
mWKKA/fabbT5g8yCnkh1eUJd25bUuzGkDLq6aZKdlztpIdSLEhBDGpyhGV17V59CCit7ybeimTGp
Qs+e5XvG9Fnc43iHwc2+H1bUUOuZf3PvLmk8CxGoaEkqB4a9JoHJrIFM0PGBeYMlmoZFRHFQyX6p
Dsdgi8zFT0cgBp+Ro7f9lLKNgSpQ11RdVFY9LDXG+EJO7eAqgqOcfseZkQnYT+njOOFTceow8et0
rX5VA2AG6Ad7zVhpM00LTFL7yA5xvyBMD+YiARQP5E7o4hGPFuolqud47mkrGLStu0yIzr7NR2Be
+05xMoSoU+2lzvc/TxWhYy2tqm6Zw8SxAc+15MFKoqc/IQjLgts/w165R7Gfp6kTX0SBF2qHqw2O
9emf3nHsau+wPudnIdDUe7TyiAQMSpMPeB2Lo3ybGKCBzNOF3PsShIStC1ASbcI+QNh4WeixJr+2
kwfWGeBNGBts3HQ7H277RYQEpuXriZXzb4arSjuUSCrM/NITabkWMXeBZrxC5OWgCWCcyY43J0/4
/i1HmN9QJIU4XNWexztSEScVH710AlEQZvlxMgDhHR1XH0ZAveBfJStK2FktGTUcLTIFHXlIw3Oe
CV1BSB2DiORgwvAQ4gXMLFd7Fzxz46SOAAM1K79nzuWMOAMwitevDd2Lvv2aieopUHzcFt7SrA1K
Gs1kuYO3c9/itEsXUKK/vTV4aMgKCgnlXZwXFCMeJSmiwfYFyCbbZDfojp+Bo/8D8LnGvys7mFDJ
OREhm4BYKpB1i3tRJVLPCpAK4Lgp6klmTXmm3FQZiwLXBD5mbT9J9UXRlBTaz/SbxA2P02MXg2qL
CAGvz27VDG1auMEgOBNlt7YcsfDxJy7BPFLDa4ZVexUnzOg3sgPtmhxgvcvVKQ1is00SPGUOUHlf
Mh2ZGJpA0SayE2JnIHJ/HWRtXvQMwNf1nOpFyShBDwPLXlVeCzX9cHbgOTieDrL19MY3C8T9ZsNY
lhOUeRFQIqitYichMGRaG8Y/sVlrTTr0AbAyXIL5bIua9bD8F7r0PFd5fomD68X7UkJzn2hYLPLT
9RUYkBUNgw35ZH5f/uMtxOyiduYemqQoDydFac/TBWFVAJ5sse1LsIdfSwtky8H/s/8aTqZKBgnL
D13crbQVAbCR5zudITixeWrj3KRv1O5qbhHSIRKnpq3SeAKOOK4g90ILOAUeg8ULQfxSJK261t8g
0F3kaGoeVh1iqXH3f1QCNFKi/Y5tNO2O39KDd2Dkxy61O++HD6/evR+W/DCc0C8SoqeZqadudy7K
AaLowY+4ze6He4Yg6QXZhgyGoEmwJQGnZcZqs9uFDKsvO0nOS64LeAZce4uMppQOqnfwO7ir9wrO
P3tg5JeHMjwLnlk/2TTFpWAVWSrw3YIjCf61WSIvV2f4RvqvPOmG8yYbXYLcQn7eL1jQ1ZF7jwGa
Wmjj1CKJukMcCSYda6of1CCKUIayNBZRlyMMH8kQek/FV4YEST7bzTR8gxW1DizafURx81TTaUqE
2Jia4nThveCsVFcLAstM3sxhglBWT3yD7RezEWpfdWlqrGlJK+tI0Kkw4qtM5RYoZFG9p9MlnCwm
wjT+TOpRNUJjN1EJHIqTzISOexql/zo35keU0RLZnQPDRwUna4nSwOLx/FlDl6dJWQCnZOGzILF8
Kartun40g9JRlQX4dOG30PAhTMcWeyujZpJZS+joEIRL99fdKtyNLQjxoOZ36jttVlD7OH3k0ilB
o2UPsPuq7df7o9E+2I9DH+G3Asks/0tPmVZjHnm7OQEgDjbEREX5lypNywcQz/nkAMN8TmXpOP4+
KQHuRQeXYcn67xZT5F1A5jBV3v34f0GFup4TWKiEbXJ/gA6LNXNeMTSZM9y6RTADz7K+/CwhECqt
3O8A/WgthPK2e+SrahevjLmabTlS8UwOp4PcvzIdOblWC9MDxn2BB4BruwfgJdfDX69Sfe6PpvZM
Ca2H4lcE3zMpSKYzXA3NPQiu2mhZm79gHsfZCdeQ1Bfm0JVXeEAzX11vac2PrQWWlxA00e/WO5Ne
1a76jDYmb8Sv//ssx1j2eUORzaEq+7avJZZixiA+KfWpiv5u/yOsSOZ67pZYkx8qkszkiIemK7HC
VvuKfn5+f4wZdFnRBi8jsc+H948RUBDB8u/N39lB2sPHWDaiLn0YSc4cQ7BRQhiQv5/0MTPh+Qbs
0xUMV4WwHr5qUAiLO7rHMsPddHQwue0Ij+La/ycSDVvI9v5rTJa7h6DRF1Q5cVeq0gzlr1DMsOUK
WB+7/IwqkqY0zuqTCdt4yi5HciydM2Durz2k6wJIRwBHCabyXYAZN80L0X30uUjIusXXgaL8QKPl
1aZvbDMJHQVR1vhoZJUklFtvbjErsejNFej6TE+hIFUkBdtvl+eqC+s8fIDDvsUx4Smco1sBn8y/
Cv/Qur/Cy88UTn7gzbt2st4SpBVwlgbaZupjQmziL5K/JjvnbKs9zh1jj9Rt8rzZSOK/Zlk1a9Nh
lJOHi3DyiF7UeG7GwwYipe0UegZz2kvmeSjlctKJCpKKqEw9zb8gPT5jk8nAtjUmUsyuGIqVI2/i
w3ev0D/OBouknVpXu8KtpTtfryt4H0zpXcT08QB3ClUzkhZBVh7NYosY9EMSq0FNjCCbNY79N6qE
E5qLMDpq84QMEZ5jIyeaa8fog70mfRCvqZSr9NV9NIwadMrWkpwWWM4iZDjzo0laOuynPPKZjCJc
KqUcuWKbkoP9nWl1iOu6zqvAIKAczx1w3qutqI8nLZyiciUQY1BJVjq2uy9qYVBWEe05hpzFYQrp
njwJcYDV9lsGnMeeQlUd261eOyBUZdRQXL1PNc7LCPT0NSYATdT9U9GxUO3+RWJ8Zq84xeQ2dvJc
mxcVBsHVR26rRbSio69Dfc5zuKXChxsIfsvnxH98aNB3FyjbTKAAqQmpjTAFhNDaFoHPbyjOl282
xL6qJ9y0SMR38yi8au8zVa8Y6vbzqK8GXsmQZK13nmGUvuygVEoHHOlDn0YRsTYmweRONYOil3ep
v4jPPsLDwtkP9NzhrlTdjYGXuBt2X2/bqlYaKByMoJEcLYIpXq8R0XjCkmJhlw9yhYnhgOLtti1z
FdVIewuANltIiYt6zGCnJp26Lrr86Gm72rnwX5fpwoqCrDNpKIRrYBBcu3DjNahWuLwfvlzpDFTj
DG1uoE/4WawumPwPXY1ezeHjhjTqMS9MlQsQyPM6rDCv6qRxjWhH81AzPeo4TuXDN6cVZm/vFYfw
Lp7eQcLzvwOC32jqIMJgOZ/WhgTe+b4Bc9vyR94zCYIMctGe361U47gj0WbBIyaVRQCwGca/LUhp
2ehcIezZRu8dHOMJ4I2rh1iMvtXfnCUd5LkqWBduESy3whUwjJ23EvV12qGPUPq7zVcaJby89zJl
c4Z2SCyU9M0nlRzTD+RovLxeZTXRM1ZOW2bbZPmWX4mpypqk24jr684/pUq2NkDvV8ZQ+e1vx/Zk
tlJ1eKvKLMH12L3e/RJ2uyILSNT1t5sZ3OaEe2EXBBv3UGUhiJm/SuvyA4dT156C/SwT919Duo1C
CmvjNeIq5c1XDzsRlc56s2nxjfTz0Il+5FtdeQa95gHCSR/Wd8pUZnjS2myUcCQLeFSsodM5R6GU
R6Jpe+ljjPgO990jPvdTl9MfNTeKWQ2TGGrIQKPzHMdUOTRiKDtOClu0nN0Qw1fWyXOCDZQ68gSG
wRpzL0KphjimWJ6slyb4DPMCA158A0HstVC87PPFJYW4TI0PX9V+fClkJ+UnaImC9pMAHGaE+y2M
sSoDLL0yZpisouJOL+8U06brTX4Goplli64wUjTfTHvao6WuvY3Q+h9cajPWHyYi6Q/qOF+pBXKn
7afj78E19FKDLD2dVdGWNxL1lkVFY471qbOnBr4npXv35Hw7Ajt7x/kcFWja7WDVV/aWH5IDtx8r
3ZE2/CpoL61wa6AW29FlHKUNj3ISMQRana5tRNL9BKOZCzMVMWh/Q1vRp0y1rsSzcSeEzq4fBJ8h
tCAVxiLdalsJHaLJzjslLFDF0CEqIc1Xk/53tQZa7cL4f8p/TEf+qL/8BsadBfkaY1HilHqFSXdO
WWXZUKP+X+6e3/v0ppnOlGYhm/sa52cOMl88XyrH38KM4pGoIVWzHRXyxPK9Y6jHRkX378kd4lBe
2GIUkYEIp6ynHte/MueKZI3OzbTCMnuP3lx0JOAErmDKpFJqF52qwySSvz5G00HyDDJdizgGME5l
Gkx1HX69qLcsARvXbrmNdYeWGt/WXsTOIEugd18h/5o5Z5Xga3nnt1zNNPvLVmEe9Karfi9y9LlS
VSap7iJFMeWFZfKfNwG/qRAr/RljBDEZpsIqVKQ9Al4H9ovOZNq0h0W9vO5al/Nl12xcMNqZqZOU
ueoUTyvjSEN3OCtHD+e6DuQINgTmbhg+5mLEDHUQd3mbLS3InPEV4YylMQZJnfUDsDpkQCx11gda
UPYl8ZUm8io0T7Y50gDz4rBlBTPDAE5WAZx9eiswZNFEhPewCQB0EAolqY0bhv18QI3DoVMszlEL
fZp7gTxflIxH8TqHOvV2ltAQdgeYBm9iFL91PBi46ymTkM3Fdy2gUbQkwEpMGFZ0VivqbV/wQ8zO
ePUklgabxAm1vpNXnZ6HfovE3QpzSIOH8yQoq2mHg/lh2jvhXsa26IU+t06vcpZcRPpqZlv0KKSp
QQ+iSuFEpac2gy/xgE/wdw5mKFCkT52zHa/AQJY1U/abayAkjDNmz2cQtfRsL3g6vdVqsvVMkt5z
H1D3DVueMW882tFtLsaah1Gwut/ZjNjV2q6qvUvj6HhqvUN1WlyOg9Q0+1h4OSlUOdxR8WlLWiLY
Jq75F0aboXJ/LhMPxrrwKixTpJtJFMzU7/l1IODDSySnqlBki2gIXQvfGvl34Ef4kxp18Zcp7WRv
gtsIfzEvNHAyBci1V1PgG8YNXNrzseSjUXSS0xtq+xUFtPSDwf7AMlIHYpdAW1pYnaoYGpXINmrl
g0dYrgF/2uGy+Z0LRDck74EHsFdl194VnM53ZxfIofPU8Ur86cn+VBdbDLJ7OMnpkdGO73u3VBQ9
7OD36kyZOa9/LI+kqhr5FMYEw+i3N3GJgxdGefPRVy5gJMTwOt6XxJ5kyS5LCO2BAMyJ5XUAnCk2
Ei04aCQHUahaxIqXs5E5wNMwDH2kux82IMtj8ag4o0uj+5WrXPC0Lt3R5a32ria8OcdHS6aUMrlN
y3jySl85s0sSeT8MRBwGhHAogR8ZOOwo2k9qx+JP6lYZGRNrEV+eP1uuOwDWzT28CpbMQpnhK753
ykQEih4so8qxk+EG4m6KL3GxtqqOCPSv4tatEvoF+a0LWTXWS0etczS3c44CMKJK9GG1oDHcE9tu
8FCccF80Bd46QlsSdXrUG6/4XgSshGgQ0YD4IgmGiyXOQceGxxf8wBohDSv8ak1SLGYh9Rk3w7nd
Ohm0gQtHCBHuTbysYR9qGXk1C/gN/1HMQJVgGRAPuyYiZ52V2ZebHfZdEX9NF3T5AUDC9JdpVG5e
q3vZavUY7ZI2oy7TFa2bgehuyBY7kw2w/reyLXy0CKmkD9VQh5Z6oFJc6ecSobJnCY9EjgRhsDQn
cnpMzfGm1Zy8AlbYofGhsXmtiNUkOu7cP23u8cVNoSW4D1dguaj70735joqm6SrptfITajt/r8Fo
7T1oFAsp+FifGNrA+oT4n9Re82oaWGjSUOdjwQ2NqLbnfxQ0KbDJ7hWPFqej/aaZV/1ZMaUeMJYl
kGpEd/AipBG0gwsNM8AyuZgB9HBapeC7wdPQxpW6RR7fc9vD14pGOwLvWhdxoVjSQpIGsxqaiCgs
2xhvzJjLtBUVOnIuiI3HzKCeyh+o+qV6L9xoh8WYfEZArr4hHf5DeYB8VBj48/HzgPzSPC2XGG4+
2m1TiU82A8sW2CxGToT2mWJcN3HBk4uz032JfrhGDTKRQpiC7OBjauRINssa50ajnx0WtJ1dlhTD
u1SQV+xv5P5kbanNcycMVlATmJaaPyuyqqtJvmsd7wh9Vvs+85w5+TMMyfxDo0O0fGR43sfmrFIC
QaJ2xQBfQDMSc4jFKC3yb62bxY1qcpYxcyCy2dNOar3iyo0Ic0qgunHc+PaW2h3u4nIiHpPxnH9t
REWwfS4LLjYtS8re+KxuFoE8gkayjhb6lZOwiP8vg3ddwats7+xkIjNCQ9IR3u8o8t/MYtyaAvBJ
GsYr74WJ+STUWBmsxI+uQtayJVxCJm69HcclOeYcOjiHQw8HrsPxLcUNbEGM3lFPHYIOMXWR3FVT
1N8l3okLb3aax6b1iRvjevY7aGgs79AJ5t77aHE2aYyYiePU//NeZjxtTN65CqXu7waWkc8IIGQz
EagbTRhy3zkY5/IR+ITTkuotVy2ZTGaA8P1nCVNWSwEHjKhBTVs/9o8TUY1nSHeGprVmw0vHv8Qe
YBlAcha/yCJah2eFn7jdPv1yGVcbOhCsNraY0H7UEN35ori0YY/zkmWuzHew/Pz6bSQJroN1imFZ
qMVqdIKFir0oC5QvSnrNxtggl15k6WuWxL/hQoo0CGNtopbMc4Vv+8lXRshLDTCbinU0tasjO1za
vZap47w97ze8mTSdwREQU0raTCRuloUU/wHExStP9L9fldbLtRKugGoeAU+nCLLvVJ4mpdVC/6AU
v7minSa6UpmiTLzxIQLsv77F5n2GIufrrrI8MYyyXIQd+ijjsvkAqT1ViS898fAlN0NVVpHDKhi7
euRmAF8WLnjPUWiwyeDFfbLvA9E/c3vGVONpYZ4rBnhqakjVTiAVukIIVpZjs89mIxrUjDVOx64J
6WNBT5AlwyR17P9bfsO+yaWSrYnpKXJ+aOaLBXD/xTAg9gnNxYwDoEtd6rVhn/v7rxD462FHlnZX
xH6ut6shaIT7rY9u2/+klBkS/PPbWiHzZ2IwWLEkV1uE8KqIOLKdDYM4tMs2sK2Y/sT0u/nig3RI
v8RZjdRKfgZUvLcNLQ8ekfrd07+vXe3AcPaQ+dbh2ZsQDulrPoji0Qx0w/EtX0OquCfYWYnRET4w
aF1YnpFcPnwVKA6Z3wbfpy8y3VuIZXIiXfBwRMtMfkV++Bkbc/yDKn6E21KbrmwUnKjTGiwdSv8q
gSXrbuKQwrO2hOZhfKvB4+qSYylS5FahbprbiL7Oa8Vx+ZMlavra6f9DZzJCIN8Wl/pnM784QTAH
25QUil2KouZhLdYMqZV25Ze0dFvg9aKGkL68xSIq1FgwkJcT1v9VKuWBpDaiub/Hp+rWjkgoO3la
OI5o53aDPKozhoITVNmHDKsetKPkmt0MR8/yL2Oyc75qXnKStck50EVqk9bBPsHCLd9YLhv2Mp7c
8TWgYxaZ80314DQK8DFSqulk8a2ISpRtrDQUvb96JGINq9QxJ8oOBmbun0Q1ET77VZ9kwb2e3V40
BvPPa874NOTvZ8qvYagMuD+eeK/dzTmJJ6zOqGEY0phnex/G1vUCpFpGtq0RaTWvgPzAAQ88NhqV
aQ6OfNaIZNTHl98rjdbKt29oI+tXUQmnYDi5OY0WkQb/mXye6Dc+Y1ZRgbR15/90VaYeZis+ZD6o
kHExWPpuDi8430JklImpTEnKhTKznl4hdOnSGvvJSH0yD/+HJj5kixVSMnqE2JelXLRUnN+eXa8K
ODxg5irDeP33xjKThDCunBsVLq8Ucr0V0Jnkz83mRyMf2G7NRRvxWHDd9A8BhxxfdDNF3e4AqU1M
hNh/oJtYyvgrF9JkWufxZiPowmQMQWjF/zYIpefgfO19lSIiaT/BdLQ+e5ImepeJIlM27xRbzdrl
gwDzxDjyG7+ksicMEEZPVRJvA9G14krNDYNJPDDrSPKv2kYhy27n/JlOjgRhsIPeVMMt2TLpWhXc
wWlCMPYOl7m9+awFidNFQQRAqMhdCr86nTXWdoTQ+TgqrcAIQFR1sRqHYpJVr1gjgWqZ16d4ks/9
mZarHHkd8RcyHuSwElpQBs1LH5fsOgSVFFG5/1+LGAVpxHH2Ujm7tOaF4zf4rNl8IF1wI9dpHneU
WXA3CU3ghGBx99AzLZn1weKXpfrgwv+asXAaIIZKNmE6t2U7OoRLNyKbth1SCYPMzdHE1mSXqzLT
F/LENX/n3QMtzGjfawqmq2iSPbBLwO6MoHZjX4NdyhzncMGpCliZXeApIzlXHhX62AP6YgdyEnQO
f3kZrmrAHV5BJ1rc11aDun9XiKbn5QMjH76ZHZrHBpUTrLbqcUWhP7Ji2ogkNaznm+7iHBPjOJiS
Y0EH0GFqeL3uxSazGv8zI14AVLkh9Hfi2JVX9PU7C2Mk5lbSaUwB1NK12x4oCLuN3nNJc/a3ILo7
1z4XQ94Y+tl3fPFAUOQp42LsbxYmJd82MGBarme0JdisxmBJzWnIcRaE3mZ4d2bpuqv/Quw+Ieyu
Grjl+XWqWpuEgRIzpdXnaugJGWwVcLgLSx0s5rx+3nr29pqL69iiClokXAs1TxD9r/V5UBnUUP0s
u3HWmFq+PpZw5/IPJC4YFjwc6Um+oyfLsc5h90jrHDV1+KCSEW7m1b28D/PaemiqRG+3idOTBep1
lmKhLpv9bVzCmowpkvCknZkIahvOCL7zXhySOU/KnTNEZ/enNjttVwUOSANSdESkzoA0g5uYjLgt
5FPtHcOzsZZM/PctAnJXuQG+3gYRvlrg/RZLOo2aU8ZH3EIHOw6Rl5UMH9zeY3T+NONzCQhsHPtj
IaDWuFJZy8tiXG+GEyXk4y9OPrkUpmLM6xwE39XGQiJ7S492aqsz2J/cx7HOT6SiAku3+k3zb5Wf
ij6qOMXd6ZPyfjyML75djTw4fQZGY8pmMzGG1xbvPUi2q9ETUDwwuZKQqt+ESAM5uQMLwbKq24Zc
Fs8yI7Q8+FrdjO6/ApMDbnyspjIcUkLwkdDyRph31TzOZYUX6N8dXuz+iNzQ65euCQXaFs4NRAuB
QAa1xmnr2oeBgeuJ/E82uq6V5J00Za2Biym/xOp59+SnK+84fvUeOb6kLzXMLPKjuokvHQ1A0Vkb
rLoFSeQFYR1aO8dvSJJWQSMU/ICma805TL6iFJENDVs1iaogrGowiISTIYnmauEUKC//mKI0K02+
4EpekzDyZRr5KS7NT+oo+q7P7b/OkVpKa8ackHALHsbVvKeWXWAabqROnzIJD0WJGapOREnyGLC3
rWCnRn2tzywTEORgwbTitPsI3tKg+6rgXEsMs/d57U5f/HWNzOnml0kIRHbsmoivUUQ5kmdnA8uJ
LmKdJwZu0qDwa6+w99145IfJZHjFemvp+OEHH68oN8LAN8ObXP+vWy/rUPhna5BCcgS5IXNDxNB6
39Dl6nVLaTVNYJZyFUeawb3CH/YWUk/IHBvduDPXFBEmht1ONReOw5ZB93EYWN/++lf1PEE6I16N
ifrB3doVX2c1N0lgoNUE35MElFb9U9ReZHHZ+iA36adIw/xt4Q04MfvFEEVS/hmH5/Kj4jDwG2Tz
oQ4p2pvLJgjlpHqlW4SwfqEE6fWMCanBmmd5Ol7cUfgl2056QSyQQW7QIxEERJEVwz8zQmA0jDe2
7W+0YSXsTRjmx3bTRO3c9ARIvLAfkak2ppLk1XtTRNK6KrOw2B3/X+agRjqIemhrbLS+FQvunjSI
g/r6xotBZkBSuuLDp3qNf/udZ0aRwd27TEHqVhXzP7E7AOHZ9DTEvBkbP1x//lC5hhtohOeboIx4
PDNtYqhtqhzypED0mQCmq+wT7F1dL6e8rla9QNJPzzVxh12IL55/lyutBBgucOemQVfyuiYRhyZS
Zv36F6qRAhzlA/LJdczPEGbj0XiAKK9T4yigJy8LbgtpuTC8kNrq35Sz0gynKXQSXFtp/k6d4YDv
9JvMSc/0xRnzhkwyB55FaxlxL/3ya4zgoCSGdFftyqTCPf0bhpB8kRMWgBLzWP/S8Sdbg8yuj8Hc
D4aeJv7l4BeE7xJrgErlFcSNFWidgju8osTfh3+3IBRfWJq1KdE7l3pad1THl+8E8UL8EfMTw9rJ
7LEktixvAvgNl59aYoQLaYocLmXqrxJAecE/c2NTsRqScNqQKeOFiL7+ZFjsj0ih1L12nwOD7zph
g12LcIuKghiXwDaBG9QOVTSNY1tngjdELiLHH1zMKF1vKir3m3RR1MSGgQJ5NCdnnWeHEJa0oq+z
uVcSsEMrCUhKfO9Zyj1+1iDSlHm3dSrJumXO8B4FPd1I87eyylKlU64jnwNgw8P0+hdN3K9yqdIn
iXMzTZ4XBau56WWOoHBhK1MyqO/j8yQYRRRAojt237cgeMNwCpIjMiOPtcc31ARmUOP8sVH7mjA/
RyFtoatxq3EOFBeMSJA3la09znUgYJdPzbJNAV7cJgWUhZkKFirwsW9PsraQkSu8OVidQrIgpqUy
1s/RlBj27RNbpL9+PjHpG7+JgyWvJMs7sbn9cUD4nVgRogkx+o4UWNx7myOtvpQh7l/VN3wPbx0w
nUK/3lp0d7ZcXnkZg9c8W6pTpgIGLrQdX8lhWulpzcC/8UaVliqqBBDTyGyPKlGGN1jqnx8FNiwr
Amh6e83X0LUKYJnOpOMlNdOE0HKT52GVgMFo0nyxWT+md1rBg/4ZQzwztkvep9UFhwY/rYuDEJc2
XjtpyrtIWmLnYYs3x+Njqh7bY0rZo0E+yuZ8UjayzxIA7cs8QGVCOjrg/Ss0mKjqu50VQefHtPd5
W88oLTunugJ/WhynOinT68pwUcC8XQ8bWOzdJW7C1o+ZLwIe73E0+xPe0BPFQLwvEOHmdQHIhXFR
tQ7jpbc8a11yYeI0tZS7zUxd3W5KYQUtULYV/7FL+NJudCskammzBtMsXy8PiY0PHtmhF/eC5mad
6DBYerKn2ZV/RQrS1OInWhOqUXIKAzLPBwG0FMS3dUanjk3sD0e/EMCCRBAyrhj6Qnh+OdGqgpIU
Htawm+9lf4KRRMCI86Ei4s0tf3e9IhW5RyYyYdoITf7NkwtoeX9gw3D58E5hEAdTsNv7y8nO3doe
mtOkaKr49OB6ySfiAAkpFyelLYmLiRN52AZJNvqng+/x8tZbY//+Ru4ImbhpoE/qxnPnhAM6QU0k
U19UXfoZ20+z/TZSe6Gbwe/pm3k+yk/iPvgZcH1SglVLGXPJ2jJufU6wDfUAjmcsvGdp3vgKSfUz
wQrJMJrrU+6z6+l1GQsBODwRC2hnSH7BQq1CNScPtymu7F6ScGjehqWsMyNUQ7JtdXuI3oZwNgF+
vC2z1juWxYOvF/pr/APmSrwob0u4HdgrFi4GINMtKN2LGah3Td7Hh2t9o02Pq7OSSZZiwl1ps6xl
6KcCdvYjTqRloqPZTKNHbL+DY7ZJOUKuxeSS67p3aJImLQXxIKFQMOvLoK3ZCs/KAIQrnCk0+O6d
KzMTL+/dldudrGdGnySEZfTVwAkvgCYmIgV3Lfsj5SZHMV9nElamSicWHOb1L3nQHgfmCpLlIx/I
NeftFf26JWPJyn0ZxGYoOIjS3OBSP9n02QU9XVsfK4Sd+vd3y6BS+GUpPSr5u384U3ARp7e7LgjV
K5H1fbeTJQ2SDtxI3uNffnFO1/IvEB98NR1YSsqS+eCrU611ppj4EGdeATO2bkygVbCroUeTFWnl
meAnsqV8TGSOO4y6LVT/YGyOhCvupqIEuIEP7WQsdF2aYgv8NezWCdi8h6NrhcRkrt5p7+Gq/PIX
6Z2XH0GeZGnVLRmit+IdAKJZjoOpBVOSym8sJohIO8s2wQ7bY65+sfR6+2PKUQFWPmIcUwz0m75b
c8bOH88Ha0lwy99ysXzH+G930/HibJ4jImFry/4wpowJh22kBWtKzxEHlU4grtERJeiHPFVmWnfF
/OTyr4yTRVP2MwidhorXZCiuPEeKAtXiYqZGmzFGTfaoh6hWMAG0+RNBZrBBk4qjSiiVmc4YPTHq
kC5GVOxf0Fv/ZY9DBpkcVvNdwjp+Qf1h70J4Wa7LIQLY0pG6NbWSqr4WI/kHgwIuPOILN9ylk1Tt
ztKpFtQD09Kzokd0hBouT6xt6jXDtEurEg5C3hqVbnvnK0Mx+hg8b78sdBaHZCGLQJVd0j96lQLR
h8jJbv8FYy4HanHp9bX32Xb5dFVWPlpHjfLeaTpBnYcWOu1/uv41s8aAVJU/lI1gPxQvfG0D+GQ5
6AT1iPm8lD0t2o4gnVphCYkCF/UKqgzDjJzFvYVL7UoTxOLNuNInrsCptPSWDNHOc+oxX1IwTRmd
7k5Wojhzg+wQ8GUhjWd8oejTCeK//T40842aYd8ywuUT+fE7dqebUU6rv0o+UnV0/hnlIaSUwxS+
zh3hocByA05qL2CoI3gZUqS8oaKmpbox/B18+QQ11IFZxg+Pt6UtWkwdQefwdRiPVikWxf79IsOE
Op//QepmXhqvQHAOENyieYd7fpxwNKpPUq6KLswO8L9cdV7U/kJ44yJ/1nsOYhN04B21SkzxE4W9
WiuKYGy4X7MstGiPrjZWF4ryZdU7HRNTY5UebFwnnh8JvVEE0yfvBWKJnU9QoNYnwPI9Ua9e+bct
wiOhV5Fj16euJyVdPzvIMiRwsctPwQPb6KInSkw8jAFGwJQ+PogEJ27VccC6R+K2Pe4wWyhetXI/
Fc1wUmC+vEr/mI+V/5l1Md1y0FraueKf0hJhAeib54940KGsV1eqEDdoB71uD/PFfiExJwxqAlR8
vgHx8PXFHeL8/p5/P76219mtMHokVfU9x2dq6AO+mtmY12F3ay00fIrRR9ho3tEzD/79gWplwDbc
7C4JcXHYoMn9YNhqIFRPeGYijmS6gTJfWFYp0tBn0TVHrpcuz2C1uSOWHUpDClu54NISgSZAZoJK
XjaX/3vQpESmDNcqVLGk/U1YJn52uiThVcq4YphCjvoE5FDz0ig4rrhZ906EG8PdvJfxTQ+vZFu+
gPeSfNLPazF/uaCPYvIQsbS4HyusnJ61cw+PfOZW8prM7IcBpnKLWs2rW1YVqbsI7K6jOiB4Za9n
VBTFZmtQ0/Io1CfUWld02u7AwlVKS3Xiysf/7roXMbUeOAi3H0NYVuQwOCf/FZa5s3MDq79nwNlz
R4jM3XQNNuoyw+Ph5DFWu8LFB5Sqd90fCV2GlAGwcPiawdWOAZw++xblSsyVUCst8FIgX4ATpcEt
UWD3mIH4i4LW+ElAJxOlQ6HSwrpGSg1rsKQ/0beDKlDDo3g+fRZw/ylY8BC0s1HYo8QagSvl4jYN
hJz9bsQcX5KMRx6qxs5uHrqR1o8hQIOEK+6q96g/DoGxVwgbnsqEpNSuC13mxevwd5+Pv70D4vLu
WF5o4Gx+i5Fp0JrWh/e20ZGxUanM1kvTc+FspfE3iT/htvm5xsjz1UfOrVXCDs9xoeUsxpYnkSUz
rWSXSUtRurNcrNLOH6QPdeUJR1JGOqZ6vfRhk6/5i/eLZMJduwGr71fj1KJ4QWVnojzLEoNJnLk/
clDIyY7Sg6hJOlCof+tT7PeoPPwPlY1pyPqIbAs/H2mSGkCCg9/cl8HV34TyvHEIGJNSbX6RNwSH
PRNRi4STjF/TsjDKQ8L7iKRxII26Q/1iFY9kO/MJ5yVbXlLXanJy+F9LJBxbqYr2bq+dpOuoxKgW
LQcxGXbjT/8RZnlmAU4foS1eugRI2DGHfeopwAgqQ/z4T8au1php2Q3biFi8NVCUZ12Qbuwlme+C
UzxGZsb9i57WjobBQbdtTRrjicsm3FaI+fyNH96Z1QkJIsWGoL+dBVO45Daw2V6nJ4Wj0jVD72vX
UucZFoG+sf2tyAuYYUnWVnPcDR+ggWDBSHWq4KbJ9/zRUonqtNhVuWhgA+rB0jsHruYPYtjPxtd9
yjRVl+GBE1ehjZpLadsnZxFN+6j1QvHhwSxvxgZY+NjTUfvu60P1J2PX58vMYm6+IGoMPEAVIf/L
vKR/4MfUQXRw8rdvqfaViX/9TSaRQPJGzChynB8tZv6iQ1quawgPYTedsihJVO+4SZuXxJo9J2K4
PXIZvAEKvjrsev0GB63RwGefrNjn8XmYcV1um1R1hYnRRKswup4B+WRnJ/bhS0pmHdUHURiFAA7T
eXOSjq3An6Q0eEGba3voclsxhXw/NuSiXdJmAfufZA2jCL6cdOBBE2WkaQvx16WdFyvkDXO2VTFb
mvl/lrZg6aWn8FPSBmSdvjz5RSnHP2Y4jexhPajTI9+BEZ9HPRdkdeVmmXG0HLL3P6dFu8wK7T8v
ztG0eufkRimX7gQEpgkK2mEt83AM4uykSGWYW2HH9eFCj7ahE3bnoCvQazMCu8Se5o7YzlOKORHx
Wag2YsEL7GUMhQBpI3Wyl2yp265QLGUulO2783OOo/AHr2dI4TMyfN7SiQInQQO3g8Oj70Prs8xj
y1OFtRB7r3CIyTWcq2H56EtjxO78VbyviAUBwb4WW4Jc6TpEXn5xck/Nnzaknjw84J+fHdpupGMo
IulkqhP953OrJaFKv+9IbkfxGGWXbXju2wZKFtmaU/Ge1Olki1jY30Y81OYTqTy1LK5ABXlRn2nr
yHLs9bzS+osLPmf5wQbhfDST06zXtNGfLU3VtXsa9udFXGh8p7HD2OVT76J8WnxCYcraZv9bQugU
GDVwdzDUkPr8Xv0Sz1RwFlsq1PGJcVk8UBf5RUFeSDfU6eEfuFMd2/XMMc5cz15iPjUlDVuAujWQ
7H10tOTJ0A5Jy+OQrZCPZKsHfr3LaMXleIpwsBOkHNqBT7zsjBs3PDHynzkvNbpzdswiPUj+7PVj
FK2i8/zjwu129+HgizIHRHCqV4k1ieea+0eICEEeS5O/hEUtz1b1D4tDLkoGJ+FnBEFkWCurNJRI
Y8vyRM6D7MNvFLx/u4JlnV0I1WHomOct1PPKWpV1xEj+Qyfd2iu9yomOUNhJcnU8ch3XiPZguu3+
WkG2tqi4J/EJpF/mkNi3xrQEDxOc92rss8H3q4kQWEspY8iE3NBKPBA0eDFygp8Bpcio0NZ6FQ/Q
Fpbh0Fu4ff114LomthqL8JNhMd1gQQAVqlpVlQzKN3RWP8/ti6N94cF0XjhxLBTZx12PwxfyCxwg
E0F9pS3qV47IdSX7V4O9gT4379XQs+wM9DYTXCt9q3VCKTxTJy0d2Fj5EFEvmSAMekfakgv0F9cU
oe7Gk+KHm0wUcchfmqJbcPkA4oncMzoDQTEABWPdeTUXivFL59tX6hAigprQIP4BOmCRZLano1XD
Jl3u2Nv6DxvsXy3uB8ssKBcm0KyfsMiucxXO8nOkoNCRkb0IQli0eW4x17Mkep4DbavqgL757pll
081dj17u3RFdOESSCBHJdCnyKJLAI6WVM0gk8jqzeg+DZo23iH63LtB+SCOKcwwkPyB6WbERCI7O
SewM+aT4EF9aU9B1FfKhC98exPoI3yIs4I7ioqMC/BWtUVG1WCjfDly9hjbKI823EcaPfkW5V63+
hQpx20IIjkCjLfd7Vho6JhREjVba5RIVC1ueLlpaOGozqcZjfrESKAy/V2kZf/mKKJH+tW5UfZIg
PDwZVmFiMAO0FhUEJwKlKRUaGatOFODDCXhkgttweFfuAwkg/HnlNIZTnIk1XGVyGwEj0MfCoBFT
s/nMBd346cTIabiGspiZsrqNbm1aaApMwFa8/FahjspmuHz/1b6F0A8N3jBGgxXVcAeY4wtnABWX
FNBt+uMufmK+eMCtc+K7s8YbBvHTWkB8qGOMXnKLSeReXxUZyqDwxqW4F5Dza8K6cktlmZ8U6rhz
UHxOV27wH0Fwx7f82laVRCyjjTK+hdOihS+TJk9WExrEEn4LHH9YMchCu2446gqy8bRfEsC11Flz
y9JlNRggB8TYBgrAaqrxmeN8PSfQbUXRz9au68zDwYwM5PYbJJcXxvMoEDSuPehvqFJIDnM0hDT6
jvfFeveL0nkPOrha0moYhXxQONwx4rVjqhVKxDTfmEjqimZXXmu1/4c9bRwBlwuOaM6WGvWCUV7C
eu5t/Ld0jBlsSXJpPQIOPfEU5aH8VPd6oUXhs8IRB9ndpJf1Sri/sgQfyucGMiukDNYxk2KIITfA
NebT0XblodvujlbugsYFHg2R/f+5a9veN1+acK48H6uX31El+GCuE95sW3fes780uQNgMlwh6ijs
a7sUAxDnEHXxFzfr7IQI+ldkmrnVtLPqGsyVEy1cOszasL91QAY2G1IfCxnR6e0QAMKPLMH1pQAg
lhIDwhRzJx9W3QusUnHzbYOyp2gcjyrZXLDtolzSG52hROKuC1kzMc3KtmjHumRT43oFQ0s0jTFg
7m65yugA1kgOc+7t0MWSjiIUkGTR1VxB9hmf/OqDCBG+tr86yAcl7fmiVrG14bL2L+YAVxzrJhQL
zuaoU+U0bvBOhCqR+hzv/Gs5JtJ/bG4tlemT+F46KfVZf+KWEc8/x5XCsRSxgioqRZ3pLNI6K3HF
TrnJS7m0AWb1bt6cmXsyFGw7UEHdHZuGXJ3FfWMkq3r3VNdNwNbkLyxZXKvw8YqouSZvGnAEztEc
51smPry02opZtk0IN/r7Vn0TiLz2BwqkbeudAvuWv8Sz/HvG0JLmEBbngp0JTfhJFhVwPs/1u9Mn
+SCCFmaKUqGusPI5IM2REzQus9k+TVxuiXI+dH6n/OnCbjpO0HqkGyOMYO+qX1YNmmBKYRp7+P69
o/IOoFppCT3Cu/ren6XjAC3p7zKjwrRcHsCvMjEqkIwnVP2JwT+eVGQgHKJCOwqz4wxNgXRNCY2Z
8+hpDVMFU3XQ6al6jyaERLB/Q65UdtpZxw5UjpjKLyP8gJAeGOccF+iXKZF4p5kmdPEW3/4fcqzy
4k5YWZgG5m/KVS8XmUd+eIFiEyTFNcjB5dLjVIUM2lBa8BycTrqv0thGI/iKq2HP6mGWRBajnCzQ
EZI4EFR8OMA156GVYneUIJBIQ7JQTPpT2QOl8gdmsjbF1rBg229v4hQJolIPYVCkLve6PuBldure
A+12MHW4i4mTmEKjAAqDRAFCDMpAJ1TDguGZyEKKPdJJFsyXoU0lu52IsPZhA8EbL/GR1LBtgvDL
3dePk07PWwqxR92ZdRJ7WL0rchw84HtZcrkJtOuo8JBNTYMuz/ImCJABxL13WVsUacMOSa02Cy80
AegldvTkPF9ZWzBVcDvuuxEpmykFWwYtYzAe6sZaWyGyzSxAXmgHbOpXyqZKOvYjweXJaQtY/LyS
BfrSSHWijlvJy3zc/C2SCZzFzrd9kVTZ6nNh+n0WZoltKFGXSRtmdPOAh5XBAJOQaIRL0nhYaPsu
K/lDjGqJaVqjyHszu4p1JStXeYeuCdUPafsrTVR3j2twilBD+NtS/UUS6QFXs6CJXXF7RP06z02q
eMzdRpR+t3glZxEq7JtLY1zjBesP63oBq2+aDXoRb7v7Q5dgXotaNOaavC34lgXRy3ilTZltwEOi
NF6ZHrllix48C333sMsEUPBQj7t4yGi9MWl70NfYE7pJel9rkmqyNBlxIm9U/jvsV1TilkHlRaMO
2+7FiYquZqRKu7tPmKHKCjhfE8mZeyiIXjknnbVQP4wzWR8LPIhyR3ixQFVzwMcz9sVIuq9RFB+Q
5o8HEEcnxQ6JQH/iUYP+QmzqlcS6ry+izetVtEEI4VHE7GLLn7Z3T782W3TL3/0dPYeGW3uXyL3J
k38GE1cRFWez4rExouxlvuLfCe2oQ99VrI0Pf6vOM+Fj10pn/52DEPkKhsm9ldBMBtN1shalMgPF
MmPFf7phcycpIP8qP5eYPCX5etL/VNQkb1rJAhmk1mJkr/kQNRrBAGwJSPFVxWcvPRQawG0O4qcb
BwjIBMq9xbCSra5fyx21SF29GS7tNCvL07+W1EQUqAQNwxSO6aDS2Ol9iVO3h0U7aCcu3NUCtte0
39twocxuwLBijHQOCei5c8nEZqmYxBAq1eMuTsdj7WtFRbywnLimtn/dXgDtFVP6Aa1POJ/IJxCB
AjcxlDWKy9LPMy6TrZpE0yOAEmft05L8JGw0HoDtKtOUmbuK6mlnnTNabDw5DqHVL8OqpdDrcRDL
MsbM4UkaEB9zdmUCBG1IHPT/jjocJACKEQyMpcbSM7ttgHuRgpadymyizWXk0RJ+aYV3UOXTqXXW
wkKDm9SPyPNmUJEoR8OyI+oRmFzRDaVQq6qr5JgZiLn7EjV/D0zMjRQoog666+iuYhm1rLY2rB3Z
OddsYdB65jJBOQveqZNxTOBojArKJrOlMD6CtpjpLq13ZCbbEAxy+iYGm09U2qzbMGNucDeurLxP
/2O9eV7US34UkDVbCileX8yTf98k/bM+eOEnB83m5fPCTizh6devhNhsRWLdBwEGwn7apUl1tGJR
PPRHUuKRK+x0TRXiivqydA01HtpNsEQqDt81wPT1BgMFKOaW23PiZW9oz0pDxd9sbtwvZ8o/eeN2
bFotDaIQSAxzUFRUinvokSiVt5IdNYCKkhEa/AOiTUGwBZFiH5dKx51QHK0OOd2ixxGjvHRxG+VY
j7FLHXif8MnUgPPo4yhgiSFX4jLfx/X31rsY/HShTjg75IIC4Ipp4V3MgqsQ8jIFn8dqrfs7+tRY
F97wDCZpW5YdpoLm1sIS6i2xLINDw0QiAxuSFvC+BtWW7idaJrgqJZK6kd6Tc53akrq8iQsmrau0
ZHx1IQIdb+wqkVm0S8Yu4GX7MBdsvIFbVN/Tod1fF8kcvG/8FMWZXaPTru0jxua38gwMKT0vjFVC
dGTaO3i6alpT6QcQPPvsbO1G2TdOX13izx32osbyCurVjNg4arvXjB8taN3LjTy53f7H1m5Z+vT1
OWN0WFtfe9kpySWMGNlWeBGyVartwP5sWKlmetR7NFqIbGZKbLS2GwflOt0DEUn3pP8DLIAFMcwq
+eUgPC99Vncw7xPJEluqPDX+Q1O/l2vvlg0nvnhqC/gbSniNuDy6je9FcC9FuFPXxUhJL5yLPhrg
72QqSnifySZ7kbwYfuNYSqmM1aSs9Zt+VqM7HZqzVsCluRdcbxVly1oyJa7N7/IacvmkrlMRUriA
UxPHb3k+oQUBkbMWpM8hrhq6JWvfmA3X6AqLODSPnoFetfKwCFUhhyEK2iHO3V2ROXiwmyIFGbtr
ZWuU0xiYx2ZISehi16EhHkN8FKa6JMwtqrCWga/ODUSFL3PgbEvq7ivjwzzjkDPYE2r1J/H+yEvb
etKXM/1MMqYSkSEDUJcuM9BV68mOIb+578c2YM/PMSDhoGjp3HIhyxLokPzBEDeYFapLcZTbiF4G
NwAlXYk9DuSXexjWc2ncXRnm0HKXwTpcaFY6vzlpwFIOhjYQdmPu/9hw0LQ0pKTKbza6sWq1zGIz
YuFYAS69L9d9vRTc8nTvcvrRJMhwnF0NK4si/7TmBHcXkxp9KHiNJE0HqL8SzkKtOHyFA9ll/aT1
QFnAiww8ha578b7SR3BtcwuET8ptJqp8x5SHDIMD9SnAptn7bpN4DN0DKuyubKFpl3IHqcDreLAN
epMCfBTVbL1KFyraKpkDgRVTuY2AV4Rd8wA8fmBfe1biELI4TVEQzg1ctCSRYj97ZW/Kp4IyAbEh
bkrFxmhYR4DtmkVFZuc+VA4Bd1IgMBJgLXtmV4otGnal8Rcp7VmyR0XtLvnSHZjLOKttwz7A7i9w
44nyGqYpJbOd8h+uxYyl1aXBHd3c+Xkq3NPybJBTO8vlXgrsHCKr4RjadlHOqUz6L7iCiT3iCLVH
SDxgZJmwmTorxEQhwFMBEA6y7K0JnLCQfw0M9ABBQyB0dtyPMz1+36rZvkjCcslftFKPZKkvKqOL
OfquV1DlVbSfOLJGMgudSgtHB2zi2SkTP7ZOqwFWVNDHxwS1bN/G3NXhUW0usL3Vxv7qLR5R3ZW2
jE22gkzLowX9xQfqxbUDwM0AFrKGC+fHn7WcxHcGH/nY6KplE7ZMnC4R8t7YXDC/I7WO1UT9W4eh
XP0wSWm2H1EryiH9DtaP/gQZo4D+xO+nXaVgbqz/RzUgF8ZBT+cqlQROaCvfiJp5qmiFIaEEnG/D
YRr3cbuqYcy7xPSt3T5Xms/L+eX9qdDsda/LsFh9Gi94kp7kWYEzwiiWRbfjx0WZwKEmOWRQJVtR
uQQzH2Wi6x8pSi418DVkkLKO1+hl78g59btRwPJL6IoYNr/LJyAGr2HrBpRr6wocvxf0a1HegbZJ
6mEIWbUYvzXSz34HGkDI0EOiXRuAnroTIPfI7tWldNHIMbCW1aiEXKJwFSWHxBCk78AX9w1V6TtS
0Lx8EF25EgXJUAv0I85jo7fNbkeO8AOAIjKZeHZ9ppmfcTH4LFGba4k+MLhdrjGqsEyOtBDZtnUx
9tOTHF+URj4HJLvcNj0hM+iZP4PNZLVHQVKhClwkmL3Qv5SD5dqD/TEIgUWdKmS73U7dwqNQN0Gc
uURjiREhLrvHysYciNLrPLY2MINWQJs0Ukj1/TzApbASotJakVB48K5tw5ZO4UTH7viPZE4Hv/c1
4k6isvcTeXgVIMe50Fv5oFqxZ+yYkWyYT0G9kob4RcGFuasgCMKPcHMS06skZOb7rF56rTVzn6Bo
0zUGUGd5OjxbWI8UnCszEnUMkoFGIK3r9JM84TqU9Yrpxiw6N7fuFwpT+BjTMb9wn0nn5RxkcZLQ
e5WhMzM/i+LfYMr5SxwgnuLXCn4JarNb5A/38DISjVBKJLSVUKl3n7AqRHFdaXEY+q/37Pr+5p8E
5orSRyJQrlVUe19uOc+EbdnYj8RvqU+dDhBbX7aOl10TgtKMyZUCY/Xm3kpQJzZuc/R0O2NwUJQG
GByGCqVPltRrzS3UwiaRVsC/wgqlEEYy/ORQGPueQVeA5xGi5wEykf15FTRXd0NpwbMhJkgd0M1o
rhHO0wZudLJtza/AyFU35S+DW63J6Rhw/LMXiwzV/eS8QbpPh5oxzLGwypBdZKSrZhC3t5CbuKPQ
JS+3nUNriRxZsVdpL0MIO0pRX6pJ41tFq9GkXLrghZnWfTJ0jNlnnFlRftCoEhjaCrEBHn2yHiRQ
6AQ06FcDP9EW7oNfAbwYIWOx+syaSZmg5Gq7HG3eocrJeWYbN553cVZX/vk/Gz1NpKJ0JJmqTu56
LfIy3R2Po/a1ZEGYriplbmtAIVJkH8746SP43d5w/nHeT1sx5pimdUg8xWSyteFTisjtouLdPhzP
17K9ZP9cFQlg6ILFVGkgqWkI5YtC+s1OTC2UQiMRP5COkQo455orKXr6SMHwwqDabxzQkB+KELIc
6ZxQvIYoBbh0M0BU5jM4Tpqnjmd7E0J0Cb3/p6/D894uC/bjzo1hXR5SgGqMyAbkEahTQ+uJj4lq
LvEtvgbc8SX1+CvdU4foi58A4sCNuiUSlBDsLKYkW8gPCICMLSjSiXctWlQ7EG9B5Cd5D2ERBrFo
KU1Dpy0mSXs0KoiYQGldZZDIQ+qAZEeSvwVUBzzSZpxo1L/L8y4XFuCscZqHpYyRWsuW+nKjz/at
OcopjlR+4FDUunyjlAVMOZEjxSWIdFQx2+hy1bjI2hIeA7WIQzPOUbxfqKtFBAUqhl+f5E24KOvf
ZMwmbn6Zx0nW5v/Kjdt6ldzwcRIVSUGR5PGN1Nzsz2XrcdE8tR5CKIxZjHcLc7Y+zupPFfJY4TGh
1c4prqnuFUaYZQ+uZ5qdq68f4v5D9j/MmdMiGYmcCkTxxf5+8ZK1HneW4c3+WF918vjkHr92lv0h
7W98VYiwpJhTxOOQqswOsLfm93AkuNmlcL/Rl2CRxsHVzi2tn424sKPVwQiL1ewlRDkSsK8q9VjO
0ShD21MnQdTFcTGy5n3Ewip5Cg7KkVAfsUxX71mfEByPCbnCvcTy1jwUnCGhOR5h6Q9uY51f9Uom
J0Xor94HQ5e/Bty1znxwZ87ybaDuI5xjP1AJc+rT/Aql2jGWaTSES1IYNFxx3V4KX+WZpOhHDoOF
tDIKm/qPwvLsasiaFXAxFpfWPXjUE6kDp/LVzs7C7zEivzVM37WSu87zfId48Ac1DG6HqnS2acfB
ZzhhJbahQ2FiGPG/D4AhT+eJn7CZUjB2vGsWY9LwbBFIPm2dmeTYoqlfDmHPMiaC2JMZBja18oz/
U8QnDkWIjL68LZeS2O4e9bYuaF6CfA028hOH/Xkt46UMPtZUIHwSDzE3v0vXkZnbD/SY38KfWFzw
/ZCjcye948unFIzquNaT+SKKlD3GAzPADQGq5c9Z2w16PM5l8mKxsiqr8NnNTiQxoLfmACztw7bn
J+vmnSy6jaIikitx0Ob0GGBHu/uyDq2uJIp0/ux2CCSMFU2NWTVjh+WXND8ePVhXW3tuhXV5ahRy
AhjYrhhJ1ljLyPqYXXTm3TRmU/9jEzjMHMsZmGo0vG6CIlfNjIn0A/Tgs9d3NgSuvXK3eQdG79AK
x3Kr/MK8Z9vB1ooPjj+OlED1hD+I59Xx46mvgnruHs3Bmzj0Tpsb5Ra+rEwaAfdYR+wsw5xwe/Gp
RlG9dXVb1Zecuy13Yl04BEhO1EgtXPOfcRz3b2BND01tXQ63wyxIaJH6pvQNAIfLa3W9os5eG/Nb
bm9VVHV1GY/HA4NgMrEBBwK9IGi71xgXwnOdlrzj99yKZxrxWLmeiuvz+VxdwIBorpkytAejGmFm
zcLrCtXNy+phwzam9nmVyGiuK6rWpLFodhivWMHU4NcAaJTtrqPkv3+m+apid4RJzFSag0iE0DR1
gVuox74UNCch48M3jlYtGfK77u6XkFJQA3ljODN1SEUUcqTB6m09k0/kB58vh/Tm6wzj3KT3bPhS
ehz/THFRR9KY64KDxOuVLCVcGK0/a0CTHSrBn3oAZkPcNl2NOsv8egfsFg09Y5cqzA1qlJzwjazT
zh0eSTfjvFkY03fSoUaWKmW4rETC20flZxvosdAUseCiHgLwa4PXF5KZK3hRMxV+KW9UUwJIveFw
6e8A4Yp1kIc3rBFqjph+uMnfpICUlJl5Aag4lJOVuQpJ7x2Lufl4qU1V7atUuol77+YwW4bVYfVE
MnXPJHVY4PXyXEslL4pwyCJhAKNm3bBu1GeVW8tmVe3Rd8T/2Kr1jhssDHBANQFgmjFlXbEjZjWT
WCGJ9c57n7+vDHg2Kcw6tZ7nH/ctd5TToNNlv9CvR5m4LQloHIcjGn/qJzZuNAVp8BVjjN6wZvle
d6ymo7Eme7GhGSVknpXm/GXYUHJxh12oo0dthCBHZtDK87l5RmYnZ2v/CUu9xU0NDgAaR7lBluR+
XplYO01COyWHnpeAJKUrEag5ubgPon0NLoH/ewhZy65D9rjDlXB4SJXtvIa9opndbszlu9kxTFQL
94jhyHdVRPXWSvpnqZ3ptI4jurpUEtJ7MxoPkhvQDFxNvfwou6kAD3rIrHEpc1DoX5qek6HkQwfu
5/a/OnvS1aaSuIk/tf+tAH8VAI3CqvC7nhIP51IMIJAThhFwkrrmHa7zdRsy2QXoI24LNvosKx7F
4gWJ5yyZEZldiICpJQ+2scbDmoVWx9BvVnGK4UuaORHekjKocQQVGl3iI/ZJ6EsSzuhjoNyrLZ9W
0/KQDoKXAaSPmOWIlvsmmfVWq7epAyidVB6xqdyQpk409pngBwqd5F6zj3fq1ySdsJBgETJB7Y6y
ndGJEtzkTD5enydWtXD5j4xJnncly8hMw4Tsc0r8Wby92twuQxwwhwE7BKZU2fTHU7O2t7sj/n66
NEhRPwvZynf/pz148eLhsUsCkYYS2KhsQLQObLLeH4+oq76Gc3gKZAIMVGfbLPNux/UgaHqlLRO1
V5a2gxBaZdrvsKSXaU4LZcphr/mVg33HMPwNMI+G3sbx9ZA/HEgW9ff9ZiMMWRc+kfPj28CTs+oz
22xFwT/DJH+pWphxhG79ekI0+zubBDnYELgaXKsnhmRJ1FBwJTu0XxmlkcNWWJlX5FCd2SIYdQ6s
cjcM+xXRT0EYjAlyJjIYVoq2eZhdmA8d/Fdipyv4bcM9MTfcQTnza91cmO9DyZZL5S8G+AKGf8Gm
RPF5q4NZqmLtEGmCgohdDGdMBbhmBBdmY/66eRSeGQqbngHzkeyL0c1DvfVJ7jO6Vkk1dQfhmUDM
fK+3tkqHeWE8RzeUz+iSJxlDI61QDRPj/FEFGmrXjpGJ1CqFka1cKRCyVJggJTmQHFg/V3U+g6gx
cW9cK4DLTELyVbte2JAci0g5a/NmClyUOtRDGn3oURqSqknUCuu0FhheuGgV4QJEhzSe2+OOIQJB
6WASvBjIc6F0pC2Svccbpy2DPUcUHrdmleLcV+6I4F5v/ZidonxidWwwtIP3LNLnpX69HkhxuPfj
r8/h8JMbp0Z8gU3So0noBhQ+WD4vPCdlkgMjE/gtYrT9iwlc/Hs2x0DO3Ab0Eh+G/lqA8KNqpJRN
2BSpm0909oV2+W6cipSV30Qw4cTV8Q0zu+1I2BgouT402vjM16U2+xSzwWtxi5PSVE7F8P2VuKQ/
IvOOb3Qdji+gRElYlfEd2s/oqnmFkuY7doWOW+gHResRp/Dlc5YrXefXSLtGxV1GD5Lfiw4pmgxj
BuFfUuwHWuK1QNHTJPSQRCWSKpZAqhE6Uhva7IrjmFQaxLhdDhwV4CFzwhBfoRQ0NrRhwbFolGnu
acIYSrigDt1mni5eLdpyTVXzkGHBabIM/SGr5dRpYPBueIbv44k09ZoJPTB9pGSuJFHB67Dv6qry
Aw2CiyPIog9hxFjxLwfdoEDdIcWIwXr6LkJONs2amsWzyG6/azevFziXNsVLco/xijgRNXegZiwU
ZNAJ8aRCWXotfbDEMcir9u1Fqn980Mg4bpThwYt7T/rnAe5FMqvgP9+p2VB0jn3D+9m5s6U+l8LH
c/auK5GVZ50VbkA+pkNMnn5lu9gELUc8kCFpRfzT3iJf7ycqvd+SVSAfvO62Wbjrl3TFnnqA5nAk
pgeaDVqMJysCfFgU+OMF39xk+ZxLqINHKA5ORk5/ps6QVPbO58rjeqlT0F5zO5mxA7qrv3W6GWj+
cL2aydtpPmLLihuPYaOalduMsCZA3w0ENPlrb76tiOxb/7LKW3fI7lhpBnyu0r1E/YDNa84SbmGU
rVO80AE/p3ik7RdzFgGp2JTI+YkWxRLbNtq8qi2VtzOAxOENQAl9PrdUvfuOa/rIoDIyNG0Y2hzB
pwR5PEA0pZFTd5NH3rd+idEa1Rm1bD4UZpv5Fa4VmYkR6YG/qGCpVqDA+VshMWJoOiBMnmQmNUXB
1SXDal0hvpf8xQmKdpKxqQmTUYwa4JeyO0c2MX8T6NPCHbM7sh4LlLGC+7DZP2nRZs1qhw46OZJx
daIMCjVNPembH2+zz7HXkVJ9z3wPw1zlAaWjujr5biHActY5RHYN0Z1tQv40Oc7inWX9bNRvmtXd
u5hELF9fveBcuTf/VnWXQo2z60i/RdP62CvtAn+DiVhM7UryAN547cDIcTiwrt//F8TEC/FeMhgi
laMpXEkWX9+ct/XgovcNUszfPMto3j3XYpGG5Cv3PEwWbwJLLIO6SrOtLYHFMGTjuktCPYR3LRui
V1eAHWRKsWmA36jis+aqz0KCvYDTp4ufNFgfSMBovSn2AfvT0Ywei1ee2FCufQPqg40d0cWr1rBD
uGn3zbxj5j62Gl80dkiskkiXr0aI/aYS0CKTE5SKwtQ2lNCVxwSXImC6DtnuYUsgBOJSrmR933jt
1IuMqB3YFZ8iLwY9KsJo3rTzaM+eQ0Ip6cA1pvXmMtFGrBCYHUTGpKjuh8Of1JgiVaY/W+6i7Gef
Kp1M6xuAA3bYHqUKCBuxTEdqolvnL3LGDaq9mn+uecp3htZLZapkXKoH3yx4hmFtcZ/dEmBeufJY
6f3cHIKCaaeOS6a4jIK9b4zrvQBiqQG58rOPtlP26ZTI/GR9T7X3wvvyJ8OZqAqyYyZmCqMYh3IN
5FuMVPvxNS+SE0y/XEB31qVyMYjfZiU/kNT9D/S/+j5/lfZ+kLejIHTxEaosJCbwJcaUS9t0l5v8
EVNTslDgvLuwHYtgqVCuYykpZNPwP8SKUlyLVjNYKTDezRb8dXXN1P6maBylM140IEOc5LauOAnq
B6FiHcj0RIjKIKIRxlDa51wsr9lWIegn6ViGHC++UJmmde8LZWxZDHOubG5jIGzVqUm1ZjwQ7Rrv
nLH+Mg08we/Rh2m8m0CO7RO1bQj1bSUrHnUrUDC8J6LZCmBBR3jh3QvO5VZpP6vYnm3X+yDcQLSd
DkbNbGNdJ+bFPL111A5JkDV7A9shPfBVgXhgQu9ojGyndknQaW5bivkt3WN4SgQ9uVcV55aBUD+G
nyo5Jcq9ZEaWFcUcl4RWdJI3yd4Wcy8BJE0MbSHshzHz7a0R6EG+LrwPNH3FadVlYFGybDMUAsip
1EXiLXXXkgL5BNKdbyH0n+lLW4MZpnIDYMx8xlRCrQoyeUIgV2VxU7BYqIf8tZRbr2kXaKWtL6vY
G0XG2g442aBAXE1TNRku+2AswL7g5T47TTD4EKDJ0buH5B+n/5KvXmKVle5u5ZhbNl+RdzTHutN1
/L/FgvPv3SVTgQK2sN4UuU/d6Y72N7EegOCc/POv+cIGPO7Q+xkUk3ookkOsz9hRmG1EiHSHNt9A
yr8irSa4eAIvGNDw3h2X2R1Cxo3VepD9YssHl7Juyh60vUF/6q806DrV2EsWnuaKGDnc3CEV2Mk/
QBPYCPMD7uHf0Ma1y7Z1tt1U7k+v7mZpuCw2jtBevm1eke+QZgdnxLXTHlZ3BXWCA0bcXYHwHjow
bhSCNKd8cyKGVVULQLnqdVDZOnQ4iD32hhAiRw+B8sqrp1dBe047d80bZCAYyZbSqQucD+f9GtEu
g9vXtBoNbBuaQJKZ6Gp+20y+yfh07biKukDjTKINyk3ku0QZEbYijxLJml/jFGtKLCPhtWc+izGB
EnX7cR1n3WxUKscfzA2kmrbsUosnydfQICOtxEpNX3VMZr+nDtKwykXpJ1CTzD1oEO07O0eys7R7
g4AILX0gYXRVAlYPmYHx72TJRpII9MGt0X5MvWOo+6eBlse3geQpqd2QqmeTfg1DBhCbQ01yw7cL
9qcIQ0Suyo5M0Lz+CcmeZvF/RAS6Lq/O5tKhVdFnLIZNITTq3PuNRLEVhUjiAsioeaU59YUm9UlS
1w2/fJSr+VgSKEmOEU9E/HuxZzrM0GfbfcxqkXnbl1b/q6qiFuRDb1TzzvAEEJXdbLPqUpol7sVk
b+LiHA4Bq/YOZpL8PSbDq/MExr2KDuaBxQmEBbkd+VwS5ushqt+WNVNNgOEjZA6vcFLCGhl+vafc
MQcQYLbgMheFkmw6Zg3J36rEnKVWMnc26AKOr8HTLcu6XsQwO4fLMtfnhJae4FwlQ98M/NGe5PDj
mzNV+01mQYqqc2g3Hmlk9+/wMmHJPO3UYVsKtJMrvgY43s7frj6fNgRbvqQVYFr5rq3oL07vUXhO
G2ffIlb7n6ke7yQVZ9ovttfq5+aMUkzOlKRgVb39+FlglnZbpJyFYF3VtiwIkUWck4rjGtf2oj0D
5QRD+y8RNaX8K4tCHWyjghiWZbK2X/Q7z3IIBUbRNVLZWrnJNRDMCrcLK5WoVz67KWC50uDkBVdJ
3gi7RueiZ05t4+L1W9L+GmP3thEruvhpHPy0a+kv41EMDJCPY1ckofi2OdW3+qpV72nJ/YzbOLX3
MFKy0HRADjMbHXbMwlvrwAIS60i1N4nbjt+A16qKPMIYN9rc24VeGXrgm2OnrkboctR2/fKfK4jo
gEMX9yKRSVZBzzgJpEEg4lNmGLszjRdF9Yq/aK/6nSi1q+vR8da/0OzAgNilu1FzObiN0lbt/M8N
xfr+X/g1d2nLbti3yqC+iW5Uq/LMotOR3RHegAcKbyCwPeMCLbmTRuOZrJ+PN3DhSBmjyX07HBSo
vh8MImBpOFGXrIeuCBTSfPzlye/6LjSzVFVRlX5vmCIkMNmhCWcBGbIvn6I9MfgKqn7d8KjUZtm1
4aUoXvI08JRF6ksPyfh4nbatgjYRSmCtM5x2tOEI45r4FxAT5u1BJWArcFUdI6iN8N2VX0kQZpcS
fQeB0sLBfBiBXyAJ64C35f01jIWw0oy4g2jU2rvSEbKrRdt9n/H1dHuXuPguG02Urnm2cwqMtxW1
bfr+QdSOgK/zRpv8fegRGCj86XQBRNE7V+tTqt2A1597rH5puLpbv+hLbD9YfwSWpz4ER/KIoiK2
xeFSo/6HZLX3CYERSdXvAyZx7qHG7mS/zPqLIOl3TKnirdX5dTI6nqPRUnCpRoNz622uu9uDteSC
rVhw44xbOBXiCcTWszWgd+YyoNWQlV6sqILcW2EXzpbjwHmUEUNghQjN2IZRq2bvRud7pNeN2Ixg
6vrnsHZMCmk3iWl84kKzf9J6Xgrk8j7gfh6xBEB8+Gk26i4eRtdShX09XF3UNvqdMFt+QzzZm3d3
1AzXlMsWDmthrTaQVmmHw3BmwyIMep6Zpla8s2gjEnnVO+2fyIkZRCWCZgkDS6ffmrklTUQ2vodl
7u3HOPJfgdKvb7T3tVDjowFz/rv+wVgd91fPheu0ClkuPzYd6sgF/cFIwulEcglVEeaxpeUcUndl
tOWTi+THVeCY257kLPOUyI7+8An6OzVAVcUfoMZtq10xcNCJL1OmW/5EQcd0Y5oVYvlobaSZgXhT
1m48dNsXXIiSbx9IjGRxPuGrSmdUJP/3ffmvSXPgSZpvaWBAuguxPQPMe9zZT+/83snjx57ZCSzs
AEJmh6r6H3zRrXF2gV8b5zmSnp471UCwnAdyE6Jx0bl9tfp9dMCWGS3k+Y2T8WxrLFVtJXfvxKzJ
jLxymaJhSQNqqvtTFhhZjGZMZqtVZCQobIpp19FYu7NVNDDKxUZqYjatjqKnHU2x5mz9X56Efzye
9iasj/vKOsXdRaVgV25vWnRTRBtX9hy/uXY2Bj0uE+vrTguW1L74B5UQwHiBwnwi/eGc7ZL9NQT9
K9pNNYtLc6LY5bkUQQMSqHNv2EJSPUeZgqbPASpz2GtavCn0Zgv927LpxzysrtFV5MU+0B34SvFe
OvSQhMwnxOt399O9f2NfoJ1iD9IWQsXfmmvYT/o7QHXD0wb5wV9qzZnBCBM/hyFwDS3m17UFI4ZD
AhdRsFCbRkaGI0rz+mq5AcblIp7064ds5skYpKe7w6BhOEPdoMBAtQOCafhCs5dKkomoVcIWazMI
p35DYpX+hNwsqhTrg8e3TfG30fUKz4lhIXUsopW6q4gUIaLsUEUKjPF2uGSZ+iTSCMXNH9M52DGV
SffWMup8MP6qISY5tzzu/69RZeeo29sHd45pBNtSSjnITt9EcqShrvzYuop/fj2yIIdEtkHqg6SD
dHVMs+ZJXFcNlmfBnS1FZr901IJa6vNNcxHj9gUaEI6P+axkTPlEYIYeqrS1bfoKd01WaRXyTCYC
DJCDWYBZChjaC8sI6RGECjfRucS9lnJH+6CToYx7RWvp2joSZYuiwGgy0TFWkVILhaT+cDeb+bNM
LKQHRerlAoY5ku+g/OwibMke/oPZtJ0gzERZ95m6+w3Dwd5ydF/5r5bH0sulaocw1tFF8mnPQwD5
hwOgAt4ItSXNiQMizbxLhsw8EkSqkBeW3tK5Ej3cu4p70DxxE2p7NVpxO/owXlBfQAi4tLzG3UuM
2MDrnBAMLNQAdiDkuxiqzgZdgg0MlmjBMBa3Q0e45wWS8ZRUIuW0WROihah5WJcceMX/3nwzBg/W
wggUlQzRBWXq7x7I+ELAy/bAZGY3CM2HWQlOdVEcdJGFuFuCwUsreVClaQ058Qq3RumldizWEvKn
U+ISH/95HydROkkD1S63/3v4CYGX3UANqz+aR4cuNVk1rVQkvX3MiH5Fpf3IuyLMBYZBNTmZydcA
QOi9IT8tRHnCn/kl4kr90X2og/bMYV/SiGypDVLac6hoXd7/MHUdGC69HVNem1M+gy0SRO/voIQO
9owQ4jkv6YK0Rb9CfIe6M0Y5Q89GU/CSSHV+Gp/0PnNcrZppckGrGo4aB31IsxlbS8P8ZFs9bbx5
m8QaHmBGqNbJ6eJoyYgokNwQcvMDbJFR3pbr+DTP5qixU0mfh6gn3DIeGKVJvQYyxtGP2gHVIUEr
wThvVoVJtcZift/nZqAJ4Q0Sl+xfrNh0X9cJYDGB5zY/5q5TFEzoDOENJKyms+hHrhzr9rlk8Knk
/Wxob0GztmNyAHiTYDVF617iBQs5Bo8WfRm3zrLXmjleSgHjqYdvFhfZcBUjyrkqEd5lyBV8WNVJ
l4zaxh8RF2Gk0MrQa/iaD39aTFlICgCCIsw73bCmpd43siCjdfmNeufK21K1XJuxBXDYFwuezu5Y
Q1Am6FXj8FIOUP69G4scLwObcSIay/EvIIS+1ZZn54/nzdUS+W3Pmwck/9P7dCm+52XdnYvYBANT
wUlEUEM/swfz7zDf/78kzkWeLsxkp8cuFRa95ap+OFbRer1k2L2MH1v3fJjbK9FSgu8v3vmbNx52
5a+UY3bIE+UCJNjgTf7JucoIotjI+Sd7aM1JSlMDyqaIbBgX1z1V7YqbhowIErPMRYe7/93l0kSb
O1uc4HuTIba35ZVHUyOyMXtNB05HDYeD4CSwAFNYmbEVr+a0zOly+r3heRVYWgLjbjiiAi3tIo3e
lh5C4MiZkVNi+PAgMTx5LAvUj8WPiPdwHuPPl4uRpMRHhfeGMdc/QKozrAK8rrtgYIBUPJEnQhLT
mBya9rE2kZ6a74EOt1D+/5mlByZJJ3oxj4aohHQq6JW9S46dWiJk0sQm+rI28nu5P1zPUCieHio+
QRHWUF8e4Vs9dIpcYNJTH8UyZUvj7hPLC7v8w+R1pR+MFpmE7wYUYeW8TE7vdZp1iY/824uDTmIv
kmUIfHL1QLE/SfyJGOH5vYNuGvBSqNqkvPusTa0hpuhPTLlCnV+ST1yX+vo/eBMrQ1oLl6+WTVsi
bfurfejv/7LABnu/wuX58Ci7op3FxVxoz7b8Saxbgh+4UiWRSnw9rRBwhtErhoJk82mY/SpdF6+c
Vc4zVCUcNUz83t2sNShsPlfHoK5r7/NWli/YNqo18IZ8TjQQBIwXO5DvHuO/jzms3tDWYmWmJsSV
lE2HMEFtmvZ/VlZngDUp8tze26DrybkeudBN+qUIyfH3nG+zvvYAEEYgyqeZfNPKOZ3Y/fAs2w5v
ZdeDpv3U56yg/OTw1xj2Int9bUxJoCjcLoXk92dvZN8RDDUt4wGYryjrH4mM5YGQt30r0DYfwECY
/aLg9QiHnck4wIUghXH9X21CIGV8MSHg/PyXVQi+86ZagxTzA93KbL6ApmZjav3UN/BnSDmcZSfM
I07VguPrKZ90ndgsvS304TP96dfBVSGFkJP0f5KFkhz09mQHJ0nOR17FJONUo/kXijOFbpkpC4kl
M2AM+cVI7ARqJs68qtQYZ4AIlMQQXbLR8ULArwdi28vn/K74hAvXefyCn6oWY5+tKPGxqBl33E67
D2aY5dFE5AYQ7wN2T60qT81LgXSSchtSyuChAXsI+bQafVuv0TCzhJU1VOPMbLqNRnXmmNXSNiGG
uI9/b8xJhu+DxpSGpBavqiRyUUN2RH+G3uaw4s0Ha3gKxZ8tE/gwjxmMjMGLgiPK56ZnLwen284G
5asD8gmn4XSML8VMZfkHSxj/cnPYMRyAe+8AImYcNafeD7xnHl8xPWfNm04unQg8j4IiJLGu+VVg
pANxaEw9r5PfApbf+xStCkHQffExqm2mWwpcAC1IOdLcxpHlYOK3psyVcxvjPHumESe/T4fbCISR
S3RlQ9b1smQwOKuTNgJ6M+DjY30EgNA2jyaCAaXesIE6gHfiQHdVU7H7qj2Pi7oIe9jgajJTT/8/
HVzJtXNZLRE8x+Au1GalETgv+SI8skuKlHS4Z/bxrwjeIZ9ZvQliQ0Ue3+n2dFblU2oXF7DGnVhF
Xkb2xXpHiOQH5eSBVYpFjSqHNIEnfQlA98wxv3zHuyOQPGf07SHWDvCk7U/HzfHzgLZ9SxsY5pNm
VdXEQQ0UyaW2SSTG0jEXty+tG644tCD82AfCx9wwAPr0oV+wTu016Sg3A6PIlFbQDydVIzld9xKi
sy5RZN7gRHu3RWAOu3a7bPUMgimqtApEMHlAPEKdKL8N1z794GjsHjXqAYYCr18K9C2oMgQuF9Aj
4PjcxZXqkwJxjZwEz9nNw1xKYeckpHY1pWC788qElZOcD98qs6bllVMU9GxTN4V9jTQC779zsoE9
dEyfQXVSxQZUxPPqEf3GHIFpVJhpuTlfaFK9/s/koeFvTQ/EAFKnlOyTtkEXLu9mLHF9MmTNsYae
rbJK0SZBR+qr3IbOBXRDtl34EV0g46etH4KTFVJNQK3MHys2m8Xw6Uxa4Sk4uQ3hbTcukSfQMNZB
A69pCCG7xOQe4CjadtVSBeeXP3HeB8yGFiq64FVUCGXbnEiIgg1mflVCaH+wwA5EjsAInsDhHKbm
6AtF5bDudRsGMAxHqNTmVGNoEk/X1IkBNzdIKLEu5dicZ1T0LDH2gx7j44AbFkhl8Fhex0NR56SE
kts6UsmJVBzChu8NTNsqtlT5VINOaDUHrXYXCRZI5UPmLUkO2hqNp7gUWyIpU4kvoI+lvfRwNj2o
xNH599P4l6dDVAcQ0qsXRVlOYKKtJoHzHlr2xY3V7sS+Ce3AelciTCKvzsLUa68Slnxy/ttZKc+x
MhDYVNwSxyb26fuPgxmhLQ3ES6SEOTvurI69cPX7OSwPGKmKK1Ax3UAIGlkf/lPn3XRCQrziqTj4
XKnPDPyCVI7vftJXRwQRgTo8SrB4JGKuW+91D3garmTJzQEYrhpykXIZ9S2z28Phr+/KL0JRiLVh
4GdgJ5ty1UvKY+rl+Kt5HBoqT0rAVMzyBEocmxwm7tFhmRrCykPUd6c1+VBhHCw8oklP7h+0vwfC
/9+VChL8JGPngTG0H4gup2Fktk4gEC0Ttp6DwpAVN7CHh+2jASYjTZVNyMSNwAtqcK5szBTGq5dp
1/LVkHCXI/O7nmIh9/E6pZoP/2lojXU9cfmSVeQHfMJQUzREcJQcGahsepH5uQz9XTclI9dBgevF
pPcCvb30eUrl6oSK5fTAWkNO2ZFAe0C0r0K5AebIUaNH06woG4yEBXTuXsF6xQMiOU0w8Ap4vnUm
fuQsXCovyOIgY+kn8NNyp+fD6/Z4Aa/LpSgtsAap9BBcqC7vu4xzdDHVNcYZUXCKfBI0BXDtjYtC
PVl4LI0KY/D43APkg+U0mv9Hti/71CpJ0cWy4QnI/JtHJMZ3cs8fGVR/tyEFS6R9C6wmUg/2E3hr
wd2U/K+4HonBBHHHB/JWnruhh7v7bY6x9qCobZPfa1c+lkvmCXQ2BcRk9dScOi45GU7xLyyDam2M
elr/yMrFNVzKegHFtrIEXnX1+2GwGVUFT49i952qFRTRVYAiBWHGBj42J3JLG/kGx2zlTze5nBl1
FiGwqYHjhIOWpL0dg4dOXQn1ljQ1gvkB9v1TBaLIvwkQldKxT1IKCVyrT06KUJZuURMGWslDb/cJ
zYQE5HBNhDvd5+6bdvOUwCloO4+qz9U54HJ0q0EFdM9Ofszyqn71wIuIbwsGaXqHLC5A0hGME+g5
VLlzxeDaKCvb6KMrk3fJFIn74O8ZllwipKlyHsozrrTfbRgYZ/KKpIdFGXkvzKpY+jEbtCdjqGfA
GKptgk+A0IC4vo2qEuzprGjloZa6eBu43HaCdBTjxph1fcK4cUOIFrBdfPzLv/IwnFu57+sJdpEz
e4xdb/PgCVzSOssI3DC9TZYXmHzMQtsl9ZytX5ToesaISYhxjNeAoRWnbAQgYIZR8q3JpSGXs3qz
l1Jpq6PrxRTxkiRAgqyUahaqOAMmzYNCmIE/tvfvQqUsA0BzVDlVmikL25RIakr6Q0nWkZ9je2sb
wZxETTL1UlU6RozfY8vn71KV5FWr/0pLSleCI0TLI/wfW0z3PQH4SgtiklaxGvzqe1qu8aYIMrlq
k6MXA6n89Isdh+ORaGxWXAAwvsnALc6W+F+407SopF36AetP/DxqUpT9aUgrcII0g/2QpZcZ0qVd
xqMVyM0gtSeyc1KoRhF+ARqWU7VVHOOWCdSlHnuIuMVFGsA/fHXNPMp0N52LvxILDaC9SJROpfoj
a7DBNpIW2w5gB2PdJft7bk0feRLS5oCnDub54F6eKh8+UCI2VxZattKBaIb9A7UW8Uo/jd8XvxNw
iQLEo/HP15ohRkFjFA9xUCNn9xcHpTP4Pg9rLv2RZ1YlEBIg7WR9UOmUHefsm1oeVAffZ7kxBRzC
KMeqOcpukBsTIb3gFKept7nJfdtojxUcN1G0no6A9gU1T7r3t+CwBMh+RC58stx/7Egcg4DFwOlD
FbjldI82m/UljrObo2IuNIkXMt0yq31MrFVYWUcpl7U8lLbNAxcIGjVM209IdXabbiLjynPdmWSF
0z+5FemMzKykUVxMj1cqB9iuf5wJOsae6DG18UEW8T7EeAtCMbRoIiImx1wfpSlGSnJjyVa5MkIE
bEkayjxN77wApjieKUi22PKDYxX8MBDX0x6DXCwGls2gHgh9nwOXAt2jYcxR5IyfeX6yvKz3ZLaG
SRWytsr2km741jL7dEV3lsvvieaLG9/qq/whIfLGfQ3C5cbupVrfDjonEa++rsiIJRGdTKsqACuB
heKk7tGaI3/G2jB7B+tF9JV22YRaVmEpgHQ8wWLHCYrvrbxWrWoaC+iUnaWzD50ck/u1Z44seg1r
gBmbnuxQkfaCZesVHQc36gp6FKLyi2bGjqm40tNA2ncDlYIJ8pEBhiTa+GXv7bIRw78of9h8b+et
KQdED2Kx5tZSzgEdI/wuYhed+bd182zRVrkzbNhmhWG49gLWNqCw/Q5BDO8A5B3+2t/TEZbWoVdi
wIab+qnVF9MWevqJsKgt/qF3sX/Q4VpmUSGcnz8gLxRympwWY3KzOXxTHOwwTpexN6o1H20dcSyb
g7jGPxrcJYgWF1H0AXCkNRVSDZhQndyeJJxS/5kQmI7hbvVXsNcIZkUYEf9UpYJplns4WVsrBmXb
ZnYkHeqltY84b1u8lFT1Qvk/A4iGOm1RAReEYplti3rnlq95ICQer3+D7Hubc4sKslbs2RUU/hsO
vV6/r+GYo0SRGYYTKvp3s7e2Ie5b3GTHpkZe/d4Y6yydxTfOOKMNAT1MINNXrIDKsBb97+sfMJQx
BelJ34g4bymPUOUJ4+NMpRbf5yG+MclPWQlvWqO28Gr/1995Z6UfvY8D68RUarpxOPFmUWTa0wcO
XCN5HBVkBJYiFkMBpvecnAPkhliPoKb4ORUSOZ7F0xxa1lDCuUjMOTXReX1Os7EsOPGnDkG2EogR
5sJsGMM2h9SMARRpBlBm1+WiUtcNggt1cfs/Fkb5LUhYtHSSl79eO4p7oG1YobHQUc9C7g5Qeq6X
jkqAKU1QDrx0Bc68RALxCI4TzxC6uCPqeXY21ijOAIJmhEuB2pVRRRXPrDrIKv/eOANegmpuGP6T
ZXnnZE/C9ZiyMm5HVGH+rM9xyw9kEQzeJ3JpCJVWcKVb8M7bSHsAHo036ZiQGfYh27v04QYOZ4UZ
4tcnaVqqwv5FtDIMan9jmHWJ5bYayvFp9H8Ug4lLcWXsx9dlEzsF1Ta2lf9RvYdwR5WdO7pXql7y
70chdpeRlVOa20mR2uYZFZMU2srnZN+1te/TaKq+cCR5G9uGo9fQOXKjHwuFk95uWikyWLUIDTMk
9T6JSquI0l2SLycJMKotTjniEWVWhvYNAA5akJsG/RK2j/4kQjqu1m6BQbgUK1rif9CwSaC62Q57
dt6OH96PUGpaeLt9UbVZDLuUX2sSON3K7qfrcUgioIocEMUvOsdlL2DACVOAdHgNFbq+X+FkHFhG
7pDAypzDbjN7AgKZqKG1qDcCcKzLQGj1WxfNeQiHJ2kb1QDSSDONpFkpQMSljefuDO9eXzCE1BOF
pt34feNg6n6HBh+1MyfNggx11wxJHJrdIJpW7/pshlm73GMBf0XZychi400nVcQxfMNlKi0zSVYo
yau7laPLPdCn4DAKQk7Yt1N569e+P7XA0mRgtw+Yp2C7Dk9tBRBNRcrfg1XHlgLOtc6AAVNA0Hmc
qz7uaDI7TBZTskl4gY8XjigKVpzHpAWIVAMvQzfg7IUS+ZCGrLZOaUxufshnfeubUoPIBJbwO+P7
3xwqCXgvXHbvm6tFqVempblTwzd4g3lb8nd0QlQqLcTmPmFkdKmnSrW8vsQ52QSEZtDvfZirt1T3
01hml2YL4VfQoHEs8hIZZetrU4GOi64+LAjZG+dEvixcKXuM8/OcpM7vikgDDAYgcuOxaSTsLnmc
3rGQDeHtc2XdtA2aiRgluLpWH4Sh0Ioebo1aAUMigbjzUrf04CaIL29mlAO26IZfHiPhrVYr9xDG
W/Nw9oHAR5p5PCXixPp3Q3vNvZ606Wjy9coxWUC8xHar1zsIkdYE7bE+6o2Ona4W9tcObMKJ6w9z
fCB6V4JPzWkotWx+oLDG+cI3V2snuqF3s5hLOVhmA9HaTOcYzlxMIAmZ5SlRr3P1vxyeLo7Mw/cq
UYkmPuxg2dFl8ydahL514MLnFVJIe9hY+zaJWCvODf23ehL65PGG3PlJcqu2DPWLcmjSjTHQIYOg
EJOiHtOHGSTBZi5k97AaUYj+1z+676iACqudXN9M0RFVOUhc3ZzeEOVacsC2L28/qrhALfo9q2IS
IHotHr+49MP69STbAG69MGV7KiGOrsLmjVANJC44NAOKhRJ3NIHw+2g6RbCAhU9CHbRwxXerH9Rc
0k/UrGxsFajqT8BI7ij9jzupdASJWCkmsZPhqnEQUAl1g4ysMCRP+0w/y2565m/0Wu+S927AjAxB
PhNHfzgXqUmV1B8KfzgLBFn7/uSg6l/8ZpKf8VmMurRtN2EfMLD8ZT0EDQv9obCO/dX8pad6LW/t
Z87C4dTDFShrK9eISj6mmKrvuhp2+UahI9J37RIAi3tpv8xkyCuv5JJgVkux1XITqF8acFNfn4BA
1WmP7S5ssiIm0sZx/jkepHrKdnGHGhpNf8fHiRCBR22Hk5YcGS/mleDRy9rJJqhY4v0yajU9bBqe
tDsT50RzZuyfqzPiF45V2ep/qRLF5N22+Qa2+uQN90ff2JWeYwCAp9Nw8g3aM+nkRfTTaNIkYbLc
MR0w9Z0M8OKUVyQQcKz3gfWZw8/Wgrr7f5s6PtcA8NsZGUeREvjyoteeK9lOpV4Qk8hQTigpLGrP
9U5jYYPKVfmQRr6OwyB5NT7xIycXVeXkMaTYFGNR9MlVKFZzL65oLPFBVgEsBcNggDeNcm4QvqQy
493pCAJ9UktM7aiVwJI2w+L8AFzEIZyfQkS8WLO7/OIK0ZAORod6DfPLHku5KjA6i1L/7vYX9g4O
+Bx2oCfGv8YrF0Ox3pWqaKEL7EGQKKiGkvN/4PQSQOXVY2IhDVRg+3MSFwpwORmLtPIqcCjl4ZGq
xfc+6Dqr1lUGr9/GK86A5RU7hSFVm6uLvbbLGVS0RfUHEgHlEPgJBjDrM936REGYTrXSqdqSdlYj
xfeQFZ/lavlP7WJIzXyFhjF+Hao3f5zfskXgJv2FNmWEsyLxg1Yjlj3ZGfgQX6WpWTOvwcAl1c2V
9J5hc2Qdd3l1R2uacEH31zeJlsaZu6wmeGVvsJycQrTfR468DZd4bo1otYoxaZj46Pv0l8Hh91hS
XRw7qoXYaVhZPfc+nEyPkUfhNcIYmdz2AuGFtIuLVaZIf7TYQsKvmJPywbFn5fD7LP3taE6/UIsr
UebVPQw7ON0ibSvYQEW5s1pylxWPwNXudpCGUf3gr6pTzWYdzh9SGB9GyGlYvz8r268cDCE5/iOL
YdDhcrYIunAyBhqCjpsLCkNHhfLkqiXtRFM30FsRAHSKu7ZGPp+GV5IWtugP5qrH/RKO2+Q6/rjE
8w7obEoK0YV3EvqsI7wPyFG3el6lRAEVYX8ZKZbcsLEx+XYeSWpXPtGvFotb1czBxIh4XjImtjjT
rWIreiB5N4cQVgfvgiqlvMN0BZ7x4e92jX+w3Fq9I7XiWPCu4evNC56PEClRN4oHWu/lIgBtomRF
tgoKd3TiD8GqepUwD5eedJJO3Ltb3W1gp/u2u8UGCPFcaULoIXB1JQ/8s2YENYgNJ6hleh2mI4kd
bpNKgAUL/onF9sXJ5+KZz1sFhgRb03a16ClNnOwQgeuWa2x/yA81fdcYZwwRNcsuKr8e3EHkqE/O
fVNBQiKaL0qftvdXqQpylrdhEtuMcCZ4j66S4IPIxzKwdECpLHddQXpMU/Woo9itZX0je+O/grTd
yHL6gCUFpyn5IHAOyreN/1ucdKoUSZku/BtEWT0yVajRWjZXMKFIdq1zuICpZJNq/gGLtBYy3DJT
sjUbtkID65xcJUW0B3Lnn6ltqr6AsWvcplbh2WUchWdkSx11ug3Y+kYxsnFXUHY+cLE2EsIcz3pM
H7Oix21ttuGKond9gFQUo6mlu8LxnlLZjokDco9zKPf8GAAXSwo0dFtcpI8QgR6P5fj/CVCWngI8
uGA8YSGICCVufI59GzAp/Eqtvo/N/Qc3AqomTYq7ApH6qotQwayN9W9MV5neOpvs9mfv8uW1XO3K
ZTOL6SrZDrj3Lkavy8d4QTm8cYCUN+dFz2dnZZ1mULUARhUYRYMz+7zAk37WhFChh3iFWKBj0P9E
hLUgqEhT7mIBKrkUpDqsYUSfeMibFwdj2OUnX7hr9fOQ4Tkbk/tnjMXJRwIFvunsTiPYb5Y1DL7M
NcSXVPOgl6vDl7EaY0nipyH6COjlz6++mCG82z5sqTe0GsAS9x8Hn7Isn+k2YQT5xIYzfjYMuMxW
mAu1LIoCW8ZibDC4OrSqqpVltXw6b9UV114edMNy6tBCgOnJVrpCrtC2zq7Yq1CB8WaYEzt0SPMU
R1vHtJumPxvXMX+cUCSg7KKIZHOfRbnf43xo+GrSRAQ2S20KFILUn/haQ0TKd3gSu3WttCD7P7bh
/Wca3zfacY/yTYElm7I9mY1JfLFMq7p75cAuyE2ixQvgwKsC5GQZWwhHyJeBCKNH3eJ4wox1C4xn
0ZCIXMawtMTeOKHl92HuBD536sWLiE6piDW/mSpfw3FA6Fd9PmExu9T7UAawxPcGcBByeyv/m2Ub
ZbWslDLsN4Y/uZJX5jAfkxP9MOthch7kZMfC1zoH2WrWVRYNo8P8LvfYF0YDXMARUy7FKCkesKiL
tAXCnlTci8cfotnLlhQereewt0ep7POCM6JyRD9B/BuIF7cmb6Y6oejyJt0ErmFEsMaCCd88Tp50
pVr+QfcZQz7mLt1rGEaUuPU5Cs8JQb5FsLvXauPrV7Z77OuAi5YVdujHwPwRNsC8my82R60PqeC3
Va+ZpTx20XDj/Fu6L2Gz4LIDZs6g9Pe18BT8QnyvfKekjLQC2lj0qmmwk1OG56eQz2FPmvfhkssf
0BQJN0Ig7YsHPOXV7Y+GtNOfNx4UPzsyDJNv9klqAn1oLMCpL9T/xoqWP5wQBr59qDkGs6ZB3j65
q6elXzCet+28ntXQt2ex5JePWANwaxPz0hkAbP/+dbeejc9D7WNFtyPELWadwrgpVl4jruhOcWjC
lPKtCUPEYU5pLH1L0/nT3ryHDCR+0dXWesWKYfC3rSCOM2PhFvu/jO3CARWC/Ku/cG3uzJ6FxZwR
B8WrX8QCPBVUkCGMVduzuIRzglxTjSoYuoSzSiEz+Q86VAUk6tpND8SkPPRIr5XFHW4vuPhmPLmt
sfyUHbqh+o3Tw5UcmxGKLkNRR+BDaA1UUM+BKOVEzmiuAcK8UzBMqu9wAZSaZgAR+8sAovs4Pm3R
V1+KW5up1fEpAjYyHYBtxjPHwlAMjnbQpszNWiGxWRPl9oqT2G5RYksNqsCQypL8DN6ouhMivxXn
mVkOpL73JlyapfGVhr4f5WanAPugpb62HBA+A4dfBlTDn5Jfnrh+YjcFv4PW4GS4APtML5UKHrhR
Qft1stKgoT/76Tu0+LES8Xb40Jz2Bj+MAy1KO4J9gun0uNrsJV7tvq0u7dIUgN7MVIbB/maTwdSv
QbhkqLewp3ulzbjhgtwRwh/sdVxjQRRm3KW/w+tXlO8OQzOKEKpDiscYIbJ5fFDp/W0GSxj6kgOh
bwPp4vDRDseOca2RJg1Yz8t1JFzRKMXRMBbrt4ZOsHRhsktebXiW0Azf8D9qgiP6qlxVgyR0oTN6
T6KRspGaBjgVIRvZ/64AmmFLXW+ZTuypw92o20U0SY9AJW1CqFQtXdoTaRe3AzwQuw/cqZlxdIxl
S4/g4AgcWkBsfQg7HZ9BrDNVw9iODYw+BPNGyUbG1ufKVb6R8OFbqP+Z1RFGXWiNAoGVj09ApGT4
WKzqBYp0EitdDLfHMxOkRtfrw1uIC6DIg4NoKtDf2VUPfTlpXAC1wGKKUIkAx7XR6YnxaEE/M9Sj
NF0pZJihNjyCh5PMfQ+3AidBtHg/RtmwYWujuCg92M8EAx+SHOQb4g+k5DSO/oD2qnoQ7ovsrQJJ
itdQ2TlbxLXcqsqGj1PFTQNS5WwEf2nDv6K3T8QMjxMeN6ZT0aKM/lVYhkAXFSuLUSxLxwS5Qiad
2Tg/2i3QOu+bye4s3Y49u1YcyfkuSBV1QmitJdXo8NV4zP+ZgM1k/pIvlF7iR+f+NCmi3Ou/UgeZ
TQ9XHiUt63B66ObW+jVO8gMC+DV7+n8nA4U4xMjl0MXtpovPXwnORW05mVQUlwMgKkFiMUNg1CuF
2dP/fDF8gzd8URZxwpbJXk+PsmFqejQJX5pIeRIHMowYoaagycgeonXMGgc+oj9NAlggPCADL9GO
aiQO+zUeprZuESRcILxpxuz/CPQNgYlMi5d+/k/fNocVmb5omowftUPK1h0b4592voZmeh6a1ZOZ
xghlqQGN2SdYcDfZI51AMYIvh+g2YmivXLjVz7H5+e6ghhpyvd9FE8fE/s3BTxZDz17935Ww6UTs
bJY1prGzMjZFJyNRP4JE1f5oOMRy0ZI2Z4+oJd0T+IZmcN6FyRscVipS7bhYpphlVG5GsqO3sMVP
y2U1PRows1EPqr2Jwz7VczGix9TpDKG8oAzrkmhYgPTvFG69BMuim/vfKCFeE+90g1v8TrsGdSFi
xU6rhjxKyLNRPhluIRKGIhCC+yKCNN4FhGqrZHkrookq88iOS92DMKy+pACGK96IbK8Jh0Jt9GMV
Zya/da+KukurU4wQo8Xauay1bempgcLh8gT1D9v9oAfs6XU0dQYtt4PASAxPQJn7By2/05aEd/5q
ktAqrsc/IEev98B6JQM+G+bDWrYUx6AmMf5E1bEXm+wPmoUAiy3wBiUpiZNsczXsjscxRnqAZwQh
1e3zrgYnswPIt1zP0Y7cYvfy+lba1+7qiPnR10wf7BrBua+9bfSrMI1TLydRtUcXIldObCO6kJ8G
po6QDKCkL1UYzIoCiy9y/ZzCLkYLM3r6vtqdrU7LnvtUKCnTHhXXwwoAs2hqLs+X2BIuGLWyTCWu
j8LJ/gvnOMG2Thc5T9dfvartc4AQga4g6gmZy0QxYJCUXGlJXPURqZHacz40/Jto9AY5PvlGP7/L
j5k1vl0Mg4W6WJHwkVQ0KUTvD0NJ0FDi98Ro19hyiV0pCcUx+Io0pYCPQnnoinnHDdE7kEHksr2N
zFxfm6+FNqepm0bKPuyEjC61IO5W7Bb/bb+BXDDdExB8LHa5HdIi5rljxJND6X75dcipzD4/DFih
CZIyXgKmQiJ2pSC/lL5cOkTydEWbP3fwJjmrMYQzIZ0oKxVvnApc5+0pw3GJHhWW5SVCb1hT/3ZR
PvxVCm34ey0gmI4rU9Cq49xrGeEejPGkzNom+eY8g/7xmj5NwwL1XqCHapZ55A7tKpbhuwINW7D7
sfECM7tz4iCgdpXYtySWikPDyspqbvgiei5soO4bZODq7pIVLrS97c+xJnaDZljsheTVYBPi1luq
lITmY8TwQUUYDUOGJ9VDETptWgla8H1qC2du8kjQ1WIELJIGKgPIjnRz55qlj1wPb2nQwLpBzmCF
fb0iqNPTL7Nk0La70ccvQBfr5KtFvy8IjETZejc/O6mjISqDKy8YDSxCm7inKiFBJ0Hfsyb85uA7
m+2PwkDlMVo0HM57mdiwMkwbVbzvEWoo1Rh4gHFpwEiPIYoASmlwRJSkDzQ+LU+NTJKkdjfJC1Mx
+rozZs9EoX0MnUUnHkYRz6hpYSF2urOTHqA5LCtzhCC/hJqtVUG8g35HJkRfzcZRhSRBVPOra1Ap
CdnWg+s+mB/BeWPpEIM43Z1rPkiKy/upgG5VYZNXg0CvbtDcUHZIKISvLcKG4H9ifskB8MtSQArv
FDB60s9CKIdce/Gh9vt4ocuuE41wuOyUZy5Wd6HiQeAz8vW68MQhdh+UULTjbO185S9t50v6jRbF
cdIR9St/L1y1kKCmPl2SRuTsKn4sPB7v3kmGcxpAYvIV17BHNu85ZivadOJfzm3AsWOLGNpVKomU
QFA55Hiic1vt8cuiCXg1YAc3uTBz4X2zk4KhqHgl56QFKLm7NaKguCmW1IX5b48/sTVAmHV1P9kg
iRQmJO0uZ2Fy+/6Ss0yzPKCA1JMt0xDPEn2LFeETkQ+Yj74HzlNHDILQHCvcrB51qK3RgodigIx1
sOAoSElWDDG5PXdUIakBxlSiUCzof7k3MYEsEKb2Paqvnlbdo6JqoncxjrTV5+lQeTORloswSYAk
4xKVzzFSSoCQO1W63NodNxU1RFSy5ayhQ/vhi+pZmnLNgqFN3EEiVtsNo9S8LPzDYwut06Vlxzj/
HOrCHOWKDnpHPakAXVJ1EjjBV8ONG65J/ahyjsqiXz+WqfkQh48tH+WXFE82UUMxgSw8pgWOaF1r
eWq72+Oj6AoAKTlelq/E53a8brrWWvsUKwSxRIrssvA3oX7dTNBozHYkGZEzictcj+tL+OBUR5WS
GZ/oZEMzhaGLZQTSHHA520eks26XpBv+7Q2zohDHXrX2PWTzKb8TKf8UM051HLt5eVxvB52KNlEM
uLp5DKMYVNHSORj8i/t2YdnnvLOAkE1A5dps+BzzGMVP9q2dEiW7Z89lp7DKSAHAezlLxRMIQDxk
xlyPZ2oL/cjWuDSH5chXBr1TYcPW8iZCXm3sS2Wyn2DXksv586WKA9JBrSEVLM74vsXCrXrtDV7b
Y81sIMORt6iV6U6VyeyZfQag20TvFvM/ALVfFmdXEWAoq+kDCQKC86E0hQ5iHIPbVpYLuZvYw3BS
nPlXCG16M+O7+tJ/SXNnFUQFqlcBijx9MYA7714GzUOXlv3yTPLDjvkI/RXFMD2U/gYd291b4/m5
zW9V/LArObWqxW0ZJfFUzG1WWRlKoi0owJraymvw0v3u2S/7d2mTauUaHUIgjbxnx03SNRKS684x
G9dGKsK0Kc/9Z5BJKa8mZ9R18r0knfG5Y05cQQIn0vAOcWDmltSJHzq19OG/fe/JYAaabtEsVPMu
KuuPDOGiYoshX0k08mE7wOibAmO10anDIDe0iz8fR5elXWaYBVz1bG2GihU3ihUo+K0pqAjT9iGf
hp5VOX59rkU5iKpBuGiDBH7EojaHxuUVzMiphqEKTBu1oaJMjg8nH6aIWm2Id1cQb/RWVGyWQ9t0
b7aWjuSWMmtRg/xIU95h97xn6qxVGT/bIAhaJr4kDgdyCkY6fhkBB9gYCky3jET2TQLy/M05vMIQ
Wwj2nEy9p0WVXaJsDxXt7WY5gBqzo2v+jkvPAkdvRDAt1TjAlGDIff53wu2O7hCilCRs+I8j4n7w
0gF1geUpyi4x7hdlcyTo+lTFQGjg3rETbkoe4bZycBpoyYga7wR8XscxAo6v6S6D66HpEG8TVbCx
TrS3uHFz/M/O/sMIkdJVUaOkyA0t1WcRgW6kBfDiLRjLYKoA32EvT0ULhCPAqRUQlEgqPKm873jU
fMAwOu2uMJ3MhIVl4VqB5HjcmHd8X3dV/ehd+T2QxB1pjqo7c/6LTF1AdnNMcmqjgroAaT3C7DIG
pRYlFAb3VLgjfncJrCngM0sWCYG/fhfGnYfW7ueCGrElR2uzGHz/kOZSXQQWZNyf29yfEtaIipVf
eZF9CZT54WElMOEf7wRHzbRdwUZj5JUy1nIpLzxBiIGGHhi4WT9EzfxrDD+U0TOPfy2tjFSDcbCy
sVF8A32qsTb1GN5YFX5wCMZrwbBVrbmXYLs3rs+oJghn4zMDTrgbflOX5t5Z3nIgzbPu5bZQzZF3
BK6/yGTLfdxv6ZCuJsdgG7HZ7Vma+m8EWQ/3TYWcVjYbRPMGfkRv/O2Kx32GcFUWSBRhqfc2a+Fp
6s1sRkBveNswUndWpxvZAz6qMsai5cEbmdBASZ2fiLrjVDVDFayuchQWENS8k8b4ScPO8uNq+ewA
K3nwcpu+dWNXuFk6Eib3eyNmir3d0CQq0468zWzUYGNE2ZXEmm1IVZLo8t5Ew7PGQ8YvKAVuESmg
763srluMy1FZkNzZL3oUTT1uTikp62fdn4uaAqWHU0ruKOOjvLlEWUyMesSPAQQknfbG1weGcU8V
ho6tvMLrtOIznsktcDbXo9PvGm5oTZIoTtk/hbce2+bk9jttJ+A7oyNjXgeLPdbJkJsrv7aeewl+
c9rq/E8SZWbOpm+mFT7/R3BZ46ZHO6jKVVqW5N6MgCZWb0ynhUEDnZLU9JVEq2PGfBCXgbyV/GWM
58rCkCnFznAc/F0lVN85aIwh8kWK3clcJb/muMJaHGAynmmysi0kojMRQtldpYfYD5qElCsf7yUh
KWP7LQ5hZV/85BCCtaoXBrcejQ5BzhnWc5nsNEwK3X4movUeaE/h5aEqEJcpiAm7J9hA86DXJNmq
LPDRr8RH+G7YNtVhd7G55LdYD5NrmhK3BsMuQu2AIJ2cWUCjTQlJY0adNLvB1S4Ba1S+tBgErWrO
6cyEq7YxzxfzFBGQnprvkRSNtHRU4tHbntBLd0kxSKgTj8zQWh1rPdVDbVL/zNvLZ98Sz2JK02zz
bfMErgLtw1NLJ3RbaGgB7IPHQryunD3HHD+YC2kA2e9+ax9Gtpylb+QU+5/GoBJ9/y1ZEQhJSM7d
yTPot54FJxcsDDkIARIuxyYFXJYW8FMaByGIOG+i4p52f7rIOVQI7B3nZpPPY7apAQyJWnTLxYhK
hnFAriSRUhJZN9n3wrDS4aZTzPsO9cWYydM+2bvU4GDQDRDMG3XuC4hfj9I0t5LHMJB4+GKg8ANa
L4618pfieBTWhD5UUh4jvTRi8HXWGGKdDGLBvJSqU85JKhU7IB8K6xcGPBHlxZE24FDs+2c4SPYB
K1RiLLxJZOyNvaCDWwzbJRH4s2OlRJzvoPG4C12vaZi8d5YXc4VodoA8a974TztkbEcG+ACmutrF
4nE8WAqj5GEp3Pn+kwDIbzDi/qIjbE9o6iRpPvBsZb8yt1O1DBxcGvRj6gVwXfCLRzctBPxIyOwy
4oem4GcUU12Eq++fHQFXkB90on8tx4mCVx09ocjiVtG/vUBePu1ZY9oMkquSxSWLsJ1RrH6aNZpe
E5BmxH7PpsrCCqdX0dT7KU7okJqgjH8/v+Kqqhb803utF/+yck0Df7fyblWLs5G8EpWwWx3wtDmv
7Ozr0wqPNuInFLSpfVjtw440e25qt3sn1H7SGeddRq4wNAIdSjcpIIWR/nIo94KGq09LioSiOSki
1mHyYAzbYs+Fs9g5LvODJjpoIcJ/PVOKyHphIVqN0AMXsWWHnd2SzFnYteUjLmoE4D3qXSyoYE25
ilsXu3F6Jh77J0+FETX8qHPzCu0IHTJC+phR3Jn8r27AY+zLXC2J8kbAt8RFqcuaAoPRyqfeGCZu
GEmZlw1DEQ3Nj57XUQVFqlsibOpyJkuPRVAUxDZ4o10bj19EMRoGBSIc7JilfEUBdOv5Y8KyAA5G
qV32X79ZIKQXF4R8i5lf3zua1eQpyuIxtOGRSf0bmwSDZ5USiSBtjMC+ggPQsEAqymCn7U90Z9aj
U1va+mxJuaMXtNvQZcBzn/whp6Ww9rE30nW0US5Z1NzibDTaZ/GihblXfVNUKvPTj08xzrL4dPxB
rLboGOfq3jDuVg9J3gTcbtvnUnVrPEWuFyZO11sywsb+8WGHOiht63WuIjzuhBqVAghlwD6oYPtr
qlGVZkHVCBow3TZsFDe2JKuH5EGI/LmzRHkCPZj6h24byTnVrD9qe1dwamfsZHP79wZNu1TU0WzW
tC43Yy/wV5U/NXimK+v+HV46EaSFhqwzvMSY5uZA4xha4o+mhNhQ+OlsPidmtHuvDAk0kKu4rTEe
Kvi9UGHz//gVgOuJPLWh5dFoBRSlfZQ99UnwIFKTPJREqECE99+AB/mDDD9MyqNYK9zRsq+5BY1T
+U8AHoA5GN7oxBwDX8wg7bOA+0dYAOJstBgJL5kvqbNcu4NGw2LpmRRhBomS/GNK3laj06QHwDj5
2SCVmh3j4n26H/9Dn76bgXhI1OxLxIhIQElkswsP1Wx7zeJjuF7KQLehwv9oTwucMgb8DTAIen2A
jNL+O+lP70JA/WazPyfwif3oQq2ZASMJprCeJeDZugOUATS5PJWt/jdA+QpUC+Pk2cQf3X7mqRdM
HpG4DGUgETYbeZqQ5nM0y+7fQdP4NTiaJH3VpRs+er41mRKamLGyVhwmGJaERMmJkQHp89fOS9n0
srxpA5CKqWNUpfsBxqhjp6uRaYQ1Wf3zWCfqzvi7ftQUFWKeqBcl/LrzQivKldW22ET4RdEk+4Ku
WzQY8zBWm6PyEr1mJmfu+E3f/U7FlZuj1PuDh6YsXhLG8MA27mxdyVfEci12Ca1WyvSGKh9GdFc3
ghIijc9sXnObxtxsuIuw42QXgPeoh6I269b3CgrDqo+UpunEk9bFfKXWNT5kD+0NpsVkF3bisK/9
+uusSvsOFzAseuyKQY3bo+rvFcbxD47aNvdgHigMpxHRh/Mc7ytsAzZAbNvuBoCem1chg1RfB65p
EtzPmLwJQfM6QulZVLBd+7vfviYcP+fRywB0ZH2q2mjGoi8DemnuCpIYm+3r2egavmd1IrHkM1Y1
h6nLIbycGRteMC2ZKfka3l22enWojAQS8ezzVYEcVSYInR/aLre5enp1H0jg7KKkeXug9eV/Dr27
inqvl33tixs9bc8YHnG6oLpLgoQgujlmVwtUXwo/T9hnWM/8bs15rdSWhpR3NAR12cqK5caOqovl
fk9WVHQuyo3RP2MM8LkDNGTgH2MGwx+HMlNkE9dL83eP6+FO6oS5F+kIN1J6ohQxe6p1FLcGNqmZ
UcLe8ZxdJb2FyfxdY94gK+RXMzyIsIUB9UCELhVS79f2yP1hT24nCjyR3SoGhhB2KHh/VtfqXnK4
KlcimQDSxhcQDGFsOPG5Zo595Py8EqfcwG+VUgjyLxttn/PrCmWPU80vc30vlAJ3cQTLXdMnHMZP
/aofSI2LkpO3Ei7k0G1vmO5cZLjwTrTfiIvc4UIu8ooy6uXqAlIAImYItMXYQr5e+W5qP+xd2b62
gJlwZdm+fElDAd59BAajLvsLHmWoqeQZ1u4z+cQkmU1TTaAuxFLW7BlS6dfr4TXsZX0sCValV3G5
PJczus5usKDH6pOfnkuCYke8BSnokFIFgoZ1Gy8Yd6344Dz0smeqdO6T/PdYxzblKtXK8o2K/3Ls
9kacP5ApiOcBtcXLtkH8fGUQxuS4t3KjNhFsWNpaIa3MyXuOi40uzu69+DdjA7hROfhR8qXjWZe/
0JKNKqGI34B0lfulsQed2BWdOOZY3bn9N1uf3cZ9L7aLpKVYs/3NPVjF9lbNTT8yj/wNoGmv0Iz+
tNYogJsjSOqqejUHR3I699PdZFr/8dubfT8oDUcqZUxMXZSoCCY39X3AscjAVPUXxq5sId4ebwof
BHh/xhP5m+Cduxaep1liXGFrXFnl5cZ2f/47W26nYa2rtBfGuLsOvmZi39VS0ngI229iTN6maCMO
zhNTWG0kvIA8b24+dIzmF+I++DS9Bj/ucMF28V0q/vyLYssZHtVAMLO799Pp3F+eFjO3RoZhnXAa
LVIxUiXW7Lkt57NrAC4O47Yiy+sRUbTnFPrpMnG5Y9pQNwLqu4hzec2qgEdGqLTLRrBOXujw14pz
qgIjifWwFxf0Jy5Vf0DE+wdP1AhmfWpFMF3PoimuL8JcWLxw4ecbJvh4pXqZNkBB2NOa8MtEZ/jZ
XhfxmiJXzrTLSvHU2GXlzr+yp49mKe8iytfZeNAaLLStQmOjoO23gFNIgkjRkQ3JXObCv2OYm5JQ
RLvXCCi3tVsQIcu4jmz4YK2e733yjQu5TdXhfAld1eebyTn9D5vxUBw8Vlqw3guDS6PGUx0+fkrx
ZmL5JwYzhPLfR63al/r64XDWhVtdC7lmL6eLCJJobpAOZXpB4DEGybSfqSs2cotomQ64gwPDbw7T
YaJIV4bUy0jawH+BaI4NDTwanzI0q2CsD0iITOGq/4m5aXxSC4Aqj/EZluuU7ZmLfg7MApO3QXeG
FVeK9GM3FzZkqw/qkyk8yRqaHn21Z4a2zQ+N0i9ka0CXg0MA/XD+tb3bFOd3/QRQIsWl/5kVkzrZ
DWREa5IZjIp/LcvE8uPv3ePs+hTORo/bVDB73Oi/EOPN+RncVjG4TTHSK9uFby+RTqlDai3Gybi5
YEm55NIUtB0XIJ069DfhGywYe7mtMrk0ajZ8C3FZmOVQGtuC424O+psUYkCLgoR537DeHQA7wr6q
REt8jpnyOmZMIYWDUQnHQqU4VXEvnXj0NabTwjfQX9Rwqw3FpWlPVVq3l/aHOa66vjM8UC5BwlNe
gTi2h9Tp7PazTjK9L7yZn9EMBr3GSu7BxAnGHZ31EI1mO4JKJyNo8zVaWeTyym3ljUMxHGTLXD9M
HkOC3H3bm/8z5wsg4C3+6otAVS7BVq/eFjqIFjWtOqGaTIvkji5AhO/juYdwCuM/sziCpvbYB+O4
iO8k8EH2RzLoeW4ea2+FmTlQJ5su1Kbv51Lk0vANi7r81Ei7nG1uhld/SizZ814v0sQ/NqJr3Nez
dWT2pIc1Z+katkB+p5ZHXvjLaCf2EeAyVE54d18h09P0TW8b3efZSrsxduVhI7Luaztu3a4bJijR
1uqQZyO3yN7JWNVGjVRVp49oqWxJMO119+kSy3E6svKWp2BzQTXw8J9yo3FUCmiVuopA591eKU06
gOKHSl0llQ+DCarPq30gYatvGHmI1DCaoR/rOq8YtW2D228EsqvSurT1wHU50+QaDPfRsRvi6RMA
Ptwn3fQPu0qQpSKFaHlac7V39xA16x3nko/IMwPn0Az1BdT0Rb9OWc4AcOTmC9zq+f8Uf5lraHG7
jipYpKFEe6BK7dcwNWS+lqJncG+WbgIiXmKqjurg9wN2tn4NPnqbsNrVJ3yLCD6/2px49KDLYwgL
/RwuVVhYHGm72Q5XxdYSyAVMyywoEEf0ZGSgzEQuIswVJdoLzEv5w/TPy5a6gNzuYQRNrAqpVT9A
l7knQ+/xCUu3/5ENCaW0liCeR0V8WesZXw7P7C67Ko8SN/CnZwT4HNKtHXPSbkKxQuR4wHy+LNM9
suaFvPoVTRmyESBKxwqUNvDX/v48DQZMJ+2h77XclK1Ibp5VitIiOE/DqpxOUwsh5OtbYgpa1M9V
5DPAeUQY3iXSZnhcE756xyj5d0NXwqvJVc0Pm19gVLQoHJR5P5UK2CD8qlnRJKvaTSsCpJ2I8D7L
Qzo9whku8URPpqiS6Gi+NjpgUkVy83VKZ5mVFO/Ci9z/4e+29Md/yZbzHyA4/3ao2nejeW0+a3xY
OzzXUVU7hOx1wPUClXVflNm/3TYiZZUWV5ot42AHhfiHk/vm4L0fAgcSQhaBHxlN7FZk9XlyU7N7
FeUZdT/k+m91ElDOTIwVBbsgpD0hR0NWmaW3DG3UQQ2dbis0ujUreZVhv0oxucYxucA7/74tHvBS
x1JS7dS6An7JRPlHTxSIHr0UHaodgVC6N/9Prw4dcPRZ/JvxtjFGryLnqutXeIEMguzeflgUERMY
SWnmt4HlX/imMYZ5Qd0V7vnCSbsVt5FRbmo8V/eUrQmVSl7v/HDC/hpuCbVLOmrO74Kp5antxQun
zke1Q8xds82eFy9Syqef/gRFb53JeEhATrN+2crFWoWOcmGaZxUMP7pT4G+V/e8h6BZbK1c4UDgR
y4CfIK+OyywSFFLsDTrhW1p7OMXjWm3+A0PRiF5LNr1ebyyrB36X4ml/VA06X/VD0XcnCh/acnyk
z9H1PKkz+Nqav8vkaMIR0gxJI9BVXbADMmp5/9mlNJt9804C+QUGEoMxIFp3zOdqUMRO8u2r27NM
IePxlSHULot6IuWabsWF0nxMfvCGYZICWLBfm2S/mf/9DHMueebp0dZbLsLS4SpX8FX3HPm25dhf
Mx0jvapoTS4MHpxhgHACZfEquj8b6oynOEl/1Hw+Uuvs0Ck89RNG6Q15zxEQNaBP1QxmDyqbj3gQ
8KfexMrInVNWiOGb42JaqY2zJZss6UWsQnH4Yio9MPPCN+KCFuK8Pyux+Bs/3VO4JFPbl7nWEr7p
G4ba6IHNE9XNveXVVXw2nENOt3Xl2xdxPVrSb+/PBxdDzpSfaZTtox3XXycSvyjoz3xfsqXYyMDW
vfvoD1Hfa9t4XUf6tjh0WQrB78scWpbp8lMeG1qyYEkjT/CMJbnxQwapKl2hqn4n9hCl+ws0jpfE
GvNDGtbAE0pEsX5K4rjsSD9SJb1IDhPdQK1dnjScxC64xz+1lxrGCjhkOhnUj47iLx7/Cc8N3NUk
nK7/YjYoclKv0IBG00kVCDMoBsJz7u91p81h/YSUmDd1Q8gTIYN7xtSILIK1Z/7j64VPjiVCimqK
pJx8qBdP+kXEPt2PaobyhkAF+WZMdP0dfM5ZBjsf1PWjd99CCN0K8ojTPvK8741yY2CRreNz4iiY
bJidRCYzXgCuogbUS3yz9RtBbqiKQYVWw+bTEST6/Z/doEXJkGJrihhXvg2RMmT65OdgCLvFXPgH
o3tu58Qkf/QXaGZhcQzPGileWVCNsXnf5yqeUewjGqhZ9MnLovvTqql1kjq8krD1u7TZ81pQDR6X
84eH4mZlny7Ih5OsaV8GKSRkAduwRm+xHbrzCNEg1zgfyE4OARLX2txDOdldBn/xhtW9Kbv089yE
S6Cc+3gYG1POigWWMWH574jr+h4Bu1rqZ/gK//GBbdIEWxV73TMHWi+N5NyADaXbjKy9yCXZ5PZ6
9Xe6ROM8FbjbRcOiFGFEc+w/SBK965REEo+swG2N7vwNqsRmt51FajuIxNkkZI1bfbWEITM/uMSP
urBCOZucXzMaDdILpJxYCjubdFU14AmuGNr+7WourbD+4RQ7UhfvWMM1aOcbfGP1ke12iZFBIgil
gaJAFB6dO2nLSDMt7VxOKzN8Ez+Hy6K7eH1ECqIErgBhKL0/XsbzXbW+DRiT8CDV7FlgWy+8Z0Xk
/1D5B35SPCd4wWo2Iww287NVW2p7fXN4IytBfgM3rdpc6qMO35zCkncDgW2k0HHjmmYSPo17Gasy
+vNhieKpaUk4H61HjRfRBady6vMWweUMDxxbSfhr9IwZsPfY7kjamYbGVk3nGtvLQSM+RX7HlqbH
AylIYMHKktS7kaKmOf1QYCP8Nt15pgKRdSQcqcyTx/gU4CEsH8CygipGwg3Sm5lS/bu2iOGF2/d8
UuerO73ZIyrZDcD1KSyNF8RENzau+pBnV6gtQXaDRUBxowk8jVd3tcCsgQSoqxIk95p26TETH6nl
mhKX6Q66FRIJ7KP7MQOP24iKst1BcCdJP04Gym0apKM8SCTWjO84wxVV0F5yIJquX6wa8uAs/GT+
XLTCGVtXOAnabmrzWETdXoVcPNThtXRuoFvnqxIEj0l3hhGkOupfsoBuMopHcNua2xyNeCdr/UlO
92GPCsciCjcJpxMR2yiWCCV+W5h986tv3l671Bx7P2SP/0s15daRPqZU0hOzoDnSN37a4aiZ84P0
veSX/bwyLUaZXO/1858X5oNnBQfszUZJkRIElY3y7jQqtu3QRwBGGN32feihBxmjSx2f9NCNCSou
1O4UCc3DU8UvGpvPZARvfR3AGGSkGOg/AQlaGFXqgkSt+AQTM1Tv1CG244kNt3ZCmY4wXAaB0YEm
mSogj99ZWZ+3+Vwrn/u2rkrk9zQNKPPX5fKG6+40xtZBFPvmCkdkozAsJNipRtKJeTQLPiPMcszs
o5GNwWZgVTZCwjAxCKobyihSRyE6tCXh05u4vuJG1n983VOUNhB3jI39MfEVtfymd8iwxGIihpew
Zhao+CSqB/KN38KZ7MPuhpi/9A4cMxKt/Kuw9BSnD+Us0slbpS1or9tc12MVIflKs81iVhFfjZzW
ZivJwennjU12wRCarLUQAHuP9WZloO3W0lW8j2g4aaTmZwXnstkncNLFFccPwswqII3VlV9PjBah
8idN+0Rd+eI0XVp0VYVIKRI0+oI1JRWW7hmFcyNVA5ViLNh9v3mNofob1vpp16jt/BYV5T7JQSlc
iPDPm9WS9clU/WhutVDTtP4OrkqAqJHSdv3wjqC4Gli+JNb9nm9nHqGincOUlBP99VfI+1Xmiaem
SYEfqvbmDQrxf78peIykzo3/7Z03wXVgUEyb3ltf/SKHrTcoXuzAsUL5d87MsWzqyacItaLY6VvY
pYnvRzpVxCQe6WkZBORNMQweFrqz8dJzp18gMlT43Bzh57SeAbFusRiUwqptfhJcC3+Dl1mRV3Yp
9rAU7tZdKGOyprPADIc57QBbOSNLMzHcabjg86i14EJNJlqKBQooYETTZXAIvvvVzgSsBcn7peZl
39ocfcw3f31Z/ni1/ZMiMFPU6rBqVoBtC+jms60yvbqNa07mgmB7cGbLYLuzRAFfplOcw3d7dRJg
Fu0cnkHHAHBJIA5U8VljEgKTi03seUNcYiOBSoOBFlmRoldCrULCUDA2zOe+t/5sfRNQz8rEWY55
cE2D/R5M0zfe7G3diQU9arrlNBumgyZfn+v6Aivz2hODu+nTo6POq+iBfSRV5LRGYwHPLH7KorCA
sh3/d1eVJB3Xf6pzgw4wKJrrrfeXA+5Fza0ZlFaPxMhko+2R7KX+U/H5Ssxz3C80ixUQL8CKdzMN
bC7cP9mcfEwniZgtpMgTdikDhoRMEcswD/cFMT5Mqo4G6XGhpJnwiGuaX3qFNoQrjgVFN0zlnti0
h0TdAmyIEdjlSr3sH4Ik8dB2uu/xwLlmZB7uvMCVBACgwcK6mIfhLwvqttZla6sYuh8q6bf8/ArE
53GPYMZRz8y1f9hgOxJbtGP96XMTtFpBZt/7oPC6h2mSSkourN36/tkmZ/LG6iQ6GTOjRZbnkdZ/
xwxuQ5MZCbw2L/VXgAnKk5lAo19sOZrg3HsCp6iNkpmM1ErkVZKAWPetY7C0c9N3JElt1Hxxp/tO
iEe4MPw3K9wtOjO6dN8dlFVJbP+S0l6KT6ysC2katY9xiiC0U9ITjx++SrxqORHOPFmZNvePPhi8
ugTIYQx3w1S45nCcDfK97D93g0vhBNXFpaTgaCRIN7eQwGs+tctXNiyiPbP9+OgYggvr2Il7BVqz
oQm8HkavVEl7Xrox+Zy1nXj3ai2xKDJ33ZbHFsU8X5NHJLT53lFV7rTjNSTZ1bIbIfFfJTJYEF7r
yr6L+Lqlhee+s0lSVB6iLksgR1Ee/q9ffHcsa6zK/9XOBdD4ybPEEyWEd4bYeIOTvtmF1RZRK5Ue
Bp1d+oUv8qolvcve0xlBkKd9s6orJyaQeDG78Xy4imPOzQa1SK7RJmd/O4b2UZLVmMPyG628j1CJ
mOKdZz04/UkPPYXLnPD/KVGAh+Z9syoS8KtG4GgrRBCf/eYiykvVY4WINyJjZr2/jqmqM7f33N6U
gD/K9+iTL3ZTeHhPAYpmMGSNukklRVRoXCumrL5r7EltrciJueso4t9X6M9lfo1hkgro+VFyKTzq
3uhmK+nHjAKCsHQ1bpYeQ1BrivhWiu0dipIqXt6sMDVihDSowXYoqKyD+5i25UOtPhxUh3/Ty4NN
UFc8eRVG1eWTeo6wM0OUT5rKDihop+PVpegNC0DaYQv2Y6xMFN3x0bEp7CwJxSpTb5JhbVEPOWEW
S/9LWqLKdcRYJCk0gXWf1846AiDsZwovwURxTQhJH6SkvD+ORd37HKYUU+fZ2JT0hzTwlAUp/E3F
aPadIKVHSOdCbjtEfgz8kWHoxlDKAx2EFL2U6vBUchK3uiS40X6jyroV4qIiVzdcS/36pFG8lQ50
Czk16sQ1nJKQDm87atm3pmQIiJTO+RkFGLomJY6tJy1xHVktMtmp/pdsQREMLYCN2qfgwqyh5uPy
y06Q9Q30FwcNDr29Lpoyt4zlLmTl5DTQJJgIdkk/D5OrQCPYE8jeQhas9K23lIkFnOlt4gFroLze
6RmS6H8xBgo4PmU5oPwh/UFDoacaNIUl/ikVrb4m5z/tlVUhLQ3VMIOjSBa8smxyLuMCNbn4c8SV
33Ccjjw2M4p+yMolQqwf6xpO8Z9fzJ1USagmWdw+I889LG8BqimPdILfIU+RXCXN2ONixYXEuN3I
mQAKI+QOUr8bgQDMXECfvBeF8sMDnGbruz2Jki6WfD4eyxeWzJe7vmA/H+wVWPsnkeP2NE+A+lyI
Ql76EF48xq03B+OzcpL89Zo89/n4CrTmb7IRX83vk4YGtlVke0DupvjIPXuWHYg2scrdjF7O9uzy
NNAx+mjl9DDj1cycQ0m2lgaZeXcBh3UgfBaSS+WLTvcjU0z9v223ieT0JxMu2oMKxo6xhs+jqVHc
BzrFWY6HCkxsTcFDmD94pr+byyzYrdrOU74Ia151IWcr8/XRxsvYqHKCSB89ltFDaMVSUdUvZOHV
+NNj5sx/zAZlRXl7ZJ5iqubQNS9beqUYrbHYfucki8VI1dBIxDTubY4+6/PGkX/FmPA9yVaiik2D
+Xj4jFqOhAkwZTgXkG+gmskCnMEL4Q11QRwCGxv1/IItWnI65qfAWrCkhLc/wdNoT7an3VgwdHCe
HifqXCWsGxTESDwYgspkVU0kwsGa5xs5npWDNtwJh8fWbVO8RWxx9ko0WpXWOjKeyjGtElIruhau
aNseBk+ZSlJYoyCoHGokrbZ43ZcBpxVdn0J4X6NZ318xfqEx/ex8bdDu/pAfQdVOXEi/gW+pjek6
n/FEDaEBnRTxp1Q2sbWBLZZ6fU2RwFCTl6kgltTKG3WJ13AjscmSPH2Yn+CYFaSynHvtV9ivsBEb
lkCMqmKGZcp6XTpdwbMkirYOHXR55s0dSd/FIFY1WS2Tix/9D9Wr/UYHeQYAt23zlzE9GNQCi6R1
vO+SyzfFT8sXNSrXSr57FAozW/HvNj0LUtWZ74Eassndy9ew3U9lrPHzA0tRBHX/Mx+840TgpPbP
/8p5HyB2p1H8CZ+k7KjvO4a3+WoE1+UBTrBF2gvbh6VWuMFybTI/YVRHsDj0r86kkGRi928ZjBby
3YJdXSgDpYVOmvTD7OcJffiGD/onHuR3S+bn0oawuhWLjPV/WfZdLlTNVB9cTrSB2txxZ71QRejX
lsqcXCh2jY0fzP3lnv27B6n5CNJLl1otplnNkCmVk61yRQgT5FlOzNNsP2+DBNQQ4I02sSyb9pWS
z7AsyUjagd9wCejX+XYCxkMd6JbJdpp3IkyVrdG8tF1hPYxX95Im4/kjPCmc8LQxNhxXDY1j19XP
jBNGdSTEpRb+62rLr+zyfnOkr11GBKQNytr7I3QTXBmMvqvLbIxAJTSji/2AmiWDMtJ7JdKlKdGu
Y0PwL8Rmc7WeQV0f4R9mcSWUvV2SSjM2MV8QfCmgLXgoF7qfiImbUmyyZ8Sb9zQWgreQgZ3etOPG
rc4FOgoci9Zdaah1Oqiu1hjz819/o3isjxPmGRCe9Sb5VOyvtR2bjw/UQvUgP6hwEqlv91Ux3G2J
PToCvZwrAZA42gtlW7iRfC4dCuHYHJAR6nrgL+9dd2e1blbR3fweR0Cm/WFmbRm5q41ESndABEkp
szie4ntjLhNu8TeLoCt1dmPFMyC6V9KazWppXYCd5rUSGOGg65jxio4kq5T0y0OIRCJyP1c8veJ/
RZWV10E8JLNcpCI/Oi3hib0ejWQ3Rq/2shG928roJd+KrwNV+GcUeahiLxQ5NvM3Q4haliaksw3E
z/EMHPYsil76tG59zDjOdFdBezcW8YraYnieb3c75eNIklpwYHZNeK5edjxo1VrV5/GM1Sz87KtY
ZrywbZNIs7VKXlPJd1wIn81NazJ/m6rkUezl7QbL7uxyfgmmnb+w7dOCPDO1OwbFrUCttBPiRhV5
684TPu3Edlo9dE1xgB6PKvRYqIQCdsV7e26QD5XiA6cRp8br9a8TPiM9PvimIgncWnNIxNMjrbUe
KRFKVTL/v1xfqeXoFHO8WNTpAuyrVuGMPT6Q/9tIdWToo6pkabnImFXzNm6pVNodl6JIEA4u0bzz
w08+U/fMjQJfCzzznHPvjlQh5uFlEDcX2xWHdOW4qg8Squ4HsPJuczeYzJROU1hIAw+9MONu9Zls
wcUDW+Qd74m7UnG73vbwt25ymc8I3bzd3Qqybsl7ARAFbYmq4hqqDXTdEvhyLQYxUI2JSEB1TUSk
qa79/KxVPQIVSCJcCS7LJSzZN98FaSZn4uh41S6YIclLUtWzMtPHf/wr6etpJCDSLn39lrplHFcK
dFBUZtkn7fQATjoedmNzAaNDEwyXCZRK5m0qvOWM+DdHuY3aVmsbg3ZjdZ01HMuKMnJZ3Ba+IUUH
tS6KMb9GiyJPZilq0unr2ta+I+BP1Ez6zMTbag6uY1RQhNZUnM6n9uVUy+KqEmaRTiDCoNfV/N1e
yEw6t8O/Hj+6tlnGEFria2vdebg+iTTHVIIGCwqudbtAt2C7f9pBSm9BV0GlneS5FCKzEbQWAOT3
XxOXag6/fRa8XFdKUJZQM7GHxlxjzWYXcXgt5nJBfHrJJ1sJggD6AHupY9rU7wKEj53cHBn//2dK
rIeP1D20zYeLXLBGhBEpn0z6S0zZtTCF62AM24bhGvT6KVrnvjsPfcf+rgvNu2B8sKvDGE9HOgel
i+daBaAyF+lxTdBJUFzm9JIrKLof4TDkbrFtTuP3XMsxoeunXtWfqMjNFcxicgciZ8bFmTqeCG00
vlmuEsQ/LMjCStVnV4z5iSmtNaFjn1puq7e5k7E1p24ugbmN6MEFOXzN4yPtuAyzD08CvQT1E/uG
djVpp2hlsqnK0qG5NfrswRDh8Pt/k6CabRYyMurEkYnPxnlx4hegm3/C6WdqOHQRl3tvHfaf+X02
+q6lhiFWXBwoUMZB0KpGJ0uvXhYiOyDcG74txTxF5Q7AAQ8q9/fVot1hc7LcxE+hTMn8JYfy4FBi
Uc3kRiN5PTRO79+WNoVkkwdqV29WOGcofNhUSj1fn9eCnWApYaBzs6ArKTIJQWH6d/WWSpyt25O0
sFT0JtkNUsus1isqar/b5BfEbC63CaUfp/0fuSU2i0c7zpaoAr1MvgHaBayUpI5rJvMCG0K4lnJ/
k3fmwNqtz1GGskAsGJ6zJnrFvUjthbAgCj7i9hp6I4rjx+FnQE+/IpRLKi/UW9eQF2hJSsyHJakh
gD5Gd0maM3liq2d9brtA9kdVxeQTwGIW2z2mC+5Elg1anZgqXakFo2aOA/MVnfAuCVKgiZZn43oP
0iBL8UdH/uyFAn1GIc95l6CcmGNFtdEVjWAhtHvQmdWC0S6MYpmMzDEFntkuJH2vdH4tCF6MjeUT
WoJiLijTjhlnm4S5WSA1tIB+EYd1XZUgqkEneVXR71lA5AAKaIg+TQpSlQ4LnKTRA6aXDNbejqgI
VSQK7VJlsgwtKitwcfI/9KBKcuJ1oAT/YPxHUiUt2oCevdmwLB8K7pj98CXf2txxpD1P1Wk1uD2t
+9CPb/PUwGVYKzMtYeIKAQ7+N/QYC9nNnhlwzwDWBoTXAU5jvZXIWx3GGeM8THxIpeiCcn72oTKJ
ptSw7Kyu8YXAkSNuqlJ69iCfBd0lTbjzQlpM0ZNx1OqQ2MlImDGLwAJTyRbsfHBUOU6jD3Nrw6gI
yf1kx0V2Uq1T6Xvw8lduqwZE2ntLkq5yrqpSrakEcfYFix/59apQIDHnDU3FZi/TDYZUTlEb+lji
pTy/oa6a9JMIGJ4GHxO4c+SIdqUYdludxsMRNUtKRlMd42bFTUVfjBKs61luij5S2bv0uiQ0DCNd
8rGSlQRBk5AKsTOzCR/w+vArVNHLYYLji4DlHEz06aXmXzSdD45KspRuz7eZ6N5/cT04b7/Kiawb
evnJRAaK004TunPjG04LGBv1M3tfwsIztoxrztGdR4pB6DrXyJLT5G/DHlzRnUCOrqTVV7RgucRY
0qZYUwwP3DwN3pNfL9C6K6YKmshi/Lxqtj7M125mYXy8Wu3A7c+Ps6D8xY6D5gThzGibFEfuscZw
KiHfeF9DbuCAUCjLRdbdauNYX84lL+oBTETS+nXYEiFFkCxYY/FXlovmlM4bi9we8obeVBX20t0n
3szAOuZozGd8g6JIThsPZwOjvd1+tNj9/qvgGVwSvMuoYn7H+6dJZ+TEPpV8wwiaplZrnwAtfKMK
6nqH/BL4S+eU9ZSC1Y8AX3+GB2hzydDQZd2fVXlJ3h/WEePLRgRuTI9xrnGtp+T9oP3IF0IkDfGD
BXbrQpB72uNc3SWrDb3SnyQ+GLPOl0d9xxw7tEsFutoi0m0DDBEk3zx1Mf52bppWcxnTGsxnfG3L
ycwQ3mg3A3utam9QkEWRfmFpX+v3Wkwqfb48nwxflMBpIuN0stLmm19QeLWcgg5643gQYghN7E4h
ymDyjGSo2CtKtbbaZHTsRS2Jb3cVNmbie52WFYMibraXAZb5NRHnF4OHrTp1iedjuQ5ffLJQRwLe
46GLHRleJdQWKTVRfNuk/w5yWBt2I/jN3mHjKqwORz/YZDgRVtAll0DCialz3Nz5M2py4aJJx/zD
dst2QhF19Lm0PuOCyEwciqj5kivMmv7E+v1DH3ORL+9d8Y9JH8/KIMpJwmGSVKMYBc1ZshmpO2sz
FgkpTnKQ7O5+o2f0VZpR6MJwVCq7tTnrhOOk5Z5xZ9ovTVPvWAxeItSozPl4Rg+M9++pSE8AWGFg
KFbEbXHmvpkYQkkQeunvGt82bINe+6SwV7iPJS4GKETm8+Gq3OevjsuJkqcgNrBTXW+r0zuFyD9y
bcLmMH8B11N2CDYmMb7c23d2Uf3nyOnJXqk2edELvMboPZwPl9+JflieolDy1S1rpASErV3NMAQR
57h4nFmZRnHwYu1msXnSQajbUaooeqZpwO7ePEtKHQnSvBM6OS2MZ1n/wTStyXWY309QndzqsiYT
cTNL9xXsSq1yXw9HJPLKIIdnspdOYbPRt7siCG9DDGldSYzcjkYq4OUiRd+DiE4YPG+JUBeURk8N
r4xnOovSVbscTCy341XnfscSmc9o/ndIqVHF9dU1XbETIRXJZn/hwdx9LXrbKqt8ndkMHGEBvX8o
Q/pfxxSpodlLZwmXDbGnFXD21z9u4rqql76AVMI4wUIuj94SkzGvtYvvda38+EfI8Z1L1EWoruqM
ZRhgtSb6Vpk8GAHrqb9BhxQzPsSB12RAZ7cwoHFBJm5C5d1qW3xuwPR9MTP0Qr00PeGgZI3iY9y/
zTPdnaTcwVitx0oRHnJgGPdKy/s0S2JjkStiv7wqdvrIcUJLOkT9lfZMKEsLp4VSGxaJjMzT0Tbt
SzHZF/4UFIe9+Znvnkqbpyt3fDVZDiS6AiXGkupBBssgwGLbjqogoJy09C/flEMzTMr+kCMJBRnM
IaL4fwyew/zEKrA5IDe9HJ7TCAHL/AlpFjDJ2djnjKcVXGIV2lZvFuxAhgonRc7mD78g77NRphQQ
BRBIAsgzfFD1lehsQplw5jV+x7IOrmKXNABfcidK5GFs+trJSVVPKGHiWBtPo5AD9fzeRQxUhtrA
8YbsPwMb7lEDEQTy9VxVD6dvi21efVLRtoLUzlRHY8xjlP/KyTHrDrdath8Rpmm/x3pQrKku+Ng3
pyiW0u85FW5fNkIpTRcCEo8iKromLYunHmBf73/wL/SdDqCe5/nthFdgS855FIM0O5dkimj/nH0V
0tJ2hwvk3C0uQQK7C7F99fnNCxR/Nm1H21+0u4matjD/+tnyPOHIPKh+VD2ERudflmSsdmB7vETb
oJuhP1iEALgDyvOAg4ukOPqknWmIkb5B9IjowJWYPKKDMPLQR8IPt1vv4rpo/FJjW+13uCD0y3a9
iQ42kUt2qdTwpKVZodoCbDcI6nUqI0ompLmCvDXFlD8YHuQmyU3ip0We+dDKTZruupVxf7XOT6Au
cADkcvCeD8guH4/t0M0T2wqPbqhNXN0lYrOYug/AQ8Fzp3lWvaTdbo77K9at+LTXYM57QZx/3QVs
fgwu560iN7KrD++vulnmbDKyeeDPYGU6udTaLt0+zr65imi+9gC6kKyQdiLWbjvK2wvhCXVipAHm
/TorsKV73tAZWNDqSMv096pzrZDds5QylE7IW+yyrBp55vhzG/ePlUwdl+vmaf2acQIiT2ynmGrm
5JMA+DxkaQxpzCMT0gkXUrSNDT40Woso1aoGXSK/0Uw2Ase/3TVgpf1MZ/uObb/sK3va8Gn8m2Ro
8ucTL05CX1GzrVXYZHGxB4WOAJgQOh8+VQS6Ulvy+TI042jUF7iDirWFipYVCns+ITH6mh7ioSn3
VrCwGtfZuLaM4A86h+mzGhMI01UJh+9uVFGRDkjVXcsEJ9LqBxyDMEJ6euf3UXHmocIf7ZDcyw2p
7NtEcuGvRnR/ddHcehO7qxq4T4O25EdGAVnoC9CyqY9vM3ygyFEhhOXztxQo6aOhdgoZHypjFgo6
fwPUSj4LYmBJoJIMHXyCY816/zXz4emzsv9rtMV1deGbysDZbYSTXhROxjAEfkys6djjd8fvxyQ0
ryY+iLPkbFmzxe/nm8BqnkS2JfPfHlh2F4mNRKCNC9yRFDYtcTPXHpREQU2kRiVFXiaPnGk2RTPh
0kBQRJfb0XtLNrN3d7zlG8O73Wn33KSV/2lyKSOaL/UFxfGs4YnM4LzQW+tpmrpSi1mrHC9u2qs+
bhxcaX5YEOtRxFOI8QzGwGQlY2UJJzfq7HsdB1xWKGdne7egHvQsTxbv3M3quW5ADKlu/Kitdaw0
2F9DEHz2GLNOclNIWFzU70m7UdiOgsWpKYI2MCW7ljtNAb7/afsS3TIeXiiCDgtBA8ZRRcJCCcEu
QJCVXE2v6c54NRze9+aeNN0Aw3x6MbodkxMHyyvL4O6hQGAXSP4ChTY2yHXC87OGCb5V1GYDmrSH
HmI9bqEihnog9RcsAWDrUi6xCcXVQkL2r2f6WNOgXhyAGW1eflA2kh9hI7I3x4/7HrDK4gQajZZB
9GyCM5yBdKTdgxmkkmN5RiVQeOJfdT/6x5vYlA1A9MHB7EeAjw5e7qrISJiWb488+GGyj0LE7VQV
ESiHH1LS0/WZgZTHPSKs6F+Zem2LKlgzGP5lrmYb0pHc5Ja7RQe5hTLNSYeHUPLmZhETTc/XZ3t5
hZZTVolMPgki2yPaV5hxAvAEeYMMU81vZ/wE3al7f8cO8Rjpafpy1pvzvJbngL4j2hPQ85QvmNMr
CdktT8DRgYADlEjkqLktjVzX90IkkXiKG/FNYvvK2QzG8SuTVOcuTWXfQR1kns/+8vtSbzHJWLnk
1uXHdmQ85bUYmhdpiXUBzVsaGtEP6XKUXRIKBC0umNFPJl4S3YEO5boYl6Kcubs1jCm98/0Ij3Jv
z+Bf9AcZbwqnxGPhSf/Oa9KfYJZ2k9Ra1cjt7OG9Vj1Dw5f8xqZg2zd/+urbo+ULU3rW49Fd4KCw
Z1WnUt8FtJxT1h8NMcg0C3F9p82FJ1mlRDVrPyQ4yNA4rZxkUUoNktJlVxZ5NqWK7y1/2a4bCPod
U7nVFwlWvAdtDMcSqNdwfnRg/k64wXHjcQRet4RSrM456oW83itFyRgY3m19KYMcp4iq44yaKguS
pUH4k+ryzXlFXZlNBN9FdVcaElaAVvMIFksRnO9uOD50myp/UEcYjBDVk/n/hYo38NAeRBIwL/Gs
ku/ni5x6HCS52Qehdp62oSo04McOw0aFa952TFVD4m9HeEQPHEKjvqcG37r4JzCrMgi9Wb4gr5Wg
s+PaX9cHa89CD1kASOipepEAJPYqbefSVCI7VUIpiOZK/7MQiK2DFm5Dq9PTdiIxruf7401fOdy5
ZoY9TflheMH1XicrNgjhK84vcXoPo+54sLAKdJK0U1dIjQafknNlKdb2leABp7qEyOuVn/EX0xVw
GgMddIf4Rf+STGa5ltC2FOEgXpos1hYZLV8K3fg6Nhx9WhZ5eCbMjVPY95cWvl0FHewywrhfsNgL
7pkCOoUXoSj33krXRBzPYGKMAOqfLJeds1jGnqKrWcAn8Qfv1/f3hSBI2wh14f+ZGr4+041rPFcL
1Wh+b1MYfRwNIH+PzLURs6j60SVNWl2fqeexNJijO3sinGBOmxzLpmE5ibwluACZtZLknQ3wj9XH
p71781EY++2Z+IhZtgZUAf9jecd8W0/lJF8hK/1Q7aBrPMwlO+eDa6mLxTmlSpxSTh0g9SmAPO4X
iC3OeeCPMuA5Aw5KSF7LAYgy6iMhE6emANSPNO1cdrHYMvWyOGdWWrFtl26ve8KnPjJnpSkUEbod
GYyxsIhYTub0/qdZp5uUj02l1ph/4y/hA0qxW5YQRovR7Xf+PLGs2BcAr7e8imElkSQt0slLt9oB
3xWUGv1S0KtKMD9M8hvAZ7gezLoeMEUodYu9mt92DGojupRaRRGIiIJMDTOPjUpTE5kWKu6I7rG/
/fvoEv13YW7RA+iSAAf5WzEjfWyCfIvyDzQuCWLBQDUfE6rG2TOn6A2RG1sE0wBP5WhWKXQI1PRL
A0vYi7KShR3JSRPbIO98Otp30EbLxcnQTjS7IFtVKRbfLWq2YSx4JBOc7BnvFi8t+gbKN1Zxy1IF
OWjZhpiQusie0zmD4YeorQhHAYLLvhbBnZAVljvp0W+QuaNQLgfZNYmXuRJCBdrM5BvfUta3JX3P
bw+XJvBWWQ8cF02dOzY6V3uXcaIzE3+/+rQlR8YAyd2dQVAZCRumZsPDdiRBXtB0eJyvi/AOU42l
/OdB+JGMAzaGWcrMLEWGz0I4iYrCts6nUopXcab8nxPZ6d8UOM5SrJG0Jy+O5n0bJY8wO3i+3LU7
JZP1EtjaZrn/382JrOcNwc/F0Vgg1SpBxQey+8QZ8hubPTypmP8EVtUToMk7qu9D2MOKGrkHSpFl
C2VTiISpunBey+L5c2kgWF0EL0/roBKUM/j71UOgiAS8uMfuxa0dn1TmgqYaEwpAlDduUZqc75tE
fHIF2c7uXbcfRvZJ9Zgq4N553mX17RFacyTYzYCvsuvfpMpIgZ8mLaSr1zsTd8F6ew7vbtsEw4v/
M2wUfOhqNwZS5tthq6HxL0WN6W0rXaRTAL2jgXjitaPoTYRVOa3wTUExrZUFCG3IG/GYp2Y7AkG7
xR92Bc+gfGakgS5E9jhATKn9r5rwtT6SN/lYRM/R//ncPadqWXQ5detwBNzf1yYqZR11TbEhVkxy
lknDahJw/nsm3b4i/KBVBrSKe6Acwqeig0My+6+W9Ptq8Y4b9ap98yjCqrTicX1d5WYPwfH6vy7S
CKdsdALg3xOmx9rOO99I/SbunwDOfpywkCQzgacq6suAq2eayg4OF1ued+IGykPzq+6c+Fb4WUOA
Jw//vuRY1LzA/3pAi33GSqkX5ChoewV0Kc/o/kBYDN8tQJtHdkCRNajnZnpYFFLhXJ2GeBu9jFm1
dDkPwZ6nSUkD1rOu/9b4v3ky6iUNuxL+ITIGs3TvkBYb01Oso6OJ7NXkuSy9OvHuCC6KECErVGN9
TFrlSgrxrY4G56+g7bGlox3skrnbvHtXH2KLe2hB8WsN/Hi0n7EShAcXFB2TFY1rFYKCGPsiWppr
5R1M/UiDTz1Cc2qR1WuaRelrurC07LExg8KeHj+A+Kv1qQW1R+jGdtP4CHIKEupM23dRZqPFg8KG
z1tlU6VGDU6C3szApY0Q/w6LdwVPWw7t6RTVA9T1cmfpF2iwm/x/+ZcDflrXaOw+dbaEtbp/OJuO
FnCUmjZgB0vrl2TtROV73MMfh/ucr7+ovPYGvYpf5FFmFp3EY7VvzFnTY+21YnWlzLRBfyq+vpAa
ITG3bC6YiGrgeAwUKWmpbxO1iq3HKFW7sVVPj+EL53sPAB1R3ITaisdOlUZCuBEnt2wTZQFYWfwz
cne5jylxtpc1EU8jW1J88hOWgdobsRG07OBK3ihG5wbmw7H0g/92vxt8L3pHRDjNJbCY+ufuk5D3
6eLxiPWMExCPaHDn+g6yNPalLK8nOM7utSuZzIyg0N4++yHvAfx9HCQ0LQzqIYd5CoTWx4YQ5Kxa
vgAxLJaLrzJMMgrtvqRKHQzopNTpBkYBI6Ftqb0cNodE0bmgMc0GVwd2Akk4BswFBs61yifjd6Id
8zrGp4vMCBm0Gv/qboQ9m/KYarC037FjG9B7FALzzBCmFI1kZEKVgQ8Bmm496yqkW7SlhGZ3XgnK
qT3jUZEqP73PlTDOsM84xOd/iIwaFrDViA+FtbWNhGkfofMkJDVQYQTTc5fjTRVAaZYX0PYLX1qD
mIREFAZV9LFLiniv4LpTShlD7xI01AzWw6epd7W7NQMZROZ6cafxjzlR6bPelGO6WkjVL8vlAAv5
kGPuhksNTNDNW3xHpXwB/oyuTwQ8CmBntczYDtos5uQqcdGaXCJNhfasLdLfnCv3Lk84dqxUtXt9
qcK68WChywtQByY6DFrtUNdsC5Fs0X39m9aiZyRhLPZ58eGYSP1MSsJJGlHtfuZGRDRlm1sYYAoH
Wh4oTOON7s4E4zZekOzKZZqp8iCATGxbqs/3Wsvz0gSiDihSggCwAPFza1Z7kmiQL4FIgnWfWCC7
0Rjy48LfEWPoWR1HnqYXSRwPYIQxKhaHFJkuOf48jbhUroEHvygdQQaLV9FzkJFI5+N3YniTISNH
paW7GIjsSSWFSQWpJhHGxdzvqh6ByR/ciqucvOPAlms7FmpX9aJnHvjezFsIThyGyPJ6jKWXIlrL
S2Wtx8wiRr7c8ytuMURu/FJh1q+tmy2u70tAT5IuG/xGVJnKhNOFBpukizeU1aKhMn/mjxX929EW
MdDvIe0timbIz7bQaDkuNlE5i21YndzcoK1COnGHYADnK5DvL8BN/i2Z36KS27p9RCyoP6D1H3yc
IBbn992dCnKnRGwL86kQvc5dfvr6HJlyrd95d/9JKloC9GLr44g9lauMgJ/Rj2ervg45NYmWHjtt
rE0A1QYhmdrrO1t9PvhKgDtoornbypr32J4W4h1nE3utp4tAbhlGyDZHj4+quqb0WIJc/iygN2Dd
6KT+q1Pp1qgkY0pSu+gg6HCmz9QDf78L20IlmO22aIoEVo3PBId///wh12xHxVlM957ZzhOgbaT3
xNDaKJCtY5lZjzPgMKu1MDlcLeBJJMEQdHYYxn0jtFCxwOyGTvBtcwLs+b7Iv2hrO20jyOU2j1/t
Fd5GHe8gJrd3dwISKV5k3SZYhH6ZQvKwhgu/zCEVOkYb3H6QlJfCxmSaXV7nOrk+R7ICYI0lTU0e
zjPfUSH2iw9aOIzpud5joY5yV4dxApkmROUl1jKUMUXvGx+JPYxXCy2wTm54v51y+9ozbfmh2vKl
1LlWM9RdA2tdHQ4hjW3W61GWzzpsACqKrUievBAeW7WboB3Pbtd/0vf6IpGCGFNKGKvIcMEd0K3Y
V0YNNpgnf2F7/0q3yPUk+XNiW+8aZI8EHLEQQGdB9bUtp2YkKPv2kfovzNgXqwedRn7Aut8xBvba
CCM6KgCA5olZbnv2HA1KoaCiBoTwW4OrFtxVblxr3Pty2FWbQbQ8IKA/397PngoFx/l29OfzCBou
2DDjV6PHfQScyzdjqD0shAMNJM95Iv/VjiOepOqNfXkN/6g6kpqfP4qB37I2gWhI6c2mlztZlt2M
56mxpMCDqgzngNUeoBkCNaQq8Nl1ZQ3Y7rXt/QHXz3xMeJhOV7njmNsZ9HHTWR86sQqqTeF/rRKe
PCmZazh6jBikFCvvxOAXbqq9mkcuoh74HkRG4MCS4uHTeO1Bspo+reyZTvhtPSYAIN/B/QiehaQj
k3umc3M2PPd8Ig/HKbMLy5khT7cGwzSTvaBaIrI3Ir8D8MMvj8dBgXKIQqF7eCuxZ1fvKLEaVumr
bTM6uw9mFt7dAJB+3cpCc61itbfogZ717MLR45Ozlq/du3zi4CR/8Cbbuh8pXo4FR1AFJ5FYdnuA
U4Dm/R2Y8OEuuVdWkdUIKwea7A53njG8xpmKnuNtP/fTCTgqKn1IgnAYkHtGO0K4ikihgBduBuNb
EyiUCVOrheSKgQ7RKTp2+sZePA4beSobFLNnGLYoK8kWyOjeotZmt0z/+QIefUF6I2Qa8WOXclPL
zoKJy7N2ymtsxYMDPpu51VaDDCtD9eBsQqDXJ6H0/H2UQ6QoLWAsDcjU5ZGkpPxAoNiflguuIeZw
l72gT0nNJu5hA65Y5tTC273fuaxGC2+P/ZdKZAsvK+wlf421WZYoT9wZjpkC+5ZqKd4oX57FwTch
yJfbGuhEQsUGfk4jbUNrini3iX6YM1lOJy5OVbC9czCnojp6UKaVBryrn4krpeBBB2uIcPoMMJMz
Fswc9keK/Se9POlnUl9ebrrPJ6P7e/XVYUDTBGc+qw06vhPNhYjTzoSp9sLHjGnFrXIr3f/PAlMt
6srCUAwRxbFk/CY9i0k0zoW5thKLbEbkPWrOAQENt/LkpRzf/mY6waJ4Kt4RpFzA3HwJYamCwsyV
FL9HWFP921bTpYwg8BAJRJFVLt8H1Bq2wGr7s9IKGddglMQGlYY/evZVwnd5ox/4fN6YVOCGtPuK
UhqHQXPH9altkMIHikflSqeouolmQZ/Uh6PNL+SFrQPbK0qsQDcz+lV3gUplPC6OfuuT5QydZxQz
6hTTNRBBVCWkAB/Ss5DxDjDL5DzKJ583YUtU7FTBmGJYBc4EfZOzWV+/YQNcCXWSxmEsXLWlVl5p
X8k0vG3yi6PX9ynhfpjb8QaT+DYcHzjNJCzGOImIGudKof6Thx/jUkL9ns2QwdZQ5xqGdi1t6+76
xRzMMxKXlRrULXmXryOHa2Ia6WIQ1rNH3IgVMRvc5acWkh7s6C9k+m+VgM5H/+m5J/SVymkcVn7I
BlQptw+riqFCrRBt6vKb9qr3ztePi4xxfhEliD34LvOUcNw2bJ9NC43MsG6iJymKiWIxcMzztFDZ
/mbArCzmWbG2HBxsblJazEyzLfBFLAN2O5so67+pgLaG2acXeJJoKmsFe0jk3ftRpI23FHhA31nq
FFkybfxojgDBHkjkBOggnXl1aHezF8N6PTGAT3/KY2QvEHilGbC7kKq9qMyzGVUWB3b5/qHX5X23
wPcJTd7ikb5v0mLzbWPerOi5KIXVzHFapSvOvDmn/qjS3fe6dGyyUV4z92phkDtWVFtrsXZmkvwU
zO3yGIlF9ZmvpQb3NUmSGGHsGthktW2HrCuuMLeS00yU5kEIC6Kh7uNHu5N63vRQeIV32gB+NI+1
XVU9N/kbRT+EIwlgDUO/3tADxyfs4ClDdCwdN1sqYzQM6jtdLt1TsvtFnCGzWyE+GeG6sM3L7VE+
609FLEH0Pj2YJcnB2wACqWs5j/k8v7zTZqCokIpdTM0xrvIBruhLpkKGsH8zBtdUXMTwzPU83w3l
NvR5ZBgKgJQpBIjMObr+tvfRnIpnIYQ9AQWTXgsH/RXVtf1RRChyK3K4LqvD5rlzy9uFKJQMHsVQ
65N9YXpliIsEbS1gCM6sE85VNXVCTY8sYoExYosvXWD9GvB/X8w6D5/D9dzQD1Po4iFh4ZOGwugp
NtRTl6/f9S2cMmC8rGAmhmOb+Z3YEYgxYB5NDgiI+2Lx2KVYdIA0wzRA0/m5oYNmD9HCKaMoys2M
xlQ9Lk06/xhfhFd85bzj7VpXVHSRf8LRuO5gmHVIzZBtXge4itD9bTD0SoFfryjeXpghYqa8tBGF
RnZtt9RnnCSoe26I8bWVtduq3FnX+h5JMA72DiuqNlnb1rGUwxm2Cd5cPm1WgN7tuSuD3fKoq+uv
4+Rd5oKns9pvW9QPq12JM54++GAe739cfx1S1Fr1jZRw+VGYFDI61gtAmPnyxURf8VPhAx+Sref/
nYD/bKjzafNQQAjKZQ3OuNLGk7T9ig1TSg2aeHwWdDpHtxP26EI1Cwd8FSyBh9QK4TW8zQz3RJJu
GGtRPZ0za7rwG3IHNWlEABs9hMrkLuZ0tjpEdgUXBizD5IEnWT1D6eEeOa5A0f5NBv4F8Oo3bV9O
ODoO50EOlDIv21/X28MFG7nj+AS43yhdQVkOkJ0i8sL4QfiGXzeaz+Kdo/rh3018Lf+mivW4joVq
zREk9a7o2smzutMTF8bbZuBe7uKrtWcNYqKYo4M7vWTxKcgPxZA6vsGxDkz9A0cSWWnRMeh9fUsu
MeL3OCBuUa8eVsN9Vu4a8Qh/tt2w1dVyZAOPTRyIozm2Msdgn4gZN5Pfiz45r+khLkOXVVpN/lHq
nLHq+dxVYzDRHRc4JxCbUlaco1cr7N81bm6NBdNIaikvErgeqSR5hm0YhCN/1Hc0hdDqkDm8lud3
yLNK7MgJ38uMEn1xDUOftUsqX8wNiwaTVxa8HbwKBSmzoi6WFpSKyJjdEqy6NACOMWE5Wh1IPJji
GWUI1pAjV7tXlgeZsNoDXY1W1o7nZtKfs3BZvCqGdJWnoK3spM2ld7PU9JdjIP55lp3zcj3JTK9l
8pUjoAhCN8EgmgXPqN7XxFHGfIg9++udejvde3hWPSueFqCMVg/U/ollpUnleGjjJo9kwpGy9Ity
C1vKd3+d+Vqk0AHLWuueU2uZ9IZuZc/D80Tfs3/Uyy8HRdGYKXfXjsOiR17xaXnYPxwJ5XNwczB+
y2QlnDMZXFSGMgu4J/ojBB0A8dW12YJtwNOr1vMI0KKIMANXl9aw1PusKsQlQRRD+ED26fMDrH/9
V/RqGmWifVnG256DBKUupLtZClZ45NBHnqsR30n5SlVDUBbNjyjDNIeX0aAivZb7FfC05vqSnLVZ
DglEaLey/8YiCiUSwi8nYpP6jPLKAi973Up/yMQ4S9i4wJzRzBwIejh8MZYlmUdkJRn2mgKMTJf6
ePQWArtAWoVqqMN5yVU4Jg6bYXs+aD1adb2tQz2JQAHLdOdmO3Slc02ceLdzOzoT37WLg3PAwHt5
94urmjKGTDnn9PZngBf+YPoijOH55v/Eeyws17r2nLz/D24XJxttDyH8aLVHRTfLKLtQBpvLgI5v
l6URfJ8Lf2zy+6mle1cqPY7vjQlX5JO9WrMx7XFtReBy8zUAvjQHg+5h03IiHGhPpBhEHaDWF77/
QZ5FnoYogZy6wo1fpiY8yNucxzdktqsBQDxTCFe5NAN16z2ugPqg6joOlqnwq+JAPHZvNRGDcv9B
f9T7ISIapbpI+19kaTAbQCK4kdFJ2J+DecqFYstnNOjFiRlPt3SxL/kcrrsRbA/qLlIsjfKk9TfU
y3Z+10Lr+Iss8HT6vTqixpQ8kFv7ulVMIhX2Aklm7u2/oGZ0mYQVFLdsBe1scFFn4t2qJInowN71
lfnWEnd1YTuA/v0ozyDmSazaUNEOOMd6R625KhTTGG+jxIqR6jDOVtfYw55BXvNGZaER7J5HkkTe
/o/OjLwEmIIICA141DUCI9/OISSR5EesIJB2FwSQeDleKQvCRxVSi4K1ppo6ng5PUa3JxekSVVto
fC5Vzf3/UzrE6HyR+9cXKWi28RtsSRsX47Z0D3gcNNpXBzW1+FSY4uNr0Pg9yO7o6PhPN0TBfZ1e
slaJios6e5INZfgERK18a2QnyE2ICFftyXzr+dzKlj4dFpCrJ8seokzMuVc5y/uv5zk0KwZ4Sczi
70I1/WeWyoEvF90J4ACf7qhpUNAa7tAZXgGDuVysmEJA/mcAhEhlnYMXHYF+7vSI3hBMcuDyM5rf
eOvlXK29l7fJksQ7dW8HWR5KdopNHKdzub8PNVX9SwGKebBM9tHQJvn3ERHV11Yd3ROx+AlQ9lVK
QITsd3Jlh+YdP4iA+VZ+IRDwbMoeEIcNzS0m1NgXYJkAX7uaWG3u7GU4HgZIA6W62j/Kj1u7rM/2
niJzxQFFbkhaRunXEA/iS9eCJeBKwtrI3V4A9KJKCCMV8mmd32xnhj7HuIb6iroUjdI6MmS69k4X
OZPOAz8AQ+hFgEwQQMOXYog2HiHSG1UF09MXgw9msOx6B7m5zCrXpx4e6pZESGGOkvLEtosp7QqA
Rdp7rU/ZvmdXAyEu6PWn8s3RwK1Qmq/NrOez3ftau4jQTU5Q5Foj2o+tqdi+uGWlpPrulxAMRFJq
UOQfDQwhJivnXX9ck5eAkt/hyVsC0Rv04LncmtkpspZ7ElX1ImFDeqGvpDZm17AXlNVTbdMiWEgM
NE3DZ0/ABRM7AFmHnR0jvbuQaEM5DhezdPKIKVP70/aVVcUP1YmKsGT1O0dKkTWInPfCfaskmHgk
ecCGMWyjG5cDKjVXhAkpnIC2n4xC39y7KCxpaqmpKky/N2O1PrvHLy7SXSylz46sbp3w7SxXuI94
hXUKpA2FtcDOV8qpJXJA2cbwURzfiHfXDyL7zV5mk2XzW1LWajINlEmPRSnNVWezG7Y6PgJPEPmf
e/yRVfiVOKIfuBb6ZGQ1KRNgMLDYviOdf6c2AWfHSBZmlmgusJV/FoYVFwFoCrkuJL9vHm1c/ca9
M8fmkteY/lPACxMRCcM3pINWMO2mRmVrc26k8es61xV30jfffZ9rZe0o/FLINLLLXPvpj+rBse2+
tU8A18n5k8WQXD4impfj3yUoQ2UKmYPTGTmk6NLXxmw/c1bPoPmPDavHT8tcrSmaM6rLOGdAUN1P
SzSQUecOLlXeifmRC7J56GDexjYieba72kmbrl4PkVuifwNljehzjoTcMT/3g8Ob55fLLvz9iuxI
FUs1m37FBCk1RxZA6ZtSuQUidEyUOxpFdO3Prbzub6aXk27UE5QHq04m5sMZLkkEpmgtzmNfuvU4
r7T1YK7qq+8FMYSc8gSKPLRfXeN/ipkKP8VF1PdIOuUMEbwvtdEbfVUKSfSkyX4EsEPdLiv7I/XG
BrrrcGG76PfzYl7bl40EQerZQFtL5UmK3eJGZs4uH7YinHKphu99uTeRFkF20TtL6T39qC+DOFH0
/iEv1GNA2y2DRrOSyUJ2EJsak/FcHgRxFWEBkDUnoZVvGx0+Fn1FpVFGV8HTZ5Evf+o7s/NkgBRk
bRku40bu8rZdM458VqfJlLyekhnQbhj0hDckzJh+jAeN+tbQraTr/QUlMqOG5cq0hYr8prOBN9j3
AqZ5yWNIggujs1o38uJ1vH+RHtmiUEc9S+w5NjNX7+ft2/klrkiKDZS+L4RMo+a7J92I5bpwiPQr
1Pk3+YEUezFWH242SxcHRbSnoergdQmKSVS8xmt0F6s8AIIIG0uWEgW4GgWIvpSWtdUWH+ok9oTg
tiqXPAGpebHa4BgvuXPjui5yXG8Mq8cUW5C963Dw4jeHFvSprJv5GyHz8tFs6xjbUDYMLNXFL+ZW
Ag1WWjIf6grL5fnyOWIXqPJ3rBDnMP3B9EHl/NQPKi0oC3IF2NNL0Ukv6vIjUOwUd4ZJP8sazGSi
YxKEE/Lznte/nk2tZFP4gvFKyemA9bnC8kzOixyfjnZfJPCkEPq2D0UWmRyLyE2gg7YH86Ccglb/
l0eK/o/3Q3hsm5rz6oER/NSLcZUQujWKMn7sEyWLmcO9ZjfoYlvZTrG2YW+2BM/BBn7/KmmIS7fi
fjflhIQWZyqXcQRE1Rt9m1Jkkz9FVWxciIKcPWihmRLQopvCI0Wwmc1HTP9rMhZet7PA/HNsSa5S
1F6OI4x5jpPLDmYUsTCDL3DZgR6sCT6qKuhxkvFLkumlcYnEe6MMo5XsLIqqDBsc/s7WNYG0KKw2
FStvL2qudCLHCh+08z7a+CooAQncLeAmIQLaNWsWgSYyhJhOZtculVGy8OQaYiOnyUo0mUGkWp8/
KD5dYzPSmI0FQvat8eF13bbk5XQVX/A6JrRFLQOp8CdXWXHiEnBX9d7jTXkr62Vwz1faXsNGB/oI
tQmbNU/XXmcGCykadhblt+CzKBdAvOG4zuJXeDQOBm8Dxigh4qfzF6T1xVBJbg9z96evMzOypv+L
gj67YMUfq++VdlX5zubdKAwxhtLzksxujlulQgXHTspA0EzqaRBeMN4v2k64mVkSFp8Wu7Oifm3i
EWDd+0/XxP0GffQVqAYooyORj/B1f9qOYg7WXhq0bZNEvbMNPHO6LusA7Q00ljC6jmQ5Msr7TUK4
CakfLfOKmwMSIuP/EvuhGFvCDUXMcJfXrx3vq2bpmaGT3dml8ZA+HbKfg1A9er03nkQLLofBQNJk
B2lIS1d08EX8+5JQe1vK9jKp59Jt3iW4jNOHoFVm1n/M31qZ9RAXNKTfXFZhYxP+k+6K0V85Fwma
0cnfor6LbkT9bN0H72ObhqG7BqvcRaHgqnnXvN6LKoQa5m6BoFh3Odh/0e80Q8pw+KvO7O/a5bP+
99/tbafE/7AVb3NV91p33Aq3SoLhO3z+/8x5+2e7SioEcE+3chaC3pec5yUGHNcHpXy3OMeQ3omd
NURJcqWQUifEZ3KuCw9e6oX0JxAkuD0ZcEu9Ay8wBV6SGxhxKGpLFzCpbxvQL5G+19NFRI5T/PC/
0cCbnmj/9darByVvh1AhK+CMG+HTsOhGIj7Zgi9iO6o2mYozP3NZievj0Roy//xuQsSmdKCl6RWc
N090NqiALJcvZkY83f7Ibv/h377ygAwdZVWKVj0wNxIzyTLeCShet3gdWr/2axU8G6wiLfg4R8W/
NgGr1/C9WzOcsH9qLNCvV3+/6Mj6qrbUs4iqAuTMnhZaA+QC1aq/WwWlaGsqhqyHcVuKfWdSO9vw
jmp07a7GoYkpC1B4zJlJGeNuYUQAk/9eYLqnOS+45Ax+Zad3pCfp+Dr1KAVi+y7sji7j0cUAkcM8
4t3gkKpI301njmi/LHiGr1JJxe3+4EKAT5YcAZo5MK+W7jTue+g2SvDWTIPLFRSjDVGrGBvepwbX
yVAXyTKfgi6mMjfR6DYUBpVaLg6d9v0Hh8SgylfoYDxrfHansSqYqqSPSTnLw6r1sqhSVam/DVSU
mpiRMxCyWyDY3vLuht8oMeBVCt0T3g8Ku7PulrLoKIJnwX2Ame8G9CpkGY1nVEWcq17XcIhWov4U
sigrQh/lEOyvQl5DHyBvsqW54X/gItUuXHuE6u6oPtPdYRgqBfC2EP+wjWTDm/ACfA7g5ei0LdBc
nm6JIbRZzWSQaiZ1XFvYMTBefC4DHzDyK2w7Sj/5H7H/GgvnRL97Zt23qVGDfXmPFH4LTpo1HCw5
/f/GqthzFz+R4HVyJv6xeZlNLZwqSkly0CW8bmzzz+wkNSTb4UJKxXqKIfR5ncHOXSJpDYXi5itP
bNOSY2mxivew/VUOFBL2eNVnsRALZhCObANqeBpN/496JKqdbMyQ34b4OdRoLMD+1WBLpE7aCFbe
VNbTGxuL3kWljq3N4aCdiMAtfXsiz0RGwaaNCbLoPopLlR0V7G3v49v+/QVaNWEPpuqOCSLLwphr
wQt9tW+7q3yfgY1XxXAOuWOcA4CtYu7I4LeDzRbM7ma7AXk5LzSDrDkFUuqlmGXi5SlqWdunloG9
2LzivdW46tNG+n/Z6xQkC1vd/yowPeFGeMj9QBlDR5VIts+3luZ9Mebl6uzdQg9JSEaKv0twrQ0a
lby2wIrp0mXs0ax7eyJHhHQ/E2uxoMwHwFYVpU1OcziSzD6Mael660/1b/DqCk0OFGq+Le6El2oO
FE+u8MPZQbTqaTgNM1PZke6K47WgR2XdWJr4fvOp8yugWLzTu67x8nmviUrdmTlVIWIUEjc2UNLz
vq25T6rfML+Nb78Ne+TOLfExskf9ImPPECUZ2f9pHB43OprVsKF0Ud73RBNpfWvSIWAMI0YTVXkp
Z0eg8AaeO17TA5NQUArVLAY1sdgPjc5Lq2d6UDhMOCHd8VPjoI8skJjMCMtSte6KAWbjr3c9iAm0
d6qB6+N04okVvRuAinaM1qQB0TkHb72YS/47bJ0CXHobya59Lpukbc1YwqI+oDewxiXyYDJtD/Ul
oOuNLtrQP9GiI/+RUlCgL0vuMiy3umMqemQSz+gVDTbc3oXCXESlrXGXY4BOdVgcZ+QO473XbY5o
3jL7qg2kvh4eaDVLlSYR1FsODJRz8mQgB/u7+UclRCAaPxF0n+rjFs+THgt4DSeLp2p9WIEvYqRL
1pVH9XSWMTT/iYIYCOy6ZPlZfIAeIjTyoO8dXVoqp3bVtPNraen6avyJYgrjhbcA5HuqWN4FP5v+
QB9g1aEMUk9Q+l26CFA3vQRbq5PYNKkoBTl/TH4zZtq+a2a97AlcjgQt/RDpDwjiozmWXWWmBHyF
E4SyIyT7lu9XfTB2Hp8WL6b+Mlzs+pbVJYi51F8YoitHWzXKmjOpteWhVyhfV0+JejN5u9iNuAwT
teaZNwBS4TOnvBIGtmwMOCaOp14itKhEDkVNfczduEtX0RG5gZqnkEp20JrchAiynKmz0+BStRCr
fhN4sSW58Ics2ryQxuxRzpFraIO8YurXAn0eN5fqYvRY7sEXhW99ZByK3JBp//AmARfUZOHJgjiV
MVdbMSAAkZD0JlGr1vt/T6vTRyTfujw/naQTh4GkZHTxrC2YGmmapskJu9bzYG9V8pziOPlkZSTK
jPihlo22Ls/sBZYbRdGjr333v22JFuRDIjiyM683Mc+rZM8/BD1uTwbc0gqkE5oZyyUiMaFH/YOm
ugSPbH4skg4tMNE8io3h71Gwpo8lYco/5XIGFJLSSglqunaA5VY0/rNRlOZsDGDu2FifEdgKq4AT
iWhkCEwqbYeUuRVrvvEJdW22M0iavgCnkBMMhvmXBbwdaUI+o419UXlDsxEDX2Jk6Bc5UA7b7EVS
ca1sN+P3wg3BgY1Dnzp7/ahJ9Q9G/YzluKM9pdwtpsk0mnrxRuJjpLuwQQkV2Xdlnzr1tU9KEtpt
qqm/cbOZIo2LsOrNNhMPE/VeGJszvY4ShUZNyS8WLtxyn9vpbu41n8WJJP52XMacaUU8Bv1ZbCH1
zTp3Q13XdsZYnd4VqgzcQcn8PWOdkwHT2DZO/S6y+eJSFGlcFr6Ejb3+nLaDBhZzgHPxhwyI47Ff
dM2iN0Acm3jqEhSdBByxAKu1tc9NgvtQzx7ycnHckFO0D24EJKUz5EqdoMTyVA38gPw7SnewOXfB
s8KZ+RCFnpS6tyBsHqtVaSnxpGYu8RTgS4cRqiB9SlkieOTIl+AheZL0XXDpEvdtkFvhttoZC0EJ
ZQOZaz+PDJBjztE8Ste4X3qFMQcpZHMbU483+S9Y2NAsPYThjrJMe1EpfFm5lF18lqu0YpYGBUOl
0ENHG060xkuB1JqbKxB+zO+30MWGmJWlQQ1t1kgVudzzZcmDEMryCttrbjGPU8Wpg+A3Hv+lgFHp
kbifnJnNX2oIuN3eyltW1T7GbZLpQ6P/QcpkIof16DpUr/cHKyHGB/uOZaFqj9daDV2CGoNFF+gO
8diocipdNZDeWzyRdsk4Q47uw2N1OFyesdgZtEeq/2Dw42yr1HK2BjmM1qZo1zZzOsZ1VnU0hYz0
4u5jUlmsbvxuzg3cO2wfUf/jTMkFae+KQUXJAnda8atsPImBWg76x+H1PvNXZArUMqVmDDXrMSE1
KqANJqixz4XoyI924jWzyXE3tTW9bbK7f3iWYatems+RkWmo09XpKwl6Dc/rNWC/F/w+8QLM7oy3
o930ZwQ6PjiI74b/0T9h+abmcBmw65QUe4rKrIUSoHQL0jVupVc8f7C9eN/PrKImaKCJVIGyEwZU
M23njfZb8bmnp7pW4V4O02M9J4YH+HjML6ECNwUQ3AXNjFLoyf/SIrDcYYR+tnE5IoheoffPYPRD
xSZk3oqYHSqHjW7Q7FicwpueVyyK8qq8kB/XZtkVSaSPZfM87bwSdcttKIsQQ5cr67B4AbmNBPeQ
HfLhTN2khMxZzx5n/lmqU/y8NP/Hm2F1Di7Wl1nUORsqiT+jPpj4rhCBQKLFNn9V+5IHsdwEQ5Br
uZG1dRWu6wiPgUghAr1KVG36K3PyAD2n494AM91iE/hJeGWGizcIL1ZGC8Lt1MX/6hgJkiIylDet
Ieq4d4KcM8zsbHdtgVOg6S/KFJnv1+3ayj82rtGX4QEShHgkk4ucBhSo1DHXLAhuiCk4gRbHlCzT
m5V9r6BAcQfny704iDL/iFWq1yjDDfVRLYf/lQrbyqUsqoHeFKjyXlSO6+DLrdcuguvQLUIG+m6X
8VCL68pJXxECkw3TmPtnVueIDh5F+lDfc4whuwZyHtseLwnibF0PKRIUnMhQBW2ZrlwWwh47e8UM
ZFetIg806q8c/gqRfU3JFCDmATY0jkxUijtv2wSfrwTJENaAPifl1BLn5lNTFA/xM74mQoLly1dr
CF67fQEfLGV3SKpebVqLH5o1sCDz7PmKKKiqIKj34vAMzH0BsBGlwXdhBVJ4YnhI2gHckCag6iHi
Xxg8YCNlR4tUImyVOYm2LYjAjf0ZTXdGvjriivXwAp/Tm5xzXVY69wg+Ryyrr2amUd6yPVvN0wqW
9c2SQ7KKFRYV2ce0DJd/MsW+bxE0J0Pm/ZryegvRCAfN9fJ1qxeJ+uBMCpajPtvhhPNywwgxPhLp
p/o+fasufD0OonlqeZ+ESFzXFctUsBjvpRk19r/rQ9Z/ww4xHVUCrRBaNFjJGLgGvmiyZ/0WYpQN
qC73Nq+rnZk1TMUfJ6j00Cxw7mm15RyOgWHUwSxSjfN2aCKafKmdqXcH9T6NN4ZiEdfOeEoBSHYA
7vNVVyvgc/3JZV21Jrw/BF7AlA9wTze28TuWKFNQc0W0hGHm5rRoNNT2aPiCPs4Tr3ygIRlI5G9x
Am+hWWAN+8UAsVUu1/XXjKvibyebfmszOr1acGbQSicA3X7pmCDwXEBF2LEOL+Gpg7On0SjEkiuy
AnMivqTSZAirj9wlxHMwuuFq/uEwjO/D1Gp2+/H08zjRSJukK9mivcHUM42itrE6FJx6DL458ps2
KhgPyWAGAPenRteWNC6Ho6MbGguxh+p95v3H0OFj8+kD4ed9KGC6DoTaDjPULzIL8BBX2IiDPT5H
+y96gGOxxPgg66r3M7WashlwchEOHs4C8zBdMQ/cGUXm9hIWesiHmjeLrHtV1icBe3TxEiNpHFoV
LHkThqxUZM2QhMYU/s92HGRbRMKjfdV8AqGgAxDDSfwd8ofNuqdY84DiMoAcb5bv8d1ve/VSOjSJ
WMsEftf5zSitn5Zd1Y+XTp8mE4SzjNR4m+t6hhePILzdHba4zlpUWpcanrCzTmcfjiwaclcMDlN8
EAGZyFngegtrgTO6CO0KEAGBpiN6G5z6sZ9Gnv5PUURBpCiuvQ+iz7r7riGuolBLJzvyHNLgc34X
u/re7VPrak3xCP80+VP6utC8/dFTOarvgAtAnGDT/xOTs7ETIzbwPuz9wyfwW38mIs8dp3I3y2Ad
ZXKWRaKkUJe3R+YrRbp2Q6H0FC3Rn1JGUvZWzWHJG0JOblW0Ygb+piSUHM2ewsfChZmx+2U4qDBE
CalP5z1HM/UOLTF3xTRh9YRce2AoWHnluJge5nYmJncS9VGruk7KKzTKfG3xBIsgIUJw3wKJTNwd
h1Ql67iEtpSQH81Z+yGvc9s2QlYrhPA4jx+pcBCuoRaoqNrFUYIsVGBMusFKKRFiqnQI4cGtDB+g
kjY8qUYMwrL82yIzNPThFDO1wAgKKlHe4r+E/o4xbNA0Y9nSpIzoia16XR20kNt9eTBR2vJqz5pB
T2Qgwt0vtH20U0Djfe8PTZazNB7HDAieLWttpQFDkoQfzbutufi98G94GkNTya/5fC2RoKRvw4ns
P0Wks8Zdj3p4GCwurtJitf92BsWwsWh3BsUdgZtD+qlk4kerWF0LiV3bi/wNi/ddnrbra9++64vK
XFHUoQUO+qti87UjLRb1QGVa2W+2A6/2DGSh5UxNB6ar/H8pXvDA83myzAQNjAAflTSgc8Ypd75n
hAXefW2bQ4i15O/s19EYnmi6nuvd66NybGZKfaQDHjNiKrVmiYqM0/ITujS5gOq8nlYA2C3F4LeY
/c3oa1CeYXOCPAgWE0qspG+gdds6NmKdeFCqArWLlYAUdFE5OUuFN6nO29EyD90d2gIfgEocVgGl
I1abBj69ToCbj+FURwB30uUeemjOvpSeC7lY1gXbEAqSp4BGrUNCtm6hlVSVsr/2BltHkSX8Zc5n
2oHdkQWiuiTTe47Ot0qNV9cLV1LdE5ugUN/X2rv3Z10x5ppF+rwPouc5jgPQCzTKNB1LGnXdEL9u
eymaQ0QLRm4JUhkg2Pkr+Y3N71/9xIxlyxlwDHHsC4ByaTFdaK62ptQi61uPn/QLp5sKgJq63YDZ
/iRLMjJ51Vz9frvkNNuNUwM5fDl7018APCa0kOchD8kWhVuNOb7lZ/0Ji5siJAm6OjXyIsrTng2m
m7FTJdsnV7zDEni0g0DzkykR3F2zbxr+zkW2QkkClKOYHCg80ZRgvmKxILGqEy5yOYNuQ6KCqhSG
ozy2anLt8aY7UWR0yASgJfYRFPoZ8HkjH7qYZdYoP9T6d2zjcAVD/AfmGZqDOZKmnasMJ6ATnJz1
27ip5NelGjIDrT8CvRd5Bwq7N8vM4LHborU0/V3p5cajwT2hllH9jMgo9DWw8JdHHxV6CyDltcTT
4iLRRPK220YzN4E5W7DOx/O7t1qeT1hsRnhYSmcvOT0HT/Dz845qOB9QWKrCuCeVEzlrEt8QOksJ
c1+8miYHw/agCdFuCE9nFoL8tWCggmV7hEQ/jkxqJIyO6IYVtXF9HJaHw7BAHnqG32tAls8bSz6t
LbKcZyUqlHgMdwEzsVZ6h1zpiTwOf/25V9H2i4WUTCkuelxEInqhsAxA8KaQs70eZXbcl+OiB3Yn
CKDM+ZrqymRrNs7X9UwSssPwlsFiQUKtZ3hd9U/nIQUFFcemoh7v2+5PY2cWPuHTWd1qFG0TlZgd
CQ6tRkL2UOSXMyLr2jezjG8oegPFH2MM5thlms7cbXkvb68Pi3miedlCfZ1xMulHbAKk3GmZaP6M
6uMlUMR4Ao2xoA5285qkyklKfGLh59+khqfBUuxhWY2XPMMUMCAeethVqbJ3Cd33PXto6VqsBp8m
xtVVwx+zYjudrMhl11hxRkiel8ZjJMkIgHIT0Qx0vmJMQpYugUUj/ECZ9n9OOW8QE08PiP1RPkBh
WxP9Fm9SacY/iQfo1NpHpAPz2bnjgYnduFWQHXrBxqlaz1uLhxju3ywl40aXJDRCZ+/AvQ3mKQ78
tstVdrBRk9awYCxY79Uae9rLu1dCj3nIP8GN3ilE6Jo9PVfblZpOqZ+5qQftlCk9dfhlvfmdJ5HE
KUTFIutxuaaYaDSA1WMAUz+66tq/d5yWIVZOOBkPIJmoC+jIjrj4QMjuFViKP8gqljqDLz9sPHAy
0iUATwuM7QgAMVSw2g3wJotZv6LWPLORIDPZm0KGFAT8WV/vZ0A8NfUKzynBw5jzNHm5o8eLh0Px
/2rIAijj7NtH4ThLmheEd/AtcqtnIc0/aSL6NLwhLoSVuTDqYANNt0ZDtIZduU9sF5d8dPs8qpEb
r52NYJmBEYgtTnWqwwjREL6KakdE0m+f0p1uWKIrmqEKls/qr5n6m2ylXr9BeFehkP4/5zDPFAuz
9BJ37Z46VY5UwLdT+/IQoNEIJSamhff6/r5+/EPpEUik/M+ErRFrYnhWPLA9QQd8/oDx3+msWsF/
tpL3RiFdWMEH2ufOx99MBfuSIffg4lIZnpDWKS5NPEkagqZTICtvGWrDw41WwwB5vwtUyyoZHHG/
BoZkUQE++PU3jobTGInUJUkIfNhGYLU9h+3PiYX3wQcyzR/xYm5jRJ3azhuQX10/ff1lE0Wb2BkZ
q7M8/0kIVPMCFtXEC9qIw9F/ToK5AXsrsh8qxjg9uC3zBZXi6XESwCfVQW2qfDwdnfdi6DkiRM9E
QBdlxlJfNlhx7yXdfguOltiwGTtgoKVCfck1DyJ+ACDmmnlgCqHgOqCZ2p7o/h8Y9JeWxLELjBPY
hz6ZVS9Ut9dpDb3WXtSOQs/5hGaCet9mGuubtRP1xTYEoYFO+Ul0xcxFyahsgTtJtTH1m4jg6WBh
9rqYcfu4GWWv1zHDjReZmwj/H0U10218TR32uV133IB8oA0Rn2ZTje0ZVB4bzgUbCOTTq5PTfOVU
js2RC210XGy2etwiTcaypeF6lpMEB2sT6yb3MkeCSFx8nH/eZGpIple2R9Wmt1Sb4DBJ6AtoTUZ2
VrkVM2GKO1TwKRp6RIUJzwVLXNb0vqJGQf87NUxxrHkBOjqm2ZWifTUK4B6aCyj0z6UAnCMYyiOV
DWCK+vt/nW78BwKTXNxlvjmZ0KYuOiiuX3qFk4NOI0cvUy8/YaVP6SDEIINd1yakYvwrBfaOzw9z
FFlR7FgaHYUo+Z+EGGhJqp/ZI3oYQSUHvXNTi0VDoRVXrk5wF1Oti478olnsD+8qjH2yHtpGacxH
UcDsciqjLSRfUeQbaFVGnN3nGD4SRI9UrouRJ/DajSE0Vz53s0xvhol3Ju5EoxSg1v39bEsoD/RW
1tUPz26Y2zYHmEhiRgGjiSfDkIC2pC9GFnEZ3/U3fBkPZhHt2iIpTMqBpITxNBmolfRpatICDtG8
+UT+UMHVskxkjjWb1o5wlvFPgAyNHuCkzHQWkoNtpUCU6XWNc4KcWHiebHTDqDF3Q0DNcrG3bhr0
YGokBC7+TMt6wSXCh36gTkcdQI09IHf42mIbiSivOZZMwqBAdOcgqv/R9hof/egeEIlNRbVpeb80
7WqNJVsai43aOZb9C63PixjXoKwGdAF4KuerWsxfbuyQDX6tAZA0cp92TkYj4LOgy31HEVXuuf8+
fZDSfsampx1mQyNq/F3LMeduA+lTtDlpqbbJNGUb+/HIydxr1twFYLtjvzH5dYucE48PPRNt7Bp2
0rzmBDTIJtYFcrU4rkMwQIpOOFkGpQq/p6c3wj155M/oAtvjNLHlc/NtsT0N2JBYOXlHl5QDXsLN
p5hUrVXrZPlSfZ2Da4hvKPkOZFTiIVSf2RTPxIiK+3GQ7PEj1Ah3To0UD37KMFjHw/VxZR7DPH2z
S353ToznToB9UspVDuaCKjA+p0mhWQ76mhmb0oFmWr4VdzQvivAR6RLEIV32WkvWI555+vLev9E8
GFWrh/1EEBt2T1NP1UM1CWMmDY1VXUoFMdWNcvCogVm94jPyfM6gVFHlNtOtPeYZKB122/dUP4Ee
3aQbvm3PpamsBgSalL7e1Vmd0SLsjY/UqwNoDgGzm5cDm0y5+mAYEs5H9nHtdmL4UJlWsUPYnHiq
cx4z6kf3vc50ZaDaEQCflWhTFGMq1kZDbhc9G5tCvaAls3H8nrepvAPcO4Unjk9apXczCqOu2YVx
9ovRxMB+vL0Hq4ewYk3ooYR4wlpeDtG/sRaoW1aIXBH4S/3vuJ1gIMscUbr17M37/s02VyITfntY
+TQHj95RKrTxdw43vEyIaqdIA5/xoYc74wBi17RTZsh9aD02KEolOwkCusrlrXm3D9F0UTapci0d
NV9yVz2T7I6ZkJd4ReXlUF/VVV0NB9B3au9h3uFFR0jK/imTMt/VfeQqRoEu4GScBGxQU6TpiAPf
aOLkF8+f4i9XJDo7tr2biBpTzcOFs25XMSiDShnp1SgGNOe9rfldGlcdGtshRWfS1XtP89J5TwkH
+OX/dpYM35g9TP+1CSMeS+YvwUnWJnAm0aNktvaJFulm2lGfwip2xki7nyaq8rbcTpFeBlCY3ER1
ay0/1/d/XqiIodg7aAYuiRqA+k+ivw3Zfn0l/WT6+y/VOA0Xuv4qsv0RMQrclGg7RrYpNHcEnCUD
7nl4+/GWpQUisQshEE4sGV6LdPuFPdX1zpeJSS6ZJb9Jbz6ygLmMM3wHzuS1KMWSiEOeJS/xTbvT
CjRR2TVbtPCWl3ixaBih6ahenv19sLtQ5CKGlG/83BUYn83SLZ3voFrbqppI0Zi7cp85hey/0pSc
9GhYV4P6KFJ8VD/JwcMTarsaViSq5UgL5MFrFpM87Fc/jq9prh0dVjVjtWjIcsOUxzNTBRw6iWK/
198FU6Lr+P/ZtR5f3efg2usQHufNF9gVRSNhZsJ4rLofUNNrVx1e4ZC+9EomPbnaYg/wmtqY1MQK
CKC2UqQ6ZC3VkJTaHxmLjPqQdgB3J4aIRaRQBhO7kjE8NZVvia2VBxbCBt6H58AP17gdoVndf3JI
+KGdSbkEVTysoqqWEinyWapqacAWl70zZCXihjy5azGacdlyl6/YDI0ns0af6t7skZue1cWUg0Yv
981eVxzv4v/967gc0cOsnGcqY0eO9/5pDR+GtJtoTp/NuurE3NkwpI/9+Fu//EMwubFjJQNhoCu3
qKVMH1Sl/t7naFfuUc2ocqtiRJanyX6Ukueovva3I3UKm1OdCYRXbszZbrkgNCfnTAW+Bp8adXgA
yb3nwaEbWJaCdHsIHL0wFM9aGeTpyGEQBbP/0uIHGnm3/ysBOiA/vNoDMrLtb4SFM6wVzSBYoPrz
dhb/FdneKf56Q/Qg3s9DmGSzQ0nrM/Cgn/vENQpmO46gjGJKn05o2VACOs/Ib+CGU2L6bHdEVFzi
SLrUPCunYQv2KMQTxyPwBH3YITJSH+xmp6YTrIkC4gY//rAw4ebBff/79i78IOPgwMTQeIx1q2iZ
W1EpSL2U2ztALjUI9igY/6aqzDhp0a8UXnpRoOMm3lKh4FlpdELwfAXoFAf5fzo5Vc4rW+oF5URa
ArOoQbhiE37mbtd8GZHeo32xq0PxGX+2LVB/GMhOQx7lSHGzu1+amfeJDwUJOXTzQw8Me2ZQYfQ6
P4X1VZAnUBzuP2caNdaQ32mpgELGH5sD70s8HJ852aRm/rEL0coZ+N5Or14Zw9WgvuYPx3b9PSeX
rdGNWUr9i5JUXVlMYNOKiBrB3mgeC4iO3aoiY4CjAeAGD33QH7WUOQ7F02jSo0oh7sZjdPzdr1cp
i4JTjywpS3zezKmiL0kj0ertHPf02pOh4A/88iHKazVEIQ7Bywo0gENcPz72n8q1C8wdwWyfRRWi
X0HNacXE54vxYCmkWf/hHBQDpVbZdhPOPr3BF4PTinNdyrDV2/4gSmk0vw0KV9y8d+suBjTf0keh
TcnSD3XfFZit9ij9kzlzK5HHfGy3sVhKdZ/qP+pnbLtnL6tPWuyJYuSo6wuX/iOjeDNTPen9CyS+
JUAy5HZ+aWW1EpkqTELzCxVMwVgKBFzGCx21Ak+A1Ma2HYXBAz+VzQ/e/DF0YrOEz+4yOOVMcrrQ
ZrswbTM3CGFkno7CjQIV2V0jjdOk2fvFKfUkj5P5Gd8Jd/JjYQLdK67+OCRfINaCUkAee5vnyDqy
HrMdG/qeG182q6X9H4ne4L5OMCAJV2teusaHqvGnIlyZjwZY3paTjRjz700N0G4BmBZ6W0J/xxjp
SecwFFbNZzOEDnhz2cmNDSPLIUktG1NvxtoEThNlmBMxo+JiVHdGQNBkvNj87XI69a7G9JLLto8O
DoYjaImM1hSIijjBZGe71WAWLElSmuA7wD3yPl+lsRvupbZJPUg3i5FHHZiW8idrn7uOdKNiMq2x
WeaG49Yjdr1xsO2pyQP9cS0RSggqC4g0TfkaB0bqA1G9OroW7kzn+0YWRtnPJN/P5ObgQw8N14N4
z9uwcm6uG9js2iPj8FAVXC89n0gZhQ4hI1FYcl6SmFF8gmhe/pu2MYRtw7eFMPAQfq/QFWzb1QRT
h6xqOjKaIePoYRZdiYZABqFunx1scKPc9XSXNpsCt+YlCsZegsTNIXl2pi1qkuSx3ihsGy7vOe/A
6JiJGjTUyrnaZUuBb8Q5QHDOrA9hgCmY6kTYNZmh9RJsqVLxWU9BodF3wsxMKNnVbWeCZ3Yt5eBw
JHbE5gazxIpNT3qsDY47zUMEVmQWlai0JRI0AdKxWwez87xl72xdoyDTLomArRD9m0GSjh8HA4N4
KjCnD9c5FvihM8/FFtrQ3y1jHK1XjlCUgLXXOMmVc8Jzr1gIZ7IBmCZdM/rZop3Z7kqeE21gLX2J
bO0GRe8C02rKwCUBlDj0wYhtX7Klhfb6MwKjl/1rimgHzsuBIUFsTUBD8bjIphZoEQKfdEL339FI
tNAgCX6sHmfbMj2ZCtx2n0FGfQZrDzq0VKgq9AQ7HLg6tWPOYjL1Xy6RhWFmk6OhCQDUQrG/06dc
31iHAEzIeIZ6PXksoBuAmdksnbfu+PhiP7/j9pW29iHwqTIs64AgIHP6mvafglyWdFQzPeTP2WRy
hkkRAVjd72fBSSXNR0uayYC/IOcjwqZdI3bIpZqc2qEk5B0gAtn8rvDD26TuXA4sgFpHPO0s/3fa
EzUxLqctv9uQEqSMLBIzR5GeI1NlagFXmE86SK7FYpulFICTGLaoM9yS6iFEi+M+tTRYiBEN0EBl
uYpv5SSD5PRyj4NUVv+97rVmztP+mfqFPPQrL4TbYjA05/womnDkDvC+4pf5xEyQn8TYv1NWsdu4
jC7gH5/mPojDjLNKEGwrnI1QnEkIQrSDn2weFIKG/6EUb/SjxPE2dDDDaKElkkfvrLr9wlQ/7RXy
qRg0SBnbKTsiQCqxMFS4MhRRidQekJuAs83MKBwx9Xke18yagcmreVOFRzr4RvQNPq5Kql0BKfwY
73k/euUJ982KrodGgohd4BcyVyuQ2nAXMUEsE3BJpesTOV1KmogW+9zbFhffeDo2hgomkeOzT/Q+
p5tW4NxgJ0+sqYsAJtURcepDI+82yKZRuNE2oeLBvzOsMtPzRTIZx1Vm0u9YnqKEBzpAld/fOsIM
pv73Lg/wv/VxxpoIk8/8wzRyqj5tSGAeJDn/BfB5P1cwRwtplyP0qAQAt0vM9qwEP7J4VjDpObJl
KjdD3QZjNBJAp764YmxRvAwjtXN5Moe3mslwhU1oXTzUD2JBPtKCX3DC4oyjC1FrH8ti2DccAs7M
Q2pST9VyHs+7RTxd4ODiCUodenbWM89N2hFfUZrmKKprWksqnH2IJL/zWyDF9tmHWYTMRmOEegxg
rTtOU7aWJAeKe+je31g06GPRuav368HSAJ/bYXoKAxtbTEtNkN6hbJUnhOLG8t0oltkBJdgT890l
4/PBNbizFeekW5CZhhYldotKfYg5y7Y8xP4yu5n8r05rN0BN34v5yAWkMdApUQrA9kUrSBmdZ09W
5z2rUoGzO4Bjhh975AJvotlzbDD50qhP009E97eqyZ5sSkOVInCK2n1i12JlW1r/WIuR7tO8DUvT
MyOXG45RlDRbPt7IXkvdg6ChYaotGNxy5KOibMzT87Rojk1edYdNZckrlsbbOD9odixzDr7n6arF
9Ad68yEMfDaPtDeANaOhuBNXXgcXHImVEe/x5HkuBTvvsJC7SUooou6qaZ2vBjFqAAaRX2FCIsHF
kryQHkRw1KjRqyTVb6FhbOTs5gffTM2mg89D/VrOPRcC8uPAyQ778y2wrPFP1x83/1IiV8iFMDyo
mxdABya70hnAUTzbDwD3ai8uTNhN/WENw2XqoFMnUmmMUcSzpHIbx2+Jy4TW3yar7ZVXBNo93Z7B
tFN9DWwGDyltiAKC3b4PdTOrhLynzIVgMlJ4n8WoHaqJWkMOdIy95ig2Twk6VayZUHlPzgiljNY4
JJz5IrEDHsBgkO0MEJBqRPmPod4SEq9oX2VgzDAjn+h7LaqWtVQ/9ZnTjd38fc/2Zw4iMOqUUGqU
6wHsqNfcGUDxNj+XufHfIGudqXGtjP9upHsXgxdfN3ZclwYJvZesZZv/OD+IAflGh8h4KFIqNw17
Z2a6UBlnxXd3wPkvQ1WrhL2uiun/fSZD2D+9R3CYGZV3Dy+1iLMJD9OucY1trbduUd7JdyAjpaRx
N6nDqfZsYWYJ98SBnmL7rnhEFJfN3Gt/Q2V5D4quo6Wrms923zKH+4WottLcOcHLm3PTdRTa1c11
6FPpH4YCMl9YFO+hkwDY3CXwkfGR4Z8aUVC6lDcif3taKRHPdiCje5BUT8MuOPjAG/JdkEGWFV9d
2k6v+iQc1ngq7M1xRWm3VzrJ3XwkTCLhxP2eKl6ypl0PzVOXa/Wsze+M5WtPL1nYlJ6qQBDLu/8X
4Oi0Yywu7XF1dq4I1w8HhZ5RlXQyN8SDl6zMg69BrgEZBTXNgPp/R+t3sX4KPaaNtWIq98Sbs+Mj
g1T/cDbveTgpfDOnckmrcuzPK63nJlYn1hrFfYbM/blqQhKygBojZR6NTO+GRuYEBarcWsdma5et
yrKZWZMRRUnhW/K+JVt17nwGYmOf9LMOzcLMn3tTqYpHy+9B3YUK4aEnUkcIcbCyGY5PJZCUR4rR
dguHJqb4z6sAeDL/4ANhQOecdYpWX8woSkRpD58/d6fWiE9ZPnczn9n7/eqHT62d4Y/mPfC+PgJC
/7Xywxf1hZ1hmAPdqvH1eCdUbGcJWjxmiBPRBC36u9Fr5Gbezz9hb5tMLFoeukFrv+TH2Tf8XfY9
7FcOA35kX9GK2yTKL+uPV6K1j1b8vE3Tbp/rbpXpUOQtaLnUlqJ7BXUdm9EWwyVV3MzkEQjQsQN3
OE7XroI5KN3H7uY3HSYKzOCIpUOJhyexKMb/8/qNoSmEH5kXCSIeZBtE8wq7Fml2Z3oCbAUApKTY
2Yps2C2GLcOdo5ItRfaM/D55XReZOEh00xcSv4mW5vYfg0+VUHH+hUTRdcgBtNZk5YvizQytRxTy
hGwKmL327YY8k8ig8yRg8jmGECx5YYFPy93jczBMTPBZGsDWa8XgkX/94NiKi9hLgPSSn4u4AKFD
cMmF6Rhcjsc/BBHVAmuFdnNLJNMilpLVhK67qdy3B1ml6OJrXOvGQLtXTGjSXmYEMb02vXQZFJKY
bQ9rrot7x+KPlhE0Qr5d5WoXfqVenTTjl8i9UkwHkBOWtjGBUoCv7yfeu410Qmtx1LRounIYW7z7
rBkoaIFGWNWw6QoPj7rCiAnH2Zon4LzH+Fwu956I9ZW9kgVmVgVYEJLKMMigzpF2l50LW3rtpkDW
qpGb0h/K74ML7GUW2MPveX+5uT1BW0TNNRiRFB6ikGst42kajP4CQMChfRL686r4vVj2qdwPgWXl
v5o5gD1Wt3jfc8nu1zNKYgjdA2Xx79+ajWjUVU+BlctWhh75EhaascotGoUfCRlmgJCj3/k+nF8R
xVa95VF+P0y/4PpMnhmjeYcdioWyuuprL3turgn1P2ZD+q+V7r96avsvfROgQqIO8dffXFkGKNM7
D8I6wWekS6cWjzUrO7Z6MHN5j0ayF/2jL0Lr/FgdPKcltkhtBpBqGXxQLCcQmOnFfo7x3HnarUtO
0hgMx27myzubG+G4+k0pjgtSk0YU31B4O5B9X52uTZxY4egHHr+Bto4X32D86OksDymRqd/3aeVQ
NiRX7xpoUlgdHG0MMVhjR3JjZvn8dRaRPvm2Z1EpGxrKFn8x28L4xGabv8aFY/OntnWcy+HE+ipN
TOsN/HDby1u0DMc44hV+Pj3K22dqp2CqWCI4YVYUUla6bLfri7IfYn0unbpCgSM2lchsOOHDRRYC
jmjW0OqFPUmg4Vx3lqWNxitonj+cRDKraRVugbnPYNTaEkaGvUuvg/UGVzlpyd22KlACIvgWeBc7
ONEKvDpwGPUfoMWERcsaa5V+2mRyRrDcpuOQcVFwmZ3F29vWfnXB7pQCvBDKct0Q/GxcdtJzq3cg
vSsOqd/gUg1r9B5wHJhbJ4C/xNlxeRPx6L9q1ZV4n8X910GcBBPoui+e09AH+gE5PXbFJy6T8mIH
DRiDdW0AhVOg2Ayd0TIaMsfasKMg/qUMnalrTCkq6m/eLB7GcdbD3S4zYg67xtknQ8TY3v7at5e4
+lJYi8kJVe6VD+LNvQfR7puZ1wW2cvSxCxuLhsKKH8vXmloMvYHWTMKY8I+eWiUPTpZxAKSbYYnw
nyGjEnmLu6guJ/BaquIa8EmkgkCZ7TwCtAkYxEdUBNQwvEs9qivd0b6ytxsWmzMIk32LMwvsklqv
AGuZGCtXMvA0HmsNZPoSYOWpcdTVZaBBWQbZaTK6IB3wb6UrBNyPVUB85DwGwIItQABF9cXAKDXT
5UC7zyUZ+3ujGWbBJ0dKbC+sCPPNOZ99ku28LHdpRaO1O9cFkzxdBlgD3FqhXFtiB5A5ZoudKM4h
9FjB8O+0DwEeZRZUvQnczMp4tIK/vu+VL8Mf1hFskFjwRt9riT7xbekkmlXxJ1Rl7qR320Oxrs4F
2t5u1FlDyAZJ45Wei/B8WkzIePQEigmjUBIUBomw0HvUmM5g/q8fqxPrOfLvtAWwD7CsMuiSGR/I
arCqSO0CB30Ih/4T7FCYhNS1yspUEk6Gaset/A3JxEwiujGM8+0W6L9vbVnjTs/2Ezmy5LuU5YUl
3opuvBpjaUBkiZzRxkDwKJSRWmqlEpdrqzmxN31l1F8Z4Hs/aYmiOeUbKz2fF0BcOZwcP0ScpNX/
COwqebHpPl29ihjIBVKjdt7s0Vdf0UMaFobi/ygQiUm4P6FOclJIhy0YV3wprnbhnKF/bZRUo5TX
mM1edS5MFgYaET+wM1XM++GNorpvU4xYfrRxyHA2fPI/dy4FrUxHdby3OsPMFAlnX9k5rOANToTU
0cVwWhGz13AhLEFqx5LYRGW6ZtFfQyYUg0cEPmfAcK4ZjRlWmTXsv2KyF0D5U3jROsHZbCyvNyiH
gtcFpDG/l5li68qshPmWTzzIKrJgqN/k/SutKsz+WX9zpB6zgOt2/c6kPdm2DhVCaYP3lmRAIENT
V/lUPvLkhUog1VYCSy2Q7mHZarCnH1aqZ8Cmxt6+PBfSe/WPTDG5BiPCSY2QAFbMDzfA/HT9UUec
gJ5XKdx17a/gygpEhjZZ4xDJj2f8amD7ZZPZicgfNdJCASmuXL+RtwjJnIkD7iwM4YRhY97+qy8S
X40JE2/f2+2Af9pk6EtCCgnUiOGQAOP7Ebkz7cuzgPQbKnWrEUfVR7Ie7uUI1dd9WMHxgf749MO1
3sNFGYH7gi6I75VED+inSPQXg4Av0XHD4R+0Wy3L7km3SwbwOGwpNIK2xGhOqAsWTq0LwIyz2qa8
0DIEgGcDrOJj4S9jQKV8vxpHTNgvt3ryYNUMLjzoQs3k0oDjju/pXk5QeIKS5AgM0zWkvz6Vrjnl
EzP4gs21MEooL4vDsu05hLCjCaqG31kHCxaqKPEWVEs72Es81MZOHyDKo3bo+PSTJ/LmSonUtVyn
waK4QkQkwpf2RFlJz9tw81loa0559yugMGFbtmUY4RrVKXL8TZLQi2FVcA6p/EkQKD6GDCrGT7yr
Hn+NKukTnTMp42LKKQH/EiwU4qaL96Iwh3mkRrfuUSwQDMhQ6UEKy9dTYK2eJZt9eJIQdDD8JxrJ
G22m8y5n9CkEdncuR5Tt+RiylCkE2d9lC0rldMZ0JxsI0yz5g+rGOcLBu9xnlPDK1Gf5Sy7jT0eS
hoU9VS01XKE0Skg3Ar5qwmoqFfOfmlBBH3asYUF8HPokd2A1rf4xfEoF6N3bHgQvljdZw64i/z8R
1p4hNDnQ12qJ+bpPN0kmFGuRcxdT76tAbAoLht/lgQsWCNX+9Ab6D3vWD0K8PA/zu1+Y9LH1lofS
yjrrzmYX0N0U8q1ForxM2jxFR0orS0Y76GTftISju+sNbUUzpUrpQ8ILljp9gjQT63qxelYj5B8+
2itJHsqWX1Fu5oIL6aHFOsKquPELBdaf9dMiAnQP5F5wMGo7SDfpJX5TUfii809kFROtMDzk6a0Y
9DqUsqPVjhYEaDLTrV8lXErFnemkyvfZJSl4NB2knAg2GVuQqToHNAoNO5q4jbZ31+nNOHV6Tl6X
GFWMc7TrRWQFodMxMmEJZPh+8xJ+6gvgmiFugcgDOuwSRTJDDlsCU9AhwEb+c7czgzEfptx6JDCS
8rFRoNLvTwzAGgTD0VG5r78ML6ifMUaQoGYDR5vxbR7rZm14wr5SFwBxQcmhBCLuACfawERaJESB
UF86lfeO4cN6ATOEPgKzCy24oqk9m87rOKWhfFZSJhec6srKHRB6TC+N+Un3NQyS8RDFri6bIvwk
u4JLOJuKWwC+/OoJThiUucGPm5lVja9PHAtgwZvAz31BRjQyvRbYE0iTIk32wSbAt9GQFmWOeWT1
09Z8tdXtFnj7q/qnuznkzNxRZrd02WAnrwmUoCnLm2ozPyJ9D4XUQOvpXWD2lAHp8di2irH3KzUV
BDS93W6FGrGBkxTFZvJnuEx+VUH6BXONHZZMsNvOK8YUNp1amTgR6sBkn6UQyGZeu3lT0Acp/Kvi
nioq4CVUds18O6q7lUMmu4U/W09ZZ6GkeeSnYDZ9xYK471xptfjEuB0dsGtsRu7FX+mKDQGpxjqk
9PQ6cYRe0Q4JhvHwiqiOhAkjLMquPGABHiscLUBx8Sz8DR61uozlc1QlB3X9RnYtrrWMy9fMqAce
li2onLNIvW2N5BvouoqfcRpZPP8CG5n9uZNw0VD8r3CKo+yHi55xcUM3dh2tNX4vB4IcJA2MBnEK
EmL50pTXlyywGYMsDJEzf/thnSA3GuULvWqO+OtcUaQ/aMgKjcVNOwXOCQui4p/DlzcxzR71Xviu
Wi8/k4IprhkEuze5K3sfoSik0gJlOy1cVrt+AMAwNo32cVFNC0JN0Eg1TfWCl93q2ir/CdrSGShb
x0puNnqJFLMVqmVYg/HAVD2yLoPVOosYv01sPTGDez570TU2MsBFPWP5l+iPiAhMScBitpgTqIIG
zzl2o4yjr8DkA2XaenltYJIVo2pVrUmk7Nz3d7g0ZzvDwpke6zyYtcbUom1q/OvEWNFipB5QDksl
CkIfHrb4kFcLB2ffHMc8OQYjrISgM26VlNXcRrNKDsFMmeWZ7MtnCwcOHTY5c9LC2bgwLkv2oGst
DjnFtvDFZDzXEsRBZeefNxM3Gi/b7LMkglaJDRi4bimacm579QPBc0bCVZqfVKx2RcWPkZG/BA0n
bwdNeb25VbKch4qLlGHC87wa7MKEXs49dBXiJGTXN72TRubcg3NWabCm+q7yrpR5+6YIL4vDS7O3
mQVhMGhcdHkh5oG8uNK1EU/O8gGP0I3VQK5eiXhfxfV71DKsFt6IQd2bzPG5deHETQiCO2H9qgAX
EhKHjzwgTUE8gaVRKW8m+AXBuqewWv4eXxifumTKUg1lgU9bKUWXSBDzxHqhjVI6kzB3ZrdKbxkz
ok7os/vjgE7QB5qKyGplPKswpdHfKkYia+zei299IrDwakKKrYqO2/9PcQL+xH9mIrM7Fv3AvX6/
bP2niVIlWOb7TD8uz+HGjiNEKVUSLCGlljizaPFvczo+UFpDlzNDD/jxNf1iR9BiJ8nq/8CbH/cr
mvTFXNHjkwDYNNmCWPIIgiBG/g0fAj2Dxv0pmIVlfs6ILQ7P9/aVMMDjCnbG0SuVVYvSWicfa8Ft
bGPRPsrAsjrhZK1ZDWrlx0ETV7q3I4+UsLQGwbdSYTfYrmrmsdOxxTjl8+ZKw6Ct/rNJyJiyI9bZ
6sygm8f0YVK8KenI/RMzcs6H2/5+7ZC0Xsbyoaw7Jm7GipCamymM5D5Lfl0dZlxmaXNXDIEKM5Ry
eRYJR+Jh5tClQTv5oFSMh+oNtFOnKlfnf9Pn8W0BSI3TDuLUhc6rdWU/X+gdNjeEgC850n8OG8Ol
V7R0oVi1Fp4dCrf92oShUBjttyd8/Wja8oBwLMmfPv3QKmgwHL4N8Sc+soOpQMozMJoR+uo5Lta4
r9qWH4t4dgEQSSw+2M9BU/pHAgTHlh9mV8p7CuhiAO2Q4MJQmGTV+wHVrKb6YvrP1BrpZRNHLsJb
vaPT0DMO98mXsaIjHr3O9fLBhN1Am2j4wSURCNQxf5xQJ3//Y6pnSNoQLeAVihRzI+VzOo95iBL7
aXbGbO/nTNUz0+GDDbalEK5K3ArpuE0zvqCIJWt6yT8qYzYmreVOIBbQbHG7HKmtvAgkSIyiXRtA
TuqhH7d4LCkjziwnHoYIeXSDirHPtUg9kIjLzN8b4QqQ+xVQWDML5peD2XGbRywdljT8NlSKroTW
EMIa4qZHYYPDnz2DTqpDEPqqg9L7qfaiKNkoUhkbYviUK8rUPDa1/40rey6qmggm17XVBUPb2A2S
8XXtELzD2V86B9A2DWbksiZR2bfPehRPL1WGGm/kThh2MM1I9adW+g+pW8DwtoFe3A+qeAlMCaIk
cceQqnDwnU3Bp7iO0RMRyU/DoOCFqrudlkhGIPXFAPnwSoa+YTAtDlCxDkFF2V5sC1Uwok2ndLfw
Yl+z9pafINoaXzBgiXLGDnaMyS9UAwTbAKg0HwooLvlP5PU0kX/D/+seIWdsq7WYTtdjIDDwG10T
rbW/VjgFjQNba20vnbyXGsfLHEfmbYqdWcTdtUZcMAZAL0Ce8yJ+HEnJTrGAcvGEDb4kEzuCUIyo
cMLkE7d8eniaNHMKYcASh5rDLinrvP0T/1VbmDeVXG3uZ6/9tHkp/Va8to2jAyOWlXzulquy4cIc
v0zWRG5oXoLCaznq0JW7IdYUURGAtIXJ8frmu2fZ9nfE6WVab4MMd028nhZy9zbpNqnUkzHLhq89
lNVld9HLSnFlaqzrdIPJp2KPDz/f8tGl0e+SR3c8KHB6Q2ATdbMQKb8szikar8d9IfEqHXqNFaHP
7tUHtejSQObBW8B0LwjFkBikpLHPysiw3FFqzxYXmwc6SAXXYd5Hjw734M/tX2+DFpEuWEdb76rH
JKUaMBpF2Lj+CcUbDMrRDrSgMR2r2KcALWbDdx39YGZiSKNb+P+tXPGQ+1lcmL+fcoU4RVlRMBRd
04g2BLdvaJXilgctvyptc7v+3jXpWyi81kw2dhszguFDWui122l0nzxlbhxwBJFEhhh++MkNx4on
Q2Ipx712EafsbfDTSnV++VA9QJ6oNlcnned13Jh8brBtpfUmYO2pwmeSz6I2BRX+THzCTRBwrP4q
XAmkSu2xOJb2Jxz6qoh8j5NwBKB3O13QnToaJ3EXtf0P04GQfMkuVm2qbY7/JHQOsAXao6fQfvW0
ilIdGWfkQmA0UqqjAMRAMo8ZNMOhNWSIhTWDdLBNWLdCI7Df18nK+2NpAN5EQmdKYEei5poQ/fE1
qbWCShoFkBntm5uLDtPy5dnw3iongIOzKVNfLuLZoqR2C5QrIluW+2dxC60eTqQKmr6PSDe3TMWo
xcxGgOs3xnMmAD0cyiA+FPMH+ZpI1Hn8ofF4rJ8fhJmUaOlvp9f88QWDZysdeipU11EY4KFZAk08
j9TIm3D1FwjkxPD4NLElnW3SAa2EOVi9diirHVf6d5FgF40Q7vEj4JUB5OZ0mQVPAfAwWDUl9vVX
yNwSDrWhu+HO0e6SmXChLkqjK4U5XDvih0/JHJt72Qzx5MlPzrF/NdtDUQqPEIUt8PPchQKPOwnw
IxQvlBzRNhGadbgxlT79fNHB0siDN5hmcmm7DxCbt8Dt+8jYPvajLuCPe9vUsEdbBtqJGsQzFdR5
ESO0Tsug74LJNLh5kCTaeLW8DpspVdAlD6+nz5ehtKoykxR6f3VInhyQrODiduIckdThrKFFlsnt
xAyegIwXL63V8YNZjQGEfdUmdMcdbHz05yzz4/6VfnPpVYVUfDAuGbAr/jcWOYWof36nnvnBTSoo
Tlbls91wgKahtaJn/xTAqfZyUvSqCwzaLcQqomeIdcJgqdcOiCpaoNGdoXT6ef+HDn2hIWXQdeQU
UeUK5lBD5RWeF8V/9SKQzKbatHe/nbQD/HNto9kI2CllBvDKKW3tVBSfwKVDVluc+08d1NZyAWYC
zXJas7Ge2NTBrZbsrJESlTRInSGHx4mLL1TvDijGsTu21WgaIXEgXiKzwATp75B+Do8NsHyQvHEd
61fWAraeaUQxaq5KC4mQBG0bKJpnOKfz5F7wsqXEPalrKwgjxRYBpBto49bLIBn9/qBrZ9xH9LL6
FuvvrvzB2xHzpHymZw511mlz3Q51HoL7zR/5zXkmU/EgL8BLn3BMW4GeGcPttPsbiVAWGxVpeS0o
MlzdWWn5DcWhy6cooALymhNluzAbJ+deIk1na8qAQvy8TowPcJrKejibF8VIOc03+iVueJODKiHt
+Epb1rnYGaAwC3K2v5XCHKUOi8dfSGdCRUXIal7cN5OYG+GUK67EInvMmACjOvAis2SIQHN6QMlj
RjvYGCRIjtAMJ0u8U18XSCkeM7r+xB4jXAnzBVQ4yhqvRWGzMecAGQXlkinp6nQeOKEYhyk/2j/7
i+cIa0vR/me7jkStg25I93I2GNJb3R6jXVPLjLlMsDNl/pgbipXTJPkmVC7X9UulqIFNkfZ9HJMN
NPOWUJdgbvhwSHJsAX7UYfGUHnCZ6X9pLTb24vcq3G+vmsV+6YdRBAd8LdURMh1F+zvZ1GF3fWG2
UaZ8rmd0JW875Pestart5ZixuxxAf47yu/hSYfTrMFVOY476J9TmyGSBF4oYOq0FJ/Pj1ep/AFAz
toJ5twssecuZcfQBDMr+3KJPjx1qqmn3jFjFKCF4UHarUMNeDA4ju+bZkumwOE5pqi6xKai5Bq4K
6nqflW34Q0idI428Hb8i6NFJbURdcP6g8REsZvudZzLBgJGDDBv3BMnSNOlvOvWZq7q4jbRZag6/
W5BHM+gT2KD6VDzmaFJRMMAMIpjJQOS+n2kFHhWsNRr0JQ3lKVS/2A3H7kAiuA6HDSr3hIhmUvra
atPV2i027nR6D9FwFhOIcO+27UXFWacgUOe9OJtxXwYxYhIdBQ6TL63RDDSFT/bxDAXpjMDFGb+Z
oW6f8Poy33XnuFv8OUlbBGKT3K5waR4moJjVGeCCEWafNf22n0nCRJ2uPrZUdoq/k9qMkHjnS7hB
LLTAix42GMrCjDojJbCWSGIwLQPrj+IQrt/+Jy9CqYh0rgPeO3o5M0U67xPb1SuwM2GiNMk20C8w
UAs4d6XZh7oM8CyNunBzqrt+jIiKlPEuzkcp2LuTmkDN/LMnW3VbMKRUzh5Eitx58AT/DWfYaSND
ygDxWfm9LNB9XhiFcawpvTaqQ8ca51cdhlD1ZdRuGl4cszFK1DbYm/kqFg3u0gS4PIGAsmYhrTSX
NIhk0cb2M/+/CvXkIOGIcBCSwOBuSheaf1sv6RLBUJKzVLnY/YNflPXpU2On8NS775aacoUzri7I
bG/xIuoxsFB4WoA7KfDrx9CbulPyK2HOvzdM9FS6Yn+hD8xYi9mXefBNptX5Fm6zf88zPWnL717c
Xgk4Bzm6skJGsq0XlVsYfd33uu7zWiqIiJ9QS7IjdFyVftWxCxjNSnOd4U08143eK2awfeD40XBw
Mm1U2vYRcHqHFwuH8lPGhwBwySPot4MeZ8JAIEC/95RXwyD4weoi0rvSXAYofTB8qkoZrShQKfUH
Eovm3zFQLJ5wgBHqKFMT8czDx5UJuGpEZgflNhltdJ6Q+2Np+RmyDuCM9pbCz4+3bjT8jCO4L1v2
O60i2Ov3OaD6nps1ROMeabng35BWmp21uwgbSzNwMoF7BEuLTlWQY/412w2GFYrGxUo0a1GIc6PG
nqhSacl0dH96sCOyrfW+nY3fHklXbAY9aYBFUJv34N4NCHNLZtU/8yAAC2ElenW1dbChgd2N1Uv1
Il0Sh2e6oSZGlDEM5qjf1sE20uzhAcaoYFON7QLHRzy9JX7BHS8AGSmOjc1L0z0FVFvA5jrYntEy
5rpC8zdmEuiRvA/P0TUTDCrc6w6GYmWm4pHYTRhrYBTuV7StK+v+KlgJxTKxp2os7HIFVo1AYbFb
aiHgxVxVwFIvZRZqeFP+zf4XW+KZjN9Q5OeR8WWit3hOk9rZ+vVcV/sMhf1jMtY8yZpFuIvU1j6C
0W02z6juIhRCdEKqv90NYXbmuX/9q00e/WSDSMnRQdJN6N3tynmltuncN2CHIALsJk1GNaksBiv4
9F8CWGlrQ66UOsgizAVC8lT9iOBnTDSL/n36rutpXKVKi93i+ivNE46a9AHkEmCFcYgGVpYduANR
7RRM864IpsHxUr8m6ysqF0SEjzJmtOYAWZXXEJTJgixfNGMBRdpK79IPw3iuYpntZ8NRMSqaFfbv
FKuHYRvkH1SkDmN057iIeOgb8uNsAsnJKleLRszipHl9FC8Q56+2ixGqYYA4uCyz8l/tZrFBXMfl
M3rgdYdOI7tDfx9bdCWOLSFDQWOOayv83zoWdyATbne+6JMk5CvDJ8xdtEanChNXzzWQlBO9hpix
+KLs8don2C74Xnm+oZGSa3YhtOpupF+ypQcXWRYZVrRW8DYLyaF5cqVMYiAwwSmiLxuFQH6zqLrr
BRjFKaSZBo/ylZ2+i37WJ4TLmyFQgt9LDnmLsXO7PFGHdyh/3nQ7roWN+z+6qrVM2xvCA+nIsFj9
8C6BGa3pgmbb0lFUQ5UkaW8WzS6Lb/We4s7FRMCMzByb2adoyAbqiQdlfek91x93SMeXqqCKg9jw
oJg/Aj4d1KbtDLSz4rCA0PxzTeLH05WX8OlhFlMW7fr/gbldJyylUbdxBrn5lnjIvkDMy/ZB6CL2
msaPHk3XS3M1qA/2sEqAM1NJnCr/3rsSgJVvvOmWWDC5PI7Ug6MfpEj4s8ZzzVsG2tqILcPjsbTN
FaZUIFSHFk0JpRYLdt1MR29yj8zmYD3nhJ+RmjWN5WqvWAYH38ryaW4qp02OivH7QZw3o+at4QuE
2t0JA6vsO3hY4P7zzQKAGScFNDy3toBRlwDJ4lEe9SfuWj8xUu1+N60aGyUSAq6+4EVX82Zy6y1O
y3KwrC7oQTg3/eYmFbJkwXHosqEbx8UJHSGU6Za+SaYa5vJQfZVNxkI5iJNHx2fyhYP1NFb6StFT
EHc8pb+Lpl/i/WO6XJ9OIQszrWwjnvpsH+udyFuVE7PlSLmzfjcQDUOECW8Yp0d7HwWf0G/4J5n1
haaXjL/PQ8P70c3xr+wz0xp9eh3Sm5MjLqm6pbC/IKWBsc3Oa18kpvp95FPGRHKvNTu8Xtbqc6qX
5bROlBlJXl41pzO5HKh3/4XSnJhHqdrUgYHfQf4E0kZ8i9nJYr+Iyq9XpbH9WxUsByF2Q9kWTOgR
ZMNQCEzZ8AGO32SgwoZURivzJ3GG1j3VZmGJ6VI8i93UrK6oRCEz9x6N8r20yjQZ9KbenorXpXwi
0nX1O4Yaq6wWymsE8qaDGjS/vP13zsR+OP5mZqqn/2odQ8Y796RNsrh3WW0hB8UmVyAEgB7WWmqi
/IcdNsrerLQijPgNlTkxltU8A+uCWengY/uJ7dagpIQ68q4aTtBkoLBPO03oxyyBb2olUVPmUohz
KjplA15AkPUufJI0E/KKicGl8P8cywGEnI3vOt1SFYU48+8CsqGJUYmGBSj+SwuADXAHU0bKWlLI
OtCs3LoU3csTW65GH5XXpcIf5Q71JGTIK5z+3WAus0evS78xa4fP18Kj6tBMM+QUesbhVZl8pSlN
ugMDe7o0/Z5dQ64fmnSaQpR46hPxYZL9GcTBP+XH7n4sAoJ7MZxs+HIeyZk9mDYx9t0M+PX0yOPm
nJVKoXFjMwY/bnFlbY8nrBxUx13NPCSYarh5w2FVKJeLcXpByIzSzfV+IPVbVKCq6prLEYzAX9Uf
nIKORUbP/unTcR9FZxlC2t5X9/Kh+1XIlkOhxGDSR3FxeDeR83hRsSVU04Z9A5jRZH/XI+SJyfrR
FAaH7fmHpJFAD/JIBne0Vexom8jR1XcLfiNT6MPf2b3DugoKFi+bZEsgOdjq/gd8+Th/X1AycPhe
/A4SeKJ1yWc1DTrYWM5von1yaEU9CXJbOUhN/ogJ24WwEvdw4I7u82IYPlAQctCeZ/XYn+Rgu4Wl
5M9KeFWm35ZwOSDjqArsj9jy2Eiz38WBncX9uvQVAFVAWynq7svhtcBdexzPkcxJ8++6WdECZT5k
dexnvWoAncgIz14TxaCA0rCZYa5vRlOvvWTfpZwEBkb3I4z4MLupCJ6zZwSNpBkVPyKAfKaaNzwu
vhtr5T8QUAX9zhJsRqba71CRspTioXIpDV+oRZV4W5UNyYWcx5JopLI4NlNsC/MvT5q28z/37HTj
8JaZDzJCo+LaYNbLYA0v46eXGCziqlyBLkJ/Bf/VfN2ib28WDUiQvqpPh4jK70A+8y/faiWRmHsc
+ioPa9P495FiMq1p5eWo+m/2qApzEH5cldN5nfi3D0xhaZoz2VGrn7xHbMuvD1RScy44nf1IKQ/E
XwtkfmGRFBmyjnOyvFdUxi6L6dgwFQ1c8/9Sl8uRm79TXQlH9ByILYVwnBfGEB1NkMOdfD1SxAhq
31TuR1vZvuw7e9cP3oFPHuvDzlFkPiTQh1KHH+xiCgXs5C/lWAn9nJbviCjDRXmN74sxT1XSraru
pIvmnTCgV3LxVZGQNNfqGQZqTB1fEdm9jaN1oA1+LTKVxHFV+cd0BdeBFj9xvJNfiH3kyXwctY8z
tYWuQHYbvzeD9MvaRzdBDnxeoxyztnQPMJMS0AtbmoIAEF8Dh2qz3fnFy9A2dO2sYnHS+Mhw43Cm
UEOBZyd5/7HPBklZZvxnlYNKYRp8LstEezUsGGyngNyzGxdkIW+1ucg7zORQbXVW2IcqfXEdh80V
wyysn0dlDSStsWesPzPOEUzxiVC249Tjgea/vzInmuwjKNAsWamJFDRPvDe3+7VeFlz50672wT67
4T87g7k9n68CCsQnMSe+Zq7aq4XrVV4EydSZL76mLdpYlrm31whd9enpGF9pcBCuUyGcOEUjYiLu
5JzdX06SGqAwU7rxI4D3e4C95vVv9T51lhyrBJIPK6pokxo6BPDCLgRzUdsxwdjJW5wN5LyvywOb
rX3R0Hte3CobjjGSTMSLRd3YFgOdR3+ZeSS97dPspNP7h8xBHYFnU2uYgnNniDhSdRDb2aB4gI4m
DgkUh07PAJkJY2U8JQcYhSX/IaKUz5rKPNVNY6B3EnKhJkuryeagUdMZSX4ceAdUnKvjfED83Hn0
CjhILukUDIa+vtGZpc7edPsHeCRGecWU2Ipe65J3SYGtqguqrG69hNFIrnnO5ywLaOdqiHetNMUS
ZUgkyjXSJ+rsFLlmnZEfeZOskT0b2KcNM1wZM8vhUwnu1KAuYy9OFSAj8p6Zq0Pl9alU2e6IRCmg
+UCtdMHIsLxmfDuhNqL16ZEsxew5K9Kfl/OLMY4F9tSTgrQLB/n1a8zMm0Boot9LOJMhM3kf/mTz
Gx+Jdmf7USFWv++jgBaH5ivvYvXk/ewK5NTtaNd5080o/po0zeiJ5H2AQLhcKi9E6JNuiWK6L6qg
sUTqKV5olZqgynM45Q+nIkkriBgt9Caqx6mRnXqsvTNHePyZ9ipkjJ/i3tVJ2gdngBG+kpAoYy3d
1Nn0Nx2Bpq7bnOTVOCSidihtYoVm/2THv/mehionkxQI9rbitGODUdpK5SBYamDWu0YcQUEO3z/+
V8xRwzBJR5o5Jg55FqyXt+WgWl0qLdSPkVDJ04IRqEZMSmbJIEI5qQC1cQDflp55YleKm1KZMknL
9q/Zwas/3MSgGMr3neTmOwAfKHvrluMHgmfFuJiMrdnJYbpul+LbEroCorKs6vV9422CLo7lCSp1
HIG95ms0vqLPH+nDeK1haC8pO1j0SMWeRJ9DnilM6MKYguQvDbi20TV5B4NtcJn0JAQyj7kmvje6
uv4A9mS/6mlDljMQHuiL4QnTboIegQDiL4Fvw2QGGuaxH94XQ0SkWnohLdp1AbQaZVsAn4OQoGSF
/he1YRYwBlZGGrytdFCKKLyjxLLYlY7tM12WAyTDYyvSWs8t04l0lRkXU5EUPs+1b2E1dOW5fkWf
4DsZM6iryCDJHU1aG1G101ZMyxcZtSoY0DAV3609f/et5uwhRS2+7zJXKhu2ucFIZ08xO8goUQwM
ae9YH89bmCy4D2uTXoePaiac1pthqsU/nlc+7umN3fPSmbUfkSjpEdnAe/4dbqF3muzUd1Mi4+xq
Yphk0WFcAjq7cnMrNJkmkFg/DTXDYVlJnRKHLXuOv3LXnlwe1J8/7lLSbJ6Tegw2e+bHCMSHFOCC
QKDY99iKZHOKQe3npjik3NJfRQlU52srmLDuE2FxlgDhbImB6a1aRD8ggmOI1di5aWxvhtYC+mxh
ky0mItT1I5y+UGJ3U1Vn3XJXMkYggMvDTUNaDE/Dwp4YEhOgdHCAwUwIinJEhQ/9DqS0Op/eMaIR
FrWJWtbB1rtQ20E3qwBMa0U5MGt9DBKoxvAZq7yOiulP6dnsvGUzO2GihpNai53N8ifo3FjUla5z
E0/u8VQm5vJlmQcz9hOmQj7ZIcJjh7i6oCZdw94r6BH3OG1s71l3ykU3ZnEAUYAX9telL1OCV4K1
nJrX71eqCu30uyqB/3xVIWKoYIAVL3YIJ7OGUWnS499C1iR9LpLaEaBQ6K14azhuLyJ06sQf+39w
1C1ElFOEg5qYdY6I+NC4cVviLOt4Ssu4NvawD+aHsoFSQuXPgBKe+TQUGtxqJTu8XMCfNOAyApYU
NQrlxK6O4sN+a3fKuxM0wWkICH939BqYqpcxdbRoUDcpAEpoO/LoOQTuVYEj4nlDPtolWJuHKxGC
NiXmvAjIolm2TZbxwWn4C/XrP9KF0TyX+yzCENwUhi3dq24cDyOZXyuvvJ9JucG6/vpbUjyk+JKO
fcobm3hXWj++MJQx44SfIZhjRrJebRsVEqsWs3HFAUaOKqG4w+6bMSbW3xUBHVPqP02VOm5Z6M18
wDWd+bYpWjDUSZkWN24X8TFAHY7yPYqncfWj7ZoNGh7OJTlHVKEF7MJMcZAq1GLugNJEEMYfDIhk
uJPzDAHpC6srgcF7ZYk2+puDDAI+FQOGnuylc024RrasPszn5+cMUv5zdfWQQmn1JGg1nQDmGYXe
bowH7PdZzamNmOJU934eG/aZ2WIVJejPByxHFc90Ju2i+PD2ZJviNCeKimRrv7I1XocEWnDTdlJW
0eCFBKkx+zoSMQKnXQqunYfYXnhB9eFJ7cUN3wkbyXDfIa9li7MFTN8GBxxG2cY7A+miAYMQatK5
NRqemQPmT6+a4u/Mw7IylhzwpgRh0LJVIiba81w+WdjJCoCv4pNn1B/NoN3dY4ADaSlDsPC707MX
Rj7G0NEE0hyd8A0Q0Z0hIMEmc0IMTdLxHykktJ/1pLHLdukFWT8uuLluHb9rdKuNJFKb1mKPW7iv
T/r7RZm0t1Rn+ptwqO3F4MUiv2Lv5WPIDbCRE7Vds4Eo8fsB8WMHmw1/xsR/RhB1mgN5KDxfhsmd
Wg3EN+Q1cM1eemIupDohyQ/qM+fKByagLThLjtVEBgAdgQ/6zT2rQjy0mlLaRPDawmHDsdRpWZFi
UJbYvMUTYRyZXYky57Xi/SKU+CnrLXiprBLhuf8UYAKx9z7sGGzuHpQ4PEYK0fplDH/yooLHLhtX
cexoNphMUBfRcyvulqTQpVDsDdhqEKcYCcZtg+R1A9azIQ4hu4XmOA/b6STD0I+TDEhRSVgrNsS+
DR1i39GGUzdnNZVYN8lA5uowNbE+tOJxkSGP1p8wyogv0nG+Ll0LNMtn+GM4z75e+TqCpTnGzlmJ
fw6O8c/z8YC1eEvR5h9XDd8UhB+VwWnXaw6asTcY2W9dgILZHJNlCRIeGVSRxiV8BRPTVALAVbYT
+MOmGllZzGMZMjvjkiC2Ph8QnR6Qx5pX3tSqDzcHvnszKei2cTRK3Se2siP+52NfMlxlIEwvi11x
y39CyNUlSVBv22xF6za5nZ/ZlPGsuhflYIbALm0Ed9gVkBL2jdu/3+Pwdl7pTLtuOexySFjmIC0u
EzB8PbJ9JCMNlW24OZ4PK4UG6WUi1rOChgaakdl7ZhixNJOXWK7WGhVRg4tP9qOXY0v51irCnTC4
er8R0SdNGD9cQJdfqDurf6KAphaACgpkxUyXuMrQAjSnC8BBh/2FBECjHc/ikWQE17pSAed4cqwY
75i7vBM4Q9mmrCwkUvwzPU//v5WZXat/LYX+/WPoVr2N+GQjpCFL7s2VmxiTSnkBNZZPK6nLsKMu
Rm19e7/cI1QRsIN5G2oTQI2xPQZbUOZdDSJWXNB6ubACHCajMQVQZpyHrr6BwwBxG3w5H3gXKlUc
jYlaXLNLhsXL/JqzDEfhvLMaAUBT33a4mBQO5cNM23KQ3l2qn/NNoYA0mDcHV7A145ilnhUZ6q9E
0HouW7nTXvQt7jgH+pWZomjZFQZHY9qeNgXPU+EJ8ZsscnbYEOmTE7l7ADo9Yeudzld2kydRgvd2
9vFmh4rwIgPOzIuDgf9KvCNCJxPQKR2ypfgsLwjEvVATgcvprzVpvz0dv7QV9kYiP/BhdVFTyhBi
98j+I/nu28YqbQ2t7u4TMu7ahu2dHp8HDDHBNigM8vlTueUnrMrvmIVC9cy6jrbjhZDDy7sGEhoe
wJLfB+3DtuEXmiq+GYGNb0/nfvKVnNIUkbXmB+pcYe07nCKJ7GbGzFbpE/i5zdhbqPKvgiCINsDU
rMDYTVAREjTLrxBGipvcs4dayEW08NB9vQN8vT/CEn76yNk94rNM4aSBOVuLnvK9rWO3/RmDaQJ7
NYPxBw73LLQ1zAe/GP91Fyu6nA2yDDDyCspKU/XASQNOOsV9DhrpeFIqTCrJH8351AkTMKC3BUvq
Quv0OjDZ9+O0f/Olcjx6tkSkZNv+d7edl0x1whHnAwk70DxaJ1JPrJu3Xk5253NY1YPMfsUw+e64
IRGnSgGztPs5r1a6UcGpgCspcLdXkOoaMxMpk0H8UA09QP5ZSwn/OioQNHSY0UlE/bNMBDIiHZrp
emdxccJ3fAnUBBu6LHski+gTc5FXlPkGIRPOl0oKus2LkBveqU5NP6dMxI/TM3j4BoDeH+FWUFRD
TwzGzREyL8rUnbC/OfNKWRcSTZ7YQ+c34/ddkdjFLmx+4NPR6xTWVhG+SKVGLjPjC+5BWORjKyal
ltyrKoRDPhPxBTUGB1boDnahK10kDjafqqm7MVUosWAtJGDfLp9dY06d5s51xneNmOdLyACTT8VJ
MRZXiEZ87vevUWlD7dAiU8wqPB0/bh4y4SJj7FN9gJjfE0y3+ehcvsyjjJZ1rASLbIIOdAYb6cP6
buqUQ9bLdajnfhkxP2FVv1MlInrbbw8Yb8CpV0z/Em1IrwJKok0JBWUIitiyteLGdmY2kWpsRVQV
uc3KldGL1eh9pyg6V62aB1+uFIqqwOsqrLIbJcNjNXRFD+aCm551b5EHHLlvNQ20BDkGElGFFwZ+
1XHyIOp9H/LxaqXmfOMCDvOti1SCkn7StMriLVImAkVa58Kr6ebu12Js4rRkEHjr6PH9h9O3qwta
qWVa1/MBkuBcz/YXqI1D9THM4WBzvhUowSfvhKOlfWoVOHiC3WvQKo4FZ2QDu/JnM2XbhX+inSqn
L5uaUw0uBEqD0u/fDLRFSFBDHLLTm2ptXLGAnHJCzuJuYu5N9Fa8AyEsuuDAnCxX0r2Kl75m/yuS
vfmioy0fF3v51t607GA+xzuq1IwFQkCFMevrsmuQkSBSh5FIaClOKPacJgsZr2XmZ10xpbjhzS29
VNpxfs3aSW6x96DGTXTeqBQGlNMtllpP/6IQBpbt9siWv8KNMhtdUq/nw43Xh+k9EIYa2Nbhb3tw
A1u0nm3upo64ubDwwA5TToZwhUVG+8IBtcFRrvWUnvLZm41cBUdcrZJz0QTAouVZTP59o8d1ym/N
qpF+wkhh2A2poUFnSo/ZmQlVkHNaTd6f6BKywqMlwlI193FXVX7HitjrgSj/wsAMLBgYmfRHkQW6
juzO7e9NqPIT372tQ/FXXUq8z8z4ynzTKMCrXNYgYzaCUsY3Rcr1NiulnzeXIODJH9jK6+9YFFfr
zo46XpDrIfvMq29/rxhFcOgwEQ4xOvR6d0T542t/G2W7vGFNs8AwrpPNqGWi71uRuUPcg0MLr2l5
XDmS8dvsGrczAMmVjQPdN6nd38wGjK1kM/m24/+x/72LHIOeZ6FB12IR/TRPWpSfxmN2qHu4plin
aqPzQqbIxVsYwPxy41sqK5GM4FjGI+xkll1l4DtrDYJFOjqkHwZgKXZdKcnlK1R4xmS4T4Y1FxP4
3hFDsqNNUQpKP/ukMxC3Lc56otrvVaC5tborC1PQqKwsRSU0o/Jik8JppupUPbB+iSMjOU8VJ0M6
Gu5/SWfFZlK7Lk0uDS9LLh3RPaDgKNU5lZsYhQUFYU4S8Ao7Q23lDPN1CYVq1eeDeGUG7S6nz/xQ
r6+gTQ9E6iaswnHOOlZOfaEoOsJXWIlMPsH33kfwjsUyMQ0co4sVkkl9lFNEmJND9d5PXcgpo1BH
6QThEKn0eBbzgKYqYriH++7oolgN8R2WI4/BX+K456/34H5Wdcl7OvKG03KJFgQd3euUYYaGOUl2
Q4FOwuztpEZ08sEZOZd9HkS7RBz7EsZYQc0NlBsoFwncAc+qQz9WY1U3F3gvzGoNTQleivpl1EIj
wIHmpfNDpdOOocKZgf/TFFhUq+VBgj2/1jWQvfhQcKgc+Z7CAoRfOtb/HraLUKWZRJGoyQ+Ej720
38OOpM87Mrx2G8q4NKwG6ZdW22GZT4BUmrPb92aHPCa1cySViZqNdY86j19Vfhr5siCQMuw4VXD5
GqCYRLR2lOfNTbob3LN+zMfuWsYKP/Xiapl1+AHr+FlMePmeFqazB8lDXTMiJ6bt4bc8Zf9CTEMQ
eG9bQPIdhA/n3lfSCpmZd+b7RYWf993H1Ixh0tSfgCTfd+pIrZpef7yhZ8RyRBbqfZ/Q/twNHQYa
nk6Bgt8N5NST8odskzehJWybU5WsOXpMQVMeSUMrH2uzgkSpUNWbKDW8SM+SFwUKC/gV63QYw6tO
yzPcB/CBJJggiELQtIcVEfs3bVLpsfjdjHH1hppgydsSplv2TTfXHUoTheYoqJ8jb6ngQji4f663
lKjaPx8ORPoxOGixE5LXvULBpQro3MV11aAL7Ex9K7J/6zHscPaiCiRiBL1Lrx6DxN38Aqda9MrT
mQVviqh8x0kEuxM7F7NKiiHWC+mqH0A6QyeBAK3OHSkUuKubrj1+8R21RSxRwLIdF8v5HHjsuAec
OiDFq/BMkbhcwkfS+GRzh+x3o2LEKS3eqvPLgMl0c5NGoRHMl7JngEBKglcow1BKfDAsUEDutXZ+
sqVpPHC6frMMv237SDZ2n1UogmZbwSlRbReKwj1pTV9V6UKkXpZ7DLD+PzwIxhG+9SizjaF7OT9R
jHpPF0cLd+YvVKQMTu5yUrajxVl0NOZEci1kYUz42ptDGCO+MnwMNthLBuUR4Nvg1JLWvD1QJL7u
2BQ8MMhTupa8COmLfiSZeebRpeoTS+Iy/fRMLnFewlZGC0HwzYkXey5GaF1xykVXpREgzMOvCkRm
npN3uNd7rl5snm/HWr8/kYM3vnoLW8clEdpgGZmcVLB9mwj3P/kBGlGgkRr1WHgHQWVR/4U8+E37
g7tI3m960qlXRd+jrTAmVIFvUnC/eGA/i3Wf4UjahwFq0C/xoQ+Mapzj61BlddMdEHxd2/zDZAFG
wzhJavHdJnjrfhQBuwJkUGaEUmIS7R2vJEPxz7q34HxxC9MJW0vTvnbKDbay2gFA/ZM86xJE1Wsg
bTyB8J+gCGd0AApzI1E85oh+R5kgHeyYfxLLl/uun1Hrsau7b8CRFjYsnk0L72FDk5fsF+R+FEnT
1vhwgNqippK3PxcaaMlb2bPR19+JpH4qyUi2GHSv0MQb61OpInhYzBpXNqf68kt6wu7TqeYoqDfy
p3y/JDxRSckXUfJNYhbzciXiLR+Og2paryzbORuRosXWL4xc43nkLA37BB2NJpagel7FdnC+d6UA
WF4zQghuHwXW2QydrgieGwbdMU15Brs0+R5bEUZpb0gJ6i6oRLrvdAAtxNhJAIRcuJTs5YlsHk7T
Fp93vlrWxAfxqvtnoBbxLEg20P/jHxvsTbaRPPZYrXiv2S1rmCWQA7WqNBJyQ8Q1LIcc4gDReL4g
IxnV/ybmVroCmzowyjqQkNGZjff9IkEYSgLKZQnMiac+OmZPSEmaz/ClsqTfjnYq+MJLicGQBL0/
0AxSbQ//FBqvYfanLzXbsObcYGftYMMxHTnKURbm22uJ9x2p401FmdX+oR4pxSu/6rah7QH+LDo+
NbNgJNcvcAzJemTs/bF5ohytd8EcLYX3V9gG+JzFU+H5ZQ68vorTgiRbUXnaGCDI0MWrmfo8PDH2
Ffd6ICXRySJqCQSYi1WMy1vWnID8T9G6ZyeyY0YG7sQ2BFyZDAT+frHmgRp0wToh2JmkhE+6t4y3
u7q4lDbia3qon6VjZfN8ngDRtLxQpRJ44xmRCGeN+RYaj2yACAlWkzZYfi71z8tGW6QhBKws/Y0m
/n3a0JHkq8xn+k2i3nZNy/lfDQImRJsjg8Ql5Fy7r1nJbhmrkMC0TLToCIbQVqo1/uL+kokBv0+/
Tyo8xXrM9uAvVdMKKh612PQgL1KwM5HzV5FWb4Y+Fp9jruBhdkO3jGk/I0T2PVLONbeGRHDcp/I3
0MvpoGX+wFhTRHPuIUqBGFX17Ppb806Jko+GsLYxA7b1yRiqDJPReBc5YEmPTeeEXnTbZJFcTxyK
GDSGXEhgNcJIrtcovwB538+0jl1qgfO5ULRW1abyHVVDf/xp1w1iqUlQ3or7eKEIld8UmVZej2OU
C2iyYVceoX8Luh+SicZgwbSsnWZqAKQ3QFD89TN8YnDn/nYeBCcQtYN4loheSUkq06LJEpwGFMD7
Mb9Hx8PJrKts12zvRhLrIOI5N8E8h7Ob5wnORaGI/1paKi5x4IXAclSEZeHZP3/2m5RjoSTKnOlb
Rz4q41+eeqqJYjSHIu6HjZ1Q3G8MvQ2hGAlya2jZVybewNhOj5R15H09TE/Ea1OTIHn5yA8ePRvr
9NxPmGXXkxmUVKWEXifkGrpYWsPHFSg7ufgE1f/mBMu7/aUJPf3tVdVAO1ONoY37sw+F3d3ScnkA
w4le+6xXzh1W0D6agwcZYaANyoX25Tpfg+IJ7iC7hv9rXxUSPvvffU8tyrax3XsXCOGtF5V3RmRo
UMWJvc1yOJFGuoz8SPTxTNMVUNCG5xst9t+MCb/Bo5gECG/UXJknuhGpQErid3MGr+HYf+0SIKrw
tQH6fFB0eL8QsQpxDZ4WxpOV/VAOtAtC0lzVxbz6++du4KEzn7Xbn8n5QSLefNlgUNARyyZyWrsA
qGnA/nGdw8NymH5bsCku0IGE/nSlnPFPuukdNc0+kjTAbFp2lbNnzhsMhkKYuZSMvrs2TkqJOean
bVCbCxRycZ80Ff6/akJ6PM+v2QKqqIdvYyLwbhOFBGyDV8X6lbuk/nTuW2OcO2jTNKWYMU7fZZiu
GZkzTDdP76tfnaJU+WBWAx+6BjmdsZPV9T1dBiZl2pAS9FL0eZidCAZcesb34enGV51dYorsxjmL
UNpnYbmhsVnLR85EPlAsItWjIOTjf0UZq1xuzA66IEw1fOLOk9Z9gWclxzfl55EEj01qXoUZAwcq
BoPA8DC4SqL0DcvobEy3mTCjw5m6wkvMufR8hD0UgbvjXblFZob+hNsvSrOe6S/Jv4y3wqPQb4ME
jcQUf4y4tEHXWp/Eh98D/0zgxelEWYHmd3eEBvMuSHoKz+yLWtYfMz3J4Iz5P5lf/WN1qodDjZnS
JoQGY1MOIlT3CsJF2cMt22mKL4hUt8AVuzgD2iZyO3c1XuR55rIat842Kmdahmt9LqH63FsDR/zy
bYbba2h4mgufA2nGmmsLj2jHxYR4yCtR0+wUgHVGwkpxlS0JCWitmYgEzyoOwBh9ouwsdw3GysLy
f2JXsWPxAv5ObSpTb36jGBLAV//XkPcrmOcs3lKi+vPseerGjFB85lQ+YYJ7ohJ9V+xZ8po6+tAB
zEIbQsoaDvtWzxkGCgtmLrJj82PenHb4eXXwpV1hRrtk6mLd4WdqqLm+lnrLN87OeXABFsxCW4oM
WzbPMhnq6955hObkyzVIOn5a0xlwXCFC/dXZ6fyZROv5VFW9QuzqJeCxNopzkxnyn7qAt+BOI3UL
H7LyTW0COjbL4MkovwdNvpzB6yox8aNnxgvMQZUdPYiVmEjTDSDcYzFuFaPeQ4msKKtMxr2wDx44
thrc8wRwFGg1m9cFa0uyLyflRSEGhLO3vH55zexEu3tFS3ZxryX4FwTLTQajsgQswOlc27PRcb3U
SMUhTLmE4YNpaBtrx+TGXG3HPjdqNBLac3aCeIQDNiDXj+qa6r38MRyMMGjR0I9ijmMqQUryhwD1
qUnRocG2sdphisjgVmjLLgwsZQNJPQDRy2JClDStKp3licTQhgRSJHbwF5F/f0U7YbsaFoVkKDf3
O4l1AxtXreLfu7SorGHb2sU8NrVtGh6D3xR02IUSjxbHZ4eWEwWjr6yykjnuQiK5XYW9m7r+3mSw
Yfbzg6YEZkXsLpTvCYSDw6nD9OhmkhFki99efMxK3IztCM7sa7wfeUy/NwMjbcu90mJQvL+/43k/
reolh5oRn0v5r/l1PH7VyHiXFZ4Kbgop9N8Eny00Ozvuhu1mro7ewn6t4mt3hJ30dPoikD+cvr+i
+lst7qX4NMtU8FxUWrNukAv+uBBTxtbAR0EFnVsD/my8Ay5Dnyr8/kfNiKBBWBxllV9IYR1MKN32
A16MeSyDlsM4+uh/XZf1ZAlcDvgAv/1r8s+/sPDcMNlYN9hcNYNoPWL8xL1tBSZASluCATjJ++6+
1oVUrXttYeUKdDLTTFXZUkAoG0qYXXZPYEMlbiQ5Kgi6tVjXb4R33eqfpM3Of7hrYCN9a6QB61Ko
tnKIfEynOpaKCALMCIwNcVRCITs1asjZpLUl4wIO++elR7LRMmxkrxwlSJMO2iuo/tUM+m5LHgnc
aoLB/0HReMqJq5RrkEoVzBksYvvE2N0/Jx6mWrwUCuSnM6JhEy5HEXRcNGEW7eXNYuX7VsrNHFc0
O/bk2tamk9o4lqnVspGF3Gl0H0X+/V2uwID2DCKx9qdVNym4vS8hgwy8vFQVRK5vN+BTJFOmdAW7
2wS7xdlv26EL07W/nHCN8+RV+vy72fKSJSe8nvkMRjsIygfHbTqK6hnQYktMF8ykwQim150xm0DR
CE7JzgMMTIeHrwW+JWMWU0cJ+NVuaKCxBe5y7saCA8Y9//m1pQqnfgjqYlAErQyyseCqFlANeHEo
IwHVTbgzuqtUFaHB5QqG1FoxHflZ+aHfARxtLNr7MyJSAzpNSOqQ7gepDv8yxc3Lho9ORt75QZrY
vFkL/anbjMYCBkuSquaEaGYPyLmbviVqgsD5aR0ksAnbjXCLKuzwLlYWJvqJgr4/AUACLiLSYQAq
3tFEFjX7aTHc8iDlrXHwt/jawcLNfx/A9BgcSJ/QLgll39DC/VT1CT8lTYTErKnx7lQUcxZlWAGC
m2+8ajnpOabyYkpPq7oPKTFRJTTXkIBhVVmt1HNWXXkHKPeJ9H+6P7wKVxN5vQBTsh0I0UeXldry
CkZxfN6UxtrLC70WA610+jaWYA/rO0geG6/ZZFMGY5J8RB71YOMtD9hd1yX7yUN8XcyeC+L+Tb6J
1BhVpCI/SCbXj1q+nxmT/Q2mrM/PgtVfsynFTg9uW9Ng0dYN3BVKEKoRbOU878Gh8Pw49PP5VBWj
J0/oUHHvt2JiEFsNbmNUDzpAbAXmFAmlEbMoCo/0v6jvYzNNW9d94w0YQfRrMg0XMSP3Tho3iysJ
HAS6NgoZiowgHt7qcCGAqvlmYu+LYO7AVOAn4iD7Iu//UxUsevqUpJybOWek/eZ9YaDoakJZyY92
Psbb4pQiF+bPIw6A/eP/CpsfGmh0dLQvQsce6TDlOSXpu/3GyetKl8kqmvnfW+2N584Dyw2zItoK
fqDb4aZbKA3VFBPeS8Yk1qFn7a5ClAwJlw/C3jC2O+7O6BzRXkeF0D+nW8HBNsYZOwSQiW0K1evO
u1exU16fu/NFQssd+2LOUVy+NMVxh01a1WzWLqStDk5rR2dKOteKiWayFow4AV971mE1UVTfM8GL
gEzGys/EA3uCWqNpXVvyw3/E2duIkAdkokNoe/6nElTlS1TejTQCx1BNaMDazXcjDauAOubyYP3h
g7eNFqe5GJVWZM7d8GIT6zYnNw2vaYbAxzn8kLqxgPoI6f4SL49B2sQstN+dw936x0UquKgDiwso
Dqm2OXZ7vjsXO7C3g3Ug4cBAVW+z8O91SRuRhR0cDwjexzHhnNLShk56xVQ+Nl8KN68+1oRfwiie
3313cSQAjRF7FXknyvjm419CHAODH93Mjq8Sbk7f3+94oc9qgzGd2JL4J2YkzDxCt2aBAkkj15mE
1QrQkjPD9HK/c6N7PQ3qmcFBC0CIM+I+H+MkkrJG6/BUf0NrdEtxFlcd6L9hzjkz0VCE96pxUCl4
e+hrwaYfbz8mIUtkFbiJsT26cQzQjM5fNa6DQ2EOIvys8nAIVEAKH9IK/Ee9e7gUoF2a+5Uv3zCq
NfYKYx5nU7bCxqGD4i6lJmh7sBjBnUjHssjWP7OccfW4YJCYtpyT5x2xs1Iw+FwA1TNXGr4ZqwO8
LZPpTHxEyXKpiLkEuF8D3yBDXNEVcZNY9DvugCunUtFoal+gOw2EzG9OnfPyIeHaur7/NaO9uLQY
WlMHn5jogr6nbb3kI3Aujsxf/BSjUi0UpbFGNa2QxLyBjgJ9MmxowSqW3dA+Fu2e4L6xLqR/3Moy
6BKWENPH2CaQO36Ctot/mzP/MztFVnlserZsRD0gVrSw3RuIiHWyJR/dmiblR+FUk+95oH5FhsL9
dv0DhLZVbwQ+/fbdUQTXguhYi7mJCE1emfCBsVbb5yXPB9nG79MDUH1RqBzJ8lXTEp4CHb5vx2Rm
KqKeyo/RqKmgIOnxmi0cxt0pdFL2DuwzvTAMT23H05uxSg7Y7/gO5pLE7n/ykGsxCIQBR98FhV/4
bE/oGZVcCxqPAbM6aske/PyPYoMt2G1dwK/D5OhGK+wcG5LEkPyGvleN1C8lISnEaXmsNBwu2Qpb
MGdj9JhvBO8i0+ulve5+jfIKGk81vAHYbPLiiJL7iBd4uNINrm3yPSq03kTrHZtCTrZhKldmjTnK
R0/Y6/D0hiXuaQgJAKWV8uzYXGJ69djjrIMGhdBviMGSW50dJ+LySu5ST/cV1ca2BJ0hLL8hGbUq
yKTUbLj+FIOF0pUumYgfwt+WEWaxatSObrDv9Q9rY01vOJJn4DCjIjLAz6wguZAYUjVs8Klirrnm
yHkpBALke/LtTQtKdofTVkEstAbO9yZFGs3o+UAAfu3Y5iE/CZsjx00wMNPjbDjS4LcBOl/cHFpN
hqA7zlvWb4qYmDKAligSWinxOVubjneING0mVEMvMtZuXrINGYl6Wmex7BNOd9AjXMEUHb2TZcnf
1x8b3A0cttkoB5m0PT/D2XyLbaYnvw6vJ1QtVhEltproKEpByNK2IhMIY5MSYdWBUr3DAlPjoMqA
ZdXex32dFuoAEp+9PScOQexHUwlRTVHamepmUR0sLUdfSZ066GdaTtk+Sv/NxSbyeDBTzWc5oXD+
3xKNq+ktHMprpfmZ1rAbEF20LLNLqyNRRh+EClcfdQVEK6OrqhCl3hNiO+MDvtXIOFN2IyYSnP5C
bD9AazUY0nPW3OvqYShfF1QCmJmOsIKPOtjSUOhicVIDQUEupt22E6J9JphOo8+bGI7Ng+8P5pLJ
jcVYcAe8LJOIQSLyWSuMyBJVaNee4QpzYn7WtOcQYo6x4Z20GxyYSQglG0F4nu/nzANHs3ajGpgt
HHs89/AqwLrDPwajeK3Gv9U6p+JHcXnn6c5ENILFqJkpjJ551HyPZ/s6EYcG4+QILz2e1/hlBblA
C23Xzt2W0moiXZCB9YTmmQi2b0MzWZMNVRCpPqRIm/KCVxOW68NzVL0iVHb+LcZdRmJQkv8Wf20W
eocoO3DHtXso+BvzqU39HfvY1ATbHkCketTPKTLEXTcNGWvucitzgk5W7mXLwreZcz5cyQ6K7nCW
jo2XKPwmyojGJqBQj3WAbgZ9eZER1RARRaFmfrKOEI0/J+JDMcKxVkSyDHtwrXY5HQxqVofp4iYj
bj+Eqcc79A0uVwnVbjJ8jh/+inzvIKDG3HE4XVRbVB6laRBYLpk3XXzpW735QiXXFEgkci2RveyY
UEWDbjivzd/MW53Ytv474gIFyzE2dKDzx+4g9qXunqnY+r9kYYYKqidkCk7q5lPKYr7XRgEAujl/
MDKezeTJJo+Udya/F0dPgM5BwZPgZ4u+8P9h9fd/GmgxwpstAt8yjL+1PA926o65GVsQ/OsMcprD
cKXgwk+UD7QwGPVGuPfdTWq338Bwc9Djbm5ySjbTYbH0BkeZ/08UJQPjr/j3ItpiVZPJnMSdrQUf
cNJP6Z+sAGWVjdMlZVZcuQScI7dFfj0cJlnp/oIM7WyN7SZQ93D1tM5ie8HACdvwzN4/A92Ix1Az
WD9vywCdXKmKUzq0oD7hoTGzXyWilKa7rvJDUxmTTazK+YJYQKXHMVX6PZXv6IekPA49jlMWB7wX
J5tXZwOfims0jDzn3A7zFF5qovNPjEieZkwq0klliY0cMLoRQV+zaz9hfJJcUry7RBccjoD691Np
3EwUHNQFByUblzH5hPp22sFToZ93lH2oYmY4yYUBEsz6g9NegNnNIHTORKhA0ZgAo/ycZkgbqIJ1
i/lIS8ogA9NvNDEkyT8/SHSnrNnL1MH1M/d0UzQoANa7uhvWVq3wXIumbxvXSWLM9X/7gsAW2Xi3
h2RSDYw1ihQWlvW240JcOsCWYG5C1+PnbNHk0OKFDq58HlybUddvXTB3doOBvmqPMmhhrRcUysnU
Xutg6nOdivDUoi8bhQF6G+fpON/6yZeSzgFKHZg6S+zWuP5xclsJyvUXWh44e62N8+qGnTQ4W8rk
jsUHU+oveoOBX5G6QJVtNyvNvtCWWRmjQx8acFmwcu5+FWuERyQORZfCW3jzVkyVVe4opfCBDywF
ODZJLv3W17ophkz2xVqQHP8SKjTIeAAcFQwPYK7jkSwvvQRzfC977rLxOfi4scTCtSA+QpXs9UfF
jgBTl9ZCbGaTzuJmt2rKkKdqBguznheTRflfq6LO07gvOa21BTa06ENcM7gFbxXJw94NZBNZCk36
EnGYugO/GKKEKtTYpVNosPmg90VvElfhknrRF9zBqiGBbbMJM2vrDy7CbiAuQBCa94f9kJDL6KiV
jQBA9qOYyOKGo5vi1naK7tkKBk1d5HU0s4314TC907KdX5G+4aoMZrJdxZRqw6pi4X5vi/kNiCRj
9U3et4YBMJpM5xyE29ljs//dRw5M8dMomPhpdIraOmS4JNhBRXfIOQ7SsZNIoNj5fuUvS2PRWG2B
JtUkuJwL2fXS9VrF0MPJPwL5tXejProIXZErrHHKaw0mCdCjwDoWYLMzweCgQs1cIKbSOYb/jXID
xaAZCm/FNKg1TvMTfcvSLZ+PiSLAd0VRdtc1ol+f6Wqq192JvZtFmzb/rj9j8GOarjVmC1sFELOg
Nfr8hsA2b146XC63u/xYyUV91LlpTFnkcuIsmwYiJ5CrGJJXK9iJMbAY62DCVz/u2pBV3BHtg/w/
g0XXMW2sDJGIBDWf2OnfFmX/dSabDeZLH4Cdb24jfZNHJaRk+8H2IgKvZkLj6xRYeSsUU2w4hde6
6VB+SdyQxbxU7EAF8puDMbfzkUogsm510UG9qnHLI7RB+AmImH8CEcQp5rJSMPIKw/nB5lMm/OtM
okSRomVZdtDlGVpASxySQrF0vbau+wYEt2bInzssJK3ZAPLLro2QcCzjuvYO6RAcicZ6Qc7Eijvu
KD1/xvaYqDp6Nfk0wQ+kaMjlW/KEomoH+/mISQtFjK1LTYXfiC1/KPaj80SYUHlLzAbFUdKDI2EB
xTxWCaxWMowYnY0yhYC5msjbwYST06qsNXn0VgP+MLGGWB8m/M4Px0VG/ozzZvZiMVoTsfEb06dq
U2cCNY9EE/0m2V5O8fmZcOYD1VfNMp2lSwmB6s8hiIWtUj5Ffn5PGgHved6hBTxwhL2qzekzjXPg
pQ1iTJVbyyKSjMClTyy0Qa+aMJlp9v5Qo+5JHld9+0U63tUABFFNO73DGW3exiXm1wDkkDscgep1
2fT0LYrZwhDJJwU1RbRle2VjKsPiPxPqxSjM0dzByn2vsMzIDuiYEfIp1M8cYccTmBDuHaTFW+t0
udraxCE/KcA+tesqIvokghvMvQ8S4WC0/+U8Tz9O3P7osZAmPXaA14/PmR9P0iurj+hYxAngQ5k2
fxGAPPsVJK3Hd0rnZ++wM4LRe20m21QmiANtMim6B4AARWEBt1UaDqoUkwODyBadjxj0S8mspV1v
npqhbVkG8AwBKyFAUA7cuwsKYMRZt8cu37QScDqeMIDRvWXojNWfzaqMaExpOiwxVwxFtqag0o++
agYGICXgGx1p1QemBbSEQ9NeYXHKr3CQ5W11BHjV9rBLhHXW0yGpFs13iebYu1evnQp+DgFkgUnm
CZ4gC3S8Wme5P7KlM4CJu6QjDX7Bt15PK1GpwT5gcoTL6mmESZ/4eii8x85j86GJ906UToYAhesk
BevvYhU4fqTpbvGaZ9hs/ow/FVLhr+9gOPnJ5AWByPm6uAsbuckGEU12JFnn8aIsIu0SA/nIX019
XhMolIoZQx1kG6k2gOFJ8+9gQYtAXTgF8t9K1qlJeKywtiJOUphKwNoVPX2uFFNOLIUldwHXPRQ3
QniVfIM4JR+stdamucruQIdAt6Iz8rmo9SBVErVGeIFNRf45RpAb8vsnop7QJPBMXZS2gpQ0RtiP
QB0Y7qGWYWtJvozank+otJuJ+LtVFd0Xh4WRdZig627kiFp6jdA7kkY05A76cOAO6vMarBo23GKg
WB27lY0D3SaFDsoZxPjWGtqSflNS9Fq2Dh7hFwoQgCMjUqSt9ihGjJH0T7Q4gYOlzMHbw084DCMJ
o+/9rJUPz/VxbME69G+GcwUWvMy3lM9l2/U4KolXV78DrSHaVyK/nxXCtd8KSQehd1sJoYKB1oK5
tvQlv7POf2YNs3Q6q4g8xLEwjBoMXwYxo/s/ARt+rZ0Gi6AAScAQerwB/BiaBjrOHyYbm/H5aXLi
yS2NdsLYdiRoNsGmCc9tqiJ8wYXiV/jshnQo+x+zdXmQXtDeiXJCwS9sat6wOg5ZfJYjOif+pgu5
ghg1C4xGhhwpkZSH7EsxOCsif/oZOXxWR6iWfx57XOTGWyLubg/c3FNd4iyBL8hr57JwoVRwtGDR
niNrUT96Bnn2b7KA1uOQFIg7JlPcCrHr+VOLhrjN1fUaqRvHCBEwVJ0eWPGhj7UaSDwUhNR7Iu6E
JDFvCmoUHrGDdugpEGRHqBDouaXLY1+/9bn5HuRvZz5DucyUZrr7ewCk1mZiDnM35nAIqrQ/qz+9
9+ewwKdP8MUDVFXCZeCHPFPn8M0feNauzITAmD2Dej+0MVatUo4gYpXW7Xyp7CBNfkGjLgxqsKUO
zvV+8QjH28jbVjSXVtiS61VjdXOrZuVAbNNfAuEH3wOVh52RqVkmR8imELj8KLoaMSkL147kcMLa
W4oA7P0Mtcc936a4E3h0bA7YGGNNHeF+Yqo0r5mMp42z2Gqq9LHyuWsR49iUd+Prdb9SGNxNt11y
5cHbUHGurZmKivhU45MHaeKNHoz31gO1uXLsE3Xiwv85nDjppCcM5fQKIa/KVaJE6Skvw0xrGSf3
XprQCt9p6mlKdrT91pRgpZnxbrFHcJJt/yL4diF+EndSMzM5EOMjcuvjyYNqyF9jjWI1gVlAHA3c
bHT4Y2pISrkqFEi2jvlkXvnc+RiRqMHmqm1uHNN5ng8j5xmTBEzRFA2IneRg7yP6l8tq+wmGwLrc
U/nQUGbYk5CiGcTiJDzVFJh24VRyOwPwT1ldZaInfGF5y6cml8TtO4EphDObZ3OpmBd6OTWyzm4J
KwrJf7Jpur6zn4IUg0DX3YTie6WEYhmT76IKqkFOn3j1q3UqW0NuPsABcInwyUjzOfsGHBbxNip6
lIq1NGf7FyLtN5to83KMTGea1t4HGIRne3n8MlSVYbNWXTo0JRW7XYzCEQ5WBE12cR15idZt58xW
bTRog9jIulK9XTTma7iVBipdieF+m7QgeV0pG/88cbhR3zuN5Pa36Lj5sBO/DbFYbEbbdsHsaRzo
fSrcOdzzhI/XjyL3tCNOpgvpMkif8G6xIGOrDMZE71T0pOlKLQ1LPKTLksLfounjpoeUaQ4i0Mbq
zqPJeRrGsR90LMilaBEurrltBSxe2aL1gWsP+46eFxy0m51jG+HXedjjs8EjlltjDfrlIquC5rkY
tCOuYXC2FrLKYKBR1aS/FZm38HrREsdQBELRAu8d2kL14fBg/AXJRxamwSbdRWM8KCb2u3GDSgjN
7Sg5xJQ2vUeV2CpsxWSNpKSkYCjtpy1jjyjwcCNS8w2aMZxBXCIjN3yzklJusfiEgXPcvfO6eCCc
y21/nBRcSChUsFOJ+y+dP1ybPfs5Bn10FNsY9nqja0cNkWlyp930wYRJoPYZLpQgClFoP17AIQUK
EqnbtO6u/IC7LwlKOU4Ux+i1QCrfGsigOqiNxyHBopYiHqK93mMY5ncVjJKGdL5Iag/OrNA9bgt8
68HRtNREYSV9yT19CF2FBRCSJM8I3BdCcPghreQubekEsGSqxzDbJ9Iypq5eGeHybXMx8tbzwK6s
N67I0tsQ1Z/gOE3MwI0WvE+Ge3wUQ1xuEIl6MpYJHpmgqMGwHr6Y+rioCuYPE/7LfWzOmV0izZwB
no8ZERMY2vOSYUe9lsA9zZ2cPNwshSvVdM9cTjsrxh+B9Rycfaiu/0DDQ+4RHGruEyVE3aYv/IBD
5tPRXT4cUzNzyNdAMKp5D/ExeB/FORRNhwY9l0Plrdd6/ppo/7pR1klPP+QcpPXjdyJk4jI5zaRC
k2G3TMvJ5HnbJWDkI4q2vlzE76AoFrL0Q5J7REgOYIj6Kf4/n1y9eMVHOXkXA6iYAX0h4nIlKy22
ZIKRkcr3Q1lsviZF6x+pWvL/9msqH6h4SYw20d07d2CU26NSPRWXKPxzlATMHmOM8cw7tQ0UUdV2
bPbmOESFvsvAaVgg8XMDDV/0bgFPpbVQNYdHcw0wF9c9GHeMuwmFnfqOxujChtKfGk7U0kvstL45
CJZKMaqUuci6Xki+MNyy2Ai3IlPjAuHJyQ5msI6uOeVIJrCqzlVAvf8Ta+AhL9r6ljrdqg3GcMW3
AqA273oanNu90kjUSlmyQAhsIYCN0mhxaGJcUEHcIN2wc1a6m3WOfI6NhaNMSY5gk6WVtz3lQi/I
plyXJatnohPXDi7WYntE84ecBJEvJNyEYbaea22vCOLAeaDIbPsJiUuPO8L3esHVuUAXcLMbMd+G
v1xx95Xgi3rnC/yKu1oX5W9y+jrJt6cXaauwj9T6TSb7ZoCACsVKpQqUs2o7LcFuERq0POZQnYD9
Wj0BgigIIPAn8wIfqyJbKWrbfMpZqAMMtMBNpdZplTFYUKPsO71SJlNWDhqvWcFKMF78Yf+36bcg
psExNuNcHzlOBCobbOdV1BBkNS2dPVjEaZEGeEUz4p/WKov1ne9zxPNzzjmZ4RZ2MHzOc4kC0UJc
EfSgA3fnSvHP6vUyBFt35zSr8n9te4YEvSkr1se9O2rcV0V4pgfScH3Wjs18Fa1loOztXuenoF5H
lm+v5w0MPQ/IZ8v9rsUVq3p+wGrGIRJTF8Xd0T42GMoxHfDjhHJEu1iDcxcku/kc96jFUeTIJ9Ra
Mhe3dBWTNIwsNn1YHWzfRLz1zYsUHwY7tz1/wSCQstc5D0/wYk/tzwBxwaIcxTmB2biUTY9eJBJG
twXt1QKUHBSue1m1DHS12YZWDivmXtqtLvZHi5BnGf4yaMR2xSlgDruhHhPzOole+xV6eVZ7RaBp
AfY0xwMjC77fkbvWm3c3RRZp1hBVyIrQ5BiSm+33Y55WurYLbRug/oImWNDkSI7zOAzXn5wN8R8J
TUOsfgjuTjNIPPxeybWxde1Ctanb5f3jEdN9M1uuutQtwylMPQpMEEu9Dc3XPGUe3ROw7cDliR16
8UzN1FTRss+mjKlJVhijHPMowsJsZjvqyPL88IPF7AiFFqmzo+ViFa8QMDoUFUFURLUIOG2JnBfv
Gxhwdoc1y5EzOelBohac/+sjxXEq4PjaZKDAxe3djJG2o1YJA4LFKDqlYYqiS2UuG31LAk+K/AWB
m8zYSWuIeGvIbsQ5gfL9eXXcPgPxngT3FpBce2Kt8NW+XYXcEG/WdL78CIMmfPIOTmsIFWYuXbuH
5qxDACJQf6gEaqodi2ixps2spk+Ntba1Lc13ZFafVPtn+4LzUCWhJ2cnmORs9EREg7qYojyxLdTK
ewYbm4RmygDQBnGjiLCesIsOuoDZJ0QRgok+IlbbWJ2+C4PWGi2nFkxFC29P/YPMOgYNK77MM3xg
gQMlTvEO7aRmWH71LUEfpxgukd5ESJQVmDYeiK+jt1eu8KdUepYqXLIjJF5z8M8OUfCakXdG+WzW
eKX8VZHItaB4N6oN2jZDdaXUt2KyfzkGbCmcvCZvAp3YR+80ICt2HroObNzN82EU7rN+8o1NqxOX
ayrWXooE8BOc4SIVs9Wx5Tz60puXCo5XgpactFH5jD8MFUebDubrVndh1MvWikKIjbn4U//b9ZMr
dDSQk5s/yg+rhPSfHSJ7KP70W7DoAtRJHZlctV8e8j2h4cTU5/q57uPeeXKb17dpMXaHxDVeBAZw
s6/XOdg7Pk8d2L0QUcX2wKF7j4vNl1q5IY3QI6PkYBLkKwSSfEno0zmsBzvKK4DXQSMzKxdIbZC0
kk/0NQWMwQitezxtBH8wA9mc/DZIuJ2b97Ha2VbuAzQhX1LbGS+4NgZUMSlVKbU0/yA6e/WMAar4
htx24Rl4SHNicb+F61ktosg4EDujU05r6PfKBHokYuXuUS8TXDWz4xj8TLvTOjdWxCpIaROo/dTc
sXZigKPvTCMdFZzUpoFmm1v+1+n13MJo4NL0wsCdcIq34DSHDjM0kw0Pbac/7YTiIdoN27U9AIMd
vHlXOqBei1lvf6Ijv+MfomDXTZHxVugbCl2gjT3yrjGTl10emcTQov8PFwGMkuHg02FzyUqmLVVr
pbydRBdCDDYVltlaST1+hOcPBZF9/e8NgIYQc+mAfilmO3gCuu/eFpojHASW1YT9xmGnBhNBLXTQ
lYOPoXWBKB6td32W1ukKoVAzIlT2TM/h51KCF4d96n43xPVl3QEqAsqAdqlUdBOeMfaY3y331/Vg
SQVvorMRB+VHaMxBlRTtQrBssqR6n0wxaZzYFNNUdFtqMTbTAi/8hZZXW+40f6GlkzxthhcPUUBw
DE/V4940eDj1VDAYm1a96yq/tvpc5WMBPkYg+sfxiMJ3H2YBVYx9aaomMeCSEE4F2vt1KgAkKSFu
bYlLm96uRffLf+1T2qokl0838pVJCqMy/06XkElaCArz9BqzV/9JhjbHeZmrVKhFqpYQHf1OfEu7
9hqwUUWPY4wUdA4RcUFj1DRe7TxWMHEvT1vFopVp4lwZpaItCF3MS5h4Ew4eZxcJHemcTJmD1Bcd
zEbbJ3rrVoglJzifjQ5o08uprvZ1sFwiekn6eKXBS0m3EJv3+aYrciB3Y1TSAOmSHul8RJXq1lDv
JB/+TzQAs58MzhJi8OgRvqdhmHIfu3vTSI8vmFNCnYMYWUbzDETPsWFnB5kTpcD/qPmIeQWDdKGk
KpqvqFl5HbLYKCQojHsHXb5QEYwtLGARlJi2DbEs7DY2uCYpyev6Nli3ItmJMW5rkPhRnL6LNY93
CReKGeh/p9IrkAFl3vJ7fXJO7LrJtfwgh26Aka4uTZJJCNRofTz7Pg6aF7QeWuYuREna6Hl+bYjo
02qcby0KUGCuxfmrRNcF/A8V2+e5oOWYrROlvMTfT1C4/GEVc1IESUUVP2CjWeWEv7Cy05orUu/+
8Hn7M0uASgu9wfABOEplCxHwy/wDGCX/cPGRtgsraajn5igxAYtTtucmLImc1PTh0QfqBdit3vDS
Wp8ibUjxN0YrX0gMcWL+RkkR0QTGL9XeKfNaGb/5LXSpAx/fA7iJNCz/tq/chfLtC0IWwo+FWVxi
AEfrWB6WEwkYcYzm3ZH0v9BOJBk6RMofsDvcPogezSXIbJWQL8C2k/fFSfbpml8b+GYJ8nMXI7xH
iPrqejYugHtIgcQLtutCxebL92zFKL+Z/wj85nSmNnTgLYMQdxaqtk8k6Z4xrzUPZx+7hCr+i29q
f8taCaPZUMxmqosvGdfm1pK2vfgudxkvFlSOVjJSpdgqca0uCk7PGxbLxhf/8AIiXshGUj454gWU
Sc58kmFEVKWTzzqOsbyOB5g0U8HTqC5tOqzK+ndk5zwAxACKmSnCpI0VFi52V0Mn974YTExIBABp
o41aH79Tsj6xfjtc92/0G7q3SxoFD67lnoCyhW21Kckhth8NY6mxehgo9ueJ+aZdrZLdutSo8Yfq
OMRLaGnYG3Yqo3/oa25vZbN7QY0lyvGdshU2M8fVNHXwm7RlCD2RwjchyvVU8cgysXsghJYuCs8T
VaycAjY/PiTYRiO0+l3nBf4THt70HTU6o4WPJvTrL7ktXBoj3iwgBYYCag9fQ3/l2MYjjdbcxc2Q
3z7u/YXKEV2QCdasKSqb4D3uIfYTChnINHTfhP+AmtymeC8kSFBjkYTRoJs2vd52GDvlbApu45tN
fECStqxGgHkdJjzCt9/MIcU5Xh8oKsJU5o19x9NcEBLyBymR/1dyElBQ0hv6HSNjDjJjJ5g6HX2B
T/yNr++oCAj5lBN324F8IS2eioC18Ra2SFW+Gswhpk8VYRhmn3DLBg0/27X+Ogkb4uupKkvSHqS0
nytPD+v9e/xEwvbFSdoxOzH/a/tkld2SPs2JUfNsFL5Imox2SmDx4sTUQwGMOTuaM6xKoX6kPmsr
YdngADFVYHrO3KNmaE3azheNbPx7GfSzgJujvh+omTUKolg9WQo298MIc5nOHNcDdvI4H14CSkLQ
T5wxWoC7TFb9XrGzbK1PFGr03ZvAeDXyVmW1rde1bFSYhmxHOe6uPPcFaDrj/gB6K0muLa73WPoA
cQK5GuXJPukujvqF2co1/eUrD11aiQ/0VyvxdCJ4eH04p2u0RKuJShXgB4kbojNkLbdoj3cNbSGK
+BKxhrJIae8G0VoRwHnlQvHJvxARMp9VgjXzjGGXxgY8Tpxj1c1Z4butDJqFy1BoDmQzjmEjEbDP
Q0a9HywB7HyU+ahW9DGXcGLZlel5Ch9EPnLqQntXQ5df9LR2ljZNubxhlXrGQcKnMZ8YbPVxF6Dv
RETtGa0CnzoFBfYD6oc0p7YRM76zfM2UHpTeNC+o2anRjqlcRL9JqMJLh5ZGqLK3veuYh7kev8SN
E0BmL+XFL5HjUcCEc+zFaeYPf3AgFLSHq2z0s44I7JFl6czAHnHSOEMf4tzEute3mtZx0oBZSrr0
qchoPbpFjeR/I4XFh0+WDpMUBHErHskkPPWxS4GG+HAQ5ehuFSjYttvXyBHQTWG4/KNmu+I5AMaT
FVBxXqRI0f+hQYhXCrHeIfcebpxTJH9HoPXZ/SIkWLlXcjwZ5GXxOEKsvC4DrBd+Byf0n1poY4MP
bM+nqlGdMJLQWsFxgeKwmfbUktgyjCINLOtxrVlUt9pfL/q+gpCJes302lmarAxDNSqHQSGZ4cNg
FZgN3rs/T8pm8keQZn7xGUeL616Cps1uGKDeeSNDYdhBMkhs6iLVyFWjcpAesPlxBrKqeM+yYYEN
XVn/SRGNSFhO3evrCQL+mT7fxBRMaOtEBHNqb6NVamIKgbe0PeAHvIQVPAC89oYDXwBCW82fmMKC
Xe1DnsOJG2VpDN60UAvN7+RBGvAWo2J0Nq97KB7mXi7l7FhDIDV5spa0cl2ZOG+4YudZHUdAG4dj
sTU9rBI0Z6pzIS6Mj9xRiwfkRldB0u2qIqHZYr5JCxs8RbvZvOLzOztH8yqtZvUCrvQqdx0T5NNi
S7+JsPydniV6okNp8JHC2VZR+Rp+DAV8+8cc/7shAZVDdExiXJviCryoRwY9I/NxjSIduY+RXJsi
chisyt+kBsNuCRsYwS620VU3PCTQmisN429UQBZuvh89cpcFP5AFJ5uHCi7HAUNb/ceNZK1JxdIk
x/CiNFsW+qL//uD7mAEgs2DokC145R0gVtxDWZI7C6TMBppY8SVsQXzpF3xjOH6tnIXH3okMydkG
eGSj8r25RkiCkrBIhDMrLEHNjR2OmJdoSwEya8GqmDvwDM8mtqJFgkwwo8JBDwukF7gcLU9FJKiE
qen4DhgMw36BleEOPszG3xCvHMeDI2jZnxBjCAFal0Yzp+Op8Ms0XOBmAvMsnkuqf4htVML3Inqi
0v06dJKiQr3TKi9oFXNyMSH63F4NO9wjw2CmmTt1BSFKCVb3vGctL5jRQjeqHDrzsARHzZp7RHDF
SfH/i47jwbpB7hyhcUItn/PPuB9JBk+IaKQKoXHrgNiuosFSD4VLrNKSrLbxU6tMnAHNob7Oom6T
lRUcB2dIs5Fft+h/EcAXXhFBagb07NsbZtsbWgo9HXZpP8f1ZF5i9dnDDelX9SE2xBIjQs2MbG7h
WUa62fsnw6LDOaHzczEsbszmTOWIv2Xhjwhr1x4fGk3CtwcicsWLzK0fNeCMRdhQV9ahtpO5gTiQ
tKZeXsgG3tdp922Lqxn+A0ETedI3hGQUVBVB+Ooptxn/lsCCKDY3YGC0dSD+NIaJif/GiYYCQQH5
DcWJvkd6EmW8JMwN0yZf4iNa5r5sBdxhXZJxfVmaAp0dHbdP1+DP+1cZqKHIN784gamBzlVAdby9
psEPSrS9AaPD54ePGA/Rvnm0i45GUyC+Dd07KgQtjRjohfW9p4ZVXkRQykdv82kTOxvIMAMyPme8
pWT+uYA3c8y5kMelHqJI6eiaYT+9pSrJmB9hxwz4uaysmCQVvyQvOirYl1CxS8t5IhYhy/MLi1+E
Hqkz+Y8Zvf8ji/Feq39Q4m18FC70sqhTfSIroFd+yAZ2sJ2IoNb61fDlRYD0b+xRIA79pPklEo7t
SkZHrGbeGEZvNruftUJ2h6SXSiqVyqX4xqqpXvwDM0BHcoGrs8kingGwIAo2DBHmnTQqEjZh1WcZ
Mf5JViulQLZFFb6wj1RCYt1wkp+2zC+/+JCdtNcrXOeqFQNq/598fyQLSLRJ8zKRX+0ooLhMB8dt
RsIwJOXQQ9YJeVE3tUq+ZquWjYKJ0neJ7apF1By90+zeSNR7kG+0+50wwhuTgmkVKGcanNd5WRd9
rwwyBDqVkDd/Vlgf4qH57YtXVIp72x1GmSTfc1VT46EXNlrhrqdoek28OBUSx7jYrsMuiQ9wa/Dq
0nXZC6/ZiqOm4lkqJUrqFDGHSYblV4WwvJ/fE1Ozovwa3XEjytqb3tbCgZoELv6u1GoJ3SCflZyE
aWwGYX0D4xY9BhGM1pvO/1nTadoGxIVA8HuayYZHRNvjHtBLrovZwYqQrJSQA0/6FmkVRTWnRqpT
rFTP/Wy64tolYILoDG7o/QXARaBC3LbQiiE/wG8bhnSmN0VbyFmJzJCWifFZg4tE1SlnLoJJAeBz
1sa/fce4kfclWp8BRasScXfHmGMA0u/utzJYkRH4tkBvEnKvk8D19Van/sJK3uZXe3OKl4VT2izv
a7+aKajsTnauGUDAwK4V8DWNjPtw4xoRjZqgzrtO659VNN989MmNsycWxmuehr8HVvOqb3G7iq10
dhaU6IN3SdvISwjxxJCPe/9oIojwhj71bV2r4bWUIRUqJnxG6sB/yWkapUzgQySsj9KXR5LvHqNO
iBX+hGI9IpaUJy1r2gfHnbwq4jhnzeyIf/U+LyHMYQHlXtgWNBR92luZwu3qAbx/fkiKKt+cdzQp
QHPmZ1DPMTpJo79eWl+L9Dea6dU9WOpnDRiyGsoQAI/gq/bgRjEPYv22FkuX0NX61+uPEJzZ/iDZ
0yeMO0vKYSLQdqCxvtkRnjuXC7+jJAZZ3d3QfaDOudRU1OlJyahZlVDNJcrITWcD1J3ioMbjru/1
uguUTT8eMparD7kkdH7fmvzejCCvl9o5I4VVd+JzgMwS33FoPcbWtcwixy0mm0IlaijQqfINaE0U
LEz09WUak6d/raGNwAcslnKQCpnRKHdamh4E03DjCtTm6xO6uuLdvost5zfOh6XMIRT68LUp4Rpw
+bkkqzlKpDKSsxJOKMP498SuwsVBIhaXRTZsBvc2B6zlRC6Wpm/aXWDfADXyuRQDzegN5MkevPU4
MPc7Cn0og2ELvlHqJQwx15GOtO47KNYGO9Zwok7NYXXmZ2VkXifLneGFmRlo2llWGkzKsA187h7Z
pFAUIsDuVQelqTJywM6wvd5+ie7WlL9vIE/2drAWedYze7KZVz+yZZ5qOmrYyS9J+OABgfvN+GDl
O3R/f0prbJfvQ/adpSD88dnL/kVe6p9rE20MDuXqbJJfgMeOsC7/NFpAzjRU8/6JLja/yC9bx64A
q+D48oyDwNAt6As4ONhElyCsI3P4eESkxiw87/FJLNWhNFCHGEWQ/ai8OIpTtDKMiCAtcmEAyipa
oMvPilEenhSFe+JtbzUNbzqntgWQdVkOfwnoxmM0flI5xpZX3kDtkYFvTA8gd789OTOXDd//AEFx
FMfzcX+4Fjw1QQRC39Qu3eNNoaAReWujSAdtrbtSLjYEs3lAaojHCAMlpPVwTAkFifAw5L2Rys/p
+6vIcR8Gzhh4HSfGAuZfTzGeYd4H1JxL5EMhraCF9lsfH12Sa2hXtY3/zpRLt85OMdHwxLVQmkra
LrGlGBD29x2r9dRObN5bhtNuzq173Rb8rjQB1G4EALIAcdibA75nfoRm1hdwM8TwAdsQdbcMb14W
emXV8Ko2VFUPYdzVchBt20lo9jMFx6K+pp9YghtPZFK9zmqIrp+OZtkWEdct28JgMagjotrLSqDl
StmGTOXWd9ivp4a+ODDrkuomzjOivs7btw6pxU6UF3Wx7glI0L/fId26h+O/DeK9va2BhIU+LUj4
tKjsgYIB7KQsKysuJyXRvsbO0xqGx3p5n8dvoKhmpzREZRaqUqKROe3VQQpbTAdIBU2SaWeacRgz
faAiGFQt17nwJtXYs3F1kLP9pXxwuYlRgrXSb37Lj/vjds7D/D8InY3/tZsvksY4cyXja2W+Tqgx
hscKmq58mUceHB9JVy/WIeLH0bn3GW0rdW5x3NQPcZG+u0WlvDhIGDFbDHxl30d6npK70hPtaAbU
fX9rjwzdonbffGnQ6eUwD7t3G3rg8mlv+0AwJ193JRPrckfA7rfaRCTtkIA7akAbe+ZQlUX6lXZr
H9pUpJSYf1u6x/jAPHOKA0n+wRjtl3uLtxRWTxZk/aly8l31CWigOTxhgxsHfbyEqxYY+R0CUQbr
uOdIVO1DODs49jIesDgKAfwWt1haAYvFQrnerNt8MsCwWvpJR4j+M2wvptCAPiH/EGd5WEiw03h6
0ME55PW2G7r538tLjZfrwIWXQ9BlIBuEYkOisIADdp37QjRZy8MNKEzsVW8HS7pEDIMkjtsMlmoM
o53roVnQbJqOJHSja9AkqHNZhGRJTtsr/BvoZgGJFOcIdFL25FsmYGrDNvo54yem6DvxIO/NB/JK
9l0eRPMxphfpOnMr0BE48gBqg64uCU3eT7R6v5ab5Mpg5LONJK5tW1yCGLlzTI9enBhcRXWnuHU9
aCK8iL496R1kVayMpOAl4EybrXv9ZDnSk2dcyfMWoVKqCM5ji8QGU6uLln0vFVs7Yz7rdbLflcMf
GV9YXnZVd52hKAUhuGcOLXasd71EHpLBYzlDs7xFk44PiPkQpClXsabE8kzscrd3RsnupA/w5drf
iFUxYtIGvBkMn96pbUpU+Ut46D3U313pgieYi66VRAl8groYrn8X8hCGiZFekSK3NWbEttN+bLh0
owFTT5NBni7KoqvzUtfSgqcoeNCTKAp8Rnpc2blUG1o8cVW5qHdSjA3duSSd7PphUiXjKZitxyHB
DY28dzPFIgl4TYiIetcIy+4wymENaaD6QaF6PaYmLWaMWzsElPQH2BgknQl3TeXa65X4pvVu/DVm
PlnCHF4z6pf3W0BB13MnWeBTeg7BqPslRHD3ZFtN+7Xhz6pw0WpPNXwqX9QTdgUs+FFqxXKA4ZGf
GN9oehiy/M0ecf+Jrv83PTbScKrrSZsLqbrm+8Nw83bOe20CP5BSHfB06TUAY2joAGtWZJUT7SXt
QSaITqxeip0lxEo5FN+G1g60JamTmGSgCOZzeIj4d6SwWPX8pY5cbDpR+3njJ8y2Xmi28o6msX6e
OyU4abHnLgbb348LqC1Md8N7w5YPYfeq+2kUQaUfm3Y1SdVNI0p0RmToJqKO64i9phNN+mCpgV0m
0LM1099PIAgLLCEy4ZzxO8D0CICatJA81SzsJH8AnbcZM3eB2GtKg0sdGm9qXeU51eE1SdFQwNCg
ar1aeYiRdYIspKVPxvY7KMTPS9ac6s0BgfeCkvkzRXXuRcRjRLscpqkgYSJ/RE2bh7MjXU2WzGH6
DmF+Zw/GanJTu7McUyf4Jh0kBM07Jap3rB+5E5BWJJvcXPJGsS0lP6km/IK2EdIDBQweR+ewtSnC
9vp7/WCHF99bfADSGir7rb2Jm5+4KzSyFFm8GNguHEB0364tUzLEKZE7FK3bgXul/nxOVh/lipiX
KTNMLobT9RwOE1lAsM1wtqzDjARC+Mri2jcDN+FF0cAvIf0vthfpLnYfOUf4c3NRXe4mbBLPKXUg
swjVZduOtQyQRfNnNZN07Xr/vrXRWIKKm5X14XcorDJXxVyEQqXBuXaY7rSWKn9ETTOZAFomiNkH
owzlglwRhCq1zLiaxySBAAeAZkoRj9B5nfePYeFNqjHWoXwinbomNeL6dcBzD8XCY9udHve8+Tka
8VDJhKjKd4UKFdvvPSVJsRms/Ts206NkbYe6krf7uag38VyfmWJOLcZScl/PjlDdaz01q3EkUhKo
wX7Xy2A0nIVQKXBTqEOWK6OtaqTRB+f9aEJOP/e6m+54DxdkDMq6csWB5LWbilv1V97wFfMxviea
6AouSKiMtC+mOl3vopSaoTlF+N1AC4JAyrTyzIgypY3BXyMChoqMZdZQYddKsdxYi32o2TDRWhRE
3vi8dPLeOsWGlTpQWZrksmXwtIqMF2E1yKSnZL0YK4pMECijoZ1agxtX6xppRFkn2gky1Q66iIuC
2tbTovg6wWZpz87A3CuMoQmG7WBXOLOzwkn0jypfzvgCyGoMu1tqCr806AtLLNEtxNBtaZyrjiYn
JKneiwj0GqllNK83eVG8WejqHaIFKb1hsCcMidFxDkSIZ2xUXtWB+rDlQ7C9qk9TTRY0/Q2kBBx8
RXWwI0p61tUpTb6C2BxyyicBHsyDUAn+hcPtc4MrMrYHgkXBiJw1XQqbePn3gya10EoszlQHqmDy
HSX9meJXEQtfmsyXD9WHC8nryGrzEUpOMFzX+qumI5uUSSkIna+KbezB0o9cZ7geUXiQ/P5FkLEC
aoLg2cKv8lQ2o/+hej+klFGe1kBshrnYikrr0pCSqQFcgyvMcVRMUEZn6pgVuFkFdf3LyZD5xzzi
DmkblWT+EQMqGZLZFRm6/B7Z2hlIm01fuwefJR3O9u3JpwFmUBq8AY68b9Iy/ulv0HC8O6as0itc
PNmqou1cAULVCHQvubCGNJ/kZAlgUfk6dZkqX4Mht0+P4KGj4m3hsdYCn3uk3odFWPEo0aWGYQsC
AuKzodppP9AahQMj4Xi0ZUyG5j9gbEMvs2iusuhgWUsR7q279W62KGAKwQvJi2m+0uxUaVtT9eJA
2HGvbXIdXyxlU6TIsHae0u37lFvfy7gtmEDsp2abh/s14Izc+KmBAhBXSSB3EUBqeNixxE+bJk8+
yywyR1Tt525wbItnPF7BkpF/njrmpUMRgq0euIalKP3gZRzq3q7nP7Sfj6WBfHfSWPXyZ5sJqR5Y
B+7ep+8+hrGv8NOSsujw9uGEkz9/KA7ZL15HrOja8ezMEzKYCnYYyiiHJa8BG29nfecDE7WZaDA2
RY3VvgkvvLtsI2KlTUT6I77iuriY6aBOK8nvdjBUXWUdBKhG6ajYZRKxNLRZbPdJmMo5NPL1EFnK
FIxqlLDfptlYdU6HtdlHq4iTKNn6j1lxGuMFLA9X46MMr+0voSEphJ2l2bKB+vuaQuL6ZnYRTgt7
qYfndmL4ET16RepkXRD0AHZ3RSOnTh3cI+fFAVXrhkRe/tKM5vWlV8OiKTcsvppSQL2oSxfxfmG4
+UdaI314gTVSQ0046u0gTvtz4/6/MwwTaXUqttTntnr42fv1QHw0J8MajtK+vPe+8Q2PkGcaGz3v
b4/rrbVA+WynUfTNV1GGbU+AZwYGQ+M5tqbdRO7EOHLt9jGhbb+CE4PC40lM2/FfPj8cbazZjb0S
jo5jzkBB3Jg57tZhyf1DXuFvhkhXwbT9/+qRicnLimmrcg0wmNHqkqEqwwzKsW5BdTJZW/b6Lbdc
RZwqgeN236h26BKp51lJv7omeHIldqiD8TBXBabuY5GagCqoebYS7NTqaUd7WDt6YVMj4uWl8v2R
c7VuLW/djJTyS/hNRK6zQ9wMPiweivRluP/6ZWZt4/IGA0NfhsyFuB1seqYyHdLWTgrzs6Q+Z8HJ
knL6WdgR6MirQKUdYUZCSeJBWeSQOKG8zjYg4DuuQhD8l8IzLtVNbzomYD13sNzZkqJOPfYlDSlG
H35x8Khlvxin5oB2ZU3Ab840HfabeIe+7Gi+NJYNJGU0ZtDB8m60QgEl2zzYMjqE2n7nqzfHbIAN
vBUWoQ16vLybMlx9/14gCWmaabCpNI//nBY1gy3KzWjC/mxZdzgmRtezWn0JGSRcL6MEzzPFwpwQ
sPMLc/m26em7ZF3yEqeBirEm5noV809h43zXHwix5bAymZ8PfDM99j1dvBSdyrI3EdhLg/LBhYsa
IPnOeDsBwgxIJvwzjTNPI/osF7jpjfA1ec3Va+rW8aKf0igV1c8OPlZ4pA1LZjFDGE8WUDH0rmiY
wmv6ucixBO2mlmIe4NNvnciQQseaqWctkJCseCILOcho58LECIxbgWwHhKQF9GyuDSATEqCsbPyL
5iGcD6sU7Gv75U2S99krAJ0tmSZpjAwddmPViJiVRLYctK4iatP+Inlni5J5v3LLRBucPwu2/HEJ
2PP95QjkReOsUTGB0CnVN2IXFKR2qZrlg37qPP2f5OAe3SbRhPVvuJVRso1doHlk59VZuaIULNns
jbXA9z+JvQDfIKpQCAC/A391es0icsRBtmn4IpKrvhQGOqWcQckGTquyTGM+XCTqEv5eUh9eAyPu
Cuk/Ub56oGkOEhVxOJLMZ2FzEbeigHErzvQ7oomTC6oRLOMQv7k2/LA/5h5dLRtuJ08/zH9vejeW
eKxcjlUlgn7DMAyEMMLkvjElzWdNC4nnoC8z03nerzQAZJl+g+xVHyLEzUCsdPgJyFxpQdOpy188
tE0NA4iHjrq68o/C6oF2h1kKP7/0hfv+U9Ah3BwaxchjfnEhym8eDtIy7w2Anu+kP2iUq2yAri7A
f32EOC0gFE54SPjWZ6SM4IYHoPqOERlnjr+djqwllHovrvMyzmOb3cAhgN3U+fJzcyCF4Cja0q1b
fL69/wd+c1n9MMKXvH+OYFFuOyIWwDqZbdzkArh7+QC8ZWkRLm35XaRErZDYfChDb9mp/3eJWbH0
egQDMuKb3ELllA6H9xVtLZQyMNUB2Fesj9krxBLjSl+CngAI0mZxWwmehSMcw3CcgutW/RUQRy3O
HAn6m8nPwUstMbA+N2nY4lFvzo3N3GNdM4rixvIf5EuOWirgIaIX9vT4fxkuqlBpJtTE5RUQYF2z
ip3IBb/+9rikx9TSp58YxIJWXHxggnavwSQIU9jqOd6KUIJZ/vB/V9zCXgZYtsVhq8aCa5c1usb2
A62cX35GU2u7d68ereA+gLuexJjZaLK3reuMdIGxoz2S9bgup4uulk3KMYTDo+ies4maUbIRcJxR
6IXuhcua86f3NBCfBMrbQkuItc0XARRXlTBM3mebLqeGvP4iMSFP2r6k7p1CKBKy5pwYvdPb+/lr
XRq51H+9+XU5I1bwe6VhQ3pFiBY46wc+ZBlunYgPBPyd2pSRVqZlhuh7z9Yo0Q+Di/tp6U5+LYcR
YYmHPB52E09Gu+IfnyRYFBuPrd8gWXeiiwaXyOC/qh+YEMR2EYl0IgyzBtPrbKPwW3kueVjl8s6k
FLhT1VMpQL7Fa8GoCiDb80BiNs7CG84m+dF2JMHeaFUJeILrkwlvAcAacF6Y81iPRwBciCXQeHw0
bm/ZTcjm+XFZ/bj79CHVLSRbDfKvZvL1Zq3jc68AkJS8jQpsZiwNJ8rxZJaGTVAHBPG3LGWTW7r9
3YwvBwPw0+lmugp7ZB/QJA6P/s1JogFtjygfN8SGEqkq5XwPUsbBivweOG3GOVEmDOT8UN4Xsz5k
gv7Pw5ykR9Qxct5OdOaCa0sYmHgc5dibDsVnjDuAIzojAggIDdOXwAmj8F/VoM6Y9K6hz8n4lWKD
hei6xmRybt+NhlieNYg5RpiE2OqdtjRpegcJ+5kROa2qi3isqnk4CNDJWVw8n8/8BBHciUeDoY30
MbZbE/UaK5l1gzSNRmMKYgxLATcz1MkvtYNIFuw3xKLxH310+sfNfmVgxgWhVnxZU0xAvAD39mPR
/FgiHkn8WNsBeUorxRy6EPbOfScZXKlCFR9siDRMq1FCYwp8lvmY7W4WPqMJWX7nax5Om0/9Bvb9
wadmGvTl6MldM+DbYP2nIhoQ5JR93yaDLeST4EIfrqovsiRXS4Y7xbOiI+Gzi/k/Wp+ZwaFoPnsu
3t2QlsnS5jOQhuVgaNTGfyF0dxMpZrbh5GOXioijpb2xVm1DJ8Y7GsIiNgVbQyaVdw96DAzEjecJ
JmVAIshv22el/wDA5lKiR2Hyt9ezwzFGfwNNtz6LHoxazd2F//E0EdVfwLOalbUunkmgQ4DUzxN6
Ef2S7nb4cHovrVrnM6MRc4XIGA16+hRjJLwQF+PgwTc2i5xo8ILsOaDJg/rCbf7q9f59av1cXhph
xso1vKBKzSO2b47agFEk1XqLgfxDpVebji3CWObDuS4O5wj667iFbKntkTaQsraBJNBCUy7xo8zU
RMGl/3bLCmRwx7HznXn8SC9PEok+elkJUa8aMM2x+Xu30fmHHcMKFEYd00YKoderXLk24Hdo5cNq
aRNEhXYhs6hCqQQVuuOExMlxkhJrRS6Fg7ULux9mQe905g06MX/eMCva4MQqggrc/KyjnQpTqteV
ttVgBDAFszc0aotk6h3T5jNP7yfnXtEH4wqQD0bRn2BD7cKQdDXnOrmEd2IlBtDRjo8VNP9xpw35
xx1wyMpOCToFRnM03jxsl0xDiI1ZhefM75okH7ZfUOMqG/yQnipS2DybH6onP83eufiwHXmqcMfy
hZo6lnlW3OafkdU+8w8wc8DXHNAqN+ruJpEshe7QMFcECuMwhV8tOhh+nrpX6qixkDwom8qoq7vb
YQWv4vRMAWvQDGq+Yr1PVcKjbahptQzrFM0joM7/8aZUrR7LDt5NrMnCn0OcvFSzak3hPPKVJlIb
R7asfDelgOqEhggD63FExOaLWB16kQpyl8W/vakGslC2D0yz4dgHdpqD1urmrdT2DfNyqsquIRDO
AXJrVTnvd360nY8hMmYgtbWbaddFWO00vAUWcdua/8oG6nL9KYR4KBLKxUPOspH+LrbqTPOk8DZx
rZhRBobPDnNDhB5Cqaioe20Ym+KPZkXLUc++eQgNk8DwG0e8GO2/CfSgK5cwSAe/4r5lJqEiuNDI
PXE5eetywj2cbI/Ov3OF5oym3S7AshHQ2KZRstmw0eip9spItgB1cW+VgpHuJ/7f1/Da9ZgQrxgC
TaZ+a9XQzTFuVYoll+pZxthG1kmhmoqzOaKSHSClKpgVqecLUHLfKyFl1VyN8M4DBl2eVaxlRxA0
DXpY9X3ORrvX1e8xCVD5ejjR310PSdQvWBWhTaKnVrdlb+taS5UhVBDaiJG90OqlbpclkJEw6hgC
WSW2g3HfP2IWQsn3Yx4qc2oTyHyutilijJ/aL3RtC60gRenc6KWBJxgIBNb8u+7bKcZ5b08EPtRh
crN2cdNVnAvQQihI/Jo5rgJJJAN7MXYDMxlvY4p+aOVhahIp6/l23YyyUb/VxampuGSvpbWrQgoB
kVVCeY68/5CBPlpfIE13FazpyYCSNmh9UpNjQsVQMnr1wcO2S1rBelvqqPKUGTC7FcdgiDnWUsnP
zc2Iw47wQQ6H4aLty5QsBLSR4JnlejojMDrpEOjs7YHEvEV6MDt/xOhST9k5ucoF8Hjw2UFB+omK
tNZdTmHUx9Y80Gqgl9vtvV24ADCtBjBqaj+4I6vNnzMKtnSXg/mJzBBvBd3+rcUT/VXBnrroDfBq
Er9wYi7qTe4IpBFtJ8NN3TGId1oIOrXox1wal8Tq9eKNoNrdZp8f7cOBBdni+9YEIB0a9ReyUVEU
gDMmoo3qWFdW+hKAC/HPO0duE4u62PEpKlOSdVqvr8+rT0JA2nSNiUafGSzE+P5VjV4ZXwqkG9/m
v2jrTCPxZ1JznDx5PFLmy3Y4b2k7121W2TD0KvSoTFT5Pmm/KpLJBOtxqPj0cSUp1iW/cgmXcwTg
OaoIR6yCp209kEAzVca++jI0L+XyNCCvD/Y+uxRm1Y9rXO5Cur4FI3PbygYWyb0xfFYtbD/FYj7/
KzplbZw/JlCD4KrAw08nrz394QNwnttsgH+AjJ7B54t+GdxQDnZbXFy0sRrE8lvJYQrCFBCa/qnI
mN2Pqs/or9gbNAFI6GZYhpUNGxKZUMZZxs8mSuZ84WT3sgzeG3ni2sX1imfJqPO29zbO/VksEGkh
vGtkpi4RLUfze8vbPBrAzANkZeRCF+HDV2pcV0WKa2fuT+25LeVcond/d8Dzik4EcKvfBJOfVG8s
2HiX5R9VOYEAFHhYnLmr2fr0zKnnwIR4SFts0vQzOzFVyVEndTvgNA00NhnrUvIw12aFL+Y3OW/I
0ci0wn1KlUeNPb2P6sZHhTBYG8ri9Iy/wjx4qGhePjQb5kc6uPDBr9gexLTNUp70jiUDs3l1LqZE
df6ou/+zW/sGaNmjpz9PvK8q28neOT13M3SIYB/ODhwTBKqs7mwQw7zxj6gzEtsjML43KSLHA890
xDpOag8OR3OIwjnHoIfd1DZRta5sAiXrBkJCSyvXzk2deOqNhHLuGLcatBEbKFmqvdsjh317CQTK
IVgRVFBNfjhyOL8kbWxo2DEC8RpLReS2+mpxnC4t9Tf3CQV/vcD5DYoXXu6xRyAuzvuvQiOca8LD
m3sz8SptPaJ9MIAXv7KKK4b+afNjufujn/Ism2hpOZCirVfx7FmA2Si6CXBVp8Us7un4HqjWz3nH
W+C4aew2ZTorBIe2kUm4Wjs9yYHmnv2YoPyq35AVFrvHUGttaaa9CJDo8bhNzaxOC95GNXQueIdf
tcgVWsdteHFFppRryRP2s1Rv7+5YWwf+s/xVq6yGMjoSBrhMVDOT7RO825WFllDHQwNx+WfH9o3/
bcJNz303mIEWamo7p8l9/kfNzcY6A1DY8t2ZOaPpGh7yACQDNBHbwkTeN3XWVVML1ZXm0W9wdpMR
PwzHATAwhhWa4FZJqjzvRwTXCB37ozkn6G0+7prDAT2v41DEsm7mSD5NN8ea0XBtG1S4UmuGkOoM
+ajyRLtliAlEGA90qqeXhDNy5mVCdM6OPcTd/0EskAN2Yai/MkbowdZKLsPF9rcuEqldKSymkt8c
uJ3tZbkGmqtQjIoYI8B6CWF9E3JFmSUppU1xGmGtvO944KjFWnCYlk0R4DxVLADDp1SEd1DCO+WD
M6TRCd6HUMQKZqkOWsrJnrwvR8hdTitUaZuWXE7ixvD1QERjhsVSNDf9c3FfBvvujf99LWIiwU+N
UEjLOc9fbOy/Q6L3xnDjoA93ObAbgmzqRDVqCVeoiok2kdvQV6Cks8UfLhzvIpNrYR+WhhnZ2fNZ
Kkws8w+AAetLMx9CaXP8MQAH8HLkSf2nYvelV12RY/X14ADACkGKDWt+kB5doIYn7RTdpYFk9kPu
lDUgFIZgpXCcAhTPji4SpYkbeZxKPN8OSq55sMDvaxugBklxkNNG9DYCXvWHy9qwllbjTE0lYWay
93ozGuUoGT+vn3Y1YafGdun9vbWlj6gOTDWDzU2Irz/RqzuA0fLV1ue8qamOVDVTtYpiAtnBsGEq
hiuGJ1pXiB+xW5/nN1SABgtNJ4nyWhr8UTRxv62sKjE7ux5aW4BD/u5+4267bfGyHrvKlFGeEDvw
PSBYLjGWJ3bkyjiVhySDDCCoW6afkTHLk2JOTLtcGhjejvu72Muqq1kgnFDJIwc3Cdq4NsCqrWpD
LEuBMw59+B5RjCkuBMmeYvJqMUzHJTKWG4R/s89mwTCc5FnkXtYlFn36/qrAzTrYkMEgeCTX9vXh
SeLnqPHO2/ekxR2BbpmHP1UtKYSCia7sGxnzGe1a33UJAfWReFIm5iy8yKIBH+OAJDS/gSrhV7hy
yo1coivBE9X3ZF7SSGSFBQTXvmuLOfe2T7pM9zz1P24El7bY6TRBoO8r8iPoB7AJJRvTUB8ISftF
rKymDP7zZHgBZfbUA/ycZ5h5PjCM80nWYB0QfNBt4wd5CMmouV16JWevJ9J1ywPd8q093x5QH/4c
F3fb2mzblVS+iSbtdkfTgotDX0bPbDNKS+T8g8z6pxI1uV61/ANvooS75tq98Rg+wUuSSMTcX4TD
kpE6hhZi0cR1zGjK0Z/dNCLsN5AIlqz7eRSmUiiAOpe6ukEiAhmyNGh+JyZpbd6LAD8u8tAv0jJp
YqLiVYZp2JYWkfsfi+QXgRLlFJw3itKLfcs27EWjpnlmKgkutck39RJ6XoVmmOJDHLQRXp8RE/H2
kDPxJzJjiyRqw2UQz6A+nNGpaso9by+FnfsTO3r9amnfOLqq+vNYJALc4quwKnkLCOlQU8tzZhxV
RTjPYH9Wr3b2JPIdJm2CxqWsmrzhzbRGh1J+QVAN1WHUJ8vFmQK/PYtiUZdW3t8HpIAiMtgzkalN
+Zlc4mmji0A04hAq5QalDTukcQZ5deJsALJAapI8DK5EaepvsPMkcxq6QHY6GlUkQoEVLS+1Cs0F
wgpPA00ju6qoaVjJPMW8KUtKThX/dyYCP8bxm18QxhpAWYdVD2oDHaZoDmuEVeZDwPbyo66uFqPC
8cwTg1264MIQKr/y8utK6TLSVFd4W0i8ElHKrp6fKSXGyUZUXdyODiJPj2tzLbESj2Ub9RWbJmOK
QZBTj4KSLB6p6FQATtjcgZ27r4o7f3cWIrO0l+vAzcTZzRS1SyxgCi1KXRVJyqFMshw1MpcM8KCv
oc4Xb7Df42i03R+XWfJfZfh+iCJ4wVYsqFFMpwZWrKgEkrml2BkXq+h7xFe5+CW9gTAk5Y/54pmi
GXs3NCeSMaPXfMRagDLBsQeDDYCcFqM3XJUJJ8vZOOOlOxUi3TOX3RInML2T98/G2X+kB94YrrXn
SDmYV0W1hnX6ciyj6ntHZ6qETnID+mf72pVpm5fM2G4CFdnj2rpXo2s5xsyRhyJR2OICK8L3WLu8
P3U4bn1VltD45q53AWpQ42lNkRPCCYKxQii2xYOl6mV6KcwIWMs8vOVuT0hMM4asTnr76Ji8Itt+
U0raEzqHDGRRsyDNsRmoge+amjop7+inHV3V83JfRiGdCV60gkMa5o/w7NEH+krUpbDyBmzNgAG0
/8c0Hl8/lXvSA2i6u1DewcQnCVHUQluuZhaxtVgwBf5DuQNHqNo5lIU88Omj2eLq9eANs+33BYin
5fWQgLsPP+MY9OYkNT7dNjWUWZ5QPtqOLE0KE09VRkT6siXexq7LPeTKrboXfy/WdT9OUAsgHwMA
XhDdYM7EeRT50XNpXz4ejfq6cU8E7YPtjW48IQSwlSwjPwD9tsAJiFovUBcMRiE9sSF5MQokLK1x
ZPHUPOUqwVHHdss5/rndDZKm0iOv9w2NAB/7FbIjxLSnqlXbXueT6E9nWfsKAbr06ISQ8dMKb0Nd
eQsXyiTeFRRA1BbvVkMrvnEVoxCh/P3EjIFn9D9ismrLYpgBrxGWIW2zy9IOPB+moJfjlUSufG1S
JH+0+MXdQlSVR57fHFCJm/F+ziH7dUCMvY0L4aQ4Z7hfZb/xwkY8IUZQHxsoZ8Tmen1Et0J7b/Ap
1ybPXfs6HbVhcce+g1ZRUMcBlasWTMdIk49mLqR+smFAfmGGmqJ72zZkpGDC1iXCbyKH/YA6VWYg
Y9wR0GPBMP/P/hA3Lhsh4nBn+RI6wd4udF0MVkLqS+feOwajkQ+1TJZi4KPDb4MujJGjxSKqI9+J
hEr3LDKs7fJj3gqMQnO5wfB/Je29P65fsBrcNmaJVilFFhOONRXzqYBxWF4Rt0ENz82l+ljdK/9T
zmwwro13KFnJsDvtyfXY4jzowQ7CvKR9QMwpTvYBo/9OLvHqBNKFB0XFfeMPwyBIZ8C9KCc4eB9H
jj2ZhUqJv1SO1s24HZ6/YBwW7pBODJMgNdZ2MZyVYq276jMcSx+7vJ5PwmDV3gbG40lDZLuq5k+m
xK7BlHU5QImk30No9kjNhlLwyfhmLaOUMRReNzhO5h7HP8EX0ZfGBZP11fc858kFkSU48wUld3wk
PdcbIPosTTFH7rEF3ldC+tHhXQy3f6n6FFfNbK7B5rLYHjRzVEWQ0DAz2I0OMimAs26Fy+FGKiqo
VJqxyA8HjWObztT4vxYWumlyQUE9f6wMZk/K8k+21RmAyoS17F670spYhRKrwzPLLtx0n/uisCjM
BrTTSkyYGndq8aEght59GMl9dhDnONcb2cMQTbJn2sQUYknN+pGeenEns2bYWoPSf0cgoUqFvcC7
SzpI15nT1wSohsPHzzOESRGarYBBmGCHzOXftKBTIJYUhBfl+n8G1oUjBvLGt++TB+YTBahxEfMT
eshaRssXnisukTdg+DNjDwYBbdrb6s4Ji9Qkoxt4+0IRVNytqO3IW5qrgf1i+JdxDKRG9SYi0QIi
iEZH6MHhmtvwXoUstqh4LdQTH8ocs/vJ6oCpYDshCl7FhdGzCskRyLGLxNw43oW3cgjv+kHWGdHt
Ans4NnQqriCXNGRmgQKubas56mLmbrY1JEM+28nG3bT7vrvkxjBwcBm+F1Fka/iaG+tNpblGg7W1
SkJJB3kBf5iPZQHmP5UnLPXquKWZ8x2+sI05rg9XqDd4iNcMzcYG7zRxaLL10drVK0iD/WqUTgLA
loFYZBQbtRaV4oEi9a/s/xFhqABBDbuqmZHRkG/nVXSKOnka5fMd+p2RKjzAHywmsVfxuMomXXvN
fBm6XvMnCQTLBUsENj8SEsl7Q/MvS03sgaB61nmK11GVUkI8AFQSWDkNaqxJxWgjWt5Q1+khCko/
9vB21ZMU8RzLGxtEh2HpVYttyEEBi6wLtyzPWiXdW84aJEW9UaiooI/uXRF+Gq5a4i0pOFxa5HNV
fFbaUVY+ZrIm0jFmwWukR+gvs+QycEESmxnMUcTnfKstgcCYIE7mcmPfsjNtKntEOlVKGWsUo9GJ
s6+oM6APiqkXZR1Tp4ovPQqfoTTrvei2YdDKg12xAd7SXlltKAzyu+BXSRntgDsNc3bRQ+JLtfAh
YSUBYDNvbLGdAY+HUpUN4H6mZb5rczwSAHP6LmmWnwrhPEvNjlGRpBVYsgn0updZbkiM9haD08hE
4TmYeRcMb9sJMA6r8KUFxHBdwUG2oHR3CVkVFNt+jmRkE0eupUEd/sHiNLrwdUAAbwQ4xjzWNJUR
KCnxW0Sss32cb+JPtSmH10eMsA87SHYIRI1Fty5GduvUV0+UJjM83JmLfVLkXhXRFg65WyGXqJhy
HnIpZ1XCsJn73eZdsh0QqQt7huRb8hRoniiQKTFjQnG1GBQpjKeSFfnsVPzdQpLjfEu6pI3cSlA3
mXGnU+Kxto5b+2igdXHKqCflnPdndBgeOg6/czEpuUOezoEtwAFlC+BiLkIVF9swBm7Jh1EwSRBz
uKgdFzxzt8JGfLTeeda9nugmq1EkLXlSGMY4sV6a2xLljJn4PGiHkAdg8MyB5G00uiQLDkc3CUpn
VwM9ZYd/AjLT79R3DUOJiU0INrN3/7isUL/zYyk3YtgtygG7B5TBQW6CO0iemZCGBN8bRa7b+nBY
LTM+p93Z34buLBOCo3L52gq/m9t4+XJV/hPMb7fDAx2jyfmeLYSS3n00YBAYJ6Du99qx6o6Kascg
QF3JbkVE4BA0coQUzUtdyC+PNiysy+ipFTdfkJ1kLwXUdxJzhLTTVYuTZs8lct7jFyJimCBgPmjt
y2hE6Cjhf0YtfeI6wQL/qnm7TC0IbdU0nzY6cqyTUTXoVFtB5seMWU9nKdaq+lHf5/RNDJSw79+s
VIYS2diMj8T8BGzW8YjKYVse8J+O7GbCmhcyxcZGlv3caST5MAUazXSY36uIpRR3mYpEQBq1b305
VC+sGlW5k1KObLJAzbyq4/YtVnk7CHTUokkbtPhsU1hkJ9sZjnid1DJ5y/AktUJiq9Z899aYWW2u
9MNh8Q8uAlDylM3WP9VJYgpIi+UpgvasxLRYOtjTb3FxxAejy781J3zAiUgEHEwkAHyIp9/I8VYW
+oHV/ZnRq2e0X6OhO4VoOO7V1FDz++Xe1kCQG4WdOQyS/Xur9SjDdD5sSAQ+4q7jrQpIHPc6grE8
jaAQQ0mX7HHsUk9krJ61cdccwC2ubXLWq/SJNYDSMLyZ9+RL+Vz2WZH7zeO2HP/EZjQ3+MQgVt5E
yafvhk8TH4SBQC/xrdA/mp/n+MTZyWXlSO8CyfNN3qv1ATcx8R8FST1XEKLr3jRclxwED36/8bvk
pG1S77AqaJwsEAaPS69Xwn0B20ntIFYlnTA/8XgOauI8Py1OP1bTDwD8jqMM69aRX8YZ1yI1TF4o
hH/uU0qvtHzzy05P31wWZXm33tIFMeDn4gJLY+/QNC9Ka8TROL6mrogNswy5HodukjcBWn243/u9
KTk/r+J3xL6YJ4LEm88gRfrMc3gdbmcNNKDiEFMJ9Obwm6kZ2P48YamGO5Q6LBQKdI/cK/UmjOQt
4mjZShOEmw+Hbb5q9OB55lHgrTAYCfp+nS0ypIZ/FfFgl5A8WWe9lLDoISI8MemOSD/vHhB6go+b
7/OX0AuRjAbILjweaCQBySIq6mW2wMSKZd+HJo0Uzz0a9DNI+Ac+sXDy+Zzq6SGJADIBJi/NHvtc
hVxk0x/quuV0RjxgOag9VR96tERe1QEvdqJyAz21T0eTrUFit5TMO229Xp8/uRZgJCvQJ6jOShL/
NPOv1Xj0PbgzI7z12ap+gD2r0U5t90N1BVCK+ZKDkSdz3Zlf82j7LJEVxRAoouleUWXYAYgbzx4b
aFv6qRg0HUsg5FzA2g0DMvtK58Mu8fvZdnrCsmUhxNDCfxslfYI2hKaPtZ0IojWQNW+bRIk+kYnn
WoPwen5nj7MBKbwM9LEMlQrIYQLBFWh7Eo6sbhXVj9RiMQjg954bqTvINLhUyQE1k/WI7qHpMYfZ
KMkHCqaEedfm9Wnnie9ab6L7lFCmnrmp9/sL5pW222QKKxkMOpwrfLVdpics/uMfGq/FcajuwBUD
jH3ls3t9dbrslhnNd7j+ydzsrOZe3886s/7gpRYFA+xchwHAIAulGXNbcDcYFjyqh9omSmvIqKGK
pZOqqNBe5u5NIQsmEEB/3X6lQTIX/mw+d9qQIxKhGaW1TDFX+6XfWpU+fuaL1FTPiMCTTzkcvrKz
rXiQF6y7abAHOzZPDHtr7Ug4Orx7baI941niIRJQZnHuxNtS8Q5KuiHORjYnbN4KCC50sd+aoz/a
B7haoKzIJA7+AbJrdOGpsKu35zPCBzjEW7JYUEa4dGrM3KK/+Qh2ZCTgbgmB3fS8/aVxN8QAQGnQ
UsdXEy/Rz3osT85UnWIJMu7p4PXaoE164eraAazHAZy1cno4/Llag8oVtKgl1i/7JijlSJ811Ifk
js69Dd2T5ly8houzFbQDUQCQDSpVzL/D8a84uhrfjD/HpexkXS6NxmsPIizWPI2itYH6QToEPdN3
0Y9l14cApvztKMNB3FqHv+8gMsmknI+2oluNFA3M0MOY9lG7GxoAaCmKPQl7aWtAO0EeXNvoGl80
Rm1sMxpTkxWU3YjnGOerzAiI6gGEgjDy6K7WUXfjg6a0pPr0qumMyOLQmTwwuajWcjFnBJiSGtJs
k3GLJn7wSG8LLseqsHoOAkPbeBxSY0V/xAPhywKa0AFAvvcowNlblPaeqFNieb8tcjPn66yYqFPj
GCDKJJCI5YjizLH765kf7a8LbJLuniPCa3rNj9F9nwVf66KmK4nEtldf1UMOqHxa3HOFCuFU/DQI
jGlvgiASKTd0tN7ziAcAdR1JHX1BB2bC0eMlxiOXp7V575MFugnjzEfxcSzejq3wC/mkUimX2Dw1
03BhffJkS8Ha2NDZl3JahwBZy9iKp6W6MRqtLxRkuowGpUna4FBWY9fSR7xbCj+87g5ROW0qaK8v
ckhf1han15w58eK9mlFEa4kREPTxvHqa5/FBQ4/0nAIPRGbsqQ9MUuXpIda751S2yyKG/yi1O20b
VYAuOk9mzBJvPuiO8OkK3xYsGg+3Ypq0/spsSDxTWABuKBKXmSDXQ6MSwatgHzOlNBy2Zb1KVObm
siUX5HyrQnIOs4ouUj5yrXIEob1Mt/2pTeV610sqbcaJsaZvVXsofJ+Bsi5KMsmMY/Yca2k0k4Tg
1U55/g3zaMEqEtMkboseU59SH4QuK61OWDjeOCWuzRR4zMTuel2+ofxdTJjQrBlDVCZjkP4zzwgf
3aqYkLp/BbnBLS6JeQ/yMRnn/hoCsxS/6ht6Ckdd1l2WmroiNDsd2ITn1g0NFzgX4KxFad4O3pT6
7qnyEaaMIqeCse8DjQSv3R5nagjz+yIhm9tZEiRqQyZhUi91M8SZ6Kbnhl11OcuGH1lpkj7jM3om
M6OpLu1af7Si9sniMPO6XvZqG2X6EBjkOw+TSerrGPI7Bee6CM4sSP6NAM/Dw2rIVZsixBQnuPvk
JNsOVl8Ti2gF4DcAiIVJFTzo0VHhSiyJ2MpGzFhndlsBS+bI7hRDPA3LPwuojQ9XhZtoJ78pW3sG
OwOE0WqQP5BIdm6fY7k3lVU78jRYKKni54YJuoeuk+EkRpwdcIdLAHZCZNeAZyUqt/BWd/TMAMBv
+nnMstC6c7OnH2/M/g9wbQy5S0U4/Zd2BpQ3i0GMijxThVmQ09KRuodwDrWY4rvVLWA+0dPtUCg7
mtBNAWcBmtJLw3N+r2WTt+F0FnfBpUGE7P1sPG4YfjBrY0Qct2OOCl/6GBoo81XzxvY1lL3mXsyi
OKGaKI4uzqZBc8ryulaExdxcMDWYQDHD73i69kh2dW/WTepcIhc2sb+mtnqQbs5JaBAGZl5nYRni
DmUx6BWQdSSofkFgn1cGjBgPBScWSfUqkm/+C1K3XNxb1Gpq62ZYm42yEhbPPpvZj4oQeaLUoVWM
RXXXI9vuwcHdFnldsq02wiut5ZHaeMtCTqhDA8ZgQrEmCPwPyqKq6jUxKbCaRJuXZiUnrYPy/L5v
EYgJyEmTJklWnLv8R5yXgW7MHdsK/rtca+2tN+ZmWObAXWkS6NVN6UnENxep/nZafKuwnO8yWWU2
5pI3j51DD2lNW85sT+4N2OYxIwIWvKI6qwpFxJ0qen/m+dJjz5Op0I1+RLR7gngm6GahswQAFGaN
b0XASjJOYqnp87vmmLo6JSLbqIRoSGUgbDCxw3S3yYUnJEqo1zjC6rYV01SHmtLCfJQeZpIO2Hne
Xu83yhGSeFwPaBLWWAhjxeGxA5sLebgL5KdlyrglY4bQJZmyMatl3C1SYV/elvdR1pbqolyeK7Wz
NIUs1LLh7Gh/puTUvCq9s5ZNqg9bZ5yfqUeHcXPxB3shNAfzLXgXwuIWcEsx/Tk8NKtds4tEyvdc
0AOd3lRLsDUR2wpp0kofLkJHTxHpB87jmJnN1d4hqEl0t2izVu1hG67SyrQH3SZkUcY5Dhqh3ZjX
4gZ/Ri+zBkQupZpJqRJxnHGuIluf/8Blr62CvnTHWLqkJR+QCNX9IKnYAtYsN8vVSe4rIeUCY6aJ
NMjaiwK2wekah8WfaOt6M4hV//tu0HonJSnxLaWJodvseVLvZ1QXyaSQoRrbfDiFjS7Eu3yAcMFp
ckLp+43nFSs5Po/XQtTdoa8+fvGORUo4lKNJ5syRqjptbf8IdHzodw61Veaog9Jk7k4HU8Kh//Qe
VwbQsZtt+bO/yRqTSSglVzxO0PVRgsxG0NNIZNLTNST/OaZtfSe1nZlJ7lTM1iI3bymFSLAagSu2
c5b9G3uRA/MH24ZmER9HnKDzV1iLYtXphB7Zq75nHJ/63g9k4ZNypJIQ66fUWC0Yca684R0rmcaG
swYLgS9Oj4diQVbmNuh+gfOpTThSBfgK68jt6ckY6/+9fESY8bsRiq7VCzCAsDOZ5koG7CEy7dLj
y0p0sSmd8GXVl9637SlAhXYBaZtwZh9Auj9wTVShCFeCSdNiy4M5qzwYycvADWTnCl1fVfKORLPg
zygouusHyZ2SmiKKpyq6HFHG9HD9hEWWnoZUzHxbqdXzhQ+Wq8fqxqKUIveIH347z2hHesydLBrA
F91kFUMZtEECSTe63TbIbAZVZiT6Ubce3w6O8A9q2pGqf2jDP+e632w+mUdCWnwXiUNItgmjscp4
cC7dUd1EU9c1VNP6F1Gdwd+0dzecqhCFIDBkZG2CVjMdnpidMIVoVHxrmUJFlULGYVhu+FG+6CpZ
Yd97aWTDIjJm0P35h8WNcPw5+f3vuWBHbczAjaLKWaMm0mLzdh6sQPuQWJCLOLhShhb/dwWslB9u
eRSrDCQ7dNfBqAVVwHQW8lAXksdDV1/4I+lYMxtUSXQRsBShFUIazDon0jIIHVYrreTG9/f4ENdW
MmK4tiHCqNXeJepuYflqe3d3rk+pHZLRRkw/mDM8YhzRoCHYYkilqEjfrK8qTFZy4VRjYcQsH9Hn
Jtx9BfiN8fMjXXCrRLjERL1Q6/g1c8kQj3j3IzzxbsDvqrGM/jmhTgI/a2Evzm8jHA6LZIh4no2H
xe0nh7SBeS4pRuFBNSRu0iKLUY3+xAUv/xiUbmUM6VVbk6TNSJrxS2ROhCJiWXt5ts34uLl/OpDZ
5PX1098fYnS2PUyV0GrZlseXsdlG+ikBgYALpmJ64pod1IZ94YyXnCYibU2WP15mMowbJr0EUPyU
OgN0QfhFSeqtUNVTFghcAEMvUzq3wQY7myLv39VufoJh2/RE8ib4HrN1hTIi19zeWpOC+3nd2rlF
Ljy4kLa2HmBendUqSh9czbJziU9w6fdrhRDDuGSVoAG1RKW8GapgHLViZ2Pzegq7p/xemPutjYjD
dVlRoHPvx5eimK5cTl+JMhPhrh63pKqM/BTgyW9a77NYkaLO0Q1m1EwpPSLR8qqVF8TrKeV+ykx+
VkZjGh7dZ/4cb8M2a7vOpK7HC9+uM4lpTkSbHpmqgGu13a2DzzUg0S9+ZLw8UhfZWGYXIOxr7Qpp
WaT9uYqXnCLp8tagq1SdR8Gze+7gl+f2I9lv1bxDxct3+hcvywb7yjPpp2BFGut/HMHNv72MZoad
5XK7TZVjy5FWsZojnnpiGFX9vjwmMBMDcdqvROnMS+hXQEVWswHhID8MZNEutQ7WNG+vIx5IImLp
4NaQHKVK2IL/Sivu47Zxq9NMbtzisLLIVpkIJFP+jTD2byB03/+31xm5OeUSfhqRmJsiwxpQbAem
puqOKE7rgRcnGYBGIyB4c+JjQApG7IRv7OFolMiVbJhE/65LGhMc9YcAdttgyn52EYUZpnv9IJ4w
ShKMQJNCZEoMaEb8LbbknuEtdbNJjP0PPF2syQNrAMmuoA/7fmCk7d3/+5eYkz1VWyq9Sf57dg31
2/vlCvyc71OzuzIHo1Huzy6P0667xmc5anxadGLegswUU+NPhp9HcaC/5kVEwtcNJ2iFz3n4fmWH
tC/RtwwgWAhbggyOZL9K09JR9prsByN0aTvfF2/mQEk+1uy7E5WT/aaDWx0iFLgR0ub4w1PD7Agc
a59+4xXiwZaMpl5+WYzJkqM9VkY9MU4l7NC+KcT8o4h1GFyd2eibNUWWkxn2KhpWgki/Aya1fBax
tGe1wLNIaPH/7ClfdqcQPvOLGd0VXjP8sshocFWVnSE13AHED7y9sdjAYxsAOaxrBVgMynNgJQht
JkzWzFTA/C1HU0Ue1gUb8btui15f4ce7qBDz66vcy1fsYi6FG96GBm0kUVOiuUhG+GSaoSmk8/gx
D1EoHWfBY8AFEul9u/xb6sNx/iV1y2yvxt+a5ZPpDMDHU0KF4BLsWxyL9DVFLXHez/MdhHwjEwol
mOJuj+mlIX8Q/GpuhqQAZTydHEHQohUKpr7rC2yQ1dMS9XoP0XtjhMM80pymCYshZn62lsBkDEa2
qJECs8V/uMvZQJS4iStbL7QPqZXdnMI6wkm+XhEu54uTmfhi5Knbv+1E9MQEpIQgfYgu7GpA2obh
ujg7WlGBGyaZX2kd1ecdfYMV6YIkXXfc7FC2+akA6p6eX5CbDdbWGWW9gTsBib81m44WesETpqJS
PGCNAqADcdReYrt6+FEm2zdcyARnr0iAhybA+vJ62Q6VhzZEm0CIU2ZAaxkVxIJuQ6U94ys5vhp9
hE3ExfvDYT61J35Uq93BTyTlFw+DijHASz+Ji1hHnGXkMp0La8WkpycZgTLyG8MPXrjms/UOwuAZ
MjrMhiWwxHMtcMm966FXs0NPmlUPnQFHh6utfJcx4PXGfJpsLXA8o4Lvwgpw3XqvZPaFln974vKT
3a5S5qgLZjqbFVT7nJzcNg2tVLJ6dkWL7zNua8cIvKy301c1yryGO6fIPjmCjf1OlhOu7jJDLBrK
TItq40UeAb4pcUsyldLBY9DpCqj2fI6mnBn0ZUIZXg/d8B3ShGPrcgA7LhrpzQa+8MrUgMX0Hxip
wWISSEOtvIY9JlxrI3x/TSgzH9sVQaiTShzw9Fl/iBNAPNAzoNcgVX3tOUDzsxBeePln2YEXBvh9
3aqCCgdODuTzCGhOpJwxjA1WIdkYeqH41x7YKqiOIT0D62fsGU2Zg5tBZoiprsH8e9Xm6lEpNon+
MyO0s92iXiA++tM/1TiGrimgahP7y8RWPtL2RIoINvxSUzXwG6k8MSOK83lplHp9pZI51QWzev/k
h7/FOjU/6Afb/Ha4jxqWjcQvyAt0LTF79KOlleqVbMailIcJ5DJ8mX9wIJ9Bu00Q2Y9jRPWoz4pD
Mq4eRciPTMy1j1QsGENYPMZ62JeFV+zJ6ALigoh8lD1RLrWiz+/p+lgPEBK+mlBmygRTUN7uuMLf
VcxCwxanfBHAxTOpNNkNeg/GJpm/mJ3MqvUe52zLvgnSRe64QcdQ3HMM7B4Wh2oCGI+wz9zKICLW
X79TXN23iesPGd8LVYwvZ8Ai68nj9a2LLRQeFRHN6naAUgIWc+47HVReuRopkp81adtYepCQw7Qt
lFRf+sQbkhI6ulLiLHo3d/KAAthfnilmKU0e+yLe8Hs8X9QwrZ8xqt2TU8xrC4dZ8NW39gPbwUv1
43/HWEEQA7Jm7VJtCWTbRdwCl7Xymyl8adApeM9aUEadHx9/jI2UyWy0xwwwMPMbUrYWT6s1Cc9z
pVLCqrT1FN0U8k4CNFakwT+CRMMCzJkeKW7t4qcM9n5uSUYDnPNuqsdpDuWfJAO6xa9l/3g5g7AY
/AZZ+8cckYo69KP6p7AkCZYgktD3Zrg1l6v9XPCgraLB9YtkO6ywxVyUNiqcPZX8DA4nl8Eqsr5G
XBO6DPlkXYBaUp7CEzA4pLWIcbeENc9BInU5uyFq6bxk2r7X97D+uObcS5R1/QONYVtaKog2RCEM
/GOBO4rGz3SRYpSHmKwejzHN23GTh8ezW0vBJsaH5iW+neCrdh3axzzvPIi6KH6HcSsscFQWQxVR
PZ9FGFZjy9YOn7C43Jc9e4zlR/1Zkp0yt1GUBGb9Bhs+z85ZYtrv/xMC1jqjRloiMnt1zN8hDogW
/N1nZqqquIF0DAjbtGIj26o/yZoGSdgbwfW4+q6OfnWNS27F5rGuAkP7Ot04lzfWzsatwM9B56jP
lHXmjLRtd+Z6fZBWoIUBr3871L3sI4/4xbP7OVuLxL3IInFM0LPrEYWvQJXvaH9qDJtCFhnJZ5ci
GQLelULPX8VmVs8r95vljlhUVvFJczlCZB2csTlm0in8eKYsmsfHUiUdIRxJ39FzulH+X/hF429K
3Jg8ZplJumpgxeOw1nbEnqbl0G5sAuqzdl18Gvn/9c9t50g3yvdTlLUwQfDPVVuP9Eoj9UZZvJNw
aDkIvN5MxfIz8zx/5Z4zOSjaCU3lMZ1QyPirPlArXIsyqTOQ1oNbwxUHXHqBDLZyu/Ff1aVbS6QP
R88ICI7TCtgcT3TEehTnvYIpPTvzudy2pD+l+figjh3ZcOGs9uwVB1tg1+YzD9ivZ/W7B4GTCgxg
Ow/RzkYtpahzW3b/gSbu5svC7OvDJfBGcyTWdBYa2U0ltGNnB/gQDCDIjao1hL/jpuIJX5soHchx
zwluSU4y89azoqFQfbKKGAIX4cEMNFHG3VRKqRkdynaqT6UsnveRWMBCnozeiAJx2vOdz6dKp7o2
RR37frw1L1C7WHO1JUEqiIDGs7wwbhgXOKedzA1XZRBYtzzfweTrwPGj3gA3SyGiiKCyzoJH1cV2
r+lGq25nCl0tshXuJJkeI3sjkd4XIZSXhv91B7j8lJRnQq85y22IOi0hwRGUHtdNsD2Ihn1aRmZX
w7i7VARs7fRQ4P68LNi5ef4ycULF2mXygzitExacVCK2cdTIbEOKzx51U3adiGikxabQA2yTwPC+
MxFWMpa3uHie3TxmLZ9ZM21o3ZdYpceUSUzn+krpRZ3TDMih1S51eN68BModpdUtZxJnyfEZswbT
QWNgKxBYNNOq2Zy3GEHLMwGsmOOfYf1nkJgeZAhe3oQPFZxa1p0R+4USNYb4PrNLdhMLfgvw5M4I
Z8+2X4zxfY9p+vpCS/eaQwSBBvxb/byMb5ps6Pa83qTH7ZFR1e6PdLZ8BM8a+TZS3zR1b/wW0JNb
ZtZhYvA07GWTcggw4xS9ZYqCkxbUZBK6x3gxo4NKgDBCmYIaQben1anL3HWbRmpg6mUwA4Bq7195
a2TDyzJdVhEL43h38YktVrHUivhiTVgrmo54YFM4EvuIGoSO2pSLdgBr5VqXobAHudFgtOCsjXy4
hHteOfAQddudyBFj7UHHJdzvGSx9qlQ2EHz4JLUybf2eeX7hREVS+d7kFuciEUI7xbDBM0XpxS8Y
3ICrNX9uLBlRd9l7ejLh4ACvwM9QpV6dq/iwtUBLhMg1HkiXtcoh25TU7G2InYI1pBJ9NsKiq0QY
AWRD0kNSD3+irFgWiPAdBDrjoSQOjYVLzKHVZ6d8ywyiHgbgVumPoLR9WN1tY7upSXYsX8viuDNs
JSg0Nic04m9EcafhPtkkr3tg5GTsyZZEPK8ohskFRmvU3FnkN5U2gu8LuQeqSA1P+S5gfdAOyQco
Bv7CYhEGHnGxWU/Y6QVjSiN0pzSC7zwA539qGpj5S/ogQdKJpAtyEs4JIxck+RceMFuTS6aeXCyL
ykGqagQNev95zdAI4aZ+fikTGYAlfyZFZVMVAT7mYSvJGwKGCVrHRF7W01Es09AdmnNhLfZGD6ut
aoP7K2MhyhxCqyV90qlVPVqLwFVtnNqW36a5gTqPpV+VviW+2QcZXy7EOgKMMmcUsiB9yXN8IG6P
9KxACVn+cLO0efC6gw6VTaVfrPGDcvAerEb8rL0WYGO2kijtxjv8HHH2gBvCbC+zzhrTiLH8Qy84
GY/dHcozQqbviKsr/2tePPq6L7kBOlQLq3MzlnWWE969izFszqPt44phcW3RYRKWnsNbLGGPU1ep
nMEOeW2Z40VDcRfD5Ru9htGny56HZrJrDSDCdZF3Hi9xdTuixf0Pg69DCb64VcTm4Je4xgcgwAnC
l79DXOHcxYpeOH0RtHdw/fHvC0qBEW4WWq+buvdwgjBzbavNRXGbGr9qToV+xUVlcY5sewN0tmmz
XpwOzLL/7gqyMBpQFefJevzWF/cw3nMZoBYPgWDDBa7JlPeiFXTvkM7XN4f3sxtdtvYAtGq40GVg
c/O8eVqBsx4kXe45v+B01v/zR93B/EDGEtS02AnaMrbC4Q3AYdr9hdoy1GRjmL3t3JuzBvagGof7
u2bvau0pMH769U/3iGk8M17A75HLVY1dXN7MZrkl8I4rgmAjkGncSD7j64XaAYSo1Bi94eBXyzX3
HVlB4cMh4wsvsNRfz7dWSQGKS9dxRWGqRHkcKeVoSKOxPuiF7ssvB4uneHrABOIi0EpHvNTF8vu9
f3PFn/tieJ9fcMQ3jmq8wlYTj+z8xI80e17JhUC/ALgxMYT5Da8Ki3K6HK1M6OiIM34cc+joTAKR
T8ZROw88lDlAOy1s5cnTETTzFdZNbo2BbK0i7cAmNjQWPVHcmc6yXtKtgPQdv9NJPVLI0ZYcBqTv
aj+jjb/L4ZiamxfXv8OVY/38RT0kpu482yRgWydfiTKJ3uHCpH8qUfaMHTLwEsKSJfyXKmpH4maU
EjznV+JixKWfxJXvU/kq3JijAC3gfS41yAMTAmQj0hd1QeF53XTH8pYl7Qx5piimYO0Nh35+QWp+
U6VnkozOMbMFNNcw3hcGJK0zBV80I89cJxyp31YmlLql/IWCKR03cwHAzPb6zlpssMXjOrddyS+K
1PJs3tJp2oRwbD/5/1II1tsfeQj7yS5BfedbM/dwfX0fwlJplbUdWSuJdaFO5rNeovdmRXsvYp3Z
EpVWlIPHsxn2wrAVUdaB9YTWzFnh5vIgnfWqd0L/56DSXwKV/3ue0xND69r6oVtiuL+/DkaBQ2FA
h4eu2g9YSDCNsSOUWoTF7UqX3KUVxWNBnf9Mu2BH+yyNBhEiLEBI0sZkw6adGEoeVVdLu+nfmB84
3Xajp4m+zYM7kJ9JpyJ1VshVqvSoN/z4gCFA/EOhl7tEpo/Zi/lH5VDtruM3rsWDP4ZlPLjcbwEr
q8rTLzKdzyfMXuYStTeXwnjSLS31i98Olmo+j46n26lWkyCN4NWRX5hRJp7xC+NZTq7QMWrwQqXj
A7CRbgHVq6KpvU/RGlJvGC5S6+ggqPHwwt94eCnyw6SykebhHB/cCHLXkrPcPOL841b7H7VuY/3J
BqmUHamXIlxQvfGTOU8noYPSRkHw1zN6+K2+QFfTOxtW2woPur4FQzhqOQOH1mRpLkDDpy3fJmQX
7/Or6lVvBwQbhxL17sNFwEIc5YoZ5zZA6T4KnqZAMGYOF+ZZZIRoK8Coc4zR3P5mPjDw966npbz7
MSdLKpB5CAX1R1riHmqAwUzLNaxAOcVJz3dQFHKdwQaowyVkshMOZ2i2kmyJDuwquNpwXWtm7Emx
IDwqsIT3VEAubYgELJynsFDK/ltPHFkQGhuloNfc2aurgo0kjd95HyIm9Bn+4xfQY/wVBeDkn/fG
7FC/uXOGLwsb9ENeRTiHalV358YChFdVHHKfNhQqc+GpeA5/ZFrM4uwlfT843zI5TyTVwB4Lvojr
lIY5A6UlcQr39eZYbNol9nZPF0Lcnd/rIMLCk17QsVeJCc/gHKIqd3hA2QGxnGDctGz6drK+ABn6
OhPJ5D3mU/ka0F031SxiaoypqQ235iqaw+dw6I4tCty1Gy1tYR9MDVUk1FzyIY8T/n7vFjHfgfiT
sXjxjo0J1XpZL4bz6rgHyXCK5lfpX2sDgzAOwhnzpbYgecCQgtkFFyNSUT24ElkG7tIv5XEDerPi
vjMZ9GwQCPK9OcVgQJwt8s5Qge2wxoTw6RslFGp0KkzZYDFqT2cDXGHy39qZvsTzm1keoX6GHzLG
j4ldzd8L87A7zYGfe9xiHneuiY/rta18IlB9KHJr18YNDYLT/W7fttCm/XUmMAJ8o8k4c0EAjFT2
8JXbC7OO80SYhIOS+ig+AT4BNx5uK0U6fmFlzLTsFj/Hy1Mg4O2K21TYIqL6PhSDmOurWLZAD9mA
p+zkpiNr3iox9we/529mvk7aa1VwdAYzRiDhDXKzFjnrvDb+C0GQuMF6PMjjuWANkiOUyQtQDULR
tA/VPQ4BsAfWGGwL6+hSguveVxj+IiIqDr3JztEzL63gfQY+RflTQxQgjp5qGgde4LgsGkLFVPy7
S6g2XF4KSr+FbMgM1QZUgbc8fPosyk7E3ZbhWX5vg1iZouHjJAgwA88FK4dOJmShm7RZPECE1H27
4sMa1Q+CMKXOdexRnyg3KMPVvJ+4MaV4CXzJg7Wk4S55b/8vWDucABUYE/13G/jYEI2oij30qj1H
NnexyZGzWBNEbUs0WuCOqJYJ/BrMP9a3JfIGW7SdVEDKPY9HB70WXXb1GWrNManxuzNN9gUEGlrN
SHk16pWdbyBKLY/SsSf8t4ieR3J0BEbT1c2GZkY+XrDa/w6dk8ziUd2az0aZFlTOeeWUFHX3e2Bp
3zSr3HTcveojNtP1h6chZKLlPeyGUSiXq7qUKP923vdc2Il3yTL4U8p26mqXJvajXR6/EWVNZMCn
E1RMt6CHGwot6xu7Prw1JnQWNBGEsSX5gmATPSZiDOdIRMzPK6bMxiljSgPDCoHO6nMPKwzGjUIK
gVTb4jvrYfEhM54Y3iEwK7Uig44UEwiHL9V/U+t7GkyN0ZwVPGz0AI11fMPfQmKdDsgwPcHet8Ku
HiD7zxYsm4lK1D63iyD+b+oV8v7DMcFHLD7bEq0m5tK7T9PHKhvuWmMGrt0cF2e8k7N0VMvpmAGj
o+WznkslQSSLqCCgQyzzPV7blFFZJvBAn2HUDxPrSYSeAgDY/9fGW07WlBNk+CxRc7hqlszbdDMt
2dwiSAO5LGYWuQi0fisOrk+ruSBS3xD4cORMGgiS1/9o9ZL5lVTrPqxtwqBx3KFo4nY9mq4kKa5t
oPrp9JGOxnvxm5kTL4KJ2FS4rehQDUfXYIqz4QVhHSxeSNWbLM1PaF8qs6wKGVKlxCgxU07IT7zb
65DUo7tmPXxNzauSchIjIHXN/6DIMaGKXZNFnXuCUPesxZqDgGObeFthOpnGMGpphhZP5CfHZM9O
fDE3cgxLmW3LzSQZJbl3bVcu3z+rS5nmCabMfshU3nvAxtKtwRYDqfzHcJrAOvTfVmwfPizZKmYR
hl0MavLXWTuXBXUTgTuEG220OjlaoAxcytcXZf3Amr7AH7xghfgpDW3XRL5f3mq4S8KZaJFzQmr5
TGg8OBllO4qVXdzIcapyYk4gPpiiSox+/eKfKFjGrwgt4kr4laxJ4pSL85WbM/w0jrAYFmFMboO3
uRuxmgwngaTFfFBSAxEcYJoTNGfbm9WaGXTEgpJkIcUjSvl0pJEJKAAHHcaI81N4SZS2iQFqWDH9
dOO4YTBjD90P1BdBOQ15HZcwE+zpgKxY4WdaIVNCN7nc7otV3gF+LCYgGek2CB0F7gouEevY2fkk
dNKDWy9fuOsCUTaoz8gwk5LCI3MKEDHD0iW+A1dly9T89tmXM9OsMx1naUwma1ydvZfMokrKIBiD
i2zNdKkyf6ns+ay0U/kIT7I9rqDNmst0535F4dgba2cayeruCqLtlSczJ+oq/O6y+XXSvaaH66mu
3Ii1Ci3jA8XrlBwCLD26EDlQUC/UdRDmlMHLuxulojtlAniLUALLsQDILFnsiP8V8rXCwbgxKYfX
e0lkw879DrbPOWYS5eT+TpyyIooN9CpiF7Y+3c68F3auNx5zNM3i1ZmdrU5xwf3uIt7xIFZyHZpd
XKVh/M3nQ1sP3YYqeEVhFKgN18afX7rdHTfBsNe8M5RS8K53D3KoTJCpd4Prk26V/NFapegLpuGw
tk7FkqVkR1I2AsiidZO8kDywBeZNq7DTJYvxC04Pi1LmAfDYtwBOiENBySdSaMMH7bRGiIv8pDWq
7LXorWe/EFIv4UKUmEci1lukIf2Fk7r1ByEyg8x23XenwxqmxCKHgzvCwoiP6NQFYv9kxB9OyKzU
GJjMSas5v6JxJBJUSmka1PZicMwumV1l+4bC8qWoh17GAS3MebhAKB0g7eVcR76FfHAoWq/yOVzB
mFtt7Yi80Dor8bMkmVQYaPygxiM+gft2sN2J//Q5RS/wVoRVTcuhpQce/vpgr9GtdafwcoP6qNdJ
afIKRaYh3UCItya5HaP2bUSf6koqpFhFHA4wrxuuwjut4cmnCK62Iq4SvrOl/z9x8qo7NJomwrZP
RBMw/S19b8QZ+y0Y85ytxV05D0Th7T4wAMrTtp/fi6t+mozv/223JLcdd6b5PfYMYiWEmxM9PZkL
GMd1ZR+e9wMJns1/9QUljVTJGcOTwabatjBzoSibqvatlYpgeRBxTsYQuEtu+eiRDbRKEAhUu814
27HRElLARIirGPSfyS9V7Cpzx/2YsviunwWm0H5CpFO1a1Im194e8mndjsqEFXXKb0xAtuRjQTIb
lqS4q27M4PkwiHVvaEnBi9z2fJ1L/Fd+7p8lKBFDsDLEd4qfAH9fU70lF5I7CgxiDJctkmxJBF8/
toE5UiUdv12+jHnmlnXwAxum1d5DCS1MYg+9X3eyC21N2t4PkPSk/XK851BulyPXN1IFaFkhj4R2
2nJlIsRCZ/3ZYrcqJxgfeW0QUNUnrGsQaYmV6Vxkp4WIY3iQHn1BaaIgaZ/boENwLOgGrmELUk48
JKssmQa/3J2oxcZSq4cawka9pWqjEzmp+a8pJgA8/ZyxQslCBjG0+O/5jaV9+L+ol6DojSR4nzQY
XBS3PoQ4YWQLYvRD0z5C6+sn9AP1NTho4ZGRIXPewtlOtPADu2LvyeZKA/vi0S4Ztpgy3M8c+mce
sJNMzBmQrn6BxcoGKMBmcBH2RqrR8vjLCX/MVGECYRSNeqUwG1nMMKQ4VHVK4oPZSghA52ATgJWF
HOqxHclLgMDuUSpabqGIOSToH/BZ9F7QJKvUxLEQSV+KGcvwKkokhwRXgo+sEEfgGwEYoMLdI32z
Ml+Ffg6OGmOcHGZJh3TSWC+DXx1A0PZHqk8W3mcGDj42RA0iYj+eAuwXnxXXUGh8IgbA8UeLYJ1O
F0z40NDKjqJMPvsmCQvqQ6TUaYU2zJrOkrIftbIDeJrAHCzI0Ftm1rZFb9G7ln+9wfUZzjAUhwLb
wv230y6aA2Zcp+sb3o/wUvq3t24toz/jILVDdOOHmHOueCMqg1cxYbwtB6rHYLiR7DH+9402Afqg
ELQzDevXDZUFpolggHdUQ0Jg5jlFnA3DTpMG/0bg8g6+IVrc2AO5Sv76OMP7LxKeB2x5PmsEF61/
bRuC9E0W8SM+S8ua1ZmeVZnfKg4bAdSHCsWEN1bgmV4liZxP5AiGbC6ncp7RnkRCzcDZF9WQ0Y5S
APRyTIv6XpUFtuBXMh4Ijt63XkPadsjOXgoM6/y/jXSUExSDBR3K1H97eyORgnv9NuLga1yfA3i1
+s6yiwJ/37YZQgVBS/iXLumufmKg+emiodWBTSi/izv9s5lEhix6PfyQL2AddgLeGouV1RfAtT5L
ZZ4Mav6GM8xeM00vOJaurwOsZ5pI+LVfQXcimrSpKBOTsDDJA5qV0NjdxZY2eDTF6pEHesItMobY
9z2KK93xvx0tt8ub9073Vo5xFW+bu1NGvHzhMgGcU11gNDgXgAWB/tA2ih2yzuL+5KNuvr9ezO8L
gmYOr0fM1AfbUsOdzx2kr7WatLHY9tc7JQDuv4HevdyLgeak38FW9wKbMZbb9cQwQP5GG6inEqE1
7T2dGtqNMbCroNAG4js4LOCECrusiRGmwPky8elGwlXeNsvwdG4hoXeMazZLCfoeJ1Zz4usiPLI5
xqXDyQG8bREx2qhLJEIzv04fENSJnW4dyWtmkC8bhvDY2hYM2OHairxvi7bsTzA84Pi1UmVtopYW
PTaJUcfb9mcoAHuOOYTVvT9VqXuzS9UxZ2mkj32peEUmxfXAuTxWrYWPURsVB+mZ6Ac3anRn3p16
qGzEvo/olbRoZqjpJyf4f9ymjayub/pWCjXaXIq+LgrvhOifVMX5skheE9qBkH9IAsjrqQXIgeKI
ZnhA93Edt0uQI+yqa8wNu3eUWXGcTffEBv75mGxba68AmgV7uMsBAiyEVg3RvqrTSVx8GSaT/AP8
0JF3pSzk7AJdGOOUDQ81E01XYfW82AFkjPI01RhGH4r8FufmK25brlNIu6cGnHbK89XZGE0s260s
/35bPAjp+/aaGjhw6ckb2tlOepoEWc7KK5NLZvovtr2q8m9WPIAk6v1gi9BBSI2MYA7GE5kMZCUR
R+JSk8esHWc/VEBG17jnX9WsVI+uh3yJIJpIyomitmcIsCmWi2gSuu6PPElDEFQmZ8DJ9nvtVzyh
qojJt+tBedVXpyJHv47uQ9uXiQoaVa+CMiMyH/cU9q6qN8+dQxfGr33cTp/lwlpy5zUab/FF8BWS
semZI165T0QaEXeYGcNFEA0VZ7bztVV3Oj7sNQf+sWMFdn8AyUPFGVm4mvus4MWJKA0KfDOROIyx
46UJsJPTkgwDsYvkZ3QjeBMu8etcaSIYKQZIPPSd76hzpDNR9RtUOMpyPL6eG/kTO/CYJZ1PMkno
DVIMKG8l8Pzez06+JL1U1+Y5WTHZuWnrZv9ZXDYNsM7NIvhhf5Fm4XGYC1Lw1y/vgbUjGmoVCSto
ZkhZXQxwCh/UEyHvx4V6vkZY5HiOCQnXXRmukYEtrh+/0Fe5T8xojXzBqrHAGuuavGzcuC+4zj4D
MiJIssDosbw2mYZaeaiUEyPRCBY6iqptyicowKHQkxpjZ7gL9UBEWlmQ0JIo8ls7X1ZESGJp0l4N
DCYrEtMvPdLmKHNYHrrDKSQL+mtN/8FUyrzjHwbU/5xhbXk7U4BP/316CDQIrWiun7smR8DFU6st
EOtHVgVl6gpBp1Wp4HGTO5yuA6fb2XYeL/xpA8nsbjy5tUR4rvRZzR+j3cRTQdf2N5IhQ/eyHb1G
SKl4IJa3A2uZYkIzCKmUUZW2EHQRfM+0OHGZXAaIaDyfCWR21qMNV7UajpBpY6/YPKBEQFgkxkxN
XX9s46L9Lb6elFhRtWCGlaKDSSiaXaGmqflx0MSxt6c7ZgK3bthTKxHwMQhOlybDXDaZyPLc8WJp
DkUrAjtm2O/KBeHSu982wANSCvM2DnqH7A4VtTdlOmFopt3ga9gfjRYRopSXx1Fw9j29LKFOJ0/8
j4ip5rcWrGUJade8EX6O7Nlmes6JfnNe1HWYUP270PBAOkP9nN4xklBay7u++XfohBFf6cboRSDE
siww16PiJ+L16ahM+4UIJzu3tXnWSYcf15ASFDL6GYjXqN8hmlhKyd+qDftseGXTWmdmmLkicYe/
DEps/rccQ1IR+htHYAEXPDgWnmSSgaU26BGyDNP7zTjoIc+aZuR8kkd6HUppUl+D/qhbNQOPuDzl
v+GgGQOIJykOhAhch4nChJjbL/d3InGaZ705QKZzeDq8iqK0MzJQPSvxGVh1voRE2tgnkHH3p2kZ
cAUB/AuK0zLxDbTEmPCaVmD75xeRo5YCJ+gGziViNVtKOMewNbTM9LcmgPZ0jZixFJIVbfx5Tfqk
/qK/uDxsNDaI650vKOt/ifkHPjPES14f6q0CkjBMOpzr9zpwwewIggg7DmWYFeHFRcKcQmwI6Cop
YeTcA5XwgWGCttbLr7ecG0xDoevoUXrTPFB5zwTZXz38OPMV8d9SOd/qZVs34Tb2X8m+J2cd2CXX
BQIvBQQq+iELF8eupiELVo58sP/X0tQ9fJka+FznBBhehjUh/nQZAqlKmfljqyP6ArunqrMvZFbs
tDLb/Kb5s0BdH2aZPjdPFdWqAOBspkUa0FS+oBfb20MIw6VicUYyXzfCQ56hi9z6MoNfR5GMNuxd
rnjA0Qattv/thI8ADI+hIJdqr+6Rhj/CJASbZNs/AV27j2t0qURA29+ltICL2Pt/4VSpG7sc2QYM
7fyFjkE6XWPO1ve67iGL/Idts4pLE9nWHNo0AEgH+kq79ZGYFW4lXF4cC812Jx9tM2iy2pMgSSUG
hRNH5BsOgG7UWM+hP0HsIEHVLNZbAbqmvAUG3k+BURsyGU5WZFz96rA/4cfJ4ZOF2fczXZQSOe2p
StIUBLWKRAGkrKr8CcSgow70n6v9yaMdkooegLlQyePkZdPJSGskDqnhLuZLarshHSiVMzy6f7zJ
QeZpjc264jH4zkl4RdEtYmPonAYHmwAglkzH4+BkqpkXXgjXM0496jeKNUdImJxaWBzId4SUHswj
3+EDr0WU1SsMnvcVJydUn2vCZF5+j7L4V9cw1f8dCgSy0bQ387Gp902s0aQcRY77spQygaj/QxA5
E6HDbVmHVuIGl/wTSzznfYmJ6zCaPJxb2e2nAGd2P4HF18V9Nt4FxAFZDW85Q3IkP+vGi3RY7jTN
4rvGNPQsxhn7AVC+fnFXY3uehBQs4GYteaHnyc8nYkilulquwIcqG4gj8lsBQE2bbpZcIaVS6hdZ
buJZcUQIw2BAqgBis7KfKH4WkjZ17YgKZ6B05pEJFye2KLSeW20EZLncjPs8VFyqC39Qyxc+V3NS
6GqCjNXes6+QiZaBjD9N1pfoj6YPPI9zIeLZzkBU7p90sDNA+NAIP7HwlnkYYQO75GMhX+o8Y7Et
UAXpd+rXG4zBG5NFUtwq2iQtZvTORiHVgBWti5DXUwFYfjFNosyYM3BTj3FXvbuK14OOTCmCVu7D
3jIIP1tXcgGns8siOO7HZK+Xix+7hHhWB48vHqUSQhQFVdO9srT5sFoosF8yMn2nxKtnD8Or7+5G
ZCDnvtSXMA2f/twZ3kb/VRuqAic3UnXWvCeIAVTXl8usgHMKlZWqbcXp/XBFrsrS42LbYlw0a2s9
YzTOXcOm3uPsYAYcnryCciRol9ySY4/7dAFkbt/wJQIIg82Rlih8w2I0OshBlsbBCbPuc2SCVn3I
V0515fyHcmZ7RareihelwBJgiLvdfr4Lca3LxeSqel4FYM8gKcSMPfPX375hQPURv6unekhV0fY2
DVID+oD6WvJmgcpeWIFUUSsqlKmvc7J+ltx+CJF5URQtDiJGV1n78vNxySZsEc/yM+MnoedsG4Y8
+MnTu8K7RksE/NCUtFtI0QRTYLqNIRbjFhUzmL5/YvBeATN4uiunI8qFqkwD8PA2yaXWIP1H5TY4
4ztS7ayZbsbkD5K+mxKdJfNrgKrWJUwPY2bXnQNCKgsJgXTvFyu7L0U7xsvROoriaVqSM30EojSy
Fn6zx0kG5xbFCtxs8Zuowt5HErvbYptAZMmABpQHZRp5VEoDa4aUHOGcS3y2K3/YlcEj6CQegKnU
FNCgWU1nYtCDPWjwsCwXY7sybCIeI/x34h1Cx/R3NXK68TNjB+b2VCapa/f4oRbp8yuWYTEaT4o6
iGAMTyLCx46jgFSXjjxYMVj8f9XQq6ZpHckJ5xSRnMV3lb29zSY7KNYW7yanDhf5fuFgnHNcPcJG
0JQ/NGQqgOEWhLqY/gUQnCKPq6yrCFj42+SKK+pMPEGKBk9Na9xt4jdLKzVECTaaDrZKLIuTLOi6
CWQGdsRlM0yWZWoR2YrXxAaYD3tdJ5dpO9AaKZIcnei+U1fCi0A16d1Os6pZrV6Xz8neHVlUEzT8
dubDHkdSUR5QK8RiQscR+/HdwJLrT7iArrKnKmoT70+dXUnUP0syaykqAcNM1VYCdBJ4PNn9/DVs
f58pjkGfrqCnUj3W2Gt/lSUbf3Te7m97xxpXvRDVvGujAQw5jusqABMERfitt1ypGY718Wu7qNHN
1fMDpZ60z3vF+2Zb4OoIDmU4wwShwgYckayVTiShPjH9UJKXrlfPU2K2IdkPHQ4fCskSnljf5CBj
iW/xKCPrXnjx+++Rp+ypf0CNlkQt2vL7J4/s6SpRNNKnqFMlsSHZowFvnXbe6ZS+SGh6dKWargpo
Hw7jq/gKAFUk1XHBBGZzg2HrNu8+btIeSXdh0KImUsZlz4/S6/d6OPRhscn2TRSG8GUOhkcLFWNs
v5dN5pz9dCZTC424GGgQR8KKf0MFTY8Pzy4Oze2eiqLf3pmaaICrNvTlyz2KFj9Z/ZjJAeyrI8/Q
/8XGru6MFM1d2mjPT+cvaLScFlwb0YH10A+7j+RUjUeML3SxStkbPNcExDS5aQy5AxCM14OZz+yD
lNfmkrAU453Sm5mgTpOiC9rbQmnnlTXk0fswNuLXWd0a5spjn0vG0q9mDwFIeDJK5rwccLj1gYJI
bKbi5g3BBW1/QkhaNO6M/imF/jENDbmtjxLtFVBPFm51y1lXAiFYjpSICRY+KPP/9Q22eZgIarEm
hNLYGFYziB3sIkAVcT9jwHq1c95ZxrPP9BubPWjcYY9XZWMXX6/t5XRci1PWqUcIPIpJF20ScC92
MhSmW1EXSV88O+fyM8okhCWTkjZlJX+JEeBP1VegxertKROLERpc56kOeTKjfUMrD5YcS/SMC5tX
ZrrUZqZ2gkIifOIBU0B/CDYVleH+ox6c1Zv0JIoHW0A79w39VV+8T4oeEts1MS1lbKK8a45ReBUc
8lSpxs2eM4Vjs6BW1s7wp6nwrxtP8aqCNgJzj1WfJiaCxrGgbtthACzK0P05SNdZ8OqAPv/wgr4x
UnC9Q6XW8EfuDvzn4j4dPmufZMIltxIcS9cnp8GoC3ccWUi0plcqSeHmN50lT26DzVSphSOtcYDv
/xvG5ReTpHCu4u2RRiRv/zS7zvhacmPKXDalIpR9/PFO8A/CjLZwEItkz/y489CKaTA1uJfL6RmT
0L5Ggy7z0DBjRaVexnMV+o2M7rrVXx1pmEYeYmiz2dS7mEJnKivS4M5e00iaPXQ/ymSMCXTsfqaB
bpyU3+ukV9H8JDQqYM0tPKkqfQdJBTnksS04Ouejnfzw+mJBqQWpzcFJPz0fMeuIFTXRhlj9K8Xd
a4z2oVj+oE++/eH/bxASfG7ac1hbo2SIOIU0nZBGffPMWG0xBseIr3nLzC7t+KWIzUVQxnDx8uqC
79ABrDp/hR8Bt8QmLS7MWBwAUsBOZacPy80+Jd+heSlXxO+zCKG6kGi6nfcmYLARRZmJHHJZweu4
cYuLz3ZFIlBqK58+vip99HNTrc3+B1st7a4FpBLgYDem63CLEJ+DamU0EiXYwSucwgB8ix1JGpYP
WnjHxAqtvOHiedQkGg8bTzusKZMIh5uvTQPSYnEDiWdn4Tg8GGL2cU2UHRMDCWg/FhPj675czXG0
j+noYNR08xDy6txTh5liAbVJ+8YdFGVZ5RyisM5/sh6Iz9hc/QwgcIB4ejcQbalfdvFiBOkMVb6A
qOFSNXnALcCtw5Ou+IMhEaQn8MN5dzs+HZF74iEijUwa1B2t56OJ0BNqF1wlpNA5ZMlGT2Kor1NZ
QIy+FDpNevKtyXk9I6Nzy+3VCSPsKt4qyivYuigYdz3YLuVB7pMGtdBXct+bXPegTxJNJmZvW1/t
wje1Oj9/3JWvviPQ7Y6oZgmp7tMRzs+tvFR80VW85fNTKLCejyR3LdHBInh59jJxZOGF4BcyXqoA
4atfsXPIWuNyB2Q5k2SyzPpagvGqVIlBKYXKEarBQqnSgWX1SDJOUnTfsMrhQgxbZHEGE5v1uj21
0okVHR66k8wlyd1xvFVfwNGElXLv66kAzS4bZF/WOKpQrRautteAqHz/M13wKjxhFSYOXRuL/6Gu
nGRH2O/hhYrmetSNvofZzPhb/zCYapZNlb8gaCepxdZbel9yiPYX4clBx3N5Y4yxROXoH5gkP4he
DlxqoxvmLsPJhiE7DYqqkVCySLa4AYG/5N9u+reB0LWjq1T5uYjYkboTDwSapdCmg+Ek3zGJPnxR
LNaMxbAWpgt6ReOrw16bGLSSKpKllQgGQnwxZT5QKtuHzrTbquz4MBnSCqG78jh4HyqoN9+TUuDt
axGdrDs1JfPuGwiMQ9LySy3+78L5uXr5EFqNom3iZF0XOhgkFpAZz9tn2vgVMy3cr7lpbOiC4N3C
tM2R3DmkYu9l+5iacF+TsCEuvy+BaNvAq07dVwE8lHqFenzFIFBd8bo2YoCmxTzOcqC2zs0ruMgS
okJH+efMG6kJT+K4a3m0SrbQnCdELj6C+Lop1p4wnd+E9s9KMA4ki3rsMlRnCg5YCw6XnpMw/mSH
x/GaiSwBnSBXcKDc1l0Qhr+HI+7ohOUa/rTOPXBnQdXzzqXlVycO6++4iQc+dCDIPGOzk1ZIsLH3
c1rvMuySHC+RomFf3jm+7Hof05sHbzc4oDwchszIqF9obsRQnQolsMhEAtTVim4bKcskfjVld6M6
V1SaV/MXNfAop4cyKb7eg4Uoih5YgIhzxRrbf9mB4bu4clU6+09KCSkvb2R7T5Ra+s76sy19Hd/4
tBcKX/T5vvJ61azQoxtJqHOXKrgCCJ7W8n5SYaJfvPlBsDZwuj2sRN5LVxFVeTKPPh3RlXy9wX1G
Lzkpdk9rWUQplh2Es6Owh+suOt5KK/Tc658I2tXKDI2Y5WTVmj87Vec4SrkGJUQ0Jacr02qCQ0RA
2JDS3VELltyrFqPjtksQIVaV6xvXQWhNxfucCtgMWCPDrs4cf7bpgdMVdP/0dFAGPkQmYcadm4lK
SvYVfCMIXJRhGqXjvroXdN5xs6IsffIOFWb8VXkwqlrJAQIXet9chupnjGfucijcLbaS1rEcksgf
BjarXHM7xvS/6TfihSaPXRHUlzaiq1oHQEAmEcNz9msmEqG3HeZQqKxeoh0ZeqcXWXld/NH8Tf8s
CE9nO4fuSgT+GpBLeHkLS1fzdsB0xSnXF44zYDvQ7GDnXrOfpsVfFI2DMfZ76I9/D/g35XwHIuku
zJTxz9xT65C9vBiaJRc7fK8KqYvrBDGf8NSSv8lOkV0QdBELFPgebzeO1yfm01MC9MWxv4Vi/1Pt
lSEKPqPE8066qVcRQCxeEKIPncNieBIYpxWtIYWu3S50GaBNz0PCtmy8svWyYTJC6040YcnVh1Yw
qJp8cEmQbwp8bvx6wqXaYS1PBgILyz0fb8eDGERcQe26Rrc1sSqPSyzPN3PUueLUWWLwfvULVsOL
7EAHGkDxNKujFF1XfvOB9Cg92Wr+5iOdbTPswgj5SUPUYY0zaYWtRTaX589hQAYsuRiG5/oaLPDQ
3MvLNplsNfzkj3TI2BvXsNeju9/fifQeJLW6B8/qApVwZoF34GjkI8bX9YVaDkGNHAaaG4Ybbfug
UF0Pa7ezs+t5USfSURliUu7Wfu7NmU3/tgnmVinOUeSsatafISakN7vW86wHffaK0cHH7B/5VGWS
6ZmMuhROxCC9oDLqfuKjrILff2DhZux1EsKwOX37PDI5Mk8kA9UA6wcnC2dZ0DslmJcNbiAq+1k8
gRM7QKE7x4Hs+PKE0s6tLNOd2JhCjFRSqqjCaKlHoFJjsLuiOAuNmBQpNxjolW4XJuTffKyB39ud
B/6NK2FRClURHnk7qJgWNNvj2+ZUZ6smlnnRVnd9XjbRG6L/bERMjCm4Jq5V0uQCt4UcnA4xFyvU
czinPIcHmeP68hmgS9U9N4UPoLW6WRekRrkzinL9GWofO48NaKSids5ONViJY6iskzfYE5hBReBV
2UiruFJnwQaQJ7jbtRwdU8NgYdyzibf49q0gPdksALFi8PHR+4trVZyCWTsBdpF6yemVlu/bVNWd
jUFKPT3hDpeJT8zqMhAYav+lpEVsKFwrfwFa3GlJkfFrnhbWbZGs0Njr39J70m0K7omOiGuhdHNB
KMfVpAsQ1duMnJyJHVdefAGU/K9Gv7ZPZjiBJLdVHCyDSbVDJO21e4bmmv5MMRQM1797dOrakDIY
mRm1WOyUd5vE8CA4U2tyi88q5BaaQcFd73zUq3M+kBJ3dTTPvTDNS8Ge21ll01Kc17tE0wi1Qmtz
K3Z+XSHdbGFOKSayGfzLe3cMd60lg1bhoJ3swa2SEe1vbWSe1YAYG0fzW+c1iXo/OJf2stHFh+J3
PSoe/eqdtE5sMd5kw7fo8iqLXe6Zi8UREEgmbZamTzw3Fpw2ilY3n1BqA0mbTO00Nn4H9fyqkyl1
BtUwGtNQyUr1YTxQ9I3lUYDZclvVWwIe/MB7NowvKYvhOE40VwYJfbVl6cgrTMI2+HMKf1wZvPGS
hylMRd0KvYzDYQ7aV5xt1xPRoKYrClaVkG7jXl7byu6oERfeNLol/0/QvSNG2Y92FvGRyqJy90aR
mV97Qbde7OMaVjw/r/rt6/R355Yvg89m+DYAmSF9bw/p8JGJcwZw40vAHuBwyVzPdaXTc8IJl85l
nwnqIpy0tZHb7h8wHpjGwLemrydjs7OBkLtmOJKZBWKOyfrLGLjfQNrq9OonPLMujModGk6JnzWs
RRwLSNQ2UVe/CozmmxNN4SfDDaVdU+utRRqp9HeqFd2GQ8jIblTCX3OSuV8N7Q3ljR2wSgzA1jVL
bPwNe0ZRt8quVNK8RYQf+hU54YRjS3U7sPXKDrkQy1YNHQFDhdG5WRGqfxggsaWy8igsnvhl5onI
DocLcojJ8WREEgR3uBG3szmicDLxEGFu65JhCCLaAj6Ld7NO4nFQaMTTs3baNf/4yc1vCSCqYh4R
uo/UjtRYotQxdtso3FeZo2UgBCu1qE9qNSnZe2X2CRZTB2yZ6Qwhg17/xfG2lIl7I+ba0XBmkVrr
RG2UM/ERvyG8mAm4AEN620I+X35QljCoaCH1F3klT6//PWuvDm+QM9vZdYhTirCS6TztC04fhm7C
BUsY1lb+HwP98PHl7fTVbh0nKLOJfTSyLdzjytwTGHfexZc48Ud3MPvxUFwe3QKw56mhCNpmvJmT
HYaS1minIhbF0rQ3FgzkyvNuCDomPmUOFNBIxvJZCRveFOeT2ccbias9qAre/V0PgN1ohfi7FQ0A
+SWvTs/gWxC8RJ8idSQSXxwQFXz7idBEIj2iCuzno8XbyWlC933lO1o6zlI0IAwgp1rb+1WibdoX
Ykh+oQzDnyNIoA9zlGSyt0FqSgj+TanCJ9cFfnSfbXKrMy0Pb+cVZ+nqPjwawqjJXBHcLN3t413r
1ksFqWvu/GxVLJJQMD3x68LA4NuxUML9wqwK1AA9EwasMDOMDsJk+ocEJ8tHDTceRLd3zHADSamQ
wLxXHvGZc4FnFRpNe3frRfPvL11Y89/BB2urN39qliqqq12jMagNBaOjKh4xWwlMhxx36IYu6BYP
AOVDpnJG3QRK4EI0P9LmTL/Rr5orvEMSPLYGx3eeHMfiAKey6uhio81STX8sYjx3nh3KlP4AzNmb
mtIRd4gAi/l95V1bWqkAtpscJqRu6fxkLZfmZ+CPpbBZvbZx+7aBvyWOnhezi5rSGfMThn6Z/Vv+
QdZfzhrgwQapK7CN+jWlk0SlsQ2px+NGQA5YjK+klS0G/spXj7pon8MFJ2iPQOiN7hSZn4niTPY0
TaMrIichBkXlAk9cOjfIgXpCLUKTDLwziNg0AM11596uu8X0l2DpJZC7k4kLpTNY2i3UzRMKXOvR
bqrwOy/EsjGmFJDaNaZYc65LiZItM3FGk0vgQk+m26kICYfojkcLEHJBeUsipDubjy/cTZmYTdpN
QFuzmHK/36VKeiD+7RRr0NwosL4y0DeXg4bhfgXGOmLKv/TMpA884LbFYBBgjlhauBPg/VWyP/7d
poEtXo9SB60rQAqNyUB4e2lk/68eHZXZjA/RF7htH2AGlMtt3Dkny4aXwKqo+Cdla8Vj35Tf/J1s
exXzHDLol1Tl+i2UaaBYbjqAdz4EoqJxArxoqP60nQGF3H5rcd8X5AsCRLX7xpu+HrG4uCoH3Y8Y
4dvZDfEJfkry8G6FncjRhWLmP1buMED7coqdn7cBPbxZrOPaOrWHP8ha8GCH5UNRLsy8VyUq12xS
z2Uzmp5nHLU23lsAm7gnRMEY7FZ1UPEJEbdgUZlVYZA+uzbLF00PIs8/JKGqVexOKfLfhWtejqYz
jtH33S7UqzU6Ig8rrzED4zQ3e5so/9Y1uHdQC6RIJTbMBrUbgo0+aaf/dq2/TTcyJbdE0xW+1trX
EEBfzvOtVCRnbepftyj/WPMC+OGjN1GhUavVma0vMWvqG4AvfY8XKqIQ+uN3+MLMEIMGQAjEH5RJ
9udKX4FeeMEGq43HtKAYEZox3UyeOdotXU2UuLmtYC0FjYFrN/xP34BmAItXUMw3D2S/R+LqQad9
Lu00liqUZXRKQAfaqOVHOxRoOB5phT2jo6Bj1g/akbk61/5TU6AHeqy4Gok0MfXDep4PloiFArlM
zayxHRiHCpkMXklOVkZ2ZeAnv8lrKYAWK9QpAiiHSIRF/v+EjjJ2GKTXn4XOUkwbDJParvUH26WT
IrTW4Rto8/DeBixgfWKt0zYuEPUR8e16GtEJyNlKq7rw9PXgOGFY8lN2Xy9N2TPoUgIU0hpb27aE
V8zhWUpVDCVIzbshwjGleVdwzUpJhwptwLkyoHX/RGhXqmV39afRm/KYvvU3S8gXP5r71mZmdvBl
oFbgQLtAP7AvAdONjB3UPaScmTZqIxDov1FKZO9g9RjUuY3ndUMw3VSYCf+YIHhtHAdoMZ+3hAze
gkSShO5TXJMlE9jyFWh+sVxs1xRGpoqEfl70woo7lAoNKUmj6Tx3RPUuc5ghfH+Wat/q0d3vEYQn
41SSeJQ12D6TjXcrJtcfJTvqrJPX8a2dXOZ+QmIhp5ab48iQmJc8N1PmzzwR7HKvpZUqyF514IZY
BP4KQnjdeE8nsdYJ2ibBdM0FzW0cm797rIYdzsHhd9A7o6FBGwZhf436qJa7JsjkZsU7Bs7xOhnQ
dDEAtFDlliosUPtEKTyCeMLkGpdDT0glUaH8FicqPWfyRSeDcSlh1ppH2jqWsT0RGCuXXJXYdWXM
Pz4p6KC4Lmv2m4Giin6ZypruEszDqJi+pX9Oo0oU1j/WDDA61mG1hbtkFiL9yVYIlQ9IXRZfSWNx
VSkWhIu1z52Z+QyhCXLNpVhtaoh8Lp23i4mIwzKpvU5NxW8mTB6uFkqt0YySwtMV7/7Xs68Uj6S0
l+rjzrSNJXpH/luEDbYqVM7GdeXOzOQjJbwofgkOxDZt3nsd5Z0R0NvbSUcTRcCZ5y4LnGF6KZSr
GX2K6m2WvvuLDpjMrw6ud9w5LQQOTADjtvB7CzVFkwcKdbqc3WUUkkfgdm6+5GnAyB+Czc2sn0aE
IgfVXuPjqent/qGTNeaxysJl5R2OP71wT5CnMh5mU6RJxt2Nyyvnxc5SeZXHwNnO38OccT/eNqC5
opC/ReeNssenF+T+9pwknQm//sleqCj6alf923uh4RzISSvnC+glkqUIK0iUXF5uf1oSw2gNIIOf
gw9PqEimSOmwASy5x4s4jTSkGuchkt35k/LoBmhJuyNOBW/Gw4xZ0Z3RIFKhZn8Ydk0ny1DOa1/x
iwKXJHXkOgTBpXYHiS5iEbDCfY5a9V2viO6LxKX+XzPy1QtODgW5dT7HouFl2hm9mbz9GSpuuCQu
COypNtRMudb5/l5xBBkI4d/X/FYN0hcY6zs3i5xpxFxsZwiczH5i0+u8jmxnWgrkJ+hfril86nFH
sBjMm7fUu/hKd1w7K6kxjB2ljbZ7/hNCFvUTDzdZ4ACqBiB7FaknJMQSie7T9ywRYYvhV7TVx2hT
BP4Da6nK6HVfqsHc7wR0i8gwPuvtMTZRTrQHnOeqWb2q9NULky2B2D3l7rz7YhABYnCg1YLB5/zK
M9lbt5yYnb1WYa/EzaR3p/8gT3EVBW+gqaQgUHYDWMUO0fCjMCBgvZof9UcIDYNm7kjGmw+1KcNZ
Tfh9cYgVCiT4C0yi/n3jUKhrxTDb2DsT/+6kTQOqHDRY090KOSHQbgWLi+PCCWuNqP21lvPT/sC9
6lpYc2OHsSAMYYSSlm2yCGmPYVzWlB115Tntai0NZqfjkVVPCuEFYeJ4DCQAyAmDLu0PkuCzHlfn
3pF730bwZcH4LGD65oKbgQZVFlwkZipHKJ2do6A8PxaU8ecUGFtTnkPuS7PHetoVDxtjbY6eiohB
HKZ4jatkg8bUG5tSsadKh9zQxVA16PfmNJ+sypDBcOZQ05DcOCfn3HN1dBkgXhFxeqyYwBicPz32
JWVysjb72wMnlrS9nRWtPiOuwCVxyfzDri3NroKxJwfaxhFr5OOxobm17UOt+nPhHado3RLg8SoJ
gX2Bcqt9oFgmaLxchEjxnzzzuXKtscsNcb1HOtNQd074P905R7eETiQkfJuq5XRdP5ivyRbU9Yty
1Khr/x4wRZEhFW9XDMtV9t3jVdWd4c/RN9Va9gigWZdabA679u96ufga9C5j86xz7n5cT0raT5I4
GE06AaaYNv8s3HcznoRMmtqHE09I2oyuGLRvplXDPNen3h5ngiUOPWt174FEfc2NY2LMpaAO6GT4
b70irHbtpTXE4RrztC5F3nxUhLu6FCxpfwvypAIKcTl2nDN/yeIs8S+nFteGXEEtW/HNHgZr4mtN
f2Ekh1/I/61ovNAiyXT/2oeUcm24CBIkz/TyqdbJeeC+ZK7nTL8/5AwON0kyuyQLa7t74oirrflT
BVP65b5ntDS5RVxRXLtLYrler0yBe6WUre0hOTyAjY1Q4vW1Op6FD4xm/VEvuYtiARI9tT3Tjf80
BDDmoIpf20aKMV9z+TM44W3B2pDoTjYDWfw4pkaF939OZqnm5Gc5AmvScwsl2lQQXDN7/EE/GHbX
lmdAxjVUvTF6IMXQHFosR4Xbi4xomKVngbFxnt4BK5eyJ643OywV2bpCraLcijGsJPPrWmvV2uze
6b7UfVLRLY/i7W5PaR8POiAfrfTp+j353E5bOlK+hqVNEx3AkRA9hoC6rGDzNOYT8KTAmpCOKOZB
7LLMZ7vf5rnSotXbyuCDsIyhTWKy9Hl9HZh66pmMV/3DfqH8wQJ2jn8m7SVJ5o01dFufu+Nw9Dh0
qVs+cdontkfISzse25hBa/RevTzhbkQBp7v7zKJfmdtAZPX5NVzot9OHJ/7zZi20zh4nVPDHURnF
vGBbBxOYUaaqU49ti11+2D2wxg+csF/ucEZ4iU1YQj23EMnmO/8GayJ3oEo7k11n94AOLTeUkj1m
jhyTUoExhJ5lgQYwdNjqRDaGVjb/Dzrv4vw3TOdEuETtc25QfiLMs69BpRQkIgpUuQw5+JqdH+OS
zqdyUt+OfZ8R/qsfrrvNeV182YJlTYAgZ3wyvJyFg/Rqt3GU+qh4Tu8fx9XbkMH18P5lYx+YyzGt
7DZQoz5SaRLonwcMBMRfhfZGr5W6MB9YR+Loe7SlwVzLfXwuG/DpSktlgNJA1pn6LoHEMwAvKvVe
K1DZqItMsQOPOhn18d9V4rwbnjzs4qcKvY/0MiLBApZ2+OgVJld3pjRXjNg/8w5QLEWvcGCJSyvf
ZGqDzeodUBI5H1/7wVslEudg4aF8Li3q95beM5pLjAhr3C5koCxqTmmq8RimPwyMh6iAS9wbabAl
V3P/d8RyTc9kGUWye9dK1BLyVcpF4xydCRXNm7pdsmqxzh3E6XjRz2Ou4Br66txNmvyFeXeuZ8T0
iZAI09444TvW5PGEV9V+r52SwCso7RaRYCwp7vYpp6tqA4yzJ+BhBUPHru3Po5u46yJ5C1ZVTlYe
pcSEPDrLDFkPPrtaCB2quH00GFeZxVCNsIK2lW5g5bd8Zv/wUsd8ntLEI639GhZGtUucoGCYGRss
3rACyHEYxfClvM/YsrD4MvYTluUc6w86anPjTG4CucBPEcmALtlY+zg2RB/X9NaVbjMd4fsnBnk7
y4RzWIGO1Boy3S/aZ6+1jVBIeL1UqW8tnZ4iriMYPwNmeOhThQWMR77fkhgm8GyGVIxotAShoLK+
2O26ToW+0zCtgkkhjB9NY56W1xiYZ0kcZLRJxBMKIwcFywgCvma5rCiGQXYTTwkg8gNbxT7fWsgh
2QJJE/gqrQA9EBQ+X8s/ZGcqLp5RgUCxSSzOt9LDfYVj/iQOCEvkX78sPN+L2Fxt93BhmL0u1V28
K3sOszgxoK1dPvzPPq9sREKUTnUOT9+S3OTLiBNMt86JpKUWIDJuRFvrrKwF+95nyOmE8WYba1ab
hrr5v4/XyUD2WVwBjMoK7YFgiYrUAW2W1b6QgFuRxGHG/S5q5PGlWc6aNZOeqcX56LorYi5eza8A
ESXMbF7me6yBrwhnBf08svFuZfoitoVADizWvwquRddlAurRAly4SyyagQXTAt6Cqrwz5SbVCVHV
OygupI5FIowqNJaMJC72iANPZY1AFF7DOeNSHV4zyK7ujO6jXqR3PXZGqYzKXiKPQYeugP11+dZ6
HD3eGhKdAIsyR2pJKmoNm675koqVF5Wf4Hn16/ZZaSplzi8axJHKAymr2cJAE+14RdyeL9AU45iX
PcUmfVPtmEyNWY60wWwj+95h8cGYeY1ikndmGRscMlHaWRIbF5l4JJnGhaWvTpcHpMXKqT8X9bb2
aFR75QRhwbwILMM+tlFSQ/orhWHPDAKVGqIcCI4F5vhit762sChBuuvneo/RDKn/Qp95oIQyUVG2
TOdV7ZPB8JwGYtX3DlzgjC/xKmiJvfXrJj6DsWnG+Cb+S/GDMDEpPoaV46ODASis2Po4bWVozCXx
Q2PpjfPYPYe9bsLVFUWL7nY+Qzv9qlblkGov/9DL8oXZbwHUO8mJnQPGejxFQoz2MUrrlerb5opN
28sxak4PMxrkcgX0B5BIp20efxTlexULO21WBbKjGiAQiGNGU9uZKEt8+x+scfyaKXLI6YSw8cj9
EKfxNXbCdcMpD+VZDhUB0+8Uf3v6RHFL/9F2fdLawfz0e80NpXU4Knnm81yryMtKVb3SBq49OB+s
hz1yJnSuABx+aoNypQNOE3Vpb3nzm+rrdBdQyBE61Fx8gbb6k2Nybca6HQUKoMpDXGtf0a2jghFZ
gek3cf7WnI0wlYdvgsMsOiVjUD7ykYA1/1miTfnMvMmhJmuPIp2m8PbAIY0XmiQwwFLPRIGd0uW4
zEGLRdrm4nPuQ12DCNUbd9bjupo0PAlI5dSjVSl1caXul6yDimmjk/ZoQeQZxrZP+ZBugV+Wz/9t
AaR94kqzdQiKJY4tad18QOzb5t8rhFl86/Nm2Sb8JBBnA0+Ix+tjAiRIpj9ZIB4HDUhZYaEulXrQ
ck0jrK1U+b5+RFzgXd10MWK58MzyfJkuXQepz2R4oJyxcn8HT4PVd7Vvez2svXmxsyUNbDm8vxWS
UIBuKOWscac+eRl+Qj77gWROk2q7MWHnKtudFMRLaHNMjRfOwLQWT1/ZenBY3e4eap/wsXiaBCJw
pMUQfsd6eS7H9ozhVwZol9FJrnGJBBn7CBCynJ6cJhOj/nHgxsQ2dH65KaiFSmz22NJ/EwBfPvJX
hD9kWyRRZZtSVJrgq9QHO3Tozr2QGSqTihuwOcFsXrTTFE8WmdpUDqLkyKK3pHTAjRCS6uakcbw3
8+8R/HjOpFRj8y3ee86qGgCVI3pBl3rsvivN4V4gLFBghYHeEC/5TBRtQZGfiSYbX3xWlY1cKpJ0
X5+UhFfKzu+mev+QyMt6yUQ99+75sGIkuUdobvLbc+1pMQiehyYEyIta2R2Cr/NKnrMHK18lpSOZ
b5T+QvChkxYxhSPZeo0RO3YmCJdwpm5vxlZ2UKT+sTOYvoI3xy3KjVdRiwiuqrXviEK8gBFrU4Vh
0SoGazHdEOb8Zx+cYKMY/54WKp0s27vIlloPoH9Xo9/CHfQhTLQY6WBTs74eQHMHOs6HixvVk8lN
IuMVvRi1pkr4IRY06KMG6sq6nsOP4ZEVcX88Pi5Udo/ThE2WycUh6/11Iw03SMeSU58t3tjnjbyQ
ajW9dM70FTZChzSg4sveTGle8uw3wLdb+pgOK2MafTPFKgwcwXWuaYGjex2nizgoCWJETAMz9zow
k1XmQRnyyZ24HczQeGCFEOnuzMKeml8XLHjlee6sJW8j4CsVbha4GPw/HbX3NrHpPdw0E0mXPlAT
FTH/qP2PuEpXM2s7EEZgg7jbly9ZEfoxvxxPCD8FL4c2AuWD1ksL1c0ROdRiwHIRmAHnqxICU8cG
ShgzEwSP+8TeM1fH0totsREP6uw09ROab555fRKyVgQMasPm20vEFf6LROZAJUegB8N5TtBkZy1j
hnCo+p0eIJv5AoF/uMUZs8qqmbaK8Z+rb0RvWGwy0r9H1Fi93EOXR+GiO2HOBN/8ykXtN9aE4Vyx
uL/J2zr1R0KQaeUfFHQef1nbJ9Ogv8RI+mbgH3wWVhcSLaq4IOFNH8E2P+XnTxY/AwyKUtdtmy/8
mhabzCmG5dEttIMZqMMkaXJyGyd6nxYDFPxterobUZs1T5olIcl2VBGp21rV2Bp+f1ihqf9207x6
AArxSFh6qvAICL/N9/hPw0zn1FilwVyWcOoR2MF9R8mFe9VeFPXwb7xUfA0D4ejc8PH53ZI3cpiR
XWDboxk8phT5vY34hxIWLfhEmxdJv/IUSAIrhra6ib9bDw+bh0t4bANARucluQ7ofLe37zPp4o5h
v91RtADPc8Ac/l8hcLlc6LOoSOgiI0mBQ9kOovinxSdSny8MnS/HktI3EkL1bbnbWNcLDyJfnVxQ
YjAvgeYFTxZJsKdn1OS+Qe3FiYexRNaIFagN0igZIe+ONA1c2yyA/d4tXV66W3753PqaDMXQpVVL
kTCK022nDBqoWenC+jqe223q7Oge85BjJH0ZSnDxTyeTZpYrfSiaazH1PVeYpnntosiTHdAEvYGa
l//rfXRBL9uGkMq+AIyK2ETtg/DGW7up321ujzizdk1ejckVUzlBh+MHvyd6j/nnv8g25oJg69Sf
7MXXWIj7q/GIMH4v09CqqcdoPj4bBqMaTZMxsh4T8s81ioF6oKSlRqrfgIjpZv97+txs8LfcqAe8
OXwL4PZPWmMP5EB9fyVDwSDsckQkMiChU3aaOTQ5USicPlD7egNTnQisqROTTwMwF0dZlaTLDLfY
N+xL8d4A4uGR6+nyb+dllmPhD4GDvP0bdjGGp5aBgHoRMcckqlsRgg1QLYamtnrPALHHpbZ8FTXr
hHufBND0b2NwZwj9CDEqQYggv0APMZDxIr6/jw1MK/wCTdLfIYZRxErt7kM0G4JRs8gX1M/hPgbt
eHdyuWJOtQ82U4aRHjzIi03i1BtuxFvZIusJkFCfrW/36U+VhpVjNQ+UX62SOKz7QxJ2dxYBgz1V
zGzEroq4sWlt9Z7ArhIAALFOcfqKZkSF9iOM5zX7Kdg+wUueQt6WozCM7UmP2QhVGcAxZKvpian8
bN6+EmkTaU5UYn34HUozeGfypaL4DojP+L/WIqZxYGtS7H0GL+9+6tV3ZdB4lDRt8xhCUxM1ZORK
k/pQIlW4+MIuwqsfqVJ+oZV4e9awVEtIA6Q398qX1tMjPgsK+fFKx1jL2DQ6oMDfJcDVHz29sjaR
k8DvEr+lSeRH4zCx+25vPlSTF08ydceZd3yG+Fc+E5T8ARQYT/NRO/3iV2vGh3pY2maw8mc7VInu
vpVNKnuCN5xq7R7so6KOK+IXQ5pKS9+bfQTyNruKOI7/wsVUQujGyp9o9SxEJZx/tsW2bkIBh8J7
RvkkbKd1qUWMr2Z+FYIVwoqRNWI2pfm/zUlO7Ab0igsGpQbWhistsNyBo5vzZudm5X/E2O9FfDDS
OwSXC2OE9Ip8TjnBWp2ceDO610j+vM0o6hKoqTX95gmeOf8uHHe5o8/GeVAqcFOtM0LfgkWR5x5s
Lbjw3YUqJ+TrYF/j91hpwZat+Z8UGpX+73CTVIG3TxWsSTb0XTXoUfuGbTzzDS+PfNd8YuKHGMzd
JF95Lf5JD4H8NCiey85NavyxUQKEVchP0ZaBFZkXHiGfj8cjCYnQ8ETSuc8HzLwjL4h/LYYe0E/t
C3QgmvVV5hcsPmmXwvbSjZuj1KFp8tUUJCzPGANiWFiLGFkAEPRpDefKogSI3i7Mj4n+5IawMf9M
JSciWeH4/jTTVuarUvmAG3jsZ4C4ytGAoXgd/fm79KIr1MpPmEJYC2+/AolGGkjBfOtfOUmGqxVK
vCNE3YBFwbCcr4FI2liNsH5bWXEpv5IEdEcN2wmKu8fbE5AtYbWaQ59b8uce8vcSrYH5Xu8nojor
9fNFFoWe1ks2Kn4/Hx5G9fYFe4JeZfMo+HsEw2oGwiO3i6jUHW1Zc6o0a1w89SMoJf3Kq/pDFXc+
YqK2YdGw0wDuusIY//vrRs5GvAmInxZpFXqmA8yjhgdk0KNqzoRh8C8xDAuq4DcB5eZiYn4UGNvo
VQQE7mcz6pIi/dz8P/Zjhz6QnHjctaNpjPUAwODZ24prYQd1gLYu1knlEJGUronTpWJ4mHWa5VKN
gwVSaoxtHbe9ygN+aFIWHnI2CaoVLXUsghRzTap1ue12OHah3/MHCs28DHvCTz1teQA7g7Us4BWs
M0+MC3Rt+WoHtcnPkmqGZQqyc2VYsjGR7hHy+tOEmnFX0zzs3XVSjiJiQMv5KMfH/clbQ14CT/NS
jdTpEL/ovR6I2nmjV2arZDlSQxyFazi9GFa2MYK63ku7KeHhZxry6EPbI3Vy1scoX7TQlAajWrZ2
udPvWbVdxOGLB3fZe/fnZM1TkbYuPrB86t0BDET3GaXW6LRILiYzzCMyCgLg4bBOxCMopGLgTh6Q
uHn1sJx9trA9nwQ3+t0USG4KKmwE4p3M5P+uu32Md57YWG2rOAnyg/vG8VOAfC21NFJ7NY/agkdt
3e6symxiN+JAtk7lATvmUT4RH+u8lWXMAuh48trm+zYvWgCIjo+Rt52+HGTwu49Gs3GVsH3byDWw
uewZtGeITLSsY2gr0vtL0+yeKRkA/lNSxnLg+sVb8qQ23fNC5CEcKsO1DJULWceLOY5jcEKXcL1t
Ud2b/2fR/c4n+6FXpIq/2XOsPguYOnSELKhWBMtN/iEkryM6cAbnTRw+Z+aAfqmWNWMMLYdKxkWY
SwVXn0aeU7Tsxfd+E6jlowxUCFP32TZmdx8qZJU1DbHMDzN8/is7Lv+hOBcqJiP9NM41atWhUykq
a8A8v4/Zo7HWGwHxzAS6mv53NttIQc0+OkHRnZT0zSO6zubrKQaMM2X5qXPubMC7XyNrzPB2vq6j
NSN8aj7Ty0lZpGVvkJfR7MO3DdxXeTTbny8NDFA5BYIzZMEAf6WOMwpWsNJHm8+BaH5wh+mZpviN
kZvEQDt2yHSBrTe95S52OAZFV1ozQ/cbPpVhwK0zyKSEQTFptV+ojtYaWoFrMdFtLNxPpZM1QlCr
eAexIxCd/4+67lpD+iv5TglzGgt76HSvjFftMzxqF12G5eZYCbdZVcQ9UtCVRIqT70dt9BLNQMBw
TiaXSzSUosDLEJwDRnUsHFz4rsfRUyVNaN6oSmdw55wDRUF34NE3n4ZEKS/9nskCKANMRvkpqy6T
2AKkcnGeJ+ssun44fz75jg/OGrj1UubmY6XoRXisDQ4UtchBrI5w4ZDzCF36cMS5hJTgiX7jBsVq
B29EWwfPtxVqyabdrvuk1gtEYHdHvYWnu5BeA78eVju4nLnfwoc3HNDo4281QUSkXmppN4NneWhl
E+yGm/SsZrsXqQ5IJfU4wqci1Kh15z8ET5wClAzAh6QG2TTAplqYhqglUEo07Da5sxVB1XZBD7ph
2YTBmFjO1WV/IbwskPBpnQsFAEN9NQNWJX5eKgmi/dz3e1S8k0rfNIerK5FV5bYMpWJOSBB2LIHj
0JLcnTyfotZJmltUJOSIXgYolKIKH1Is/4qYT/CdEvWoxQglbe7D9PYBvtGD5pBKjPpQbwut8+KV
jNFQqfblFgSmN8cX1sDNx5RcxCBtmO20urBoHvSzkrKKGA0WDaVkYtpsWql2qWvPzGIqTZXIGuvF
YUXjnnjCA9KdgPG8AlBQ43Rq3qst7S2+goQUaPQLfb4bqBDF5L2wHCXXPuAHQ5L6d5lekKqQET4s
DjZMDnkSoJlC+0y1Sq72WrLj0npwRO1mZryXCnikk13qsjYbnB/9IcYY6H6oaxlPFoZ5B5qL1vXy
MBEeX1/yFwXVOmZC5a77A/ZqKIRzF9S29VxtkSsGqxeNIofEWnPFqwJ3XLp+j0emsJsVxSSo43HK
3Ing7LGYYvUE21MfoMkHAoL8Q+6V8nBwgpu7HewOXFeg1KAKNPrIzuO+7XiZ2O25p3PvmMZyYZqJ
iYFJGW9aMpa6WT+CJ+TsgJ0z7xwUXv9JoCq4eKProrjsRGtJgyNG1ekaKzun2IqIg1qyUxlWX6hC
DzpYh4VBmIRQiW8Ef8FIxXGdTM4kJS0nriikEEjbhwnSxM1RP5Rj/f4DIMYD9MDs8nxAlAfnxZYU
YTVH9xowO+rsR1cYWJIhY+/9PC9Oe6mcYOzNItsa93SEBe+QOEGW8+5NKZs70aiMTfnHPzTkyCqk
wbLqFLoCD/vrIQo0eFAxCaKmAVWY/OSZ9F82HUiS01IBCbuyuhNZynvmM83bmPZ17nwwTei5jwIv
Ydy3t2ps5UhCxfdEMlXoCmN9I1bbcfFRL3xN37Pis6QFbNWMNIA66qns/hJa0NoCte0rYV54rllA
j6+mPMa+zm8v2S+teaywAGYqzIQkRQoD/E0zpx38kFiCfWq22VTwP+zmhEOctSsWb3M3dblxFRpU
4N/k34JBKs2YS7D0EK31r450KvJX0lJSVTGf8Oqy7lXhYT9qwN6AWTbrhI0MzZoWOCEf2oGGd41v
r5ILLlimI6fj8C/dgp3aQbV5lNhUxgy7xca7STXZlAlsH39gxIYJgCGegr+3SGwbvmopwrAVvRnl
/G7U33W8rjEmznjeLAJB4Sizx/5uL2Q1MgO3HUMLwxjo/VLq44C77iNPSboK9l2oMJDZqOLMjUIB
ChJIjaNRUvKO7SmWgt9ZNB8icwZuiqr97yTUVdLg9dDKJd0AHoYwsqnkbmy2HOj8y+fyCTcHfefi
GMnydZqs4uPXqlbNRK6IlFVmbiGdEOKI35Ot0spbDk0e3LH4N/jfJK9K90zFfktwPwUN+b69zjEe
V4VpsSEWxqe65E3/PhN+ZhzSl9P8Lfptbl70A/EgSBm+Xc7M9GWrmGKz6a/LHN3HpZd3/ZV9gkug
oC6VMUu1JMiQbOSvA3X1YmmSpBrVFM7JrKg17jOOZVyc07MR3WVdhIOz7MmuhS6COmlyiw0RPpze
TvlRgE2UY84VsUaQoQM4cHIqWj4aF6oGHhAFSQxbqcnta/ubl3GN7mIBquSGrXMvXlD4TRll/dNT
Thy3KCXfQOIuY3exP3c2OUHTF7NEAUxPkuRskVWFWKsSnjypVrp0Que7Ult1hmxqQJlUF7HeEjkZ
B2HiXwLc5V8r/vGf/1QI0ysSRYHYdV1GVe4Zf6bBcaiMkEAnvM0U6RG712DwQrbTUVTHTysvu1eE
2SNaQnPV27Q9MzczO+aYZaRdQAxwU2pJe8Hzr/vFRGZxodusCsleky+0UpnQLDFKCBKYNNW/IkTb
D47uM/I/ckNFN5rp5Vm/SK5/Y28ChcY7RHhPHQGNjdYB4XZZffu+MRvNpmNXApe1VbfwCc75E7qF
c0LPbOuvtOxlMu77kEOQe/iS/Fn7DXtF9bYuaTrg2QeHuRszRLJktzDO/QNBjp/8I+zdHO1Hu7Ag
RFlmecCufKc3G+loRxFbzTPEJy0Pu3MaNi8tKG0K6DQsogp1rgGkkdW3Q+6rtf9ABP1BU3ykvKkk
AaTULS8NO2JMruBk36ptr0ABWOm7k5fLhCxkM7Gyp7lC9EVALWNl0IIGuvqTNH8diTm+i7hh3jRN
/9Z/d6NP5tpmSe8omg6Oa5ZItDzqhMnMw64TaATUmCh34b4IQc/EYIpq1QsFpTmcmD9SwDSh7tOb
n1/ZMn/h8gO+bHsPS/qR9vrL2b52fECBEX2MABZZ2ySIm8J82+YHofOZNtPCgBwlRjClbzwA/qWW
hhfGUFT8IDpTFb3LmXvLyzxVPLfDwYensY2MlpszBohNxTjApQnuLKg1Maf606HEYZHoxosfRIL/
4ZwIgfHEuAAkQXRIvmGUDKnGWgOWYo8N1tb5BSDYicPPlLpte2n6xjGjFeKOqsuyISowkEAfkMgn
jRioInwy3kZZX/0ibgeFuSHcK1FKC6INSeucJxfYJbCI0x+D+P9TaXABB6dh1GQSrs413TeisSni
4F+BBiY+QaAvn183Lgv8t1WBKUBSLlUZJmTjLST2+CmM+tyogdfN6WezPylvZjjIC/FXZEQ9cMFE
gvrC0TfnpUGCRLrlVTW8UgIjai8nIkn5EiAOnE3tkxxwx/PlNiRByFndnz77cDC8PAMGuKvDcTXk
njTa1h4QNNBPAzDfsHzBGNBKf2iVQvv8jkJObGPkkpXE2jDPwEmIuh0+75FgYsSE43bLIbQVAVkE
ndX/wFiGoI6ie610IttScXPgzPUoSTnJ4EejEytNya9vOwvWOYzF3iKzwFgM3DeqJ/qNxa6OSqoL
DOycAeSa06d7OQmp3GoH0ED9OqZVv2T8po2sNc9yBnZioBX+Bdxfi+A+AlQ1FxRMyGO7WVwpDhFr
4nVQgqAXAYk7QLGnekeMxWLGnYgoNpl0u8jCeraEc8rjn/RPjGtVdyhlv0oYOG0KlY+6kWQHrUKH
jvp26usaFFA46Hqd88k5nFLhZa9AtaNJgrgg+CIaywtBUMDvmTv8UlFfSRndOWDjVucmdAAUqu2E
+VHhPvr9hW/O9o7GPnSYwBaYI80n8bcZ2jm/Tg0iXEdijM3D+IRM2M4E24mFt3+u7VCRbCbdYXwu
C6U4j6z/5jJhUjC37Mrpbc/Z4+khS6rNDSwUdJHNblOt50+GDeAh9vt4y+cPq4oQ2uJxFS1k226e
g5VIxUUuuBDcw/5pB0nSizzeNHAfNWvNI8tvOiu+s2qp4u6Y5D639JmQrXNUlwyTLFpdR+icLgmY
+n+dhL9wx6PVpV/idq00yNnev+0chsDjdd0EFHOu9eiZe1Y4/m5VcrP1xVJ6+gQDF1UPSNYV0CPR
vqBetCnOy4dmo3TLlnpm9vWlt8TqD7rO0TRrZoUFUPJkK2znUXQ8LgZyTneh3qw9ulj+p2ngY1nN
Yyblm6hu+9A/4LyXZt6+dIuzugvuCqhsNW5pi9sWcy+Q2l7mY8to2M9LT8Jxrc48Y85Y61XSbuua
jMQS46ZDyofFaQaxeCEm7+DeRn1jlsHjOCGQOdHy+2HaGUSeXwf8Jk2D73HjVwqT/CqcDeOXgmKl
u5z11iZ0dNzaGYZHlQ6RxPGp2qBQFHbwoxiKbqf7wrRGNRPWcA0KO1t/Gk6YQbwB7En6COKirldz
MMdoAMp04J9URXzswxbuNnvYH6i7B6Ts62UqxIzdt72czhPuPnth6vrfmCEdHKjsz74lwnmhJt25
n8ECfoXB59YrhN56Zf0Oef4Tqokbb1gbPcrxvFpiMpfV/xjajdkymnl8PcyaBLsxJ9XDJBWQN1px
x0ON1RdmucD0zoOZQ6Zr8zczoWG4KuimsQZxYE06wAQrA40Cn/0QWzuVWgHcxiruiUVS+WFMb+6a
rN678ayFM3IpLxZh+ppIN0/UOFXzzQ6KEv8bjb7eEyovlQCl8kryRQ+XI5oUkrM7Y2zUH93PSLnU
kQkveu5MkWcnS1f/qL8bweLcU4f3KnmnjsBg1TC3kLtEsVbjiKFtDHskkcUW+ijBKpVvEU7Hy2qj
UM3a+k3dDctgbjzho+bJBRd5zOSvHbgGNT0dWQwkuIV5/54szY3NkZd8ao8X0gkmgZ3sQIBmL6u0
lC23tqqhM9PuQ39tEsJyG0VDmzrbidECUfG9+fCLU/yXWoy7Of/ZG4Li9rcTRPRju9r2Q12lUqJV
e5Es8KcrABSLQNYT0vEEGMFuMOMsYf5yEc62J1tYVRAnXIBiqtAHSAx7v9ZeAhmHylsJwD+boBbI
DKyRl72BrqiHGIxR0C/3DxqcKYcg+3HuhP8Vh5LaaJ3/aF0UFFcfUZ0zWJNjAc7K/JvR9tVgqRYy
vgaY9TDs9dZfRSTKhSGIorZAvRlwHPB1WL9/RedwJAS1pjRzEXgiQx0FRuEzIbNfpJiOosVSKleT
2tDsKxWs8p4shNlDP2DRXlr8cnscqvv0i+iQnEJmWN7wEsHhux4uPWstLB6ZckNqrBnF9P5CQnNP
aRSEcMH3YRkhUKDcQqi2odBRiFk4ue/oc+/e/unXjVVp4zFWIiG9c1pdZPEz3xc54YjB3Ps4nR6z
u8eoYh6EWIn9kGIPmX3+ECuygZxKVHEWGa31KWvNDGATN1mx4XaYVYIW9lFH3X1Ja+yjPngXLe86
/gNgyBGTYRLIZbMHijUJd9EAGcvXzYClKw3z1Db30Z3dYCBa3ax6xh4BrEnYMmD8vRs6YADlpnUu
yrGXR4IRXnCLf/2vJCxd46zj1pyARRdjit9mTpuYVJEiL4sFDcyItb33a2cxCPPOk3F2BYGwb7yp
IuA+mZh3Rx8pibLv11aFAlFpKgHRFyF2gX8BUvYzsX35zc+IMAnegWKdPhWBdRo5pJa66xOx3oFE
EtrsVU3n3sgah57Obbar8+2L++yMzq0s6VD/8jhpoKHb4M8YHbh+Gwf2+r3/kcBu3D+GSfVqSH3K
CFkbT5HL8Sbgc5/mag6ZGKujYAFVbHZ2lUhTH6V+VX+mCdOUbFD4c6yvXVNh1bGXYZru2gzv8rcx
iOpNn2QBTLt+XinQ0S62USJQc9DGawSX7vHs3bsVCuSASBmaXVNyQHEH4xEh50SkTwqOXGF5Nmxz
X3OWFd78/IlqjpNCfbjaX4HNRxU9YiYLqWiPsSVizxytlhsCN4ODZfxl1c2AM5FkcqZQTNPv6Ioc
PGBQDrX40KVhf3Rd9WVQWxS72/7hFS5eS/zZqQwS1QcwRX1PxjeWWGb0a0tsO59TEJ53AbqL3xm2
AJVIqy+unwCbXh8dIC98WSfG5Y9xLtajVtV4vpvzyiKq6cx05J8aTBrdn4h7xQC83Y3EfU8j1Nn9
wvnZer1RYbM0tm+ZWkR/DjENsfh4k8Bn71WnBymYNTQuitfpK6N4MCyNoebdMInuZgivEZxn0js5
T5iCT42Ps5c6YKL9F+g0J4K2bMazMCl8EnK2YMlKZ/R9WGY3l7nZA+efKewRK1HZDUU3FA/YVS7U
UtuQieo8hVyU1hKpFR15w55IVWln+ET33S1qBIMfvXW9YlxcXP6KBfcAsYct5ACAbsgXjs5MP6it
KpVaaeab7/s3ys0+unMfQUQSUd/QMVYjh0w2pUs6D1AUkaqNLeQmdcuRhSxogtoQj0gWTio64R5q
A9FZ7xZmF7IH6BBJdRUZEsbZ32GaNE3y5kJstXT84j0sBhJg1JYndkQ6ItNaW+ivmJJJkv5uSEx7
7RuPH0ORkOWi2uHfEE4Le7WiYHIg3QoUB5etG7bFqHe1aXiGqL718IWCn5/OB/OCYKquakX/LiIG
f556If5XFCiYk9c701sP0oMl7Hh3/4oJdffhIow5/nBHSIglkBI7NkvX/vGrtsD0yiMphc2z/38I
YCaZV7t4y8CAgQdUUbrr1UruVY1O5x5LmLfjAo2w/jn/bQ2sLeL3TlrlAdbJFI41SSa2bpI7ppHE
VADtiSBN8ifJyrYsLu2qHKOv/scejtSA/9mljhsTZkwl831RvTBcahwBAk9wi/0mTV10C0zY+rGL
MWJUSxQb3QIiV0Pi1ub9LoYhzZzCVhDf1I3KaDwH7us5LH+y6U1A7k66YhE72lvm0Srdr3GsnM6G
lFt0abFl0ZAMKdF/R6isrggWT8N5WCpNVj7Pm4vcVupmGXrxRy/9XgaK2HJFzWl+uOPnRZZG7EM/
K1hS2ZJCKRmiC5GtLxN7Afu3lSPLkwr3oOJIeOzw+8fy6Kk+IHHA+ERJ1tbJSUxEPL1P+dUEZqbY
CW3c3ileOY5C+yFNyUw4M+SVUzFpy8PyVrdEdBL7H0ZjN4xy0pT0NhSqM2vMpGpWnwgeB5Vdq/qU
Z29+BhSgM+yQlbSfLYPKOzhBWi0I/vpfy6CYEs65Tu4AiY9NIdYgzUZytu7YBjPb6soK7/8NqwNx
YZvxOwvaW3oA95P+65oM35ryNfaeTJuOMrneimGaGH9BkWEsTKMe7DG1JCtx1nmCqW8Dp9FyTp0h
+6JTZ3hUvXxbZGr0wbKSkvWu02EuH0UAHqHp9+An2+yh/ANLty7wxHLo7NG1SH4HzU/bGghJGEW7
zy1+zpJgFWsNwG90mfupCwh3QNDuJpStGLEHstR2za+3CNIH74QVFRgiFthaUcaXZoyMKBRyllUH
s92f9u/JvLdc4+HG/o115WpBSp83meD1VgucSB32TBjCwdYo1vBV+Kgd60nPXjpUV4NVCLN3VEBh
QshUB7msQlh8y8RTigc7WcgA9RbZrBoJwQQuVFwcPi9eFpOUeJgShZd2NracbqlFDZHQzuLcONn6
BKbWSMJ0gxfdj+cD+lkTltIKwR+yC73n9MGI3+p6Ecoosj405JLQ6EOQ7uv6UoeYQ1hUHV8RYxnW
HmDrJY5znViLd6bpdWRfqkgSWIaXEhxI2m402uQ/EXgq+cGb/KmBFsTn0t1ozIuSUTaqb9bP0j+v
EVNC2I4jSusEO4PoprfwwUs/osdCfOfohxfMn1Zc7ghMlE3KQNpC9cJp+LuVIkqo5VNToK76AKfq
VpsMh/39o3pU55oa+6VKM7AkF7802/OvQ+YImPY4Ra0Y+OwTOg+VB/IKL3Fg8kW+DbOStx9Pqqql
03ianjun7cipCyhONaJQqi99vqqtcAN8fM3VVJE4AgupTGTNY05YYSILbMoiATPg7fGu1NM+Qfb7
P8isZxp4eke0mX0Batrh8zXMYbb2rYk7ik+0xPE+6bX4UKOvYEKOxWD6x8sXoewutXaAEaw/bBuk
E5hdeC7qsqb0zdBZKTJKL/Tnm00wfzGIe3orcebDrwLxjF9D6gMDjUu6LqxtH2B/JVgdvqyzhWIk
eCbiMItNJBuqMkdjHm6baR0PG2mySfJ+G+z0UHH4ek3y7wuarJqpOycSMfOtWQJJxdDv/l0r/w3C
ukF4zc5PkrnUr7o1PSIWRKiiQn1eb+Hji4Eb38y2uAgOpSLtyShjIfrrJG72puzyatRC8yIRQDgK
ovy9z0YkCVMu3bHoX6ulj3G2Wivstlv1NN4NStCLHED9BR7RciuP3AFb1xjwVSRaCvFBsQXPESsa
STo6yxOf3kfLxm9v7KfzkHMwna/ftGc7IHv4XJe3mBH/zteEjuUeCPG4PMWtGFL72pEKe1xoNZGD
vTXzd+/yPbLMO4P/Akut89QZ4s0PqTDvwFnLL/PLnPv1S67s4Hf83/Kse0mxfxYZmjQtU3gv/r+t
eq0eI/AhcIz+e4ZfZJadRFxVuvyPJTRJk99v++K0+3EaM2cEtNQ1CsHYgIrErFO1tFZ7eLT3M6bq
2v+48zgRPMWNHfbCNf9RIxLyC8hyDWQk4kKsESQ6kJ8vRydRBWhfGW/oG7m8L2TyQRqa5A+nz30z
EWaFgV01xrV53XLZtQPApq6NHOLN6wu1j/KP6/saUah9ZJBciSTsZQ1qYINKwC/fFZjJuFkPq2u5
a5KI9Jt2TA9q/vQyKQOq9ewGAzi/3vAR0sYj8O98mVMtnbAGbD6LywAm142B88a41cMroWdN9I81
+mxIPKukS4Lx8Pp1/2dAtDLM/DqmO18K1nACXz/odg3IeWc3LntlAqRNwD9hpRGn+pAPYlYzTWYq
C2FI8PDQ4nce9vxsbKYLVY05zYwHGLMEYvLL2Thr5A9fnTlOy2UeQrqvhq/VgPReRp2sL4h+X2aH
ZaSs+rfQksHcq1T3gNtA8Iagn0XTIeE0e0VmTsHRo/L1OHXjSmE6BZYqrTLyp+TLFwvDWbVCwqZW
jyTSpnqqsF4NEpxBUpb1fI5AF6eZETXuvxSKAL6hkScFMjQN4pL1Q1bImYMJB1H1cyvS9GjgU1rO
Sr84UBDw/FuokC0E88vy4wKHWRArWKAn/40KL6GVQ6S3dPZwePOCSFFepcO+9opNY7bnlA3CG5Yg
dcB5Eph/LoQUcNXft6mZhthDtHuAt/3+BwkERsOioZhX9migtGSilBx1QJcBTB9DAqUuj3jFxyaL
uW0YZbDjWHAi1SbYmwJ+3CZsiwe2yeOdgQ9cO3URWh8MHOIdwpI7qQ7cmz7UvGovOopnsBdN+x5y
bf9bhNntU9c4QrVZSGfz+rabUo4OjnaVEMOloSq6RGXSSN3V4SDZQ78iA0SybOXRrnvXZe16e/HS
KpYY6qfey/LQIU2jXjn3mkzSelvb+/39k3S5tGSYMGrpYM45g8FhJ6zXAGp1z6JMjA65sAI+8i5D
CNT4YPFl77+tRy8XtrtiAbB/0oqEpuZfaNBJxDyWyW/XeQUF6gRlrPTV7loA2FnwHiVqp1n/3Rl5
5IZTBuX0B69/QeIQ6Bg0fZojnANcPXwCfI8qtvsqU1f/tK1ExayIUyohcJgYR0vJ6nTZmkmKf7G9
y6OIdpBvFcFF9wM44IrJ2pOR6NykjRQIF3ZeCcvnzxWo5vUEwOBBzPt6+Snvy44GyrYSX52DsdFx
5o+3ThUz1xC2Lx52RhG1QQ6AF5zIkNwaAvBnFmhlBf7vNaddyfSoS1hhMrzFkvvMf0m7R5+HFoA5
aLC9onW92dwHf30+ZGtWCpzE6gAn9hcH+TvZLz+8U9fAKgilIFPCe7kRNZF4cCUuvVpHIcEYGV2i
fG5HGVvdKcBeDSxuAVaPRRil9ZBblorsD3PXkqWZUvNuU9c4fr/cyClpWAFNLd1uPuIFvn08pr1K
PWPxMUN6wzz2UbqX955nG/nmDIw2kmJl6Wwz+JSVqNbRUj/vyyIZtO6brqVRjn5VqPLFHu6fzKzK
0B5z66NjjDMqAuqJMs17/D7iemoqGmvcR7mgmBPw7VFKfZ8LNUjHCgRHtOMyNMO+vb2X9d5FppNV
Y4IT3xJ5oZIlarrOsm+kZWPI7xiOgc8hCIMQ7SIVtKzNfxaYyqzRfwvekvfKfYqor4En/4qDEoQW
8w+wMaOwtnVHBYpV6QRJmh7921cDfWgqoo2ZaAfl79p3HhpAG1p6earPldUvcaJd1nz3DIw5UpTd
hgSOmbO+utClI1QA8HKuwqmC0xjmvAN5Cy5d/qtZg+T1fjqxCtHWBRi3uR0NMLglnd+bmBQshk2l
Tt2Fg5Qfv+XOTAGuZKkTzMD0+QR0NLU0+RQDUEy4kDSBBKpE3QvFzg1+GfO49D2aDC8QxQY6TNuP
2uOc/Q/9ielegdJi9WrAh37CdjfQCXGgbq5y0ja+FZ01gp6QTN5TSYvK3nBL5SmJnsyPRwOOWSsB
2MRgj6SV2Aya96h2wTgq+Ude+wT8ZaQbEFhIYhpQIt2632RaqKqW5GgVcM0BqYsL8m+BU0zczFQD
PKRyIPLsUNzrM3Mp7z7w8hwH8hRwHykedoyWOh6rtdF8PTQIToJbBGEy7VmGmprrcE5xN9PYPMsa
hVkuONRWW0IjdQJ7pi3SPsva9KorqKEFD+q5vMpMfGQQXN1jCsIb+WYPXvfwF8kdY31ESSefPjOd
gbV9c00e7zG0wQiN2LedkWpI0Sdwgb7NXxedoj3gHLs2XILzeNWgUmlnKQ6r5WGc739pxn+IwlVR
/S8u77gABhrOD05EXragYUH7Wa5rbyCljZbC+QrNZ4E/jfvsJ7C36bci3y+pu7iEcvRf32n0T+23
MA7v8kVS9/t7dhIayvo9UXlj+wxGMUPr1krVifBC+6qKRCxmZaj0x/YpVuUyGLPmqe43rP/7Q3NF
nZvfJTIsY3UNQfIabnoRZuCKM+MYoMkYoUPxQ9Y1xsi9OejiJkVt4Q0M/AbVhBi2BFFb/y3JNFv7
P/Y4pYKr+Ofv+d6R7ERVS/juG2r/ED2eOKVaA48MqYtZ+mzGO5aqA7S4dKr6bqnGHJissXEC1W9/
OhQ2jMFtIXRh/DExVh+B3FVG4FGdoBkaW9r912DdqiorJwMkCyrmN1lZ3dMXlc+nJLOnKeULwnmb
Sr5ebUDSq7MUMeVjjdt+lRZikRybV+N4D/X5va6WjRltpf+8kqxnKREwPlOpToaFUq3BHEO28qpZ
mIm9NYfkEXEv41gSJVIcy5imn+IQlsg3+O1nyf604BOAKf08wdrvbMY4q7LNvgmM2Bra28kTJY3t
PaDfGjgG6hwhunXosYQ1DLdaUXPsFc/3gLvAypeJ79BFH7AlzWXu4PHGXUcYBUbYp6E6oiAnvHcT
WeGtRINOYbKKAuhEbsolM5PO7UFA/UlfxxAjsIJgqH1lVkIPSHuFO1GEobM+e8LjOHiVFDLfXMhT
PVe/V26PEixGQUFa7eL9r9geDVeZd0sBEvHkbt4h1tnvPrCvzY+JZK3cfl/AWaQQ6hB8ysZI5y0r
LWQMQr14R83a/+/xih4hgDErB/Y4wnnbOesiYKvnIrpU4om06O8kGIi2WDEHWYwNvFuuomfOSNoz
T6HvtHej1mA/2Pm647z3fBJKg4a/hJPMvnbKgdCbWUHmsekFiNtY8DtD5P/32DCrjuXvYjtyUaVM
JcMF27q2xsgyG2qMHR4fuUNG+IsnqL90e8z+iTEj2XCfr4nXE7hQWjhpTAWdhYup84fMNtK5VAjH
aryJTPnPw0LVYcInKySHk7IVKWEQSuWkgew8uXVbOCwIFLnke4sJOAYOyo4qyn6CfulVLStxGfSh
0/fLQWMtcmCs0Q3OCqz4syyIeNaJDUSC7cHHrl89ZqaAfScgNF/8pBfsFdtrQXUwZy8Ahrjcki82
rkOfqErhnmi/8VWasNrFzXbVLEPjgkKqPhREY8MoK53qeMTTnCUtYlVxq5fPkUjGo/n4N75IDsbx
6a9UYaIHSaU040INv0lKB8JcZXqPON+56SIdj1kpkHrYfRxOnMeO8VlROS6Y+mP1BKo//5UmN6Qz
hQRs8C6jbg9kGnaSeAo0yvFVG7TajDURm7lV/CxSsx+TYWmzdzhitpIoMvcpvbIC/ZnAs2HQrf8i
t/fGBCxlIGcLV1QLXxxhWjgURclaA9P1o5D8SBRy2m1OltD/TBRtYE0+awIt3qpPf/YGq4fKgQqt
8mh+Oz8aVDWqJiwK3M/WWrntSmbZEJdRnKfHRRjgM0HO/Sdj/TPTwmLNqxg9gs+e/BEixBhT8o79
Buv6N7qVQhRLYO6X+zJUB7KARK+5lM7zGiK1AKeOautylRsNc+BiQRNh5CEQwmip5P9mUZbmdvTC
pwk5f3lTj0FUqtPVnBFRd0rixfNHHRCaQy3EINHXEG91WS/1joUjHuYaWWR6VXMX4qFPjHxupkwp
bWVFH2CtLsZmiUA3P6xdTJkyFsTSbl/4eD80KxAmvhT9fM/zIxu0E5R9vt09+GSfCZjzs9HscdR6
98WNnCQJ27S+eWTY2bahQyEsO5TEG4CypnxgP2L8bEfYG3U7cQb9q9irYsE4DVX5pCZbYK7iuJjG
5GpwVyr3IghdaLJII5ZrzndQmbXzz8jzQLwcBIqWF1l3cYBS2/JfnXHJrBLx7tYYpc1uVipKZcfr
6RDQ8xc3YhbyW4hxavhHsAA5VkVL27OBnjQleQdUHC41Ev38o+H+sop28sNC+LgiaDIvLzlI2utk
XlSlOLs7CtWeVuoBOyMvsSUusffd7xHp4fgM1n80AGNaNhwZD3WtpfmzTXQWG3LIJTZcE5OpoJ0L
0qlLK6mqiraB3tV5nu3p7SIXcELCJf5R/Gw4gcPxyPlOqUhyessS76+c86WEodP6CqMCXfM+RYvi
7L2xiFUo4rZq00BgG5hCrxGaiphHvcpUtsmjnr0jHaWyijC28cZW9YwpEE9wUtQiImsEpxroAdFf
Mb6deUCRc57gIb/Nv1tgpXrHgMR+8K2Ct9VYALgGnuwmik9bHrolbvhP+tAT7rMqjWDFhxcjugsg
2O7CGjmYlvHgHoQ+Yoit5BVJ7DCUknduR0JXvzHm58B8oOXvQEXv1C/+KhxV7z0MBZ5OjfomCTBh
xqKCXXSLbXag7aPUNZ++YdOXGBVFVN8F3ujvw2FPYTy/oqcUBLl+4lnAshVqOPi17PjwnSc/6OWp
S7ZcDNWSsNuT6OOHrt4KtwTsG194ZU9u9ONg7Cs3SimEkMi2fUZqdiH9+jdqdxyLMEEfbY7X3E/b
eORriU9JMKFC+oh/xfoKsVuqkM5yohaAP6H/kiR/Gxsiip+w72+SzmH8J2YqMlXE0ZGqNf1U4UuD
A/tDZLa0ygPzvKu3XpJ2ffqUn4CAzTKy5M7bkrDAtXB5zMTOQXg1tV7IXsa1YxNpI8uF5unMFWcU
SGjJoRkX0/UBgnS58pheC335hnzw0SC00BLs2dk7DNo1KmfDl3zAfeU9qaur/OLpIJhshprZZa9G
ajvCWu5SgW7upI1qUJ3/V73RiYYYscph8sU3fJBPSLBwYh2eELMq/+Z9qQqwHQVIT8+CY3CseGT7
3cA7AwVBo9ADBqNJVk95wG3wRi5TOD3g07MqkOCYgvJfKjAk53zZZMq0Nt693MkLysmLnWWJNP49
PCmMsbTl46V/TDjDAvGJVAGIEOQaNeJYI7yNfI6aNlEGEY9OvkA/pgEQm/kIEKKcer/0818bKHEW
/YKssvuWWq6O2OKs+cENmyhdT/GF1m838zDZk9mhEkCylqiFzbP02SijXw1eSQ3ZtbVbi2QtBjGK
eHJ4iP96Py6WHba9+R492G5pmJxFNScmw6fVUSNdlGfjZxF/ji9billWOQAAi0piZ6iT0Raoe2Or
rbXHCUl/mkooaNi3XrZIFYFgSU62zTIf6Q++r5mdgSriu+dUd467XLDhAtC0fRs2581az1zqIEi9
QDy0cxo8FMpRmCtZcIDlJDxBCsG2Zr6MuQiOtGZsR8r5VhjNevdRWxzQlMYcJMOy3I2FxDVQNZ6d
j+cWYLhhSsfB8Conued7s1CbPZoImK1xcp8fObrHyadb+vwXWJHCWbKeiV8rnbMIBFlji1wezX5T
KRNufWxD6iMsIX7lT5BeHgjGz5PkPXOGJapX0h33BkZvj6pTYGRHUmHWwktLJFiWeJTr5+IP8U0Z
Hk+NpWooxzlIWGbnoj6y9z2yLN+3GXJK7uBvODlNks58rZmcji7FriqD4OC8i5z+Tf4CpaXK1lEq
CBRJTVHqRitD16Nu0fOes0Bt39AE5eEij4jkLCBKxkkV1fn10XW1NL+VTLTX3wpEmjvWHFdigDij
ELdutGvV1PCGIi2yQiGruv5xyzht2o4G8CdcwfbS63+aUVgVgXXRf4Jeg7P1T84POKlaf6NkAt3f
50Cmd6hTYW+pX3dRCrhw9v4KzZKp/xFUBhuyQQszE1IK9o1+F4Ezj+sBFOLaLC5BZW762lkIMGXl
CdHaeXzIW+JtGF/qvJswzatRFAlZ07icJh9QlJ/wt3oIlhIWAjxQJVa3ewhib2bj3s/8t+MweZIn
NZi/vGFvkRQ3+wv3lq4jZJF49Op1XiRqpstTnT59c4g7WzoYkNy2okk/mbei45vYqPitWUV8Ny7H
LLm2Wc/7WXMUhivss1+LOFA8fnkPWoSiUpOKnsXnnqGq7etH4BwW8pil9I3raMQezeig8sOEdgy6
qRCiMoEKD6W48rKjP8nLknA1GatLudF0TN1E98DzrqQHOYzwtevX180SJScv0K1Pb/cAMiOT84SC
AddMkzvlLsLTXlm/5Nof8iNi4996HLXmx3daWvIm9jdctbHdM2ynl2bweDnzJhLYyAdueiZFB/bv
SSjrpjVJAkWJiNprAxNruVhYPf7slj8R4WMtZyaedFefTTIw0+DzbaWdLoS/6yYpzqviEpYgX/AG
/1YKasTmeQPIa/R031ulNTlmqmwMMdK8eK0jneOGEyf8z/+CaZDpTzsFC4l41nlH6+p39DIOGuRF
1sO9bn7WWOFjFeNQXxQw638WaD67ewf5WpWPi+50HWmJFJLhIcfXSI7pe0wSqlEEMVg7B030k4Sz
kUwWG36P/lOys2aVZCTyAyfWHA81YKoH98k/reJOlGOZn0qZ/9X1HZdVAK6WSc0JyUDIPHQVS/H5
hdKFxAuTOOs9mLpg28JOF0CJgJLeK+Sq2fUmVai9DjmPs3jryaGXJTPWktCTO1u5L6AHx05NKQT4
n91OEX588A7sP0GAmrjVF9L//JrE6FAgOw4XjS329wqd2C/Q7wuQnZ+dV9RMdHbesTw0A1sZEN71
kNbk4U+mPrgmissHvA/yzjGe+vMV30cnHyNV0NHX8X0qPgxqxPLZpMTttock/w027q0KI8Y0x37l
VEw0OwdtQ5yMSeAuCZKmqhAKHntnYZCzEXzcoyJ2LRcIVCe3NMi2yJ2G9C1K6K/4TiBeCpyQ65yG
/dXADKMa7Gpv2c2L1GCD3HzWATIfxsu9vzAtGqZHvY9MwWezx5doTo2YXVFgCstffBmn5A5POSwp
KJw5h3WKTktfZMzg/Ht1WsQNdLIwayTImc3E0Ua+cMvhEzT2j/zIeNNbEm3XU0ZjSTe5RqImBZ3A
TNlT/ISVppcZjaUTBe/3ljlTTj/P2gnykxdmGEptFmrF499lemA3t+CJo/xBy8geNDt8PZqdSkpv
qeIcfOY+9dtbiTNGhTv3MtxuwXCIGQ7lwoSqE77n7tdEHJ8be334xpcw51oeqom4HIvxH3hh4IWC
OEvfyQHrMRKfzBYbi2RRWagKnZ3Z3vV0XsmGg1gNFbAjtW2AOFdSCO8axVrsdcapBQ62MsgLn3wf
jlpG9Hxzyq5at8zfcpIHXiZpNnvpUZyeRSSzrzICE7c3+dpytO8VN5xbXhQ2/9gxzSd2eSqLUxOT
IzMktnGbd9uJvbGOWeWiTF3lF9cUnkJhV2pW7MTrWMLeLnZYb9OPKgEb5aZzymZ2FvapJKIlVO3s
aopw1z1n6QRHzuNOCnK/baK5Ae2WkBYTi27WIgscWmIP29KHm3DbmMM4MjQ2J+a5u8HBAvoqOdEd
GDaFkjN9xcF4Bnwnh2KLJtn97oyLnGz31yHbEf78npBgZ2h2emDY9qA8K12MszmaCP97pUauggbW
tCmjBZKT0cIteM1agwfu9sajf0g+1tkkVB6Xn8xSlXhbyfScuqLyAbOQXir7PcvQPJkLbp7XCRqE
DFPyDSmlUFTOyMY3yIoMsUwJMepAlHCbHs36g59858QWy03Ps+Rign9zDissFqT7ruDCw+Xv+lFr
1l6dfOHKALRGa3al+t5NOXjEyMHwWuCJ4a5+ih5rE/71KlWQ0lcwIYP11Cx3pRkgqb3cXtEeIkJ3
j3A6I1yAtxTjiY8QpnaiYI5ZgciQEVFoE6qFlHwAauaN8NMU5YhPnHmoO+/MoiVnMY1UYdg5817G
756qkttH/e1pkzrUuplzUmRCGrLf6N1wIemxfvWZpXjj4UidOtp1J0skDTcR24mqmIJ2H16azxoP
o/DjLIvyma1vDvFSsRJw/6NNXZYOTyVx6CHikRtIPw/Wz6PZ9QCLWZswIpWRZrnRMu4meMvt1CZj
u3xb+yYqR1tdwJGnVFLTn80V+SvhIwnn57G+Bla/lWScY3YFrhXODJpQfYXaeYJ28Lw0W//1HJLg
opgRXi3kLR+EJ03v3IJP5JmGwaJoj/vo6Bj3DNgTlEGq1S3vQfG3fmGhfg4cAIJYrikft2xnjcU2
10ew3kEcOHWXXldEahBD5mcUZSe6KITPzfJuLjfVGzUI5F0inWt1zH4qcs9BAoaLYfHy/puJFfJo
XbOSfPFzWm4w9bZE2vlDfQdV761eWhVsWSvS4mDBacyTdIxiJd6Ytw7d9tQP2eK6FH9haFNueP99
Olib8nBLK5MkXgk7/P21xqtOg1VjMMjLjZNnkSH0Ird4gYhXwLXBFMEipwZc1K6Z31yRHjOd/DF6
1yFHRkpMZb4Tz4JllgvXD1nIPJWeTVV0h90CfTjEVkSQ7gRKcpgQ5TNTbztBqxMeyOHjPAp0Z13t
1VuqFLCawgCaFxLISlREqxQsblsZ7zes7iS2/DPAd6tjTQqrvWt9Ehbe0AwLZp50j2DWdhmAdroF
fLEljEiyDCpsLwB2ZDqhz5DM/gszkO7bINZMKSR6PMJ7Ke1Lj4A7oI5kUCfQTc4VdNdOcvT9PMkH
+TA9Oy1WKjCuMbHA41oFpwtEsFuCxIF5owPmZO1JL7h2Det06FKxsyuv0InI122Fri+/JriaCfYq
+19HLQKjheOZdjRAwdCFLZ5QQYA7CWOqDljBlYQ+LZtqinWXjzgsJgs9Ia78Im54FqKmR/USmXal
OQX2YVvQq0XWD1ak5sYZPC///i8Wl7C1Y/nmNTTupYzQKyRy6+U2EpntC/CNIWc+kMbxYyg8T9N4
KFEPZ4GB2pSm0B8TqEb5UDBlG/pKUjthPg9tsOM6eXZrSfxsNyCFiUl9qjSl4SxyOxxq1nw4W6Zu
yzO9Fbbb+JvM1FibM0g4HqHkQrR3KlM8FQpXDeQ43Tx8K+a78EhlFnzsDonUXtyH3l9vin83ZF6H
HKSVj1bzt8QtU9lgSe8nkCTas1tfh3p92O17iIFjxT0UVF3DvQDaNh/GXfz0ym1yMameNnXXxGU4
AXjuvKjbBI6rbokGriCRJ1A0ALG/2vUXqghgzvmfRTGHA4abOPKTz+lhALnudktELGJMMWE5PIlE
QDLnax4wER3kTdxQlzR2VHALSnUQE9+VVBL0vYOLtu3W9kBIGr+p7vJ4opmlXv0qSS9RnyB94j1g
sTCUy+P6zLO2uGDppzXot7AH1qpAeb9d7v55CkWaTuPVyk7ot+disIBKG8Pqg/Pi95JA89HZYHfO
EcpTJowCrownChArd+NPw6mGavtfC0M1isWpKeeENTp5xFSbVo3O77oY7PRhLSlcfCTOJVTzpl0B
9jUrFo56hr5RhjStSveetsHGLSwt5prluZIBs//XUP3IWXE1OMx4PAcF4eGJ7TRoG+jrI337P+ir
paHJt11gL6wOPEpQrCAB2RBiLRUkcmse8BcNA8Zbmxbr9WkI1MeGPmSD/z0pJOO1msG0RccWE0tV
GNyUHzpIg0jAA+mAhFE6czwTExEMNZ9pWZuEmIBPz9JlhWuhqMjYX1NV6edFSSniQEe7u60zrAeW
HBUg+Q96YVkXrAa9EHQ3fyO16Fxar/tvbk5SrdnczsXPBed8Bdj4A3U+0pxSKLJxkX+oxTajMbqB
dlEtg8iyZLr8RUu7kTcptxnFgt6npWodqffVHxsi78OAUAUQbnd9R0cWt0vp9H1sv/9YsFk/vjfZ
qgDVWyF8TlkGqVnRheMlxglwVaxykVUiz4ddW7dLR3DyN0B7RffbPvkfFJulI1pwjlXqFcTwKZ5V
0icRbB4udgd617lgZLBRJLY8FtqWMIhgSF62dRifwbv99W60d/HZtHECMTzsbRG5MQNb1FSHg1ey
gj1Rtip1ZsngFah+u9crp9q6SHmtZl5YS6mYP6VHS8dzfeQH7scUjLVNnYQkkwBUQdWDNvVIzL1C
e2p5m14OyTvXHbaChWIqfcv+WkBYaAEZhQ5v67gqms5B06Mp1vouGCWSwhUpxK96n1Og7pq+meFO
qg9kYd1skmPIe6V4KsKf9afW3nY90AE+pOe+TnCuDHgIZy7lMCPInwtc8qzeCYusa49ihfb5Itel
Ef/zESR9kcDEuqBtkV3NumEgaGeXPJH/du3q699dXBRYUhmgjIN8J8K4QKvfQyEw/8Lpzptn2FZm
N5Y3ZnrHxDNlRRaCLBr1qrElbeMzsl++Ski/Fgc703EMryR8teDDMUZJ+UCtfhZQcd+WUs46whcP
1cItZmU4m+2Hu8MHnsOSf31WNrvGrgMS28spACFSW8N/EjHL4QdfAtVO8+ERO4Uwo/0LO0XKiCsX
d34nk4qZUuOqKr1GRncmQxhkWIw7/YXrqb8uNKs8gGLIUwv4s1pHZvf+RTelQL6bTxCdibfR/dfb
+LJEGBYLDo02Yy73ghQ9m+GYmVZquFy/JBwIInEtq8JbvvLzmlXe/maViElLvlVprCZ3LR4uf1Qd
cBuWkjR0lJGKtmg0JfTYc2dP3XMKajLdTDTq+Lh3IioMTP5hIe5N8QImDU9hnsxENHpV2sIF2EX3
L6ZIkxIyIj3wD9PURzNo41f6UaVCFwVi4XdrOPaExRwy4kBtBMdvARfUglQwyN4SZcpBom0ipf5N
p/01rYlr37UykdQPhPJu2otnK1Qq35PKiwtUAfpyy6ficdwcbdI+jJJScSUZrZbPNViQv+p9G6xj
Q23a5cBfqvK74m8ghGbYSzJnDGCvX++c96GdCZzzzDxb/ge0F7mwI+Z1djWTDDD9ebRBygcMEFEF
uCCnQM6iBOR6Xj6vH9/1asJH8oGkrTPPbTzHP7e0Q+8lp2pc6HvNFbY0I9oWZSLCofUDcuRsKIz1
vDbbeRzWnMcjWz+m2c+7X//AxldW9RH2goHC7deCeK1oP5YbHAhhvQllduoxA133tdv67M//NLnk
AKrjyuMeIs7hkLI32rdxt2O4nvLoO/LND2r6G0uHtbKHrKRI57YqjU/i/lxqDTmmHDg10VaGMvcR
7qQ1vzRymJ3YcnptXWecSTnyCm63m4Zu8ZnRYb9LYrl5UeNhvASGkWsMJ86VCaT1MdBoak4GxInM
21B7S9j2Nfgzc/AFijgcuH/wyervVV/XwufVYatsJxRT/ddKBvo+PpI8GaFqbzWn6tXx+XLnxELr
PXMpBlF2V2ZW1jZaflHhNkjELw4X8tD98G5nPIS72OJEOBIj7iI7EJVMyJ0x5ZMA73Z/Ey8RUd/a
7/q6R3/1oZkNXouixNHdRvHNZhb+vaF0upFBTFAgmlXN/V3T1DkT8a+M1xkYlmwzHheIVyTHY/nG
8byDAfbOxwnWWg3IvPsP6gvxVdKozwAqMvGWF5Efm1akN1hV1OqwmE11AhRPcodYXa2RZ/gmUo5K
Hbqyd7TWl1c7+JDrG2OSIdC7bvAQ4qBQ8Pvo/REgpHBjWYxhHMLCZzI/4UsLxta//ALjG5Sz9jQI
liFxJRzqF1wqjlSQXmzIeX7qVSeEWxKRCZI2aN2sAXDuSu+YooaZykRNufon9m81+qLgF7AS8vwB
nwHz53VoxHOj0Jn99Pa+RV0eA5WTOsCe643n5es4f+T7DoC6iqh4ZQJWHjpAvb5NlM6NSo7kR91M
V1ajKb5xZNYaDuBj8uwm1CRDwOoDeCut4VjL95xuAOcUBSs7xzsacz85J00ZUIUhD5WCEV8uWr8D
dFaPD13q1IsDyWAYzwQJi8avv+q3BNnoNqwAALtRf2bIUCF3/1ZF6In9+GwmYR+WKIPuipufmNBb
UBk7vqXLN0Q7ID1scON10Id3Gh0bVw3uzrifyAeq5wzoSs6n6LHOHT3r6kSgCp3ee0JHvErFALIE
o71KA8WVy9W3zyYvaFDTgPiBzW8hU6+9FGg4B8iLTOylRsUj/mB9ArJ/mWa1y0mObjk/u2bYaI1G
kMI1wZVh0n8S7Pp8ravdp4+QKfhNNaPGyEGWboaU/E6balb4pjLKY85blvBuW3iSBb4ZjeISRGN/
2UfvaO3RPkhlJDO7UsFIgCvKF5yU93McoYCS7Y1klBkEvmDe6wEK/TQjz1alzHyOJGsQr2zqeqOq
gxuAg9+QRrslewhXZIe/Q8ohxa0Na67xadC3v/yUzdzn3L76fWI7gSrUyPLlK3KabmcbHIqjozwE
5XWXcOwwc64Fo0iQmT+uXhlPt+Oyzjaj0duHVgW3PyA0h/8hQmWEkAAl7se8R/cydI7+XgTp2suT
9Ud5VFT/9LD++e0eBLmkEGUcH6rA3ZI4JloMz9j73OyZq5DZ3kY+S5xkmBcYNy6zrWvQZmJMZzAD
XTVznrQ+WaK3Dd8qHoAZ3fqimKs/TRZEh+K/gtX7B3AqnKofErGlz9yjDRTrTNQR98NWpJbP/mDc
F9OYQYAaxbSBHM10k4JXstKV0O2MKRwGtKBrgOBO7lqH3x6yXEPd4ngpcId3K7JXx6o7p5gn9C7p
rpyIaDeGpmsYOIYcbrAJoeFwXEaK8+wBG35B9dVMEQGNv2BBMqSCITIudrTi7bx3v/kAFtNGLSHd
Sw+DxIJPhB7bRB2NlayhccZZTsl1meOfmaZz3xitrjr1SMmX2+7RiHurQjkzpXETqhdcBhs33ViV
OI/dwHzL3e5cuxdgB5rlyuIs64a7+9ZH+eintYlEopoIN14kh9PNNxN4u4x56z7m2kK9rbDfeuvk
4gCVV+rWSzxZO072K/OFkOLUcufWq67nVwwaYm4NDWjxxIT4sHYlKJPwkfusJKi30hfNj+A5uY9L
e/RfxGaTcJaM9XMpysrybbHEQbmHG4BJpATQ2ElSm2bIroEOKLmCVfo4/RFlzS6Mq31EoGjEvigU
IeyxyX7ktTcFdV1yEFICbUzVBUDXhD1tMPeHUEvvQlKegGvsUrvOqniceCRt1LnEkfT1clovoYG6
Uq+eXPy0r7gPB3IOGf7JF/bjTlBuHVCVAIDmssVjdjWF24+B+jJKKVj4mz3G+zO3O5+j8EjNBpiI
ABmj0/tIsmWnziiYaZleTalFmSH9IRal0643kHW7DJPGqeVu5TWlGgfsHfuH5YoiQkYl32RLSoHK
VTn6v/ZdmoriOB9FYrYEh60MyyLSbI5fP7TFxQZWI/T5Iw9n2AA8ra/EaxMrR4Sfn4hJ4KnzG8Fg
7QWbNwGgSOXYXxzXR+m00nMgvcwJxvclxc4vxrJv/PRbyH31AVa0lOcg6GtChFTbxbrQKBndm39g
Nv92tPJnLbjiKF0JIYHyn/PRxb23S37YAlswbzowpBTegfroBX3EqZfj6OlDr7FsOjdSr1fvcxR0
ul1pbozYPtwu6PuxE9l2mVa4L8ZSmU1D7+gFRSJf41YQb02GS6mPI5+qhCZ0S4qZwlAvzG0cWEb/
6b3PUG4gA1E9Hj6+4jEYPT2Na6vfpFD68l+pmpAlTPgxOPE33YU6Is7pE/8eff8ajWuKcERu+jcF
L5AQdJ6mi7/natWuogZpyvuWplfNpTj98m332wBzD/7UKsAHEYvoXsRg+eXd8oTUsotlIkkXRL+L
z2+Gy6l0tLgzYPGd4NZEQidYNzjSLWs4HQwiikDFcqO031sfNYgc8IZsXYP2QZIq60i4ZLljtYeO
U+rtsh0nvrXXQdeBb0BPkwgm6iq+wqAcy2sQ5ZqkoeRh7qvb5Q7EbhDYa7C9vKWZtULzhmO79MJa
KP2Mf9KnTHSC+ySI+B0CVvXeWqG0LQdPO9YAQRuPDXjsHQbzUXCOXJzt94gEw7QdVNmydPPLMkWo
1IlZsjNYnDE/y2OON1wEH7PNXOshn1bpBaSpRWIJiK68k4T+LoF+rsStYeyLwMx3jitKzAdegvAz
4RpUmiC9OztoEhE1y2VB7h5eAIS+lWC3kiBO/n6uR5GNU1kNKGBSymFvCDVvhRVEMs1JcGcRNat9
n4i8/SniQlkXXnvEwzpQGj2hYb4hFvHNBX1CC82Ig5iowC3M2XjOQR7BV/bA0VnZu6DKCqOEsWJD
/fc3nId0IG2WHz2OwEfkc3/3245IXwtp1oQ12cQanE4W80K2KAlslDHSY8Z3p+jKjxa5qt9sxttY
2DhoRY4auDKdcIWNxkPZzlP9BK+6KVSdaF+y2jq3NnO+bskBjpJ8vhJnTNzHS2cgwfKv8dZn5wft
BYjXHR5KmwbCgrB0tGOgcffsErLptwBU+9TXtMMcDM1BIwTZyNBvTS+NqyU0Ys13UjhIM/2XJNPH
nmHwOc1gXWCbSDuJRYOxXOdr5Ka1WKOPm+85k9j6ios3CWe+J9hv8hFM1CitVa0Gv3xPbEAEpsy/
gUSO8F6grpiY57MfuG6qT/+eRiNKOb4smE/ZkpEGd8eBouevVzh6FbcZsxMP8/ryhaaR/pF4rDI4
9Ibfg3H+pDWGN+ZBZXkBje0blopnZKuDLDiGj0Ce3/2CPZQdUFzfjFkYFG+80c644WHcHTP0pi3o
0tQVQ3e4CPUTn7rIHtzgxvn7jVfEU81oB0nE0jHaKqPiK3pc1FfAzY+CMevRnWsUbQKCNKR8m7/s
b5H8vVRKjrTvAxFsoa6ICR2MrN775vY0cXAWAIpcCMph+aUYC6NnszjVHBvszSBklvROixvKtU6e
hrzCOorle/dVyGdMTgYUoA4NK1eJYYk6dOvwIe6gitpmCXSx4gLSSdbJ2BdGKDNUncqz6GxTR7GF
2xD8dzWrnvIIvNwhLYIW4TZKY39cwd8jKtqvdoKcGOrMBExZg52f0w5arxk5oVi81d4a2D+CW4CT
hSpqdBBSFDerJprPHMtYbChfcmpOePP5oLtXPcdUd6Pcnm4c3bKeBV3U/3xHfWg9hai6THDMKq1u
XhdnRmL4QH9PbSDwhJcgqZdOyfrqPxALyvWpXdNTF4bT9u5HVN1dLrlzp2HRPSUuJjEmAXvLQ6lg
K4dTGhItzMH33br4p0aJjeimeYRQqYK9FOW3itU9IgTf3Oyy0jSNl45Wl7HNaFu5XxmJC7HrGBqL
uKnWAhsI6h9ormISC5apUpUd9ikk4tBhru9n3ByZbmOICeVg4xP6LBbnkHfo986pRVb3z4o0Ucs4
M9VWeNxxD5yy8BIlKQb/JU8IsDiNEHRGWSNwAIKnhsvOr06KngOEhMXVKO0ui1wYwmeTY7v0t51J
rcB7pn2kYUEuPOrFY7OWMakA4YITij7Xe7dI1Lt1pe2AohJZVadhL/zf/i8/xN8a2IMbUm8fx6lp
YQvAhK7+lwSLVgTRgtevE17jgqUs0uYby/h0lD8daDotVtGlkCzywwWCuzQtfoaWMRkLWxQsYddS
NisTDlEHXAVrd5Dfcjwj+dm041WALuvmQjOVI8kNmm1K/PQ7EXDgWxj5HAyf+frZmUc0PJgSRUrQ
ej7pyMzVerAac1mr+z58nITF47etU68N4XC3hHkR3uoISRwUznBrg6JNtpHI1u+2CC0YBPiNBxQB
cmHj0MdYzVOmNTPk8fY6YLR7tl+B6usGX/2KETu1yTX+k8OFYifaXiH2sPKX4g6VAZ/P/k/H/TkY
lAJlJnBdpw/UIvWtiiCV1tXydOfs+sDON26dvyG3qtdZp5NjRpnqfp6+Aw5xTyTNEb+4KZIyfWKB
u5YzSaH3EoPomBulECvQBJ8ltBwmSWi8/w0azjz37ELE9cpXe1LgujLnQMxxNPP5HlrhY0YZvKMt
+MbReJLeHOIt8vlqvR3zHLfXvEtN6y71p3I2i5syibXhUu1fMJXMm48WFvglexX/Y3caT3tbHW02
5/Xh1P9120zt1JqCnp1RVqU+DnpxsVPQdy11Jnh+y+0mgUzqoPsdlbb7FF6oU7mSoybobJOAP/XU
z81V+J5sE6TANRMBPXYXkrs6a3y3J7sEEZ8Qg+pc6JnsfTCqom0mc+UVewxHnXDtHOZGoAZpbvIK
Zv9c/kAykrrF53OVouqnoNiBHrcfYAdnuKX4YB+4ZW+KpGRab5UJZq5FXtI/z3IPt1ePW9meWr83
xmijWwroXATWW56hc5oC+xdrKhbd9kzxbECKGCzv3/7NNZE4u3LWuQflqMPZNZBIdob2BbXs2xF/
+U12xa1/WG12zaUB+JIh/gqghl/oxRDqvfJE4lt6fetIY5xFGo/wFI6ozblp3PcCn2JSIozXPBDe
hzeD2XrwF8fSHFt2TRzrxgFCc/f+AJAFVuopWw4ln9+sAV4BUM3BKP4mXUt8c/GhQ1Pbs/qzXMXv
g/FpIpX699LpoFms216L8wmZMCwLjDXsqT9LHAt7Fr+XR8Xl8nIWd5IW+e8Y7+oGDD8VhPGzyebI
9UuJSF2vc944iIy3M3TvYr27K+bvggWqES3/A5kYVKBuNvuIWapwIpq+hyAv1qJAZo8mGMdeSttC
0M7yNLCkHz2y3AXhlHDcqZZ8MDmnP1zGgBc6MZ306J5sNPEW/RY0ZyNwsnvbqMuXf0BXDaXMqxgV
pUuroZHi1l2fE63Ibf/G8lfa5U6mpidA8XhymGKpYetLQvjisWl4msgzEnbYcoDe2mjX/3SDjyns
mFF3s0M8FJ3DusJFBwiadp/duPb41JcP8k5cVSzs098l9j00bYs1eRVgCCHVTGYFYvKrPAbFEJGF
T6khXl1XOfZs+z5j7E+L1nN75YUNmYoXzgTFMuysYASlWUM1O9CGkcbbSEhGugQ3U0jw7e5KBGtF
G1UcH/lgYZBBTqxFkhhcgxpgS/Amlpf4dTPoMuBJALVQHwW8elurwQ/r8R+/gHQnqcw1uiFuU9eN
tNHNf6gRlerQ5pOgXyr0ZIexV/Tm6zlEpNueFIlCO4TyUn2Dr+Bsf/fLWzPT9xaseCPPiahIU6UC
n/PskmIOu1NwHWBZElCe1YuXI6v5WRuD2M1pSbeZu7KyCfze9iD8CWvRZagll6H4ZYYJ36v/t8Sc
7H8WoXQ70M7L7xv/DzFp4iHAFXjGQhd4bIqpcl+cCCTMKPWbH430tJ8atjqP3vwPtgvkv+SeMhrS
5SObyHM5iqi8v8hLloV97x6u9ZpqiJScVe22p9jaiT7fX4rsnZR8AwU1BxInWOjBic8P0DMK2/P8
GSEkOziVoWH9FLdO8FAHE4czNhErEiOz6fmzhPUTxz0wAzRmN13eNrxJzJxhcMapQg8rj2gltr1E
U8Gi1iUSXFPEoWrgB3CUkAcyg4rxwF9xLXV4Rzl5AZnINwXtze53DjnRkXEukEijowsiYZYtazYj
HtZpL72F75jpwPY/E3bq0RYTBoNtCqSAFdft2w82yL+AhKTqL86rSGdQLscTpfOX4FRZiVB3VZ4l
dhJYsm5hykkH+K5CSTjSwe/jJ6cJe0ldxf6IPp5cfdxOoaTzbJlVPn6Hal5/UNGXTsny0GecZ0Vg
9FnbS7GEAM6jlkDYLZ3nsekzhOHnDr3Na2WlWGMKQzDFbrlN2d9S76ubCGaHy0lrj0fnkKjaZWPv
nx7sC96xo8PevPc1knleXU+eY9/KAwpIZpFnDSE/9ZWQQJ5pf+xfu8hhY4wSkcod3D3qmPmCBLNA
OSVWPEJlR59/F8FMSPf14EA8wG7qqQvS9grKUD7LcFZKAKmqe4bZHt9WlfD/WJl35xsu1+BiAIb7
/ateInNb9UPYLt9MxOyLSOvtYL7Of9xzKqVgHbDcm5OeFzrgwfldIFf7h7b91xDvrLWOsZWHwGjX
RF8D1fE13+mcJEQBwqKzQoxhl5IPLafPRzZ8khCWTE/CqWWWUK7x50Cez5YNGegm2Vsp15yci5Xj
P2WkwYwInOZjr0LTYTqorNu4RU+nQyIVHtsjv4IeatmWIo+ku/TBV5ixJnaySvL0WraJr43o0GU5
cFrUbAWInBistwZRRkvAlojaA1pqsI7VHtJgWrWicZIlLZTcryA4/fXxchXH0+EcbfOOXrESs0RL
d0M75Aw12QfYNRY67n3TKkJCEk8FttGsySU3UyTN+b+wKscrk7V1dn4NPyZeYkyfhYGyyj57Xaog
jQVIfk7mP7t1ScfAVn6RghHkbDUjQzRxHF109pSKe0H6zAESujKWuybBc2oaSWK97KLr4K0BJDYu
cc8A140UicrLoyNJEQiNGUHiom/jLl3XCy8J6MA6+QB19ZqFNrrJoY1xKVzOxs+qlIv7aVhWT/Bu
Vfef36YtYUFxGK3G1h5R1r44s8knnQr0n9iPPsRB5wrOiAaDoKFxN49C2LS+4IuX4Q4aBDK4XKzm
1psWnC/Lg9iOsK+Smtr4GnlArTIATWBGwGzxy2zFu7XJCsXHCGCgy+RF1dY4q2nI/aDIjmQhS1C5
z4XKPdNqjo0AKWHKlc7HiZf2O93RVrDbB6XKcsuTvTkqAz6hQmy81EPPLnD+v62jL0EH1gDmf17v
4ixAv5dRYxfeg/SISvqG+fjR42YsiK1UV8e1kj/ev9BLnKskWUdoRYs14X2FmGuQ/8k6BvRE57vn
/RGUdPrYDjv5v0lpRW62SpX0TYByGBQlVavaX1oQxVDWWWz2jNM+7z0t8d11ZZadk3gcUFctMAIh
xR5RHa+cG25ldEMr3dNKZgYmt/GlmZeOo2D7HDGOlljch3gDANl11MvxXFR6djFn9p1tEwMK8ct9
L3XkdIOnLjlpML7VNhaPbRemNUxcL30OdSQb9wwWnGAM8oIyJUnYZVmzkEaUfffWdoeFvCgcDYL3
ewJrCyG1BgYC6EE8R3KE0xo9/YAb/XwoUQWrJTpmKsbXPn0PEYLVMa/EfKAsvAfpphe/LUff0vpl
fe4znMxchFyUG+t4wCs6i/xJlmVNGd4xzrClxzruGUrIVENu96aFdU828eVLqKxk+6WN0+iCuOee
aJXrH6VVzCE6bcp/sB5F7E/gdFT7sKt2Q2ZC8mYoWLe/tW+X8Gsr2S1wI801kLcRG4yO19pFgPkR
v5YAcRUVrBeobHXb3NX/4uVOo2LAyaeqEQwh+/z2r+qA+Go6blJ+zl4RErXMY0L3AKBDSAhcqf2A
Lx+eK3zLdGf6LFWBBORrkVjhzUPd/u+3lagSirl1CKrsh/K2LeWeqBAUyKmxRUo9dAsSsmiL01dh
XPzkFqHx5+bh2LMpCvexuqMEbU4UQ/1LLqsfm6ACyJO4NlKUe0hhF5YST85SPDPfcSSg3TGH2Ey6
ZnlOE31IQvBNQKdD7dB4E4MYLMjLaICBpGpGOdTLy9Mk7sQ+zac0c6qfMcedqN7qegZOGqK/GzHc
0ei4AgkWxa0Q2QNPIeEEoBF3Vl/GxB1T4Ca5Cuz21m8L/fmas5ZdoZIBOhcjkJuXcRGvx4XOoYe0
qBPeO4gFw/T0u79qYR0aB2zwft57NRtBdyaoy+NMcloMRfDqtQoINtAS4FEliyj+9TC7ci+BvdRt
2jvDHwtG55Y/ENMVDyjmTX/hvY9EEUgCXx14S/2Xgegum7Y5ksIdEYshYUpmMagVHYV97HzPZBcc
fEUPrnEzHsjFjC+PQzpgrbaNdsYeszNsC//KtPyPqZdxtxjzoACOA21yhX528Ssa4dTst2sz+pV7
znwRiG4X+GGUuklNUqetMH33j9KWrHnJ85wQL9d7ZL7hHSZC4y2BS/Z0SYY5ZrfoUPyduzXyrzEU
4oMMG0FddgNMm9Wtuh9cfpGbX9gNSz6XSZJhpKqU76PssKb2hl1LiENTd9dY/pHhgyYo7fi4k7xB
JnrYeBxl2dRnQwNGlH8x51Cw6vb7R3Aqu8ZpEUKjE/hlJ3gJYXSaM4W2/3n6TcRKj+FWiTkYzWsW
kHdkJb8CX7mG/VZ59CLIX5AKcJ3P8Oma1Ix7+oqTukUaeuos0qayoNenKmcpABW2KkosOqVgiS0P
+4b/Ttz634yQhb+AQANVStCo5s7HneCRMyfcFgu2/F/h1KCo86PSANhLySvmye1kKmsbj1h/vhxy
F58noxDQRiAWa35/N1J7rJeTno+iYsAZ9/ZdqdETVSfrE+wvSwkiAHuFKekXo860+0m5rgiHvoAp
iApt1VSq/+pTErXKCohJuzvBrb6DZ4on/JHKFulckmjyBpq49SnE0Uyv8Hycg0FEvGBZ6dsh2V2I
n/oNo8UHz5R2S2GmO5N2rGNoVUp5hWftoh/3E3xU8zvgz169O9NEWCDzBSeIsq/nldsnOoLtRDKf
SgGL0mM6138rfo2FQ5ysTk0GTs25NRXExdQh9DLsNf2ft1z5kCQbWP+8A4fuqqDDiuhmn7oCIR5U
5uGpEHqIpIlHyg8BFJE5RpOQ8SQXxYxiC6fQcd8KXa1z4CAVG8M/Ocbdb8Lw2/kh0ksnupOOuglz
gSdbh1qR2xPE0iL8H+R1UQA9H0sho1sJKCHsVB4+BNoWDvZFWS/3M2+JJwB4UsA608MiZsLAMx2Q
JyBKEYd/WXFliL1ZG1K9e3AVAnbHIfh17A74AUqZJ9kfp3gFDwhjJN3Vvo+ztYGyZn9DX79UzBy7
EAmKoEXGNcWJua0ZaIHW4maOa55zGBV+aE+mK0VfgYGGGTDwirR7LrWSkuE3WoXM2vuAULh9yFMx
wQgwyp6dayBMWRtVDDQdRK7fer1cCkafevVOMeWC8mrEuVeX8SCDTgoDc8KQMBmKwhea51VxOyYQ
bHwPp+DEUoru0JHPwPvO+kHAinTaNgpJINk/Be7QRPg/P1wgQM5G1emHO692wHR0OcwxhYa+VvoQ
5g4unx8xQMjJog3mCYwJbsUkcT28etQm5ozQiaFj0325aPsFNlkd4jZ7M8vJvOUXbEqIKtjbuCrJ
QnPFxDD8vu5j7nhwywa/4yXR6vijZLRQD/N8jrZ/F1ELf9X4ciT6ZanJH+ZbiLy9ctUqFMmpnQE0
Tsv4BxDJxYoIzQayZ3WjM9VcM2drkDvqz6u9jxgKyKRmtiI5aer8IZCt/vjsbbQWskEAPYDhv0SY
TjvpYZvc2Inl20bcVGBYkMoFgiOdgNwxCPkec8OifT9jthFSMp9D/zPV5ycRZyBiTt9BI5y7PsvK
YIYkTORdTiR30oVQtNeBczAgRQFKkxP4tdhO74E64bQ4nL0JeNYZ7eqvfa1aasfsU7u+AKnSPAR+
4RoTyCwuITRZPHiDKgJh+1IdGpj0nz7RtG9tynPokC0wz2H00EcMG8KRL2CS9qXWT2V1nnmYeNgB
1HOycY1388u4h7BgpQzm4BuFl+48WTNWg7lrZuMDbBKavr35weUBnaAa1oilCzhAgwR7T+LFaDC/
ED3rfxMnf6/b+6uusA064TePwBZ3pf5IoseYkLHyDobZtFjHk/teWc8pXAitmKket/BquwjJItTq
vlHTZQJPjm94252LhF+DWCc1QTCMalKPGROMvLqILMsz1+vo+nNfzI2GsLhA2moJQUGVTIfUwatx
BChitCjDF0NGuMcW+szi2pzSE8R+iwTBvh+LsVTa06BpKMgWvgLZd2oHJPUuyL0/QUxkp2dYPLl1
pKMMbGsvwYxLiJZHUG0sL5bHM+ijk0xjE7gjsJFDjtJcvrCFlZEQhCaoF7QH7OqSi4PRUpvr2Mtb
zZaMK7AGyGOp7Q5dsNmsm5lrCx/Hs952z7HSAI+KQcIdS6/H8zlke8i+R8b/qzf7vCSuj2AFEXna
LZVIraV9/Hcxb5Db4m+AQKgclyHAw3f7KZWZbxxJFgvkKp8nu7MDBGp3yxzLXZYHwlLbRi2+y9hS
rP2f3vTw3bq2oy2ulmzQnT+TDl0WqpxK7SeJSEMjipSl6LzS5PXeFMWBF3gwLOCd+bC4r7UXsy9U
IaBNrknDorM33KY60inzZy5EGVIt87ajRkYb9z21YoOm1hcqySvmRHSuLDVsKJrc+HJq1NsMZRwF
JV3zT1mHgO0HE+MGjHwF9lgGwoCle6kXVMZZM3OntjsHC1HBwIekXX2X4cZzhMk3q2eJcKeRK/DZ
h2/pOC1HQk9LiR4etZLXlShkV0XxW5LQtPjMNuzQWWq2jGgXtyqTqLXQAeczEH49Su5DdviZTOGt
o9C4F7w/QcexINHfYT7/htkyUM8NeVeqFjivQFvpMHutxxqURdc9FZ5qdQeBSddTxKjiOEScquwJ
8V6peUvNQHrwjhJbuOly231+IdpP0nIp4pwQ766ZyOyhdydDQDfpHZLBiarBN90JM35/61IF+1fZ
9tC7mO+80xPr7eA0R9LRhPGR059xBkd4aywn06rlbtumgX2gV+OCOyIC/CA8c+7fTaLF8S0+G9dj
ChjXPRvF9URIPJM6gOdJLTp+NDLUgya0FnjqUelBooo70YmzLe9WasQrz2o9zacw8q+JMlLynL9U
0Lvlvff0j6oFlIvb4lmZv9v6Ji/wliWoIGXhNssPxFrxgdkeyBzKv+rPcPNafwINFV7a5jpmtI6R
wFfZic5ar+zzaWfll29syV88ym+kYN4TR3/L3ihYUVZQQhZ5XCpfrrjjcsCIi5izauHbmWkuaAV2
TdNHgzq4KkpH3Q5NBvObWa172IFoLBdZ6Rr1qFo/n8FGhMhS0yPuXklovk67nT6H+sux0bUp1NpI
UCDpK65wcgixJHAN8qBk32u+RedMcjWW5mLc91/sKMhM/Vibu+Y8Ip+BRavExYOZpJUtFAa0HrAO
5HthoPCVaVOFpOX8VsSKyBOkiB66wCtul0cNr07ae5Dla460LmsE6Cb363h8U4KDn9bjFYzoeh2a
jF2YD+mjJ/OT1/vx8LZrGQMzuX43f+MvRZkDaJX8v/opBYcUT38q9J8lpbpnHVBdmt3W6+HTW57T
52NIEdyKldYf8tbBbmFJQvO+1XzD/zor33RYFK8y85hmsPGgx11bvKCnLcWxxO70ZEUUVGUtOO6x
WW1RnIAKUN7iqhYnjlHYqXo/z8HX7ehXehj7SEDt9Sxjs+omB9te/GKOA0nBTbJaMlR45a+Pi3BE
zCnK9Rh1h+UPWafkOIKkeaN6k3HeBtamhTjFDIemmj86cwyPUSnm+vLDqkhEv//MTjPPc5KPyg/U
B2WyZbtCc/KcB2UcfwEL6JOvucF7HSyS/JV5ZGfc3bHEqoiHNSwx7kP8cZK3pDyNMRun39cCvA0e
6MYkaSK9VMJ8NzxvoeY+HT5iK9BehGGrY8+zDKmykYAT0TSkyGN4TBwLJz3FBtmZKIVJMvhlhGF8
JYKlVPZrL9jVSaCSN1NEsobKuncMZl1DYKngbDgR2VIljiA/4+Ncgd/Wh+22MsG345h1Jt51vYR7
ILLmjPiqzTqZPhh+SHg62o+BKJKnhKQCJtOtSKJnC0eEM8ncGUXmE2YeEjIt/vWYbE5bwfYWZ24q
xfo8aYGxYHuglsC9McLYF+i+92ZpRkPHXx77ycf2ZqdJoqRpsmEKA/7Q/EcDUOuVcIQXkn6MxHEz
GQDI2/YiSI5JpsfufAWPljN/9i1YX0srcXM6GsRXghaGst2RTI7pZEv7AOa5Afjd120sD+Ex6iCY
c728CR1iX/I/S+P9VxEtXlGhRoYS9da3QKO13dOQhkitcT5IhFko4DDJQ/gnI08PR8BC6FEhbBNz
0XQ0bSdoPvW+yfZ7wIIUiYGbz1OVrqyJ615xoredsC5js1ir3+MaL2GXsvllybTpFBsGJ9PFSnrf
lk1F4UMKq9YHqlWCiRgwh4tk0Q1ZZD15ktBrOn4XWMr2OoOs0L2DkRygz2tPjxdV7NbJryCnXY0E
Sr9ATJpvgngprpWQhmY2vSFe1xK/I6W3TyBLndg+23J/OUiDnrD1ApoYWtxpuWGCwRz+IVjn0/np
LX1ydjKSeJc0W0MtG+c5HeveOzMAetkTKnpsm1shqHkWTAKeyAhGMM8jdsCOzX/d45k8zaJMDjbn
cDPMSgWSJ5DveWMEA5FgVsxdZXeSGPJa0tnolvVhlGrsRQ+G2UaVlOD5SYPIk6+LMcsMflHmTe5K
Wxt3FcdJYc03z300BeiMYrvQo8GggzUwK82HoBALjbZrFf3pR40fOUgjbvTHZ45DHPLWUJVZfN8t
RIWuPVs72ASKmG0muCy1xAbupNB0YtjyRSH1LVAleJ1JLIF9zFQKwLf0ZpG+eB31WzaR5JRD8nBI
wFJo2Yj/qNfMCV5KayLz8i0DZfJynhLb5s9p0Go8xD9Dt1WzcuXpyVLD8Qj/DJssIETgJcs9w2+8
aCSU09eeWeIH6IjGrTgi1vZPhMuhLwAsETQ3gqNM751AwHc/WASmUtFa1tQ1jJWX19USkvLRPx1T
WR12rwhUYdGhcU55Iav9+W+GM/IFgbOs/SACM6pLjQA6oXc0legXSR9m7+G5cWqaejd8zPoX5Zwy
x3v9eI6FzyVBmP3qmpG4BjnQTzr0w4dJlaZnU6idwGcpNgj0J+v7KJiqT4mBILGSqbfKfyFIU9z+
DdvIh+j9h9sTszWhcb+6085LZIbw15KA4KEXpD9h3Bl+31OiLU9y46p4cn2xE3CoqX+eB0uuLIE1
RT0WAhRph4wGOoMkiYFWtftD1TU9Tc+UXk9dkHawT1ABVF32r4kHcCnns7DNbgb5KA1N9ZMZnZ03
WBc+CFXCaapLUF1WcM5jEgSVwqY+p1yr5DKsLGQtmbq6E7mhI8Q1CB8G1Tvp3q7zi3jKEoqBhS4z
goqiQ5VOvJjGNfq6/TkhEZugDU4a7eM2F5Yd84K4wyIVXp0/2sJhkPjNCtuDr7d2/Ta/zZuuWP2s
3e5g5zM7JSFLynfb1azaPL5pmuWvcwLcrprnREjCt5WZtEGCiFE2hJdNibhq50Izzt54oJIwcAQK
/PtxZ3wv7jzV5KtfwhD2tqD/Jvujw/nougGr/SIvEnGCGSKAwubxy28QyzLjFTN+7iigzCTofOch
+A0iMzp64V+gUMvZI1MpPjlOnS+w0GSITixoCH9hCknSTcDAmKZv4uJXbt8LyGmnO25D8JP4CAKd
NMw/g7/MWkqklPn9e/Id+D710o/SuO2qFNteqD1Q5i5gJMUmUc4xqa91NZWjd5+a+pM0+wZglbLq
DSa6IImIWB1oq4M5Zyl00s5dcHdmMXkVebfaXsZUAAfQ8nDJOHsLQwGiV7i4O2ZfkNZSieXlcINb
ukOjod+ObNecezduD2eXNzLg5JrvDkG1BYdN78qUF3XJAzrYC0NROVON8xOjG0xrhhyCADv0p+Vj
73payOMTbOabAmn9OTf0KpgkpDoBO7EFnZuHS9uEFEzS2gM6pYrkvNlKCNRLrB7U9Xzi3we/3IVq
njze2GcQaan5O1/iN0hMrfCMl92diwHIUWvXMUHFVV1HzjuvTEsWs767B+ksubJx9/qnHysSzjX8
HYEtCdIoOvc2Wul0zba/5dM2vVCXPRxwQNYngI6R4+qLuqxtinjIIUAhqUdP36oTUlXwEWYAkrHy
K5wXpJwAzbe8ko0TFhs5x273l4s4TwQbW9nG7Ch+W4JYcxU5itU12nnCep88rprTdpwDUB0pCo/w
HqogoVETWJilEEf/T8Gw29PboCIFFTIYttdxvQbbl21+CYK6mbmrWWEj2DDXd/2zVIPs76vs3pm3
NWYFHTbopg79rAag1Kky+TPXzPP1Oi1cDj5CNWjWg9I77pPiJ/cVHPEaFxSG+sz84u8mMEtvdBk/
BEFOLAwMYKUmXZqmh3f05DcDuWwqx7FVFpBmy2m8A1eHR3a4LMKzim9CxHyTJUHC2OZOMttbjInv
oywMJjZMcTo+P47JCI8r5R4FJJ/669+bWLLeF1A0XyX29eH35Bfktst+xKMhL8jmKiyo3hVBo5zo
vt1inmHMPvncuWs9qVM52hOEaLJA+Vk3oAA0B1KNJjtY2d+syjesywDqFGbf3T4tRDFoCTmTF9Cy
DkzNJfeshMAjk8SGFfA2G0gxr/q8jf8ZYv4tDgqU6fW2hYr6NZJ0xrCSZr0TNsmwcE1GbXdWR/l/
fFbXH9cBEAevzKo0RfPuMGmD+QTOs5UB86gfsq9JprU2tVv5HAYwA8a6WkdZMvofvjFUnpwnTvC/
fXA6QjF/JcYCB7piLAS7SQYsAKR7uHVccYNiT/cEJXaZTAgR1CVf/7FCRo4BrcQRxQ6rIsumFhwk
NyPRqNvixlLHWXelgKykp1jiLSRyJqNPvqU+PajXnL0xZ+LVNzC/vQ9N2WV9iqZgW97Le+y1jkN9
YGUw9ctQL8OiEc2huywn5l//fvE2oP2CNhl6ZewNLz88xRifUPU54PYUTa+YLfdwSJKXcrv9KnSC
VdkkhMLyA7lFLPF8LvpAOUDwVQrpN0lmOl+4v2e8cS/sBrI3mxF1oknCFEDTd5B5/LtsQNNdznpJ
7laald0v9kfuVZnw8v8z5CEM6UTnFvSP8ZU+wab6S6HppmCkgaGVDiwoNryZEKPOcUXM1oYmDzRE
cq3QtpEzgKH0zAOXu2XUxCzbiLLio8e1ME4Fjti7IPOuln3w+ozi5yaKO1E2erE8hMsdtYQ7Q+S1
B61Gm07jTPO7GxlYnejdUaXbMnvvme6OsmjG35DaA9JkwxaCecaXZjl9ade6S/nhodoOVkh4ITxF
vJDL36f458Wj4AJVRsABznddQtfHY8uNPlsL9NidjAkbWSR6Me6FCi0Aed0c/JAHmaB+PHqWKnSW
jguj0wArPHrabKaMsi1Sy9vHV5wCRLIM6g1G6RzyxvAt3pvS+B5IGIEW7w1ms6z3g3p90ToygBWb
XfRx7rfelA5hfvqKkYg6ySgMCwaDGbxECA6VuBprzSU9D/zg3ATifnHJ0INgl6SjGZ2nNdbkjtd1
ngfE+XZAKZvI2LADhRokTwy9CprSC1W7f2fRhZ7V7Gqyoi3kMsSVG04xk5HXUDTJz8F1sSIemRxv
yzyYMPb1/2rZrYUyqet1T8fcqn94szpEowTWF1RZ6nUoIaL3g+gj394z593Pkt1lkPvf4UVvDSe2
NRomoDBcFlPetChvTjUpwTOeSA6UVtlzSRwPSxMMEd2lnX3SH0R1Gx3EYhL36TYzFNFy3GfMBqD5
4UjsFNiWQEGJgX863CnaALA9wn9gw1DskF2yTFqucftdQ7p2C5zh3Dg+LUVdHNqtZDbE6t5Ac+pu
GVhk8+wsIEelbyoRHsN12rndpQNYsl45JKukI3DZntfBLNPaBuwckWLFzuuL60KSgAujjchZPeh/
metJb6tiTHVfgBAgfRJ/vJsvQo0o2uzBxnsk5N42HXDRq/AaRz1d+Z1wZ4RvBKNC5tdNTgVkL/Ac
1S8pyDHRYtcF2h5FcVnJct0vtaZ06Us3WxSizu3AJuVOQOIXjcShaqkGqin8XrstSM5tNvhVQ+sx
QJYCm2QkZnbtf8MJEytq3WcI8uPAgZYZ+emWl2drebS4MUGTh8EXvCM9BaBMuJ9nLhtye+PM2TeM
3xM8iGaDnPYeOtrhlNof1h1CIuf0dCUbW8IHloTe0ctjBNf3nIv3rTKG2KFHMqEFBIIwZ03n2jky
Uk0yf+hZmZz+GjcoiQOeMSD/7W1BebhuWgnXt33EzQhNgQ8xBTxkBZbuMdquZpoNHFZu+e9l/90y
+ZSdHx/zT497nBJ6Tr9INdc55NOE45lom9MMF/6LmMDQNvVhS8UQYAdcvKn8gTd8d5XGbJhEIGMn
5RgqvApMCzNIlxG+q4RbK6qm8Vt7NY7ZuHQKjYVM2GjCwjlL6+SZCA9Jj/dg5qT4/XPjqiKxhEDy
Qvcf6W/4aX5oGO6yxLzBW60J/UILlqjTMYVSQ6CsPHEBcXiEnxGVKBmL7ywxJUphSDOtGEEhRfvq
Wk0d+eh/MkrWoDgBfM5fn0ZXz2RuFboHeIlNfd4zvu5Ugm46Lvf6g/iV6e4+UDzFK6vID+/WMdkc
WSwaZbXfDBo5vTdFuBTwSnCLw/sqOy5MchB8xHeXM8rKnE9tRhbYKeOdsbfV8tpZXnV8XTv2mJzK
MLL+lkek2zLX64Wij6y+LodX93KH1fFca+fQ5rZ6EvFYNbaHGqtIdyiszrqTpBGIckqA3EJK8pVN
waUkEbafx69bnE1LzkzdJd0dyES+JyIP+4fbI88avc+EEMo6dY+syhsC2BRnoE4F38nQeDdFZD5n
G7KNhl+xEvZeeXjFsBAzM/g+GJVvjR+aEptccwsd3qka5/zUvfgsyuiq0K6RnUe18Q9ADMUQkw50
6G7xnZDF7llPr2PsZxAnXFgz7EHzcBeglTOMZtGjhygixsSVp5kW7+vXFbRKDawn/MTo6D9UVtDr
5g/RPj/vvpz7RApSd5nVFqBRdCfpmfPhN2c5WbQAHIKuNr82b1ttbIwXtoI679Qe4PJY3WhE7ywn
c2gNwnBEpv3O1JhRNPbB62Yj0zosFbV/rsllTOsHxkA0GqJFroa+CVUIsM06Mi+eYzFfBiIEUtMz
igi4kIlCOlW89txqhXqevpZi48nHjCBmPddxxJoTMv2jdasB8eqV2mFwJf45XjFw2aNcMW+L9BKL
HQYGcoeV8Qf33xaoYWE1iEHOCDEJzfRn6PN3zL15cXQ5zfDboye1A5fbNOHM+K3EsjhxGrujBv5n
sdSZQ1uKmMZ4VsNInexKV54sN0aKyz97ByjVQ9Tufbck2fhLZZZJTaDds3f2PVGpMYXt3fdaddyy
Iq7hBgsBmw00klEB9vVXiiFuOfTqhlAn2aPLySHtLluGDu6ACver4eCHdgnj+BuZTW/ZD8o3OhOd
uxXUloq1pFj16bQGDYMYrqGYWpgYX2XuZmENamu1qcRMyD1N8UNJR+bkDhlvHmz2LKI9nuM3DGG6
WjXHS8frH/3bt8E3u7YmW/UcpN5A9UIStw1pyLxzOXzphrdpeXBK3DzeEfiHeR8TVVeKI/eypOw9
V3O4PJtdxwIb0oGtBF8px4cjbUkGA1WBGW6skeA5BgV88kg8uVSqz1wzaYDcu4UpFHa4h6T7jrvY
7X74lObomsrbC32e1hb/vU18e+mjmqkfw+oyy8akOYaJyEaDXlj1E3B3MzNR13KdZb4sfBXGYsd6
/T7nXU2NVtW2Z8D0QOme1RomMl7T05FDT5IoL8QxaG4Pr+0LTahDQSDct5w8ZGID51GfXraLX0HP
+oZXYUHEqNo+T5n/xX4qkiR9yM4x2+fH6GaUhjdEFNdsJENmLzlx3Q2gKGh8UTO1dJCcKhHa3eUX
+0V2NInL2zT70yD9UHP06JPHqfhV9ja6wqADRpj9xZuZQ+R0qagQMAMnfb2N7Zpob+hmLl+O+4kj
PkqcRJEyAPv5186efMDwPjmHaIAtwR0ZhSspcbGCoo5802TermuSwNxS9PDmcHAXncQd8+n4zXmy
tv8yMtDwcgz1JP+V7mLsqhCK/8vw7N+LB90qV1NYILLCThIs2OYOC0GuH2cjquOj26h2XIiy0ifp
SZ7iL5exKMSHsG2WYIL37X0YH1pnwMMCWP9TLTDFnLm9wr6Esvn6ehe36aNJ6ciDFUln/bjwtXzP
g4m9nlqHmeiNFOCchd6RR24G+ZPVi9vcdHRzPW9aLuM5/l1QHhExRSveNdclDyxBaRvs3FZreVoi
BZca8iZfPUR+Oz/Vpdk8M+QFiu/R30R30+N8u0oVN5yZgP4DH4et0JIjwJfRPwubrErvLT7ekumb
Pe2Y0ZgNRa15lpLOILndpkFCcUIjuqd8he/EJ6AJL6XUz+a/cAD/F+mrS0TViB0hUI2PheX14YC+
UhUr/xmFf7v4hK2TbsWp3WsjKVBODJ49sEsoSD3jNTPdJnpVas5zvJAUxbdjCEOlUz7rejaH6Wey
0+YtAi0nULAFWYNJPOuNNO9KNYTx8+iMQmQQxyEBE3zw8LEfZYyZuqfinlIu2WKuaEuGTIEhKOZu
2y1R3BlOmF4pFB0t7BjGd+3uRub7+DGwaIGYNWHBoIfI38LXn2mLQ13CVkWII6bnHMSC/4tOi2ju
akN8EDICmMgr5Ph6sqJE6DEPcvbBNLNtnzL1kbnJV9rQCCzx7RL8Xr8Ta0/wLS5oa7gcIAIMrqsU
q9l4ApRUvLy7s3MGy3NOrvt0up0D7MhvBhpRKp/HQ/zSGyGIaTij/Owr7aiffE0Ygel+YquWXbzA
1tKxzW0dweKz4aCy67ECje2GPKJ/Y9LviiClO3GHCTuTHq5wTwd3/dpgVsY1Pyz2m/UXbDQ07iR+
aI+H+YMX1bxC9oljfkc8iORAMGjS0M8TA5Sjvakg5+HYPOeCifRSxu7BCn2uKrpWXRg+zX835gwJ
J5jUKz0x6PcJg5Nj7uPcFzPUD/Wk4IP5YcGhvKaI7Wa8GnjGLb3KRaO66XRG5MOKwRmY8s7uagK/
JNnS8C5iWMUHEsROzZwbJE709qy+IqQp566cDKYzAiSMCcYRk5NuqOTRuFEU+HgNtx8fhrYhe/NZ
EQWUBGTBhajlNU9qhJT5jQKLtYlIxTtUWDMWAO6GMvn8U2XjndKFR+zrtpW8+1fJsgtkjuiQRyp1
F9jKUE6OLg2XT730VoLrdEGrxH1TqWXN//8EFP57eKVdwmFcka0Ptb9DcQzxtZVbCWBpj0vRJO9a
ydR+BY1KuTfJyt3IkEV6LOBX9QH6xpkDWRhLWf3syrfsdZmEU8jvYaiFbzgOiFSvYUog/m9c2XD/
YXbhu8jZiE/T+6eoYZFarM7dqt+LpstvZlC4oyN9srOzhL+P0UcO629mTwB8nkCg3q93cCzIl3vT
qmPXCMFG9SssgpfUm0ygvy78vOTveqnP0fUNeHaFGXjuLAVeOUs5iVo0jvyPwuI9nVbCma8JiJhT
FUw6bICMxNOvOEk2fdYmxzGcPaCzVoqMYH43BAHHfiabiO6cxeCdni9yVetg4MEKSHN9eeNTI0tR
4Z4bhUeHrh+Ni886sIM9lvUi82c+S+r18qUSSbZ7VW6nNNb0XRQM5W0cidtAr01Fd3lS9/yNPuQ1
6FJPaRGkSyTxirbSxi8E5GP8AbtST7S0+Epa7BYMVHyCapNMHC09eDpy/uNCiFWaazaHJ1zywpx3
sbeWdA+yenBpAyWnJPKDnOGQykFbaWbxQyxeNspmoRoCMOEZ8ZOMghoo/UWx3L/4oHce65pTw1GO
jV0d/vss+UpEkhKZBT/ATlOOUzfbnv/iok+LHda6ZDhIckUmqBUHi7QF9zusmchZzuGp4KS/8kMw
ieY77bLCykdYCz9qss1k4dxCC8Sem0ihVlkAtWomO+GrFRQrg4pSC75BkIvX0uA6KZOVRhb8/bgQ
GRWzM+R2NMAaF8TBn45Mvn+C35TA6ctIL59Yo3VV5xjvFDWpCpuMo4boTkSCcYt8klVOF8jBEIZr
3mY9O1Bq8u6vauZkUxjmHy36hl8zlcqYxgKeEPqoFZryMURf5TlXYqXBqo/MvQ6ftZK1ydmvDhLA
nCTWUoz05stC5fnO+v8RunX0h3wS7OlU7o3jX1VaK//mhPyHROdeQ4oIgRH8aTWnypGo75Jeqhtr
EIwouEkIZEWzueHMBoCjs2Cim29xFsOxPVVrTtUo4Q15JdxBhWI8wX5nClSQO3t2fckfR9MCWTLA
hXqBR2zNrnlOgnaJADRwMLz9raHGEBlEaDUn+AaPMM2B/8G1jRPrHV+0ctcEYlWit0cPr6VKUxCF
0d8XSRoayEVHhbrzz6e620vlrhakqf37nS0yX0Jfl2t6SPaGdV7HzIhfQ4g+1OHZNAHNpqRzsGZr
UvrgkQM1c0ACKaC/dDyAQ7IhDERAZ1dIgorgR+IogFvxiBCB2KTBauBY9F7lGTsJqAZ+uE/1lLEC
vqS80FYjOMpNL3Na1oQDLm2XeiyEvybtEChrYWnp19goVrdOsbXy6aIbzAym76P09s/1E/CN/5WG
HTkOFgw+1fFgl4VPsgqBQ+lokECLl5YypcWdlnkTJioF+jLoa2Obt1l3idSPL39LYFAE0FX+pk6k
j5puC5S2wYTSjYOrXN+RV3U9MHHVFJnB0ZGYDYQ08NQQh8v4Ft0TAuKkCvgvXRUMUYAPq3BJ+4Q6
krGqMwSgMjcZX8PdE/WJ2FYPURGMuJudEe0ef0JfUY2XvbWtAFR0FnUs/t/tHVrds8ylL+OMfygG
Xx818AcCEgjIg/3irl5O5fTMLpJO+/fVqhBwWTu0EZ21QsJFbbKQTyCyCt3Qi2A666/01icshKo8
Kd3iYV9jXdCyAGbYT0umHqTJy4fYqF8bMrhymHCgz+sxpoVznqkOvtoZLJScYA3IiDpwRpXVxOPy
Yz1kPqx/hqrhGAu0o2IDjXB2CvdraR0l4GVpe018Lw5feFKVRwq1P7zQo+VdsoVamTdSEB4OGzMN
3JUTMuWGIm4mLSkcqmC8yBBFvtqpskvYkIvxLUh2mO7ijOknMdBl6OTLhuAyjozJg9oNVOUGHPuG
rA9B7lF7LkYIHeshl+S8GoekXJJT7FzD6L9Crq0Sk64PvX01vXnFBlPiwprqvxp1rREBBT5JWCgm
7RqenHrid89g/UIHmgUvpGsjiHsPpOPO+w3Y9Vy6IVw0oTMbvsH3eyFI14q6MAKtVLkkI1rL1tUU
iusOgcyvPC2nFAagzeOcayGWqcGIisJLUOZN4rFgoDz3HTMs6BP7IRZqxQYameHQqeZjhyxN9qgP
l7csdFS7W/Ts8+6708FCCeWqrzHZCOsyBmNg6LTibJg3iCNRkOdqyz1NF7WGcDTo9V5hGpdF5h1e
9B5p2kEkY1HjVPebtDYnUEuAYbqD7ndt+9AygbqTTUUfS/+okNR2u5EccSZJRBB/KYJ/EatKZZeC
VvxowSj1NKhlnl1dp4aynb+SakAtfNYyadNmyFrXikVau08Ik2S4uxdAlUwft9dacQm1xifsp4aX
DhxZutJ8g7YEj4LTFsYOcklP5AeZ5sea0Z3ZRXKR1zJAKQ5EYYFjdz6HiXC4r47QU0QWUKeorj1l
r47ojsGPdDJsJAYXQKyWmzA/aa5tYpfwQxIgiGW98Pf2HcxRVY8RnPRQnXkUcww0Z5QeF6O6Cjin
Nbwv8+RZiuLKQZgUSJpNwz13F3NpEjXnwufqQNu4Y5h4nwnL29GW1gRz07H5IctY56KcNhp0qbxi
BgYjmZ6bp+0yoc8gTwWgAdr2w3V4rBs/kihbBOISziuZ9sUBRiiTLcmRs+jqmE1PkIJWKdzTIJE9
FOSRbk+pcAX6ZfYTXdiFALTSx8Sl3IojBjNPA9vzetyxVy/tc1Mi5sPCu2OcnBpTrHCw8mihxYCD
s4ocD5zcVdRgx0N5BUb/dnYthd5ERVOoipnItufrGabfd0Tu9x87BbSuaqB74pOHwEMiP2Zps90y
9CSMA8MS6OVCD8DYr+2habxMgUzOX1NyrIfHytxvaqq6n20PEdCc95rRcQy3p+4wCkIxibweDeCG
vU09T+0HP5gmCmqpVaXKbCuzcEb2WFB8LaPKvNwzm9aCBGprEbtbYLgZG7ojzaX9xOfS95EU91BU
ouyogcmPRaI6x+EnZtCoO5uod42dsftidinxqPBRmwKtN6CH0UOnnJv03Z31QnBhG+c5S5VgZg6Y
T9WLeDJtRB15fqQbbjFkAjp+j2ZmnpkOv7vytFy1vo+V6JsFxJ0KtIV38Zwa3lBuOXXfBCy17qSW
lYBveyRXHvcP3SrirYt6l/+qr79nW8XuCS366BFaUG3nzvRyN0FuZeTEbzW5RAA4SjlVeLhHtW5h
o7ZDXc14SLA//qSLeVYJP8lzt9gJuWw4PhyOvO6tfJ2Ds3hRzToStKw+GoZ3jmJdAu6okynor6dy
822g1Oth/tTozlh95pD7XjNkWujVQ8NyVAI3s4A06TqG56vx08haR5xn9zw+69EZ19jJNsqKAg8R
bs/CJ3mvjorxhrIzRzp7uNBp9rLwkMYkfmsm523+EtzFqSdOr/0uC79RBLV8cBxAOHRrv00znVxD
IM/nKsMfmbpOMo0HO2CswwmOMxrXb8tI3NdoxXpmLey+MgHgDD01bQVgMupcnO0WGokr7lBW6RTn
f/ml1GNzYsRzcvcwHf2Nz9ZC9Mx4DeeBXr6z9UqvjcxNQoO49H19mwUgE8ikgFyWCjmHyvFnwQV4
++B7NnqCevS6DkJHZ1tOkkfFp0o6IoRIOCA794ysIKcqKUsKznoTpfkpUdCIufRfR5IHGLKi8pt7
FuFY4WhswrazMT9qXssZIE1l1OOfavRLvcxCG8bqOUoAUODMGpDRhxtv8bpmCJ08xrJQz1KukwOy
QeCvG33NmdLMw4M0W9Lldhh+4ek64CTAn+nFQ7E8cTxtVJhTiiwWwmhwkXm6uNrfnw0sX1OlLs04
rGUoOrC5VuL+yvVwu6saIgo4iPQ6PkBs5/Wbcv7jIJ7DfPG9VSikV2tAlTnpa2UTg2RHV5s0zKDe
8UVfLFgucnGE/jayxlNAqUfUgRdrXwbKeBbJS//x+pwXLEPVpc+JU9zTFcF39IrYKRJk2aNKZ6r0
ZPQWnQrWNx8DtRI3pYooGwo2mjoaAvSmqcZNnQWKqFqAkU0m6Yg3MRG3HMRiJ5PsJP7bre7BPXXN
u1hlv42et5MXHXtgLGhof2hTjd5X2tTiOWEEf3qXzdKQsvHEbcbfVr0gYvcfbXfu2Hf9ueKF+9Ea
jFCh8P0lB5FAgBu2OyiZ0kh0UJ7US1SO3mYkNOUjrQHyhw8PD4s3Z2eGRL7e56LbQvh5BhH5xOWx
LjPg+8JX9Z67unOCilLD9ZrfBLbFZ/gI/g8scQM8vAQyiBbPYdG8c+8QEu8m4l189JrPwM/qMobR
z2bLD7kmJuMVNyPEd0hu+eOzxQZqxNt+APJzZ652zhO9s4HDO8q2m2mORgjqhRIKwSKuFovDACJx
Ba50TO1QCAEFxKo+MPOKQl5F8rVQuJkD7gCBTYANO4IV0xK2khbo7Pc3v3aCbn6a5TewMpkyHy3e
oC5fimocL5IpR6Fiv1gvbe4Jl+/Fxtn1N7A3jklzMFzHgzA9SQrhwnSgVFlPCi4bqcH6J7qmPLMf
P7fIC7RpJI5ASYbLi0jztKlvNQnJGq8ywlwDO9VFBk2wFYeL2qdhtgJcW3sBMbuWWJZDBz+R7F7a
hnx74HdfVK+JC3q0d8cda640OBYJjMEhN1imDN+jdNp0zZiKd7F80lz3EbSMZvjZ+iQWqOUkKKCP
OGuHS4xF3+uJWPw/SCSn65PdW1yunJUVe7vQkHlQ2FG8vEdJ28XrweJ9+4JPCT2GWEMUo80RcVfP
aUuz+ErmwmgkHmd8mWAQ+cLaJY9xlyxV3m5Z/6SUs2nYqh50QkBcY4V5feLrbqbqBadpEFUHgTbp
z+/dN8ggZq1kWkAs4dxgN0aERHH5jb4aQJ1lSmipiYPWZhMgAd4mhpGEeAJovYY6YtezlntQT02Q
NnnWUkAUhgarRdvNXoarHW4w1cpM+1PaJ64XT/pjm1PnOcHZxf2wL/gjDCvXKxXPnteovAqyeclA
XfgbSN3UUcTppJLdmFjHKIK9GZDxr1KwmTzD7kHkR4Gaalp7WiVCzsjFDdLzeePBKvtdOiyphbe+
EnaoBtMz5eISQkMAeB8/mSFv3O8n1aOQfZc0QuEisQoeo4V1grQkeoEnK7FCbjlmfqySzjSjkvdy
9QNYFmVCAlVJQvijcFcjbGGrKlzRCfPcuEASkj9uo/xk9lVIO9sdeapkZFR9eH5hwMuuGdwIbS4B
FLJOxSR7ldx5eAa4y/63nXNcmlGUCFu2Q2ckKZGXPrLDhmqygne2ZvSGb8WJ1AZ6AHonIlXIpUjE
OX+IK7pp6IB1As6nx3cbRVvYfgi2Lw2OV4e0zvUvC9xGnF2SH208GvOp9ppzr3X4MZk6VGrJQNrJ
YpsD2dblrYWVKE0CmvpBbMJ/KrEYGlCS4hqJMISHkYtFdzdnhNt2n6xzmnWfm0EAYxVbQXVrTjOI
emEquOSZKH0uS4ituQYPKBHl3g6TslT5zhKU2QpKI718iwP0IS288qR34LNCnI3rVtHAuIJIZ6rK
wFvvpXZVwz9qjt1D3tZFCvJ1Gl/5Fshu9M5RAJZb49eCw7Lx0YhRQKdLGgHRkzvxtBObLwYZPNXj
dPtGzrViv9jlsYawu+JHdYyx1OLKhlriCkrYUUxL5fUgRMN1g+35WldvQXcz9XfeQx1Wn6UD0YsK
MoOe0Irsd4c7eZFxSIILn642mmW+rpHKPi0o2s2c8aiR3WxNAWSdFDGB7Gn/02K2384oAqkB/9lJ
zYmMremWH8nG5O6wWMBMzWj85h2Se4lfs119Ra2rgFTLULJtD+Bt20WY8lTWoOQiFLkCKatxuaHK
VGs2doDYFL6Y7V4IMg3rTbwR6B7EWMNdEHds7CeuyTfsmDFDmEyKXfdlNh90QaTAYD9iT0t4SfCW
2xebSHQbYCCqWtBS2zyEILBrcwvQT5MHZFc5E7TVEFURxZbOI+2cWXy6SezmuykxdAOp4a9N8AmM
BOt42ofU92t7sp0trUhlJ5H/K8RGpjv3nezXSnsg1OdTeZTCtQvmQcakvGL4ctgThIjqlFSyaTZd
LkkuY0NwpLbRaXJs+T4ZBgWJiuO0jzERK+zT1/2n9z0gK3G3bjoWY5Fo8XFr65Ytu4mKE9H7YOi2
HKmNvSdRGUySbh8AXUwTGrmy5iHGURiCBRZQfMQmYm5FOu0eX09vJcRYzRwysZTLNyKguEq4kLwD
dAa08WfO4lnaf0ixp0rluQzn9lKOjBz4ujGWBOXCr38H2aK4noSSu+FEtG5E7hGoc4JIOnan29RP
NCMs0OXDl1mJgBpPF9MwIgAxCB13MchZgB6Sr5K+GXq1TH9aAey1nW8HOMonWX2zKbnIrhwba8Nk
fc6KjZJrqG67VVMciXsovJdVQSwsihyCr8IbJZ2Z0izhslsAHB3z1Zxif/dOB2/gnYqZbH/vi2yS
FJdWTrh1VLqVYZORjBr8SchmYZEQG5SDKiiPqt7atlaOBGIHJi3oxTQeWB3mkU3qvRzJr8xVYzI7
5UZfHBg8NSGhorpZiyrtT1PGyswX5ZKkzDJFtdslYEZCdzcc3Yh6f2Nu3xDepjQnByt521u0LtII
4SQm7ZNjLAfDxiBNOqSF5JPvrZM9fSqv8BcjFzASk92wNK/3ATRfSU7HSncAnbhYWY4yRMttR0sx
9sRJXi1vdwJXIOSDy0C2nVJwLn7YWe9inGysd8Zt8D+4UX2RvYSDiz9PYIDFb4SZ7cDVWOWF4C/p
G16Vhwevjmm8GNTIxFfX4tvROrz9+3UZlkdxq6Cg2Wix6zfh90KL7gsHd39GGG2bbSDfViE7L5uC
VJwEwmvIoHRQGK0QWL5bKON6leGYHrv9gTes2+tE5F12WRucQyA1TnL+f8p+ZDlZvNS6x8ItHfzx
6lnQBKRLbXNeLf9FzCKM2TDQJ9ZouubpuL7ENnis2E5JN0UjYfFRe5hN6yTY4CHRUo6IbShJoY6m
i8e9DSS8ywn434c6Uv1cgS2jiM5+dgyMv1F9IZ0YV36mR4VsjwzbY2MvSRXruZHiBD9aE/wAblPw
KYENCC5ctOKyQVfN8XHJcLOOVQU5y4FHdUHl5gInTgIhqxlCM0G8XQ0c1yUaGug94CD3kljWA4lH
65FDhq/9nKjubIbXdZIXLbD7uWmKpgDB+XxzZSqbgIVu5SOgeekNBDvQRVNLi95+n5O14Sxot3QD
xV0yWem/TvXFDRcvUTcBKyBawCJy1ZjxqpZ/l8K1miQ4ZPMVWwR3pEqSC1el7CKsNIORgWCSPmby
jBYZJTk590pAYRNokmZcWv1q2+0IyZNdmnKW+AxbYAaaz7KTU549b75HILqnHCLmzYXfIarQXPUP
n0vjmUaU0aG3Zv7H8AUu4Jj5QWA2DTl9EVYNmfKzbicaVDKDHcK9Lk2ZLJNJO3N2GkXOdMnG6A6s
jcQULd5rnsiZdV64BJ5ilWShK7ggdLPRrvuQkibQyIzvGu4oMvw/w27L8Lgg8r8d+QmWrAFN1zzy
CQj74nZvR4zBuRWggW3mUFSU31Cqj47hl6yZPzYW3/du/YB7t54n9PrmtrzDLZbaHhyAZrPort87
cidaUCzjU/Cpj0gKvF9xecDM8eEyPlmWb3NOARlIJqGdMWAn8ef5yOkRxv8pqjank2za/3w8FUC9
h1rL6UjezN4M0irdOqrVq5JoFAz4bdlqgi7KlvmxdVNtj1AGW/86BWuAwwYMNd2bz0Fhxw2rg+Gk
jMAR5VQR5ufqThddvawFHq62JykPVnHTjsayuYP+W01zfW4nBy5ognEX8oJH0OYmw+DFAFTzQFy1
bZYOZqFZ2DL3HT5zSO76S7d6gvHfj8R7YaZ7zMuu1kkUH+Wp0mTkLn8hgm6qIZMGAKHr8FwH1YM1
3BNia7wqtt4BKl0CyX+WqtUydiAem3bCt5atBqrGKlySVVa1DdH8vajfjzPli1Co6h3fbt/Y4z+R
xruSFGg88ZROKQkG9cnKfxLMtU2TOScTm0kyDeeF1d5K/heZxbPjb4KUwuWlrQoSdTLvOCkN0Oeg
DnTiP20BgSFdCra6XqMEkJs2KC8PlJSgy9ZUgr/bJ4dTlpLEknHKcUWhpVaqbzAA457uFP82rm+H
zuBh463PLXcnGJyt6dbdMnvSCa9457Qcp5dhe3eais4iTDpaYD/htOrEN7M+4mSokJ9fQtGwmktx
AGVOWtvHlsCB96UyeaNSrKfIOtHj+IELoUgaGTsw30BewCruO7C1cfBrp3YvBEyRULa+d2x1Jkkr
G/DJEDxmBBjigNYsYEMtdpYuOrNLukE7rXRdmFV0qBwPIObeNwnvJAL5qVQIjR4TLSKiOlGt0bl3
meSrpSvvNTEi7JpPciEjv1xvzuHuhoDU/6XxxbxzTgaYQFClBsSjMBVUlh0m9cqoMPxdmXkXiUi7
cF36Wamq5k1tb5pAvw+QXvQLA6D56ffRAb5/uO38mu3O2Qb6un4d+0zC5d3//aV8sy5vA2ltQqGD
1WgCiYVWxVhL+qM3c21Ag+CkPn5nsV5RxLGpFGwuP27871wGX20kFtWmOjM/xfQSHz0Y6TBkwXW2
OileasmxqcLYhnDD1UF7ohsG2MQh/Ry+CNWSvVlBNSvx59+1oczIB50O951M11+7bYhy0FyJLHnw
H4QVkic5/niXjK9GOi1YaPCplKJn+SEvW6PquegGoNnE25bqQ/nk4MYgJwjvmzKeQnSyOtvgPRXL
VxzKjfAjl+LmavB/W528EEeM+mED0Rpz74aRdteUcevsLZ77j2x48pUMBAmFPryPN4h+qJQ0gRXK
0WDAHzoEcQGvzwa2lDIi+JcMkZQgcycI7ySNuwtmOeQT/HWLH549pZKz0LYjUQFFgm/ZWPCdgOis
wdy5f8hzCdgfarnPQI3HSgjMT950ybwmjx9bTPtSm5gNZfj+Nz6kjA5Y2TcVD1wKOxAtnBvWNzKS
3niQVdrW6+molTaz3Czdd9k+PtIH/M8wHTFNCY+/FFq9OGjSVLZ0Vz0ULg5fCZRMn2Eki1mCSXgl
cgCZKUgUvb0A3Y2QJ8FWNcW/6Ss7jadiu+zZy+nrWxkXwpQephzG+axQ2hRNA41SEhX9Hz49TxNr
A2ecOlgZqCMZLATMJe2UiO/FIjs+y44CAdPZk+mN2eh/60637dd7GsB+0n5IjiJd3e1xFZBAXzhP
QiDi5vIBdtj9EN5EiRb94imzZTMxhtSbJu7rClSlZssmNT71Ff3HqjRvimt+yr1TOQDZhZnHf7nK
+GII/zuQNxXvzbDRxg36bIlMgcxcNFQ9mOyXRn44ZUYpmBa1VOmdgxrTGsV8TCx0PYQCzjbPJwRT
FRb3c4v3xwWXv+G1EJuHdpAMAf6b/VWgZ35XKHIaB8ZfKq7lh4lpze1IJQs4NXanxua0YU+RQitt
PZ20igahmqUvNG+lrwsXUnSvcm95iywG4MfgbUMVwdzjbKJIPbVugeNW9Tz1PA5Ai/N77X3i1KkN
L+gKJBS6CSfCBVJblmXGTxBIf24E8EzcsBX9sFMM7lAx2lXjiKMVSdI+jKkN8vMhryvLpGHOdgTw
2kB47PoyKZ5WgHpYNzu03n5ddDj8tOBpwMVdKzDhGVzYr6xKb4FyeghSdoihdLBePLXQX8qETKyI
9fmg+nwXHrVzhnGTMZ0qYEgSZBLp5sLfkLtSoJDGUsZWH/I72/u8SRLXY5VMWHuwVOzsJN+Yvi/n
YYZs6iuELlWjs3Kc2sPaKnsv9ytXBp6/XX+LLZuGgqBGZedaLvhToYkPNeHrG8dYy0+KxO9a8QDV
bYpu6Och1UX+40mnMPAPA4x0fBOglYeThY9SgvamrTDPHOP8lYN6+Kv5D9+EkUTkbVv1MSumGLSp
JRqG71yXYzZ35DI9ocmVmKhcTeBxUNQmxQ9UNbUe4eB35JIusoRAu0Au0baD4y9UHOuW0mnkkbAJ
Whjll+nAi+WoKBzws1Gewp8urBNtoOr+I4SBtgEYOSjiGJVsuiTRNPlunhnh5JVipQwhHdYsTM9t
mnBLDT2ier+rpcM/8hqzZSf9VobuPa2+4jf1pS+sm1mDFVil1NnUq4nCTX0WLWoSZZT1qMrpy//X
lGBbzjSR+KyHLY9dYBBc8qpP/ggb9Ls40502OLNdtWfbdOQSb5g9RrbvF57VbhZzDo1m02iTjAgS
mtLDiD9vxTe5DKSXIqZPRdXeirBnvAw0TBa8tdZ4Gf6MTng5kmNsnKYQu7DJDG8KndPHgS7zTzhj
+8tOAoHf2tQxL1KjcFY1uieSEk7E3s3Qi+xfb/o3u9PxvxCqsBpEuQSFc3N+iElBqjLZNf5WgU8p
kyR4tYo/kVXxIsWfTdO+Te1GkJIJTwF4TVbJbzeCdE+USd6ifswboVkregyEbQZ9juZiaKW5oxeY
UwoCY+gDrHBWnu14MWE7i5X6k4t+7j+jRvrFz1kVShmCRG9OF29lCJuqYgln0yfVcSAi80MQjNTN
X7mXi1MB+jmTa0k4G6X0Yarq0+T9eHutn9lZJ0sSPEzCevIG56aD/KKQ7MFyYglTso9ncy8Vtvjq
XDUY165clBWbuT7z8DgKsIBj1w6eV8Fgp6Zjo5j14pLODEBcXXfYZSRaZJieCgvdGnR+vOETnP8r
nUEfcb5+p9eEBCLlFdX5g6SB2xG9xU80Aqt5sDi+P/WG0b8+9d0rDlW2sxcnbQF4Fx0gF1tYjZbE
ZGUlbScMw01FHfwW+GyC+k1Wqa+XYV6r+utv1/REJXfbP3uR0uIkIxwRaaAhl+pG2Rc5lw5U+kyA
MdbgpNsBGsuTINwezukPGH+VdgmTdDn63AAwgUVs3XEC0P03i7E1f7KStE9oZlRzRnphhCepUshk
wzuosts33GFscD5f/yWTM+0wvlyIcLkEXRPsOAVLDEy/J/8F7VfhGX6HtXpeYfc8i7sxznb7rOGu
Ir0JrldsatQ5Z76DPohQcSyvdExrWlOYY+l6+OXB63A50ca4UA1ZJSGe+9FQY2LEJqPP2b+e5giE
gj0gSrB+K+XodDFlr00iroIEc064spJshn5m3YbRwug57zTZb6LoAfoBgNi4k+9frCK0TY7P4sJP
eR1tbAHZ5CvA4aYKuXSoCg3Ff+6Px1S7i0VlGO44wXwUVpx5TRuJQPY28WLPHrwlgBApYL6PcjYK
EFmSQ6MMoxOHUr24JFTUctsy+LNtsOJSMa8zjznL6PyT1/U58vDWFysvX47+3IeYihvtEwnAO2o4
dW/cW9nOvDPLgzlDN3HNuFbcW2Nsx+GTc19CKjbs5HBgMxMhz/an6Fa/roqD4OzcQ4qmBAGVJEBP
mfUHA8dk3In8rcrP/ru/YcaV7BoIzk8Hids1RDJxRlQYSwiodrHM0hNZgji4UHQrqRzEw+jU217a
fsjdf/aoyDBzyt/ot/Baa+FNnV1mezVgac0NJoayyK1UgKW3ENxnYTDwlrtjAawTOGz1Rxf4xY47
cudsxk4FUH9vCf8uZo/QFKxyCV99oQcnJE0MK2UxnH6nC3WL4HdyXpm5e2+Sp9P4mBWpMfcSjMyf
JRpFm1HPWzxwcCxyKZISZ8shstQhO5fNIQDKAeiqA7n80RRkrvYSjVNq2EST7+IdImpFOWKWFSAY
eSw4Lw3lX7d1I1s0fCFwkJdsXL1Q9Am681AO58LV/BKBzm5yX3ql+11bZWBYv1ZJ+ewpgBLa/G+3
kMFXCta6sGfZG4TWZdU9DgJSmDNOqD79FBjnpoR5q8VCNM9T3dFyzqYo3u/Y46CQ1/EyLARLZaoh
UhJELA1mO9vANLbuc+iJApwN6NmkFG8IpcaLZLf0VzlblvI9e9WWN6kxntrRspKjv5RpC8rL7iCI
sRAfqIkvRLmIR9ffIskkO3OD5+AFjY7VkdX8ruF58QED29xnNF0pLlawOy8okByB39d9VdLGP8WM
kX9zsVUxZupKfhXfD+hfCbPeAU8tsBUGE9CThwkMFrhfMkZ3T6fIsgIocHLNaZiU3zwg0INiMj5T
sizArb5pNfKLxdfpI4rhgwP8FR6clKUeOqhuP1d5Bfm404lqtr8dnQKCJNOQ5JRqlKdiGGd2wlm6
Z0ULg87DMcyicBDV4NByecwykgAdeJbWdmLamEe0Y0JIA0k89uNT83c8jWAXs8R7zFc5KEEID1dG
VRdESZf1dOvmb7Fv+vL1dth5KsbE4y51or+X0Ma/umiZh6xtDQ8yp+97yEUae4nTCZZW4cFVTMa7
DxT10i66Na8Nvd2Vy+pR1RN4UvUCkuN6qFM4WWCfopWtrYIj8/WwJ4WM8OdMGf4VXkw1UdctlNw0
JQKCqxPFlRxJC4p5V+w8thtz+8VXkeAAjqmNZ7Jqbchd457Sc8ZR2m2CYrMRFVGLCqItIb3Q+tsp
22rA1a/GlNSBGjy5YiCpX7/gZaZAtVUEwHj7CleFJ8Mtb01MoGi9PID+E+2CcTdZHveIxuBVuuhJ
bU3eoABsAWT6wyyEaURStxwwE+GhATIi12HiYPStAiIaUOxK9wyzbNzzo+6fqkdRpxLZdDkPnkUz
nRKgWHZjGqW64Hs+MgPjD9wpizhHNNKkPYE961nWvm//xTnPe+eEqVhKwK8aFpng4rnDSmxpsCCl
AkE+SqH2uIZJjoDmksgYZBUsCI3lclesYpH2QKw7zKxaD9K18QOKf4bfkB23woRZo+92oyHUO1xg
ez9Oktkx0nEBcaT9G00JcfTArx5xJ6GhrLI73rT71PgocHYVteRj555h9WGG2oiuaN3SEMoZAi+s
4DqFomPyi5qCXMHdh0hofwdBKMl2gqV66She6jM93XOyWhae662cjr3dnAvNobZGmtHNznqQbRnw
at3SuRHjokvjhBbE/lAj4agwGGmfbx5q04eOt4bGu74WuDa1WWn06uentY/KVXeK3oJnlWFr1mbU
C5pf/mf/UNfXSCitdGvDHLVKK8hG+BgNPU1dZJhj4KWL5rVAaJ0XZ/JVE2ZBzC07I83vxAtrz0Y9
5mabHEQtAFE18BkGtTobbowd++pFPwcwTzo6CyMX1XVoY0irhRUEYmaelt3W83hlnX47u+d+al3o
ULPp6ZSrWDFtQUuarbkH+SWBiRr6kpZwat9zdUm9M6XI2qOUe1Y8WW6h2ygMGWJCPdaSEL+VBjwn
iZ19ipnAmUjYuQoz+wRplrsiXeSW/NU2pRWstzAWWS7/ZYxD3882FJv6x7wz/NCSkMyCPfRrpZjI
IDCUbkH9N/txLQdxOhYTUVOo0tmlyMdVwQG2hlGTJF1N+ySLw8eYfoYO69DDEAnEPw7TL9NmvUSB
ZUj+XX4Uj90+EKHx1lmQUhF1qzWBlyHkKuX7vTIHJvLuL8g62K2Gx/p6wwF2WIF7GLAR70FPMkFx
FLjPgatSUH/MSl3JhwxArCLUjN0s+wI1F91kiqwML4yOYZD7peB73e9omA7+1B/oyFEGT5Vbiuo1
nMjStyPWkmYiT0hpGiAMcCF9tg9Mhas53OHozs+pmyx9Pw5W9lFz6hNzjX2NiYPN/L4oKIrCmc4m
mhYt8yNhHgsKrX1easynO2bwCzgTddKXRYZmRdobmJPV9jX/f7bCxxqI/eG8xTopPp1ibsjlsCz8
iT19oI6r6rWzzb401B8hIMzyvqggJLPQvcBYIxPs01SFKKa6E1QRW9p/tkjZpdJXKG5pceiQJ8Tf
gtJr9rg9n/nnJMqyHs5A26XYJTqUj1mBwM/vqmmUXMtQhAhBLsXbJhwFg0V2g5J9zgYRdbTC7ESL
Ody+GpiIc0vwPbTjErPO+Tsajo2hEi8KWv0zDB1B3UgwWuCQom+o90SUVvlNWqA//KKT0eo+mjCN
8MqCL1RoyLj3BnWZP2H0BN0hC3DRxny9/IomRPUy5I3ywYh9b9YytYFuhZOSuRkp9YQnWo0bRv9l
GHkKZwHqA3kGOlZKRk5oR94PYKwZnriEscYXr7nOQNxne0x7U1v7FqXpFWTiRjjbowIPeOk96Zl9
/tOAVS7bjEmgI6e37IjZ0K9omct40wz3Oh4qWnkzdoz1H0vUCqBFpZ+NoSlC6AWph2FuJgXKiJpL
M9qQAKXoudVGpaEz37k+v9eJ4Xr3Xch+ioFtnigemaitWgBVcFC/32K6L2EGJUMWJkioqh7H3xLa
lnSxKYWCaaQ+VcfUbsnckunIJX78ZZIeCkzmgH+xKgAaPele0fkaH4n9BLGT3ttiU032Q0A0Is0m
gP+vcn1xcqAy8QAKjb1NmR19k70Tx5doF3bifYlKnG7YuLK6Ub161w4MJqGQ2Y7VxKAfzwLDLFuf
ybgN9Ta57pQRcK/V3JOpsRYdKnw85u8fuVKtRmD0II/kBckW16wnHMzrufWrcdSp6ftnzZJPhI95
LtWTAFHFemP9EMg4IGAx53d9hTZ/t9KMZhylZyYuQB1yD6ba523fEpnjcSNrpUUbp/n5/EW+m9b9
Ij90MdfdjHIchp21EqQBJh4ziiAwOM0lg/aNsMsLGwf0duK4k6GIH/AeZiaZCqTEcRGZyl1KALTo
oMvLkz6etb93PuWHB80YIuDoqrzMDOECFB/2sgkml3CgEu4feFu2/GgqR6ApBS5ZlzWXBcDVb6Yb
oAM/em8lYMuZc2bw2uj5jM2o3js32sZJxP2Dc3esByVRZfTUY8EnLco8n0biRJwV8rpIeSr+Gsqw
fnrugbdEgeLDrGM4XWsZpXe/JNwduy0tQCShmP2im5qWByMxXtKEMJ4IPMx1+yniq38S27gOW1ab
pY76vRvYet8Qtj4+xXOB+Qff8GncNo1l9yFu3MhMcxJSaNOpjHMoinHeg+LgG4fmhVHFfVCvhlvc
bZva0M4wPd+W3DoCQygFQakToustkvu9RJBzhVQj8a0kmN2FU+lCdYVgObsG/HNFmLBLtHTczhcQ
66fdDZZ2T0py981/reZg88M3rZd0ixxsiKyBd9eaTdGCH2X14oUWV+b6STeF1Y4ynxuF7aGCff7U
F4e3GS3LEH6B/qJTQPrWGco/M3mrS5DjduK2tDQDKTEZ1C4POHsXIDlnnPBSjggKtX1kyberZvEs
H9Wz6GkKXBj3AROirAj+CRn5g7nQF04LlEgLIHs6oHJ2YPDiZEKLtkWxRmzD+nhSqN3oJ+PO/YCV
WkF23RAkvOuwiutQw7326IED0+SbT7WLVU/qz6SSW51hDJNqQTdDQtnp93UXBcb8vDlpuNtQCSy5
v+8Yb9YfTQ/y17HtEXrAgWWSQGyq77E1McskE/cVAXTnwKS8cTCFke6f5WLgTE4P4YWUtfEIhowZ
wS5bD6LHlkL8o3CGlf3a77bDZNsLjbuqBLwwmjy1DaHDwtuGdUKL2a4czOhLBUJspmmLZXG/2r53
cE3QQ8Bbf08cd6lTqNz2KOlDhXb3Kk1APO9FpplORp2Wr2S3htBOLgk76bY05Y5fRqLQCgNWviCZ
HU3E/jDcfZ28ruAGFuExy2FGL58Ixa2p4tDHdyB1kWeOesT9NxXWm2gLRvTkPv59Xa38xuP+dQer
Z7iGCRhNoTmPtWT9dUNd1cRxSqUIb1Nx134Cm/bW9Aiwfi/Pli5Ngt1Z79lvX9JvP5pByXM9XZyn
xYwArR6UVRMKaYRe5WqxglE5pXlqDEOIxKaOa9kE0QMkDeWqvOmR/+7f3SWZV+1xCVyYlAzw1swg
DUyvpxIpiv5A4BRgI/rp4HQRgO/Su+lWZPrIYVeinuAAJW/4T5wIuA29UmS8rZKpz7unqLIoTzsE
aMjIJyPBu8fdB/1NBEigWqmyqSIkKueIq0IxUib+j/tISYEDs79Nq5hDPTRtumYpsaksfZ3qBta3
xz6KmF4Ppq3C8aLxTem8+JG9ib8UaERNM5YNf6u0l+5TjuxQmdVqvC/pZyF8Gm/ZW0xALpEUx3Gq
T8UMeCf0cUSPpmNukvd3v57+++Aics9qNCb4421pIaScQ9x/D9BygPskK0/Hf7GzKXZZejMFB4+9
1MMsLAkgeNZfFzMDBft83bbxfySiFXb/T4EGYgAKvmz/hReyrAkJm0rOMBwfy3NA8HTHGPt1A4Xm
GsRhtzdCGhpkhfyrJBDrAyU4CvJla6i1RMYpZiCSUlur0m/3LvdqH9qD7CgOxPUw4Ep/Grk5PH1S
26KpSKytPlElO+ZEGzv9SyTgiUgKOnCzJNME0ZHdkm1Tuz2d5XxRYoBVtkfX/Ud9N26C5U9535IN
dEcP5L0DHfR2rQVCdvxrwxtkGLPWg8eX1bs6Uh7NP/U5OpfnqTJk+/EvBtAOrRD6RsCioA/ulEzr
0w5jP65ObiBio7i0mYpcOSfdpDqXzljlpNuMpn3ExAzCYnGlppZ0R4F4UroPCfYXcuLO7HoPbhS7
Svg3Ex7fVJK2S9u9Ad8+Vqyr96IJKgTdPRCAaV1JE+rtHptt6u6NICueTmLPJAczfUbzFaknsuUi
SVBo7xR/RGp0EJsQZV49cn8K0xB2B7Ovfp23BbI2D+3UixeuiJNxiCqDcJbxyWxcM2bIsBlm8FMV
bW7U0f21B1M0o+OEG9BT1HmNltCL5RokfjpNQh1MbcrwVimcu0jlxN72p4Q+2aOQuvwL9EA6Bu4T
iTAvrsxoZCI0Vpcbc3YdwxOBat3e5VUepD4rtvvsln9LOITr/a7li/9ZjYgM2v/t4YJT7hyz69kd
u60O9HP3iCNcaVhqqz9ACt3P2QTWSxXLQyC5tAhs6YlwiBdmXhSiOqbSlwahtmhWGadJEB2+L1l2
2vv7Yz9FrONiWle1eEy5EJu86I7nuScE35WbDKl2mylHdOH8CA15zJ5FkDkAt8mc6SARwBjY/cJa
ORe5FlNj951eXh3wofJiDcFlPB6yh622yBXQkuyehKrp9DOuzHdU2bwTO826gUJaiNnbAzzByWIv
85VmsToHqy+Mz+1YaX0SXU09S/HsYigiKh8tGfyrpWk3yt+qoFZoJYRMV+Qdyz9SdHPnNz6uJ157
dbrrnlMaCZ3XJfyrsgHW6p8hGJ1RBpjdd8RTMq61lIeW/BIxlWX1ePbncFAV/mKBnjclAhw/xbqO
h/4NLH2ztoJgJEPSdvphoNbQTYxNEVx7ntfaSYRV9tPrzdP9fsuFHAnScCAw8j+P8xCdBCRNdR0Q
tNEg6m+Azim2svlZyaJP9Dl7TICQ8/q/slkU3hu51EXK0wJO51uy5DjDWWiJUaxh83mIg17YuBKc
cf2OxC8Rw93CwTkcaM3cx5/l9r7qxapEZxZMrA16HpZ+oOXtyLmFcIojphQoZGhJUqzSAy3UT5SK
5064zG5/oxYD93gejsBglFwvnHB7L1LsdR7nK9nFbNzfoaP396/jJBwHz3nJrZEP/ywUmN50YdMY
oDp5QSZHAldH1kwpt9F95KfX9ZB63rbxAh9gWbkPjfSN5lkn+dXVeTZYYR01yAMO627hBR54U9Qi
F/qhy9V2k/z/DZIlowMXRbfIPg6Lq+N85OBLbJbZb8cDuj5VOLFVlVJKZiJ3t7gNYLuAh0z/FvwR
D1EJ2kDfMqdoyh56Z9hD727DxxYqeH3QtHLl0YvfR4VcJqf0iaviJK35AYz9po7O5ozu0xbCpDob
SdbeC/tTJF69UV0oTQD0iDSWL/PpJtEn63nPAT6xRF5yldWN9mv2PiO23OgcnVCwsBm/1DFxrEqb
WlIs6w9i6zOVKsRkBA0pHYUTeWJ7KCSi1ewUoKYFHjFhjNhw7M+tCo3M7A5bg6T46GhUt3ywjugz
xvLsdoUE5B2W0iKa3kJRjpKRebTLhi80h8KoXYfFC0Cu2WpG7iGrQVQXHZ2Si1uF9ulhxQBv5kiV
w21guqFidQ1drCOuBleTfFd+emKbLTZ8YUytez+MmqyieLosqj9V9UohRuhK1whAnbsSKBoJQu35
2URQQ6U87H8lnedGBk1w/dxqGPH25jKTsGXuNlqOffOH2fbowBv3EDgwP3NLp65o9bNO7CdH9WZ7
zmnPa8M/EQog/XsH/VyjVWetVbNFiviKrg+SFHUqpQcLZbZclJAvn8lhsF8Oo2y2WBBEBRSt5BsH
smdgAuxmJ5wadxFYbK/U6bCSE9woSibdcHd50A5UD7KiVsdNo2AbBGjJ2CLhb51AB7LN/GYbGCTK
dFa3w1j3VOWBJqnvhQEOOjQmmaRLOgg+yIAfkZPwOQhrzd7AOGPMU2igrPoetWSomQVI7E5TTIfN
JOPvNY7zwbvzMF5y/7uZd9aq4LDzjg+P70QT090hGIRB5e+lDAYk/heluvO/0qIThy+7eYCtSw8n
RpbYadBbQSWwuELOhMqjssXclzj1GfqSklPZWQ96WqMC2CHqSW4OJPNxXyNf1CfGJmYsdgoW8no6
A8zaHeL1Zelpg9rd7VuJtZbhuivhfSUb6b7XgHQhorwqpOC1O6uj/bqYrPR3xPNtlNjD5RE2T/zQ
t+cIanbq9Ha0Pw4QziTDRIh0ablnBDzBK2bSH0xFeD6iOZzAGs5ttJj9vCp616oypjU+2nUJmPNt
EgRVhrUd3H9kOO0QDr9n6JUf1OKE1d6kWMCTJmpZQadc2JOmYBatb7YSL9i4BeSQgp8BPq66LXds
dal/W0oTnDXRXkpEZB0nG1daFJZENmQ9tjIQjvx42b6uJ6xyIiuqntuBbA5c7Pql9y5TAn4fo/T2
PNsOZxm7ujd3fbOEMCdAzexBk5fMXhW//tZvcOqmy+FrFR21FZF1mY5Dmqj0eKMIwWGBs2uuHAav
LbVJTdhsafuMa+S3TQ9uaCEGbQRqFwmumm3WL5ltFz3Z0ya4y/2PpmERME0bHeTFDD++4SFk7jx7
t0GK8J/NilGpaxd/P65Y8XayI+ZYB6g1eOklWBUVir6wZXdAA5XHOIAPm2q2gvFBBWlCMTG0w0Jc
E6o0i1OpUM95RFaILG4TJ6QVseYYF+NbO6HwFudTdFgzhxLO3Jp9dOMtuwFsoll9nC2UD4Zt92gF
ivIWHI8eCedK19xx+NNQxp8CxGJJUaN8JF4HITllxh5/7DJ5rrwXpXa+5432RyiGmB7zOsTvXXxj
cbnjHKeh3hlM8E+FR4DbXwjGDSWZXzbbT8L/k9zzIXxgzpJM6lWtRtgI6JOXdKSS3urMyiM7Etov
CUboF4ST02e/aoWpUSGOSIGqn0YBR9FtP/Ts3/vKBFee8Gf6A/lcx0ybQXAn0ZGb8yIPwjAmn1pT
zB1q+15ycFpXcMBX0uiS29wC3WsztQ7uE+KirJ+CZ08yT6TqxtmPJ2OL5hoBuUkMXihD+2LMQLTg
hXezOHCLwZLHffhgt8t3pbic6JlqDLTVLt/C0Pzh6ZRGU37TZIYgTwW8p1y9xhR/UZzYfDfgIYkv
P1qe193EFOL8CY2lQDUHCV/QSb0jgRowZDOaAtNwcpRt/9akBuEqwBAuAlt78hK1ixH2l4YIV2Rm
MbP4GrUIU0SGTjxWzGdr9/xkqZsGFNMUKqRg9KIYsVnWS9HeaFF28NMUcKnvyyLRlGNUcPNqBLNI
D/iLnBTXQmmQdEaip+iTbSl/uBvFK4mJGRZ69OIaDIKBO9qWM0/Ke+k01ICyT8Le50hTTj3LG4qM
AArC/oE0aMSpbp0TeJPUF+Uf7UvHC1JmbY+ttKB5/4Ck4STam7PVRAOeLaOM/S9eoHr62RqXIXsx
swQIkvRlz0IgrCZU+3oLj7Pu7Np3vQY9gjecejkhFHnAqbct1FvE9BelJgK5f7U3YFRoOlVOAhvG
WD0MDcoNkVRzZ4+NGWccw0oqagpK+TRHEK/UtxdUEajzs8UhmZ6Lgfu2x4DJTrsy/82zoe04PPEI
zfX3Z0xy4H/vkk4oEMeWUfqGl6rCMPI0o/13MMcB+1zk6Wgx3cxeZMz0Vn55ftel4Z1LKzBC9PQa
Wxp9jO9/y79bE7zaMSlW/UGtsab6ECaVzMKVHn4mTw53GqmpUNZ+X5Twbms5j8fo4Uywkw3ConYk
TdD1yTI5gyKz+3KANoi+qswkugbvlhX5IK6IN1xyqgHATtpYN4f483M97kDJpWPwaI7Rn0+Gg8WZ
Si0CwydIL4mrmfjGcTqeoITU1i9XmDwtf6YqYHKwXaMxGGTvGJ3i85s86tqcQZP6369vz1hLX5Lb
4o4MfdokAO5EKw9OJ7U86zNQvmeoOnknZKHOfOFVdmzG2o3LkmmDNw1xSQudobrJAxjGxlxS3qS9
1kmJEgP17rFEWZPrc3CppBvwztt7gHQVxgfx6ke+f8sSOsxgvwJM6hL2fzcr1XDFkl1xCCeBnDRi
uAWqIJ3ojdS+vFXe/Qfwdduuso7kBG0Yflceunq2e83g15bra69rUCwmDhWbIFb3yR/5EIxE3GTW
25D/OyATqJFtDDmmaMKDkrOL5tYxPTXRcfB/AUGNzLYAwCCJDlD5cRIGt8OttVpHDqp1GsOxHKGA
KWrciTSr2HC8ZG4kjmvwStQa2/WosNO4GarxWdMpGfas6BVK5fuopYKydJnVHtcyYbx8rI8/TXRG
NXoYiTRvhS0Js1lliCm8x5tz+BJk0HjO2QUBhDl2Py04GXZl7ZyUiAIqs16XtF5TZd3datI+yScE
VpEzgwKiqj/nGVprdZU0nr5jZG1kA8GaCdcFajDijnkPW0bEMrjLaD52rUAwFjMNt/fGveplnhwZ
AJXcnHuDGtA77qEUd1aA5ieffP9gJgbyDRMYplzT6PClatBXloynnGFqnrGR6t5MkcoxiuhuIHko
VAnMBVUhKzM8qSYzwrXvSEzlG38rUtjH5l70rrCWtroWxZBftAzm+G2s1kMoNW18AzCgwOS6Jhiv
28aZU3Q/VExemrOI4bsrdqeXzt0rTMQoGEvBpiahYqFD8lw/aVPOZlFe9gSN96cEWMAX5KZpE0Lh
yBrKlv99mQDDxVZ5e249AdZvqNc6B6KDBF7G2RtNfuRLOvlF87fd7RrEDox1jPEwM7K5Ne+CYapN
2swK6wk5Izve0q5fSXGPdUWSXlw7dV6s7/YqOfKn0eW5TKEHRgHrfq5vik35jvzgPdXAL54AjEBr
gTF3vUB1WHlw7WoCDYbNwNNAdb9UOTWhH5V6IhjSymCm/SwyN1h/27LYnNnPAYURLRaDGb7X7zZz
vdA2LuaOLYxkL52DWyfT+ZBp+hmRVT7HVMLxlJH7JV5t2w/5FtxggkQsDOYLUqwc1tN+zR2wM1CE
Qdg4bdzMaL2/DKF5EWdFLJO97yjbMgob9TkQAVZ3OmsGvlvec+DNUMboIbEWCYyNMkK2wgyFdQxf
QngmA3lJSXNpn/rkQtgpnR6wq450n6Ask4YuyAVC16ObaqqGmJnKypYILXLS15SA9jHE2KDEPoj7
GIwLcRGx30TZzMtCO2GyW2IAyrh3m8YYE7Bb542VJavZW+gugqxottFG0Q+BRKVDKxzbCiNVWbTu
+YuaoCUWharlXRCrwSJskLFDNNdnM3MkttnMYyj9bYp3x1+gwyXXkAws74CxwmWJQbETN3L9K7/2
Z5+Ek2NPcBw8qgdsLIj+QOwHyGqGLEN2Syy7o2KU4jSiNCIKisloYUkbvItXvFwEWyhlWu0J/VEE
ugYWVplqeM/AuAeWxOomhRxo6L9wNpvnWWVHC+Uatoz+I+FozKHlc0WP9xe9Et/w6hqjkxR9iGkd
KL0dcDqMwIlgwY/g03pQZspp7YPUbGAAavSnmJS6PwXZwNolGi1RxsGshy28NeeJ22Ufs5rYarFy
yy6B5I2arzhXUFLkuAwo2si5RsH98e8WUq8jWlWusAfQCv10ZUAPrLmhagJZwY1NK57DV6nn94xE
FKRSDkx+zzRvJgARP+Qk14pdsK0HKg7+BY/aoX59myJy4VtCsK8EncNprRCH/C1RsiLLG588LUOi
qCVLVTcy9glLdNTsVw4sXGRTh5+yazyeB9JfHe05um2/jU69wYUo4bSX43eicVm9nGhzQQZMG6IV
dN11hR7utiwVPaaghhci5YTK6zV1Rydr1mlB5fZnIj8xGgenIm50F9oTfgSzhzYi1Pei+Gs7ylUo
wO2KuGY+pTZcP0dUMWT2PZ9clOCPzUOg/lxDGysntreRylDZGQRaVj8fO+yQwWLgT9ReqJ8Km9Zu
Yf3DkXWtBvbfHe9ngIEzPAEdlR46JhEOdCvTm6JovIQ47r8IF0vChLguytcmWkasscs6aDl0fVDW
Y19yiEBJAZoin35RvPdrXQQdYdalzlkvpwGUngweQy3230eRm7grFPsmURvL3Z6AMd/BXm3d6mOK
THXO7qq+ZrI/y3TlDKvwHNc6hJLxh6jPwaNCRDbUbsnMdsMH5r85KskH7ejhFEEEUbvz3h4Wcg4Q
3vYyqJdeKFxmk82fdpiq0gskSh5/7TrY2vqsIorvBq2lPIBTplvtUdB5w2GdCpZoz6qs5GK8OSsO
WibgriTRjHf2tfGSZSuMW7V94UVf2Kxvu21ZfrhQVk5xu663MM/BxMR7qe5h7N8u3CcCtGWdPTa/
sSS3NFlZKd0aFdM4KRxomlZ3VPcEK8O4HofdN2h0h1HHaL8f2XzFG2JvWhqGJkXuejzDy7jQwDCu
oQE8aOL69H0nR13/2PJsMXoM73ezVA+17Bzzc3LT9fYMA+6KLLyhcKlTBS/44NsLQSr5EpM29KYr
TA8rv9SmdKQYdfZ9UJOyiWIUzV8lOh4LCPGLDchn+qzG3Yk2UyW0F3jk4HzcrhO9/2D3mzCA3Dpq
XdNLTNIw/kKocKRvqNcq3IB6HvgegnlGfQVL31sY08wVfSv5UmLe4xBicy+cTIeBPYSa+wBWV5MF
4+vFQgGAZMstyEVgY8VVfaQ3E0uohH3HxAg+0xkmKoTbzv284Ac51dFU2agSSG3CbPjpkoT/K2ar
HOJ/MDvDysQ5Tc32EzYSUI1WrYjQPa94XBJGCdXilS51Cdl3QFw860Lz5jbg8UuyyK38JMgnd4QK
k69tSub9k663z82P4NWQEZwZhMlYliQve3QkevtNgAkfehqr+NET/OwQ4zd22w58kreW5rk43KML
zZ2u+v+k6+liw8nKp/rJok0LEYekYTxMjGYim7D4xwb5GggcFUJEN6eJnSIHS5cwlmkjIyCzKzgL
/gIVCcb2zIOpRGEz9QSl1+YzDUqPQQ2Hj5PEt4OXB6QAnpxe0IE9uwuSj2JkQxkMmZ56/dkgiYAR
oYepNo8+vHkQ1bIhjXNJWQ0a8JA8F4kyCJIpIkwIAcVaS93UPJA+T2vV5hdC7G9vswb16gxOQmUR
yPGhHG2U3FnkMk3ZuyKX7dJRPVPkScEPL/aUDR7ly3Hj/sJcZwaE9Kv+6V1Tj4vDujcpNbaT+G6a
3YzqLChN1/JYzf0/m83S0f7YPdpf4pZmoXUVNi3B2ebMU6sabx5uMAO2SgfJZIlSdKKYaVcosQwJ
ya/UzJksIMZJV97/bypkdz7a08I372rXWwnRHwcvrA62SuvmEGEcCJJA4j/0o/SOfgluOpZOjYIR
+ZmVhdG+UBNVFv7AQjvurPq7pyockGAR4RM938y0Oj8Q26mbDBo5s7LIbeV5vStvFPL26i5sxtUH
6tW6VfOs44hJncUALklkiLUjIcjpjbhtHawL7HyvMBasCQpmrcUIcYx7aAWMJOFrxJstfz7h9Ott
sEjb95HJJ2HsM123c97EhDtq0FbjCCsKxZK5DudQod4fq66l6qAWvHXsidCOzMNhpWSsdULfOwXr
hzBlaLJjp3xpZj+T9L5lwLj+mqf1U6ufI62D2piAJQnFP1Rs8FsrRpRHLym6EdrUySovJBiNuhVD
W6+xtPWFKEiWUU7oSNrNZd1u/+t1UjxyfHMJCqbdQrkAYF8h/V0syLSvreQvb0U8ywzv0pp9lfIK
UNkfsD+hbVuNmHNxBmGMI6g7glLL6IXmaBaL3EyOqweTJgfOGGjju7EGuOaSOnbGszkO/hHjHjTH
I3UA7f2X8qYl3SXabrrc1RB4aAcYMgcxlMH/IZUyJ3951xY1NZuU4mgwlHSEYxOV8qYR3tNCnB8c
e7DbUUyIBRX8ityeNCuWmT9USbIwQykUAQ/0AHWzSe/dEcTjxvNtA11bUYyKAirkDq1RXBO8AB9Q
3GoJwABfz2qE7z/7OiT7b9lHaQu4bdIxjLybDid8d5gy7AfzHSt5fqilAA2EJf6AV6X5X26PWmuD
b3p0ATxHEGgsndY8erKyZSGFD3B/E6HWvHdiS4hSDeGQftpKjLpWvQa3+IgFGmhm6M8VURVtev9W
GXtwibmK7gYnJ6JHYMHHnlcwoJDbcyJcLyZHPIUoIYvn8HkQDIpRMuXUhhAqJuurkYDx5kDgpKUu
FurFGYcytvaHwK1vApnICj/r09iI14I87kBT0fdWASE5GEXk3zko2OXvirP82s0bHLRWre4o4+k4
E0GHabA25Uw191OhPJKGRyYZRW26xV+zZ7zTOBZFY27WX410RN0gG9iUznY44YcU6lQI9nR8Q0tt
RtkH9bTtHesYBnK26UQv/IsPdQMWGvBCP+t5o4CNifyTOd2ilgIXbitWlcMi6Kpke/4Wpwvch9Hl
mz6tnooG4CV80iLsKS5Wyv2s1yPylwQwYxYZlADL9wAo89tqKq+p8d2gTVNL+n6bAFX7p2xfhqnq
5bnLj3zQ1U9IAD5Y1Pt8bNhZ7HXGY2WGgtGTEtLzMCyKkmT/TQIHVpK8XSTxgjbtgmq4TFeSb6xD
tPiazok2PLN+iPJGoMJqitNcANLNo8ygROaElObnoqqip2IpVSEtYCPCwu+L7j+ndNRH/BMBFKgY
mkU3Gj7Fko5+2aLkkxabYd1VD6N2b5VrvcIssTeLdOJCbgEz0Fv1jMBERFwMQSZIsxbaXERNrWNV
Zqb8ds8xeLaQUc/nj2a/TdTRGwqKVsyaGiUfir3jxP8/C3jHwMajSwco1paHdRiiDG0LN8Q8RP6e
e9LIatfI1kq37LVZKMHODPZwKCjeV3WlBQBNcsQ+rjinlTpPeQQH/QabZ5dzkwMRcxC+YWbdkZpS
9n059OMk4PsI0Y1yy+wUguIWPg2e1ymosaM9WkEk1k6JrPwMg+dBklm8D3g7zb4o9r/8pHk2hcon
1P7OQzKdNS6O40yJW2DEDZEzLpn3GWP++JoY2JOlOVlIfvpCmCn8u+/9W2M84/yTSn/+o3QzJ12J
MWGrQ3rZ+vW19B/ijdeqxanIjVIomPoKnXQgrmm0Qu7t7mKq3YU1k4AdweLDrHTLdvD6oCZenR/5
5y8+0+PLDbug3/Wgcr/3xAmFaCwBUFv40OUEl+Lj7KJUVwHaNMUstkNYfgkYYhuqEKYGjfNf3bwo
esWtrcozabHw0FXpqXwSv98m73xwtcdFiqIEcQhuSAWb5dP73+QSdgHGV8woQwc4goFsDk/+delk
H9+FteWhYKDKqdyM7YYABQPvN2YZ24hHHBnpHgXeBS0LR2yj3GjlBudbEZxdaugXUqcTe7LY1wFY
BAKL/tEqm7NMyCeJ8ww5uFt7sdlFmcK3PX3XDK4l4QeCUaMZSpAa5bdC5q88GAV8StphuZZPR4om
SOoYELRj6Q/YB/LXGlpPI7pkuw7Tb+ih2YpQyZwJvtiWlcG+k+6JOTmqM6vfnMAxjn15Ss+pA5cN
pKcWdSjGAzBNjyf9+dvrFymJlXKWjiWBcBqvBKxa1bk0IUTHcCk4NvciIIQU+IFkJ24BQWz7vCz+
mi4/aekZ3IcviktXgpcLEGF5OGrwIDmtVPsiUtvOTBcjyNNf04HNKfUkxfuNJd3eluWUnqq5tD8H
H8YERo29nGGiGYZiF/MRSzMkFUyfDxY8Eug+gjK0nEP4ImrbMFe4xsnYjZMk2G48B1k7Ynyw35jl
71sHxjY7lj1mLAgadmba7UTpyTocjPXw2NLzZ2X5aVovSLqSLc5TUUtdGgyBeJXtbSAeNaWT5g3/
XR19q26LOHuABh8OGM+SQdCyAqb643RprEjztE5QG3lZTw9RocHScoGkcxDPfymNnmrPV3AIMiEe
hauMmc2Wf98EABIeb22axR7UknB6DEuiBafnWrudwv82thzldV04FZMcaHQhaQx1Tzu7ENcDIyMj
F+dti1WbRtxOCtwdm2j8FDMMlcMFqlb3YGG/5TqKbGRD04jN0R6RIslkjvpRgGQPXiFAOSSIhE+K
4HaGLvWbviwn4aHrAyBXBTe58uj2lmm5eK/L38no+WrK9GOTNDLELuQWMdkPF+ZY4cC3/yH9yFfN
pZIO1AkrbNyDaQLKAi7irWS8qKyl9PYfgZhhamacnfx3ET7Rdzrba28skD9Sv31xtQ1BXZhCylxl
xcsmSnUdi3I4kubLJRyZeqlNx0ovWapAYv6DajqbBXuYdSli9eyQ87Xfu0m1zhuBJcxv13F6GffT
NozdR8LuhFuYsU3MiEiTfqkon/1UjEkt/emWF084WG/V3aSJMno8cOLdwf/++Qa6A8KTZURH0hfe
pb8rUlGNAsyUwqpYroyyyRbORsCFAK13xXpn3TvHARK4HLb0jmC1bwOPhW2gsk1A2woJSPCKu/Bs
djr0oUFnQcTwpKQchDcEdqSvNXbxX0NM4geU5OWkYj624b2uOqLXnI0On+XhUXhzPn1zlsUbIHwm
RAZwXsAFAKVu5IzOEckWNPzszCCSiPL1B3Ptqv8WSA7wkx/N3pbaCTEyY5KgPUJNplWV6kfVmaus
umXg2oI/z3riwYRpDCWKWxLjvUfdR8LHBwk3/Tz9C7OOeLIdQ0cQp79L/4z0f5u4umbgE5w8oBny
8pBehVDFZmeuYlQEU79JFsECLMfQZzvJTUbYnZwMWxcWFo8B+cQkJWKkKzfiZIocSzQzo4e68Pmk
z9KlVu0UjX1wTd3DGUPW+IgMJ+H768yiqg7Qz0qqT7Q7MTMnQeTTO0+NOLDbXy/hf6D3FoEZxtPQ
2aOFs/s7EpBTuErvQ6k1TXDzH//6YeR74VmjM1ctl5kUey5u60O6HddqSLseGpFmlto70o3sA2Wy
s+8FizyLheK77KTC6aKfVgoFIdwd38ynfzza6xJAd56EMiXzlkUuALL1r+aKXJEQSH1QiXMcFthN
LQxP/TjY+H8hDmj5nSAomiajcY7dicGYUmXcyvI4lw28TwywacA8fjRyr9uW3OdRQaL2xADU+UCz
qJbYOtWDsUMWwdFySnztmFI5+nH5q6lnODqs8kzCDpElHwjdOMyS/LdpOsOUThVXTGQ8S/9VGdZr
TgVlKGffoS9Ni0WnLVBzaLwhHrGq2kH4Obbx8pSO/A55JJAF2ulH3PSjwzWYk5vU+z9CTcgHEaif
QZQ8HBS2UuGrH3eWBp88mInffIekX+B49ChKKbcRZNPYPrWlb61p6N0d6QHv0mfKTeWcs1K7PtiF
d6gxtp57roxLkW31EHERIEbYyTcvLUt0pyVM6Zy+dmtisf6MMjAruDUpPfcBAYxcLE0e+WqAwABf
8pjQPq/x7YjW/1NMcTHXLVU6GRg2vJyflK9QuTFGXeaEgfA6T9QADpFAFZzKuIaG/XxlnLVleHsb
/czYqKCdQj4iKSJI/UyVZuyR2JCOjPp/BZcfwwa2kKbd2NPB1dXQFAQsr14IhlrqhBOKHg0W9xkZ
fRkfAoQrb+cAYXefkPUuQ+C0dxRdpoxDHLHcVqAOSFjiCmD1TYdveVhibhCrJOJcuh8n8yt+U58Y
q2kdNmIoj3uJJ/ghGZxdmB799tp4gMQQM8fukhqJRWUsY4W3c6naC1V0yZgceRV5MzlDCJci5oH6
0i6Fd/OrEbXp/o0IAOvHK293h+HtFxIpE8seYix5jXwTEMirTjcWEhxaAgJrojuhuomRtXv6sCJp
oTB+ga9ZvfxVyEfHc322Pd8kVA+Z7TIibdFn56t6RcKHjpkm7ib/mWHh78R/HC448JsdJwIQzILs
sfjOq82+4YuQZts2eTBtgOjD88nuTdSODpKCdOXwmZifJ4DyCSdpg+tHd2vm2wocWVfnJqGsoBXy
eDm38zbC7i2w+h/IcOEE5dTazJitHNqibrSxTmE1J/wBfKhRw6GYO/RLoFrqInZt0cW5scupROah
Tq9RlVRXhRftfrIe3lZdapR4qylEuAtH5prz0S/tGghXx9j7D1Q7UOIwGpvwwG/V7+r8SG64JBms
3+STJgbYid5zdkNRleyWIUgWMPVhHMp79r7UgtIG8YK6JQ9GbQ7Kb8UmJGzbZ7AzQ+pmk9yfsO20
ZIrkJnT+Tf58BImzxEpU9Y2f8H5C4jzXhTdqrXAeqXGzpBTjH9mw6A/RAtqvYOUk5LScX9/54N4j
g78j1Zd1T+Bsq1Wwu2FGl8H/BdfpJxmqk8Ws6BeKD+3bUOeadzp9/6PuElTWkN1Vy/DnCNxwRUtZ
Fyq6adCtsz445/06S5OsFmClbHonl4o2rcUTxw0BAdraO4zOXASY9X0Cp/u4nB86WVaTlTsPw8Nn
E1tsf8za95YkjWD9x1anKoeUCQkARTK/b9/i5MEZP0uAPp0keX19iX6ZTVL3RHHska7bhOhayE0x
5SLlYHRPtv89hGtIHGBAXMS0sXfr4K0cP5CLWsZjiizbRib8wKOzhkXW2DlgV5SeADMpiRYqGsYA
UCrCRDybFeUBW7AMyL1fBMYIuZb6cm7mBayypzCnEJVScBAEEizND6EzOOgQhxqLhaamBpRrbXFg
9r3QkUBQTJbwHsoIel4JxUSjtjXEPGl3Stu6omfpqAdyQglUWl+kTiHe0v+sqlbfc46uRgROI5Hk
+hWa9MUe8btafL4WwI7WhNhItRBzwVPbZQl1tRdhJsIggHs6lL5wLb1SqYGjISiU44N0L1k9Q1uB
vUHmWQEjV6UL60o0DdN1k0+mBCOSXInWlu/qETWka/jJqqa67E3IQlfPs0O6bogG2yJQU/kHZ+S8
y0dA7OpaiWywtZzfWv/+yV8xpHqKYUldSbObedfo9btpBK2QU45fnebSaLv986+15vXDs5O5TPoI
xzD9CGwHlIa7RAhr4DKkIMyZ6B8/H1OBd9pz3Z5doQEFkm4ASEVS5mDJar/I879JCuJ/tC0OLVuU
YzoM3PGhf9Mf4hbe+lnuXAaXMYxiYD5hXIViy+o6x8kJUL/1pgPDgF71gCFzQRG/RxfQS/MOyjiU
xyZzPeZhfr4U89bZ7w1UJHyVgM/uxgQk6uEwFca33TOzC/+XD86UBrDQm72AzTLGRXCXjTZJF5t4
MnOKlOvHyWT6D5fW27sI0BfZ7zj00ZXGOZM6dxOe+ahvmRYR8BGnAaVwWtX1GDDJe4bCvSRyOI5I
wXCHbwQSlGoDx/6PuayGpJfGcUaoz0mxT22b6f3eTlKoTIb2MA1brlvt5ZynqbCJRJ1k+ziZkj21
c+HJZrFoRSQXBNjRJR3m5qBdoOAkYdWrW028zovo+sLVfdjWz3fNOwXEXDEULF9a2T8Ox8xSksNB
Ckl/HUOzzWYiTbSLUtf8vhow9ZWE23IqXqNSZ1Q1Agcw8/oFyi/k1uqJ881Gv/ofPKVDRxT70D1X
SO3ceP3dxoxBUcq7UA5fg2R/J6DFK+zqwwKLeZelbOzwus7qtSITqgHHIIKiOxff9vtxRrv+3/yf
MIH1qP8ivVifPpLN/kYfy/JUPGUkTZSgbx2paL+yyaUM1TJQm3PRm98U1Cxl2DNbFHFPB3rXG25v
m+/ZwRTMqJlZhD2tzeD8xFJf0jFbN8vzcny0ASkGGN/OnmiO04ei6VDHRc5xTL+wO+PvcNZ4zYK+
AUAFF4NLfrRQo61UV9YUBxkPHhhY/R52vjGZHLp8LyzBfSAUSlnB86dyzattcYhckqq0JZlnKUQu
Bn4ou2uMrqol9qXwaHMrVqspJxL1f67/U7MF/v5SYWRGTe+erQelbTfv1zSlpK3oI45oef25vGUy
bmP1Z7+KXL2oX0fU+tW70WcYKjTJYvPZnVS/q6W30KWJQaUABBaEd4gCMNdtmqbNdn0MzxrBZ+3j
aQk0dMMtQOnvr2ynRYeXBt88U0HTgrzC0TvBSLDSX3oTC3pRx9Xa+JFIgC3AHlMZSpT9ppM3qygr
9QUwBczu+TKlZGjiV6bIxnRB7p+vGqLDiRze0FZPTjVU9tw5UouV66PHGJD1sNm/Nrt4qlXycUsx
mHcJwWPA2YJRDjXHzyLTUTzRGWQ1ptMk6Az6HT8HKbd8g8vOOauu4fDYrc3IfIYb8cmfL30mXnxG
BwnC2wwhD6cPUGP1Fird0E3rN9SMnItoDfvQf9nZ8A5DG6r/gSnZ9fr5pyyhMUsvi9nbvdPmwr+J
PRRq7M5mleoOHingkS9q1c6hfiChY95KrZR5f3jHX0I2nqjjj15fur59IIHVqx5HFzQ2JwissrFH
3HYlLYI+zfo1nEzC3kjAGZr6pfY8nNnRCrtUdoQa9u057OP0H3Xo4od4UKHa60Dg1LQMY/7ytm89
hpAHYjQLHbfM2Gr6nRyccxTzoyDTY4m/txB2HW1EJuVtjsk1aPaOrWDk6whAd0suQa2fg6dNwrhq
rv8JF4IKsEtruzEqXBHW5DcS2pvFsSH6bG+17dV9IOULEJCB3dVpuJhUT8+wyc1gdEPBzdw9uekq
vNKG/9jgtPKfSP9sf2Xh7snxG8EbDRIJ1QM2oPh+sm2q+OtdKsUdUUKBbh8s8+KwJnNAlXiAa9HF
SE1nVr3oNjrSebB8eKbZ53cGobRGDM5/pbpZ2HL8fc/fBlem9kzftyTCmaetXvq5gvdsOIb99KuM
tK1xaDWTL3Kwv//nCHfB+BSdmSLtHDSVi/nP+Cq6NKL0w4DaVSROfsTttpx71jM5TBTxE4tf0uPA
lFsRNYjcF4rupuSHrr6OAmMH9hRdKMuMfKgVaOq6xSCNBtInrjzqs7E3rFHppqswNBA7CyXdN3uc
kZq+jokwNNAfSmie8fUoMjD8xaHx1MlckNfAQp/Hv6l0VCMS8rIJxe/TqafrA8JeT5UVsPklmgJC
Y/DT3UGb5vLPaMP+Vjskk9zJOZhAPjjBHuDMBnQ+hWf9s257eD3wUKlBtm3DeFrAROTsx3F08+BH
QgcmOGz1Y7YLYyovqlZi+NALgJNyKsg3vxMUyXtR/1q6vBFElzoxWBKZPTAhvK82bhQN/SzjOJWc
kb9q11bTvvF2zYZR3c2KNpUgU0aszKZSk1BRCGRr98CfWPsDjL+GotMaUHQj9lUKXiux1Hh+RJ4a
3utSRaheLF2mBQHRzTZWp/E/WBuCsyUK9pigQQep5QSn+D4TGcCIcaGXNJtZtKm8ENvjC5VIR/IM
OGYnL0wS08+KR0gT/URSJ8WBjv5tJpzPYKglyv2kVIp3v+oYr/SvaqJ1KwFfvyElZAiok398easc
DGkvjblApz5hJScMojusq5ycwzNq6j6w3Gnlx9zDMOxrbB7P9ryR9ofOhYluAmYG0idgHHeNPTb3
gG92caotnM1rPjCl4ppsNedIk66pT+tOXDeGrXQ2SqKAYK5I9mI+Q1jBqJkg91PmtCKs+Y/eAV8P
jZC8I9ZFhd9TGE8upmj9WwQB7QAaDPDTWG1fPuXpe+LLrYvviaGkfidCLJmTR93LY5J69bYtyEYi
Wv5qAvHbzVO6uB3vNEl6U+DbT0EZUiGU+UnDBrHvo205OCN0O82Pq7Zesp3faxQufgiTlCnNvwZB
IZQe+eL6cc+mE7PqCgXKQA6FO1ODux8IgZbsk2qNOr8ss6NMDMzed08KiCEIjo69jJih6tTGFqZ8
Y3aqpAffJbqvhy08rLSiHoFjg/lcxj4PhAt6S0dDumUYsc2mSZIPZvgfLckX8Sqko7rryi7GU+84
JXRjsH24T6jZe5cbtdmTKrg59q/9ObbdXE9Zx7ALcyiJ8EiFeRpMFfhMRSnpyuJWFesk9nAoKdOW
okZlupywRK11lmljEcbisbesFqfrk8ljXrWPzfOqspbvunAY/mjlke/rURqw15V6CfvNseiEkbt9
A7/DO2SzRpNkinFnxFHq1jNhAqynIS7Uhb0gGjFXmu8/Ri9XrVhKyBC1R1GhTgx+T6VuBv9+4Geo
u4JqbxtaYcWJ6mAc/Gw7lTp1xL37ErDK6TgYtaXPwW+R6zjawJ8ariSVwffO5/TQqlNwZPPA91CU
c9Eiq2udJ6QgVOpgSTW4QvLQGOBHg8UncG8GkNr+uTyaym5mX/BvsFlE3ktMOqbda0eyNfFmPK94
p0owcPD8FY1nfdbINWaD3cWrq85vE7dzEw6pJaB80sv7ZPnBVUa95OpvA0qR1VrG4M8lvAcj/9sQ
mNdCVSZa15lsSR0GuqXR0WYJnbVjr/D72+ctC5foh17vMEijKLxS5tisWUJGFYQxK6G8YB4K+mQL
oiWGj2v+XXBGVm74XmxzjlkeIW3k+M1vjbhiPKRWcmGjFj7DP4UZ3BuNJSWQ4m0X/tlSN35Am8JU
4EJ2w0Innw9fSmCJUwwzKIegHr7A/Ru8za84bvr8WyLbFIBirQJHLdfJjiYsxpjZx/M57tXHj9E7
USDX177hDa2I808L8FZq9ajZuDyWnXFzP0NRw7NsN9P1yJSAaJ6kUSj7PDwImqvuaNmOb0vjIuwg
VlwVqFlrY7HWywSCLzPX34iEYmx2SFuYZsHJh3a4XhTxM+YL0gQBukLfZ91wGmQBUiHg3ocnfQ0e
BJ0b8+nppYG8JDeDitmxR7sSWHJfiy01aiWTtrSc+fk2LkaM4PVH1WeRw1BXOmVzPZTfBMZtJHq/
aTciw7QIaJYgqIzyEQx1kh8VDojf6E0WU/DMEQYoMiQSQnhYTpsB0/YDIqc5PKqN501YkcPZ5Byf
UNcwhW8jJQHjHCq7ovoQrHgZOHuhXOjpPZjWUTSz/CKPz8HHv5j5PXyffPpre1PKydSmfdz9uDty
wCpKuje23TV32BYbKHmzJVkgZvesvvgIVz98GS1b5QTxpuoYnmSGfcGs9IQvNsEyHbyXI5LlaU9i
AuEWhMel66JcmZzmLsUVuIiC/VOfkY0FNPC8AP0cyvdCrqehr/p/2TiczFc+Os8M64Od6w5qMGA5
kFdzEOe+q4HA77ETefxFr5UPepqDyDWFAN5+pQ4ow6LnC2+LYYP4nQ+sycXTQK8rjZhjxANRTEl1
fxsWhwZMYFpgE0UebPn4mUq0bsOdzXRNOW2Y8smPkEJkcvaPZ+gbTeo6JdVipJnzbMImUCrEh0lA
xsctLumNdgJ7D6FnozUVMjmfdfXywMj3sYkO6pCeRzZ0M1KfkOfuSr+VSiF35US1ptdq36mWLBg2
5KM1Y+Nx668V+ziU6/tDyU+x6gurW+INWMbxMwPzSvhXVEI0XRLDLp7qB0/y7c4Vtq1CHYz6l/mL
F6yn+ChftmQeJUIh1uLcLmr6VvQqVtN02bJ/1zi3+nDw48tdUAKRMHhaPyD3ytP5NokwMnLSxEyW
j5ZPv20EazlajoZ8umgDBVTQWmC7E2ApOXbGaZ7b5lSKLXzWqE2YMagl59dT0BdRbeln7zyAA6/K
fWnBt7NPo34O1c9cag4Z1tbeR2xT6q0tRd4+BICD3dZDtw73d6krL4dmwMy1U7N63e0aIroz5cra
qR509bVbdweZksb4tmmgiCPaBOQTHZ/4KgExWZZrsrOwzVhFx8h858FFTD8fh9JoU+XIhSkpAl/+
wKwK4fd2gk1RRCClW8Y8sQG9f8DcRocCWJNWJDN++7zVCvBxXlVibF5VH04BYMMFPeAN9PW2kHVk
uwuJusFCb6ItsWpucLjIvHTsZO4my3bYneIXzL+ndf4fU9m9RusgtmEeCJ/HoglyohZk+QwMvqjq
O1F+/EQZADk1ALP4G6WAZN6P5eoy35lpT/tVvgh1Uy2spKo4mWJL8sq2Zt3W9fiZu0X5kgUzH8Rb
x62u/DKW6G3vMXLmBYrbmO/dSj83c8xcm/idYMMK6c+xAc6OGxQNNH1yGZ2X26rC0VqFFSoBlp7f
q0HyUIlMlkEhSPsnTQ8X2ALrbEhIvHnmk/t2Go8B7UhiLVQGqkjmZJQ/waiMMol2bjv8+xyXgJko
esX8OkrNYezcSrAwXNmCRIMWPxzw9Bm4Pj3pf6NhweoPK24mdFPxot2SlStRRKbkE0CgLoP7ldRD
K7VXjkGN/QJIob0yZfJwN99RZjdfLcyBO+scWjggfVTILRQBc5rKUNhXfRnphMHaEJkR0E7J1Yue
zg12UyG8cy/M0ApoJbHxS6N7TsogOOoub6Jvg2rz25cX/4zzcLefxQJDlVmwK80p0kVnapkuMNB/
z2EBUMm0slBCQRk8Q37C5ail77+E+vjXi8ABPRVjnr8iD04GGK0+HOMA7bKjuj7iIAxHIjKuKkRY
Rv6Ypzz5JCsRl+FewvX4jHhw27Jexv9bKR7VrZdqeuMMZR/X2cvauzfBbIu5jJS7sgVKV3hbaVRE
sTJCr/xw6hNRceGrT8eXfI+ur4/5fDvsu9fJC2mvmR2Q9O4aXAeuzO1WgRXt1NOBle9eegYLYHWM
vS0XOmpWF3pPaTtJolh7CKtNjrWLxPB/KG44zzAj4/Cy2jHAflYdAwAvS+vFjpQWISzEfsKvB6VI
n+vhK8CESpmtXZ8VkyqSQ9aTnUNQDpehrs1NjKraYO8yIvS9p4uYTAs2Hqu1aSahgzjxkkP6BlzG
NOB+50bjGX6z9bHz4vbHIbmIQJyMfdy1gopU4QFqy8zaZyzcKn7py++KoCHx4MpjeHqpQPN+CePJ
XZijsc/b96lmYbaA8672dSH6M3hZmWvpyX6MyKqRHn+ha5s/7Leb/10nnzYvxagjFcmIh3uk2wGp
+hXdussD4skmuGELhWuAnQqD/BvuymqIL5rEwgOOuiIJiv77asvHdV+vmKtX078I0rV+AW5tbQwT
B8unB4ZbrP2rs4bspOKDwGylapavPJti01rlBHbJulHnwava77oehzN0EWEOSNVtceVKTYn8Eodi
gfkQeQ3H30LQ4NwsAe7sMSuEG0ypd5G3SFLILf18nK6schNNu3WDHN4nlEtvbQkMgAVsBpIMet0T
pBPbDlFA4PrnPGb02FRw87MxPy3CZ3VFUkvMYKDDah2g34lxNbRrvzPw8qliQetcM8qgqspTRzuA
EweJc8XRd68jh9f7kJSn4UlRe36XujLB72SqxRo74TuyrBV0ByDZgNa1CPO4fQgwPr63CUScBotQ
S2Def8120bORHa4XyxVdNyNLWVhrWjs7OV8e15eO9ZHE3NkwIl9sK95a37zWoO4Oz0Hr2lwZx6fd
/9ssYUUOZ9TFqdSSreDRQPp7r/W1foh0wiuKWbugWk6CG77D3PGh73UkHDWg02ZR82dx4nKKIs5p
oI9sQJQNc5bYqyA2k56Vk+7WdLeB84xd3Sh11Ens5LYLk/3gFUR3AzJ5ucBxlIMfO6lU3URltgLm
VSvvItfrftyVlmF4o0mTQpKJbNvcyCVfMw8/wZoG/YUuSrpCQwtNY8FIyM0B3s7wkX8zwPe3oPb5
2POUapJ255E8rqURuHWTJCuoT4ESROPYx89AcIOtg6WEGnaOtvILF1mBQU+YHyy6b10Hsdl6mHJZ
vXlYtGpXZ8kTjcoBrO1KLROHEZGg/ZBMKqRpp7sr3KomN9liohkTryqq7OdAihK8+l+p/zj3kzlh
a2BJh6qoiIkA21bAG0iaEaIzTuX8s3w2p/J55FMYmy6ZYd/ZkbAD2XjS/tHVa6yK63l8zEv40hyL
DNqOxTwqLH3Uun4y5CRHBzviMXAQJIDalQjAjfARVdqMMSUSFRojkZAOSvWMcdE9/Uaz67nZG7tq
QFZlxfmE77WiTZYLVnPief1TgoPW71Mo3+MUCvYcaI6Yh/lZJ/9XU0jkyHVZ9wBljMaWMM7/ceX/
fEnHLFRkEs7L5p+sobm/hOIsuBMvcUERcH7aj7jHFJ8xViHJ1G9IUZugx/3XHlY2NMWt7nzJ+lJo
7FHoO2rt+Bg+gGCEuyyvA4fPOYyHW+jzWY5D+PmaZtSBeCniGo4rSGfCccPPGdC/Ltzd6OjkmUmK
isrm2RWbXF1oc5iL+Cuq14cIOGPAvX6GDVQ+1BAd1zKDg6Ep3oQX/KXkhXV1D1/y9MfCTveywFIg
RFe2GwPsQZAxhoJ7Tg8WYiU2gIYVFejgLIGTDprH3k92sMIUzuB14dRf2/m0wpoZ+qnuilcI4tKr
m58TWXdP5JpzFbNxWWKHnFzyzzV0+fQZNNkMOYr/uhjfP6oEqOW0TMP3o3qFzhMluQX/t/YYmkVF
SXmtrJvzaWwYt3mDU1XO7t9qimlVJHb4CgwHQ0Iyvobfq/Mkz6RQd9+0osKxHyUQra+OpM2B2TsR
PietcxKikmD+wTtv/sR5IU8d0QhlhPJvOI52LkOLdFJYjqvHzhf6pCo7o3yJWTVT9Wni6xeIu4Df
U+GhjT9fJdvvdGtzzLbFc6wdkDcklglBbzhSD+ifK4vToNSKNICQIyp6EgKJP1vioUpQKfsaow4A
UUWfvNb0yRAFfL4HSZiPY2qyMby1AXmfR8DJ4voPjnWCGoorJB4Nnokz0cJ6jM6/8R3Kcc3FLboh
8lMUQ5yJ3waVZCtNGo/uYgkT5N7+gsfW8LUytFz/x9eLZLQfpS+WMyjCdI9ugB01jiZdKBLakI04
WyGMnPACRCFriDz3T5wzmsVIu8iw4jjst85nLBfxWOqG3YBH/14qcxaXAxSocEyQ71nc2GYcCamw
oWNB7t252xoieRPOVwBnJShJixNr97DjQad0+kTEm936aToB0VUNaJQjhsM2s8VzN7giuGQpz0DI
3ByEdkrS/4VSG0zZEsLd8A30i2VIbQOr882pPyInqok+pytGQ9DmyYKGvbQZwU1XnPJF6KHLH5/J
gvIAP2Nd7BbyXcXlfELN1ykUqj9NjHarDZmEZ6eCtmbMpQSJvJUnBfuiYlmM9ZvOLV/e4RxdNavF
TsuzgIEkj5hO+tdzwpVKmEF5t1s+xC1ltusQCLVKJpE35tmeiJUWZTccaOzQ5P+5bCYn5gusxzh0
EoQdgKFGrbFwf+nRnCzcLgtADwnE/64BgJe2zKcOafVOpr6wcCD4qKrHFuVZmfWbzu0Q13gehyUo
flIQjDEf0FmOBjqJEegGbPavFMEc3HXG0oZn3TQkwHEphHuY1M3FkZy4i1ztF251UjTv1ZLW0ejs
JHB89t/gC+9h1prVHBesMg388gPp0l7U2J0kOx6+2JKjj8HD/jgwF+IFwQu4bmtXyNt3/dBUdbQa
RVbQHZzjgsqUJbX3X1FH30l0DkbgUfximnCWRGvIij4seGgKqXqqkfIf86OdCt6UFVD37FIpjmd+
ArRJyNqYHAWdBMAfssVi3lXwVHZGnWOeS7wCBX9iiGF1J9P2gaXk4yGAJQhEFsyDFi+Jc6IVPszC
xVUvask/n2USdaomhgE1BHoe4kNthC/s1b7PK3qQ9lenj+F19LEoqveBtG1mn4HMU+0wM+VcCFsh
8o3uLmF4qiAk05cAiNaauxA60AjD/zKWNo79zgns9nKMgzSBlhrQ0O6pI1YAqMeCeIX4pCo8K9Io
BzNy3+0XhKsr/mrHUumymwsUe0RP3quzgmSd4hVhKK64imblHAa3ypnMZzgwGnLSiIn9Dv54Wykd
SxLWuZ6HPkmRnR+tvl7yF3GSjt64RGa43a7K6IWfDjl/k7/kp6l0JZeBsq5Mr0qhYf9pL7kvxMXs
j8DpBMUVBug5akTWT78q6cwr0PezKcejx/bmxpyKzikz4sPc25yBrrYAzrdcAPa5zwa2M6gSy2nq
YcCZ6+5tB3p88/1aECB6I8h1G4XyAyAahQ9H9dhbaEfO02H5ATO8psKIA+fQZZ96PLKC/WF/Igi0
5mq1xz259JCK7N0756RCWPNw1qLQfq8T9KtowaGuqXHhirhgt7Lo1xnep5lLoXorx+cKbOpJ/2Ob
wXeIzOWlmr0UV8Zk7rD7ugxetm00TVcogwB9CARpQjXsNQssGb0UY6rhTRfP6C788RPjj0Xe+8+d
MyZXIaBhI8cYUo/ehdzHB1KB2dXqwNnbHgOFtbtMiBhKuXGEDAH5wAwWcDODqoFSkOiUcAynOjFt
qgMOD14M6RfyPUyL7Sqm4fnt7Bom4V8YQt06Wd7+caeBD7WweumjyBa564yHIEOyiSgQKkAbiS3e
NIoT4g+H00lmJC6MxWuwiyet0CmB67Mcef4cLtmmwmEqfaqOJJBpnvFfQGNaoQUb+iiCphmntwnb
IGr/KCHIyS1MO0WpPMFvnqYjbc/0M/AWvOWW0j05j52h+pgCnam3qsYTgIaYDD9lFusE3r46HJKJ
53JUzxf9DCb61p1/FolAPdYSDg1zFOxozaVZTjJOs8xl9K1OnAuzx6QWcgY5mKUM3de4kF2n2JfR
K9o1cbEzRzoB89csSZHlI4/4q8IE2l1gJCUr6BAlsOkPHFuD4XEmlEgCHLw03/sI5c2SaqNQp+WP
lqD0qJ8y8zFaVgMESdcPnL4bv9ypr+wE7wcs+DUTWKw6jlzK9cMk+nquyRR0KxxMXq6dsrhLEyVo
IRoUMFyTciVZqgD26dKViVfzJhsK38sqZjCQx899ZZ2C8A1jzX/Qm6Vh9HNlZL9S1s8xsjy0K86u
EkoHyypBs2wgRDAza3+DoeXO+mjqKj0YDybiemfhzxshHDdHmltXGRZKTG2vASHf8oBsUsC+cSd3
zLr0YKsHgtMBCHx0Oas/yhonScjdlLuJ4mBfnxPOJRYFMJHnTpgWZn/L1MrQtsX0OYc2BxXVzhMh
JV6OojfbGoQ2g/U0GsiJMAtIK1U73eMEq8Cx49JO1zhvUun1Zv0pebLmVQkJG9fTAS60ZbwF8auC
lXGxHUSnQGZJiD8n6mpsIjS2+9TPLLO1gH2ZUotkNFFICibVK5nUGioxs3Lh5zO/OsOWSiPSjgXF
j+j3Ovz1Eo6T0mZOZxxPqCx723ONwNkhgAR9T7ZCwyDRQUmqcEz68Zs0hLP48DAsIscSNm20CtLf
qQeLibm1aeNQcXJblL10K/ALSXCwrJ+VW1ZmPYDkYLq/jtQfnaMn57uacD7G0Q//QS5nQojhU3B6
ZAW07Yc0i5x31oIa7nVWCB8ExskHpqjBYBRhmw28KdZbnW3P2d1Qu56lMOUJj7RadLmw7DJkaGtM
hMfpcmMRRtT9WhCE6OFvDCNR/7Unf8kY86MwAo+VLjAFv43LC9oUEEnv4HBZYUTg/ph3Qq+jvXNH
JwR3xmuvJQJC3dmgUTejVvlh5j1je7os0n4nPyMyNaUrQq81CY942omZL7tk/s2DXRhArnBVenOe
YI13r8mOh5m33F+a5U3LckIEEpzuFx20XK3whPt1/FR5UCbcniRUihWcRcwwRWD0JAhKTNE5DdWs
QwP+ZdqrWP1AH2aA0snfTOPbODOGw9lao5zNPCGK5bjPwywaDvdxszPXXdEXB7LO1139iDrC3kcj
9vyci/rBvOlOpYpb5eetLKw4ofBKbiyIeHjzsJ5CJHISIadjt/N402ink43o6p2ZIkvS5iX2rLvN
5OzJnJWVlICjo/c5G9wY/HcTqophyswzwY0AMbQBF05Y0pPpJetfkVjkgpy/zMGiAfS9fdSREQn/
D2nmgGTLWkQZGZg8ymMRigG4H7Nr7NVVaygioUYQlkSTC+FKl4yYCNvXxZUEF1m/0j9gtE6Mwqv4
iFvYyYEowEp0+7pAnRqo/sW5Zg/Cdo/EToqBD8k7N0Cafv3VBMpUJQqgU6+L+Ewo1IRHaDilp8NF
Gz7CWuQ2mYKAx6BN2aU9M5gRwyvdPdEfr29NmK+pOtLe227MDOnPQmJKL51U7YGgFx9wYEwCvqjm
NZNdLKI9k0yz+mPSUQ0pJxP+1C6CEyXnWWSkTnsKArbvtMS11dXMYr6I8DXSXGx2CXL7/YEi4eGD
G3kaa3bVUB4pDtLL/1Ql+cNkM4KYDFRpULlq8NP6+W7eZ4yN5iNKjgz3N8OW2pH7Cv7MWkkhw4DH
xLDV4KqJpxXS0s9GVAYZHaxUuNOREWIuw7zR3crl/MwrgYP3/aj7H2enY0V4d9SiajTPgq/5TKi3
n8nw6kfV5JqTCBrLGg2yp1GggssFstyMbWL0hiaAbcg7cVZIQmdJrvGydv8RLnIvxzESxTbqhkWb
T3nSAG2bM2SeyB2xALKOWZbL6y07m01GONlQK+EH7XPJAcZu7VXjC1PpLeXeqIEipdMicABpjkI3
LpmqxvF65rN47xd5cIb4IF6DX5n7bAVP/ExSuQREDe9qKOeq5hJwPxnoRKKZzhy5IrlLVJS5X3mF
+K2GIS5KTU00pB54a7M8TCN+wnKkmw5fDHpya0VBA+X/MGc49Z8+W+rQLD9rJ4MjdiK4TT+BCxBR
vvoszJtYa4V9PyF02pMBzrpm2/YUu+VdAQ9ZVJsi2GJg+JEwOPwuJlDgiSZrVv993qK+xIcx7Qjz
W9otaIsNwOESaYfEoQ/ZhzS0YCx0rSxIq3g/89BenmaNo0ebjuJiAewCu2X+M3uF6HhJwP91xpHr
adix+y8pZjhpE2uKEJuioHoI3ra+MPP7Hh6SO+3iSqaC27pVtjbaRcfgBI659DG6Jx2+HEWHtQyU
mvOW7AOwBYGAj30YYWj0IJpyJuXs8+D4t7czoPTSvT7RffEIDu+VEQkYN9PzRRE8fp5hZuyLjS3k
m/T1hlragjiJrbTODmFZKBzZRBzSQ/z/kkpodYHdv49xWKpw9U3QT2jraKGFRTPsI2h3DQD3uVwt
O1NGK7jG7tdbEPILBFWLj7GwWSjoAvdGAZJyinFBGfsaPijzOBuqs7FvFpYJ4AuikHnSICLlYT7f
0hJNTtwah3EwF6jnAPCMOfwWcMyz+tCcDnEOigAQaVWXThkL5H5UajwScOUrlPuZa4EUjWJyDsr9
eHSmfKmGwaEnkecGkQeoq6H5LcZnK6cOoBDgPk4WS86HmHqg7vc/AuQgeyJrEUPNEGXa7k8OB7Kg
wCWqB08BFZ/k8ETRJkg/jbMYMC1un9bJCz7O1f1++Ke5KktEM17dQ17oN5MrJf+qYwOvRJm/gQ2y
g9/Hjh/ANX8F0AccL2YQNGb1oeBORpQSyOv4sLrOyV3rZNfSnWjRdh3s+w+lt7myPofsTJEyH8DS
NuOdf71J37TrNlslalhpYRR+OGaNp84advSJNRPaCbMzCU3bpAAhkQTaqKqCP77iekVIBzxgcHmt
kNEpzSrFce65hIrWIGT0VoM+Mf8RJLkpzEze7WiXhlttrfsbgol8pvRekPNfOtdSPCF02m6rFBjI
8jbP5wN2TcHqCotbxBY64Lg1303DKmmtgDDJnOoACJfd47rGdNMl/f2fqVtSHIyokgOqQHWa/ZRF
K36ATRqZOIq+0evwFXll5TJbw3wSDfPt+wqA4/LxPjTFLA4leyD2TGu+VlUX7CYu8JesAC535zWy
5JBS/ma9WqODixLaZYahUVPElX9Scf6chrxNvTsENgTLWftQ7DKImyv8hhnuON6wFRdlIM3YhHPO
+tTrYindd24F9oLfZM4LcTov9TMiQCu3YAjBcUFoVbQreI3OlY6FxMXe/x7bHUHq15NrzMsnWsPQ
kPxcLpyu8fMQDOI9pRJBqxICtjiRQ/YsLdeLFSYudxO3zosK1L+j5ASae67WM2B3B8iIBaH87noz
lmHNv7a593in/X4ShkrTtcddFskK+s2nnuwrtDwv8/ly33w75IwO/vWhjwEOIeoeZFXueYbgd686
AUwt8A8mcuLpHRLD49LcYtBN5tJHZSXqe7h/78zX7YVUDRIxsYdd3kgRyC2IitZGIjvwKIar7pd3
zPRi0amHS7dnUSny6dH9OuibNNSohxGjrcqnypKRrIkaEhPu+B1SaBWYp0AD434JDgrmfDOcuOim
56B3dmyJePMkYjl4/ZntXkVIbgwjKBR6LVBS//ZccZQ5c0D5hGezZoJOc8eJTHo+thPvTLvLzPOM
mvLEthLudngH83YPhBfpw7nxjBB82HSCImcz4NNOcg5SVq0HudaaSs0Fqe/MZNe38c0kjqCqtTGG
gRuzv9zP2CKOFTJRQ9+iFk+8UHQEVLLrslDzVdzQTEvGvs0R/ZexM/N1hyASbI07c2oM8hQDO4Je
uKH2JH+rNSVvURBvSljkpN8taLv1lRnPT4npZoSXqgGkChNlDmT9MvG/ZmFBtyrkouW+kXLNeqTm
+jT4tezcXtTH9cr9ekopooG22279e0ok4fQTCTR49v5jZbkfLjFCazsvKrvlJOOar9ruvP90XLvH
wvTnRhyhqEoA2j7GvcXe+h3vgOIc75nSNzpUg/xzMy2TZgt3FDjFXmHQa+wLspR3J4nffeAwfrk+
UKpqpRmL9Kcko7rYH+dnJE3NmRSIrl/ZX2LXGy73xS7iFRQeTq5h7g/s2IlE/UjvmCu7uHkXrm58
g77/VVDTMM3CuNoWiuZ6WRPShhU9IY1AlFzIwOCGjzjPsVcWfQQ7SPnqQ26AN1SvYf70orCD8+v4
R8qt+gzMd8bjfT/daq2ai9qCqLMwwAEi7+bZ1mjUSyTROq6E5B8PWXyPS9Oaa6bDTk4bIo/5S61/
rPMeEScoIX060TUkxgc7wJYsAf2uYQxEJQn0T2wT0aQXO9GJYH/Yy8nnQxMG0Hg0jL/zqJRqsR4s
o6Xz1TUxk0P3cEWB8QiW42KxyUOj3u2ZFwGACloMGfr930Y3TethaOsqYd9oZ/77uH0HZmYW4dfX
60pj1dgcZBednzM25R8KEhasOK+MwlljwCC+Nt+QZ2DhCNK8Q1ajwP0S8JalLm1YVMj5IIY0gdoT
zMwAzWASqGEYxRYMZGxpKZPTzbE8t3CBzRA2+4YzjnkOnu0H+pAj2+QB58GGChEseQeyZn15Qg+m
fZE6ktqK4lp/Sya5UFEgHrGROm+SnMLy9+4B+vkPkODKILzkvXLLSpBfygLrff2h/YG5xbATlGGn
NeuB2OiwBWEtXoW3x/6nHi2STqlfSSS/Y0165/ozm5k75BtLs/MM8ntHZWAJM8DMxoEIFJpDq6Yd
WF/Se9CCr9s2ZUY9YqrPyU25crUUfZhRD91i/RQqaz15f6ibnAM+9Mn2W3zW6TwHShFu+NIKt9a6
oWWaZsSkqbB6mMVxaDj3XC+NzX9FxESOUZP/qrqw7GNsREK21db1GqqXM/X22C5uAkAvsx7+4hJ7
WEOjyBjynZNTZrS/asa6/BTsD1EZHHfOsdapZiXFp1sCYMKwxMojSejBAf8TlAjzeF/G5dKKRt2d
sBNCqqZ4ICmoF4+QgbGjk8s1+zuYn80JHhKcfefAJrnz5p3hnjk4AB6D06VwxnT6ll+xvIY+HP/I
2u+//LybwB6MZaucE4LQzFRmfxcTVkj7RFpR7kCXD/y1wC/v4fT3lI5aQRrIrMPBRDbuexXASj4y
BAypaoECpHnMvat4w3P/bF7nJA4JJ4Ry/ut//XZqiy6slL86fM/C2A8soIwwQXKhuI5s9/fmdox/
TpErnr6rI9Qrot+agfVxpIq2ocqLrXvid95keKUlfUNrODHmln1AMLYeTnNKLIlKsjZcFSirGcCw
Mc1v6KhwoX7r6N44tY1s4twGOu1mxmX/qh0zLQMkYpKOrhZbaT7mpWGR3VR2hZXf9xzyRy29uqHY
qYIDtOp0sCkNk5VMPKBS3D9lyt9gIqc4kM0lSHvMFLAXGWPVXK78wuSqn9NZPEREmeMsTFytSpGa
1/HWQc0W6i8GXrQIpXlJiVtq4q/IZvLk9RUJfHvkQ7wYhiYODOb97baKti2ag0pHi7MJVGNt/KnI
orCeQv9tX4ElanHgjh8HyymOK9biIlFTqLqRKT3f6Mpn0GzdgYRrXLLXUF0NiEt65C/+Y74Jf/9a
/6qG+aVOmvxqnaSAc3ThtJFyOHDsoXaXvFo7mFhaHrDT+Q2b1eF2MCHUt7Dt2cKVa6kPAKAJZAnR
Q0n/Le/c7yIXc5ynY6KQ8e9GROnwcv1DzuAE+IXdH7PQEuQpkeLBnpioyBOpSI0wl3OeXMRXDYhg
Y5QfxqG5sH5/A27YuwxK8DaY9eNuTmLu/Z547nXegSA96uM6Ymt4MYONs4twYE4IykuwyCIwyzKJ
Y9jMke1vB/fr72LB5pipSm7nEb2unjR7jori3+bW60uhTQ1oSL3j7Zi5YBRFEIw2hPsLJeQ2JrtX
ktI8AOFFAbxxm0mP4BbLiQEyYdGEGUImM28oWleXzQ+AsUUxLIbw7u47gFlQ5mgibBJnIuoYWmch
b5xJ86llyKWJfHIEB9vp7UovrtBdteRcXTYb7mf760GsR4OBB3uiFxHYgFKQG/KqBwLBFK6gAuLy
T89yKa81H+nSMQFLrfsm29fNxhCzj62R4n/hJLHOC44wcUYqgb5wTM59N6z/mI7iYv3uE2HlGxx7
5wvNNS97sCwDQALQ6Xtwxpya5vtFXnBWgxlN8Ssh2o1ydq3PPCo93PZ88q3b4EhizPbMqZP5bduC
NyCCdm3eD6/nst02UObqbc6M4KtNQip0fYlJ/xyc3zHsL2ZYOh6J3hVaGkz+14KfbrxYyNhzPbri
W2YQQrBUaMA2PE7QTX0PULaxwurPdCqfNY6pBPxQaaP7syIq3hsbPYoW6oFxxlp5NeSqV3wIInam
YiEwvi3MnOZa/fUNYWdgNfYNOcy9ixymo9yxXmGKs5FQrktCo9B78+nxDXS6UDybktADvt3h4xqv
tn1SqAxoTP4Co/bmuxNTQXN/KEZPkVF6i8/SYkx0N6Tp3tvBmaOLjkTedk0Dp+xvFbEGe8NMvTiF
YUUQc3dOgKYKeqsMlJAdzI3PyWOOwkzj4NNaUMBsQWClT6efQK8NNM2fYxP5rN6RyGZDKX3ngGeS
VRqBFNhLOqIU1Cv8W79cLcbH79HulpLF7XrJENxHk2SxBonIv1mVBJSz97JrolsWalfv+kyYfFCp
X4M4J86xozRfKK85XjVjjcxiFYDaWIfSEbA31met6hjJGf6IZWEXOQOyd1EQhTwka/Bo/w2uaZ0P
j4pzuibF3sCPki+y6hDC3krrgJtOgfL564m2hRkoE4sq0pftQbgayv2f1IJehuS4D0g6Pr+4aUcv
1/4p4KwKGyGAuZSUsEjHcLDJwuL3mkeQozWqmyIUiHy3oJHjRXLZyr2YyCd7xKjlmxzx8xCNi4YS
IsXtDlGQrF6cXtpn+rRuj0bNbuiEScmPx2G05wonXF2GAeiHbLRKhK7K1YtuG/jDvB05ZaGUP/Lo
xzeew4PRNbaTNy4yLyXJeJIEiiMomaoxQVzRmMs8cBMPtu9O32kDNJzp6EEeb9IvM1vo2iyKsEdd
5wMu5hCPJeIRltwCYlCSq4uCmTJJZ03qxkLzBV/d+NwKYr8T1PLm7m6pXiZGewIwfPKZCtOvOBYT
Px0tDhRMhhz4aRan1diNq0N8CWeWddWO/d8XZrZT4twRWUxABSRFEFCQ5t1CAXjknSZURXI9irDF
zke+jsY696tPbEQukaNiNvaxlodTv8TofUWRST9IXy+wklj7NWLluxhf2svi1nQcaQPYBKRA2dgw
xPPEzUui49I96wJiXPYGEQJ9NRQ5S7vtl9ELLRd+aQ3Zy09r6xj1c9VST/3/5Tb0clhXkP2PPqiy
0tFaUc9LMBBO/v2KD4v0/edk2w2mvtOC1xH9LTcbbfU2hSiz13yspllGybFZH/S/eQ/9iywdawsc
W18dtRI6YR2vvqSJJ1qbcMOxOxPfs5FdQDUrkHDl2DDpBlaHdYDPrt5w8Cb9eSZYSZhg3A56ix5t
yQfhcrw9hPP7p10YnQxQfZ+5VmHuZQhVnfAkurOcEGCflkuAvZCGH+Phc2+eIfTgw4vCYeA+fWOo
26/DrQQv8F3p972BfLcO4fUCOhvvByWcGaR6XDNFXbBGKhJhmCkRsQ4aeeVo3QU7vbcI9sFXw5W3
Y+JYx5ok44We5b6ShxLyS/iFQT3boRr6ZH406al9DQFThHWek6yrRIwMHLcDC/LWHqRxiMGCa37Q
dDYXv4ocPy5e9X9tNNmj31/ZdQj/7hrn4AONjxL+LP+RhMLHMD/yczq6AsESTleOjRXgIN0gHcBK
ZbC8FYctuZMzn1F4v454jXL8896Dchha9ehm0Cnc6RZxOnpojvknRV9ZU/kxH3R/jYqaKHlp1JkE
f9hQMW1jSIigFFzkV01IXKHWPqe1EEeQ8M8/sbEVlERNHZyYyqHVN2e6wQgBsMreIUUkXl8IRqyA
uWM6ju6oZctxlxr0sZ9F2KNtu8EobSs4/70APGLPgpgBjW7VFhQWZlIAZFzJu7Wr8MaeClFgdu01
oYLkn6t7ICW25jcmkvF6F5pKQFt8ZFhHxfXRFs5n/t6UrhkY56Cd2njoMo9sQl/XyXWtKTzd/e4X
I/Ftw7MEowm428H6TBL3GIy6OGPlu2oPbT6KwThjPatdUssWs2BoKYbNl2LXiPXOjF1NFKQJ/Ybz
fZXTD6uX8aZ8cBRpWbDThWn24xxwCvrwsquG/Vcf1UczbAJkmkOWm5iFAAJ8QHvhkTNk//7IKw1A
qoAvdR0FJYAqkXEcr5L3bw8ColYU6Bfm7dO30QDywNShmFYSKYs/3I4kwmqgZQNVGjcpmVFT2s1E
4PmMhQevV+gJSOai38/c5e3suDnP8FNNqokuC8iXV4JY9x8zwhqhwAGu2YBGzRKXQrUC3k902MKu
xGaV4O7t0bkMydjzIPOFpkBrvxypEmvjI/i7ZeEnql+jkQCe4EjDfW/vWAKklXTW/7vs6Su3X1Of
LQpXtr7FNmbpWGXPS43eeSPl/zUj24n9K7rXGWgNWVmCJaCH/lD4pWC+g6Xrgesc+GFyyDz1Gbs1
ii+sa7R7y3gb7rZgNH7V+hNUVTV5AYJ5qfL3tburVBkSbWK097lEasWAI+hWtJSWxPpmo/TK3tA5
/lod50LiY2rbWa68NA5qHXCdzOVETtT7FpbY8AuecKu25OqrOWFgLYD+CLjzVupQsu+wnvYe1LgC
6Jx36Cx2fXhXy6yQVgxJow5HYa7/Ik1SEFqb4FmDQOzP2PtzbMEYHTPC8MiTggoFYRyZNBP5DyDC
3xyevCDjemmAxVTmGTCXrwCWeRWFN2Qjm+yQohMW7ban8MByypZ3QGFYJB/MEggB2XmkK6DMOEC+
76tv/PsZ0qQ+6KbEU3UIbDwCBJ2EgNfvJ2p1Om3uKDj/mNA/bsF3etNRT27VxwXisgmJJHGFqydz
NZKcKXWPI9lDUsiANOiq5f/LNcUKxkrNwhHVrozhY7SdqvsCz2XdWetHQBXA9ucKMtUeD10aa/ci
jQVUI2GX2PHqcO1aHBS0t+NKAtFU41eGsLUaDHp2qC7sl5rxNra+esozyanvod6uaqyNBO/O/C11
9fkeAUEBef+3ImkQfSfCoJ8oLFP0L0sBCAH0LMiW6xZSG8cfRNwm/bsbDLprwhuQqu9wdP78cEgt
0BsXzcXWcW79AwkDTJg+7w2OuxPDhHdnF6EfFQE94iebqU0GSbQFeL1voax5FVc409D3qApb5gEL
qXKt5iDin5fazKRCJc2ZpSYXPfcIk5UpQQG5DqkmQJ7QDRrXRpjwJzN8fMPZkob+ro+R97txHTMO
1HRToJwPoW9fv/znsbwJ5JV7/1PlBk4zO7+4m1cRoqnJLiSLDdG+Zr18/bLsMrirekD++APyGaXA
Bs6WOajpDWw9Ll76mYvZ+ugXe2CWbRZQlTq54VaJ40vXjTuEmpYjMblhL3fb9JJYBHua63Dl169D
3jh9dOS9ikcR7INYlg2hH9gEM1fRdXQes9+2rN+nA1fL3cIh8p2GpyzJHO7Acbc8CUut11qtWT62
o8mVODoHwZbbaZietlvxucu4w0l5ojrTi4DWRxiB5t9EkKYmRnybY/j6+KezI0xD1J0R0grOyazo
d0kboiT61LvSiQfSMRIeLv9BwjemxJIjNjGuDNNHASVZlfnHXtioP9ERBXXrqr+9FWZjWJU/pixI
dUra9ZmzLLmLzZAbglH77ba/8CZINfJismrDBhTe0gZdFS2ju7q3nceHpt6tUs2geqbNTeULHABJ
evaOAiHgtynt8ZrSbFExCxIBc6qVv2KDwmaxqalDxQManD67GeZOljHUvtxn+LnVhaPbN52zaLZR
f3Ax+nuEWCJ3lY9ghU8lIV7dcUltvmdUVNCAOJ1RFfz2ZL7goyd5J6T11OQBznFuK1nnRJgi3OpU
XX0As8+x8TN7ufX6pEPu5LHvILx2pqLaGN64XDEpy+xdYvFsDss4g46qgPlOVWTNavZti5AmHdbn
6TVM9dxaE3HvhuYcCYNvdhJU6bdE5GQ3dd1h6rkhELNDOJcvOUpIEfqhvJ848m3u7zmEFUsVQw3G
dVgq0Ti1spYG+ZWqRdCNpFNfnshiv9V6Wl1OzN/jsgqLK2qCmaja6TMb5y7Esc1w4+6D4mYPA56g
ZGuWAsNaUs7l1Ztuswrd0wI88w6XXqTdiqVih6yJAbD6YkU/FzOOVhHOjR4VTMky89XMW8sgnRy2
Zm7W98VP00FXOL74gjWVVpCAu8tax3DvxbqOguI4vk7pZq2XQHnKTZKsd2gEF8cvHWWr3WXSU+LG
vSplMuVwfZbfimpYZ9Tu9zj98MPXhzbWi96827CgKvZE5nuDv/s6og1Peke2R0jXwBTRrgy6pFgQ
dlCv2+D4P5RaQX0ViATDuIZfd/XTcr9QRJD+XeF8NP5eqyl1mCGlMUPiwIR8i1xfXSUaQTriF1cC
eVUUvs2jg+QRSDy27K8Ucyhf2oe5tSgNSvaCePrx0KooJ3glXxdsucgNaeTMFKHyXvKa6dUNHfZR
LPJPvYB3wOu57H4ZA52xbIrG9to1+goQT6jmC6fgWWyLYHtBxe/tCItmWBhQs6pVpoYSZfp4HmLV
9xF/exP1AxNOFjlzh3DxPVa1iC/EIfgkNdPx/wBAZSsZH+XkxCRz5FKunZO5U72k3D9xWiBJ6HeL
iwXjK/44vVIr9nAlqJcl9p6qGuH2ZaNG/XQLWMeF4rkVb6qK+hdniJtlbPP+36JLc54JW/9bGBnw
m5dcezsrXugGxrrih6P6InGK+9lHjdvZcWaqbArpYR0OENLOPyXsU9/vC/QUJISOVc2Eiv3xuCGi
vqe3w09xQf+0MW4yKGpWT7P0inBGywwhlNX2GV5GPbAhaW6OYLiCuLpMnq2ic9Q79YZkuviRDC4l
pxvSy/ZLHmV1jCx9bXbH1pGP6O+qH3UnKZnzkjx/uQMiCNkAvI57tKeNEeshdqwDUC6AyJcCBpEk
hMN7wjTIpVKj/A0EhA9I6ojlQL7WSXCP7w63p7BIBvQm4BGTo4JmO1t4UlxTuOoxplNyQNqk85uj
mjCQnQrJ97KCpxztXdlVMU7T6XwtD5m3CxlGtmcYMzXf99sEn32d7Z1wQ3APZ+Il9RBPLwo6aAGE
5dG9u6c8AM+YTX/7KDB1yt5Yh35Yier/JrOpe8FOOQFpMFZ79MuX5skeiAezhyWVmRovOH3/fiko
WAp3xI8+ccixkwNE7FnmKpCUQFZyAPWAOwu6sNv1AkVCKtm2azbIc1paqblX0C1iwefx2Ldqhxmj
0lbGpknDTnIT11Jh6vnNHw/TU1koPLCKds1LL16rv2QXy6mLMxyhYjspt6z1fkkwnOC48YeUX/GD
yXwBrOjTR0/iOzE3L+LMI3kz5cWy8buDBgQ5G/OFYgSJq8beg7OHYNyD8mivrm56EXFOJJRllsqn
tQcKYVqZbcXYewz0oCr7jMztE/9ZadHlfjiqVbjK59X0h44NvsTs9bCAAYZ0ZqCsFLGjJQ2DUmQ1
3qx+wiORVgdeyGkknRO/ykPRTVJ/Vvy4AITbZdRTNqpAjS9+N6OzJhimmmfkjZAs0t92UYUQpRo6
YEgrI/TuUKraXAcuwmjPzmRiyI+PfSIATrF2N5kr8qYiFL26OTSgC1hSfN9uH2gqTP8qSpKDWPuH
i4q7wrxGBvd28MOPsQibGM8AKp5TeHyEtAXumt8CZ3xwv373mctzTwegAJe+wwKWs0wJgc+JtH6c
hfWZ7VpSx/dr0vxXoSNZBSl13L8JiLjkqoHm4Na1o+nHqjfJm/cgqPRhMvkSrQ15h/DYHNo73Ywa
hGoLnEBhpy3M8gXjn91dfQ4DiIYEKHAYH0h+QUobPbI4uBQMtdhMXceO6u2N7YWN6oNlgr523o3k
2tTBvP3WBDpgp7urwVjoxV8FKSYh7Bsfn2KX8D9UGW/N3AkgyM8gdgIH8nY5C+qoKtgS0dFEyzmK
faJIXiDqpU7B2rlewWSWX/E+3pObeuTUWskPAIG2amC1N59hkuLFNsOYKudnpAMrqJchnjx8syG9
Wsz5iS76QzUyxb8W//V6MgQeKKRPlWRqHP3KsI4PonArXkt1tEwfHXietuZmUEN5UfqrsmnwG+XA
r7EjCCbK2qO1bJ7bQO9Y3AMCNPQl3hcKWefFj29D8+Orz34xVti1inmqRbLPLaOcH121bLF7VlHY
rrQrJgeksCAA+mZDrFasKccvnAt6qeRKYaMgIK/yxfrEEdgcvN7DZfbF3UStux1EvVrfL2S3L8ck
EPvN3e6nWjf7axCfsZ3LgqJBxE0jORtWTOq2ew0tpl99XLKUVMy9Px2G74WFb9uffg+B1kb4NYUb
8lfeQdrm93+f5zPILuQxDfrEZmIP9xQxT2KzOHkxfXL9I9tcKhJ6pPpgOUzwimb0ikK5qnhBpxk5
KST+0G2YfBp75veXmCTqzLeckm4xDR9r2gAxJ30skSRziqR/dWRGKhoM2rLYAPvZ9Ctd5VLWTYyR
gv8PPLbeU0lZrghT3CmdstBEIO87OunL4ctIXxKc4I8U6+hqpADLZYJI4BB2j2PH8JwdzAwYl/WT
93oOt+K9rb/uJQp8HdQmJuLJjBcFlQbNh0Bkr447UJ/LbU55YTqE4ZU/L+k4QSLFTsKgneMglPFg
maHGiPtFlzvgHG68G38hjVq/yEIw8PmViZoZYpb/e29LEqfjxU8i+C64RfjMUUKrtZCTCH9MecK6
d1l3AoVQGYdEi4geBGsREWNeYzk9uLErf4RaZ8WaMjNsHw8qxXd/yrNLYmeHjZ2RsqPqQchvB0eB
sQi6KEuLv3CBV8EKEBPfwQ3Df98mlRk9VAfxWyKeAQTTmFbZbdi/gmLv34xwuG7eKWtAepbqQ0DH
NNgspkttf/yeUVMqFT/R7KmpU34b8FrGz0rz9g3GgJyXtfBHWobz2Xuw1Nls5+LbPiGxqYlsMYf2
vtoPvCnS91dXe4Nvp4aVfN+jj5g4Dy6+RCog+6VZGJ4Ebpswup9ZotODWVJJcpmbatuWceqCA9rq
YVJwInKw5UmMBF5fCHHFM8EQ4hdbUtMZ87JBNjeK/uMNWMyA10hm+ssrXUgeMi7UDNXJu1zndl6o
Gibhd5D9NXDcSay5DRxDy8QQiD+cqUHzlppMtzoHROOmG+jJ1UMDszc/xpuqorIgh8CgfAVNdLO0
UT/wDuo+fgVl7NQ1jjzC7Retae7po2CMsg4OvRHf5J7P2AXV+xditM8oIXXUkpFSPLw5afKdInkE
9ja+k3YWaL5SnuWVOgrgcYp2DkiWtVX5PKXASWh2I4SuxvNfSrA97E1xZwp5yJBIYCY09bZ3pEj2
52YYk52uUb23saO2OjMQjGog5gCWeaAWxbdYWoJjqeukCSDXFXCphUuuFg4xpIHVIT+NMFAxxWkZ
7csxmBX6uHN9B+VvyeUFCobkuGhs6t3tNiAQFW+fIV4pdQuWGPagCCmMf21TMMYY6xeG+ZqqLLgw
eCaFpx8FtLyN5l0ow5AoH2BKaNCNIpn33CMr77ENwmqlvXn9HV07CqYTmdmlsgfG86Y4F4Pc4tEL
Q4nNGmvyptmAImId+kGmXZ4It1/beosvRI0cwURoi1OuVS0a445Hp74zhkKohkJDZQsR3y6LyAiK
FpNHLp5+Oe2b5yga15185jDjhcmg02RXBvmum7hQFaJeH/nOfqoLl+fj2+0Km3PfWNcFbXxdm0Hq
s3yKg5jlbQnn6/GCt5IC3a3AYHaeIT4ZU5ZYVTdvtPsBqLrMJWtOltZqRhfZEQyLReLlnz+g6Vnb
JOYrDibXF2u6ziPKRmwpNKt36sqv7u6hZhMiZgFnNUhhLr7ixGxEXKa/iRLv0VYHCeFHxe07C4dT
eWuVGvKN7adEX07yY3yDKJcMy3nWbh3aCpWzUeVUKaj9lOuWzRkSLZ6NMHDQ4Rn8X+WUgxc8Eo+T
Jg6LtnE0esTo4qfmxWO0o2VhxnvGYbSC3IghGAeE3Geetij1Qif6DYnWE9qHtHYeBOJ9miTAhUod
IaHKDqu/zdy6Dqk9gJfTVOs+M4Ar7M+v0dgEK2Cy47ng4Wjpb3FKifjiHOPPJCr/GI0/BtQfaCAi
ekgwFMpbMiVXsyXQkJzXrmqtXF9uQPRRxXCPI7uH2iIM1+LgnPQ/ezxHO6JCYJEL0sv+Jg+BXTDF
b6r8BGJzAsZDZH7Q93pdcB69FQ9pzLrVQBysxpjZWfECLbIwDibo5P3f5bCYpjatBdSqLcf7s+B3
1awvZhNEzxu+G9cTspxger9lmz9zQ0wLRM9kFmlYnWsY5cLMEYbNKz+dwgjt7fb2pZ/0OAOJHB8D
JolnFelZQyQMP9F4+/BRipIxaKmyDJvIT38+wyE0dcBtcDbHtrxs4ErbJK4HaFT5ZvoBOwB0Naie
YUgTgZQrklOz5Dg15ytk8eZUMcaWzN3NQdPrXi7diJawoEWH0uV1VJgf7GljMWSfItslHwyGkK4S
wf0MHbNgh/oiABA6g4A9z3GY6hMdRZJcyAJZ4iTKadPfxUpDZdUbtw8B++W+xHEE1IL9/8GkJk30
mE1msTMpCXAaww1OGf94ZU4niBJpzhn8hc0gqG9aPXx/1Yf9Kd+GWGN0QNVFRA2f9Z7SJz1mgk+6
POAXfyymy831lunDRhfTBT1Z3LR+Rc6FvTvqgcZ1RuPqGcTWak8t8L80mHhSfFvmclurvFKkQ1Fk
mJMNBSSdxtzDPdOzTQ6I/Y/f2l1nZG8J1rfYBx04+DV52/nEJpmohCU7oJDtcoTEmm1YE2VAYDzD
R+2edEAYx172dMCMGGMOs/K0nueQeyYm0tfi/vHHJI8m0hfmasfDQQ6XatlIslRNYaCRpH0mg/Dr
+heyccUfUVTcWwgE7tr8Q7ISQginHdiAcpYqkZHsBw5SNOX2Ss1eFM43a+L6Kjckjnn/r62XudEH
q6GSD7e2ef+Q1yMv/3wovVbdeD8r37CG1I+HSZrRjNoN4wvAtbW4kt319cR7Luyc+aPIf9WpUu6F
8WywwwonJtDqrBkUayrCVv57hFE45oZfwQwr3NottPjDI/DMXVb/wsc2nZLkMi1wvRGF9bqMh3Ry
rUjwmfe2Np8jIKYNJy+6XdNBRbyUYUc8/ztUW3f1g142tKCl0E4UxTi0dPUD128EhuX6XmZ9pIGw
pt9vKDsewnxBQk2pSiX+YAY5JsQftbEJQj+N4X06zIIY9Iif3aUxV0SMYorwkd+yLQSTRkpdcTyg
Q8XRh3oc6Csyrn7BloLLciqy4QdENDQPffY6XFPQUHo0FXp3tQ73VROEaoy/2UoP1igqBtwp6j0o
oVp7vCiT2N97AuV/Fp1srbw6fgkq2rsw33kmVArgFqHCBHkcagdmE2LKcuZ8XDaX9iTS8QkTNWrY
q7G4bwgNWEgU3g7o3MsbE9sDUC7+jXC6QlK08w1PWqFEZAJMMCeJkvfbOJtz8D8zsWinwwQK5igG
Ja1e6fHCIVMVaZ/KZZYBFqa7MLWtA8czmQqdOKkOfijKeMfk/MMrt0pAo8qe9W8nl5DdONrbXOti
jDYbT81TpTqMv8rdxFTYbiHLjWhp8THeOWGqRiTJsR6xKA92TfpX0j7V8uEv5EHfEweJTYY+WmBH
HULTJb/ZtIWEM22lro8UClb2kgOHrcbrz88rgP8dXftw0b3ksmORlRdWuqKWCt9I0pVgnVFMbqta
gEjyQo+QS+pBnuUvwVjwoKMzdGZY/+MiVMT5THfVRqpZdpMhHWsrCU45SDcyTNThHL73ExI8J9Ri
NIjVFOfV99Q0gkXFHhGoevjPrVX3zhsKkkQXJosyqgxq0YErtWcCh8SWUwtXkdT925u3b6RF6rKt
5CPgsscDEFvij+fEGxzHfy7e0w8azQJ9dmQML3Fxl8DVc8dvlKn8SkVCUz8w9uW01Opzk4VV1sql
njc0lJVSa8GlbORdHHk+MXyialHoptdFpfGjhYVvDKnOFZJyGwUgYl7cHBJ9K3aKeyQP0APM/dNC
+oBNUzQceFZZArA/3pDb3JyLf3Pb9uNoNIyZlJ5HoQP/z17qyI0DWzRVuA0r5HsMYkNYBUqWaorD
XqNSwXAiJZv42ZPEBvpc0yODHHYdoqaYnDf61FaQTMahwD9zuGgQJEko9CpeYoRf/dpCRwnUJsq/
lVMOGqzc+5fogH+bRMu+507Q9RW/GDQKYjUnK6Rpcx28L4idgg+4aX+sqXmv4PZ+fZU6D1La90UX
aIPP/lNLTg9Xk85z9bwr2x07XZ9JbdtCdAcG3ThTYKY9cdVfBI0acvQsK0QF9UQ5jZwAuiDnBt5c
GjNrTCZtM5wECdqIU4KAKjtac9v6rGp+KJ+BhZV6pTsCe7ZFMIRYk6MW/OclhObo36dhAR89IyoM
Y05aooC5iLpYHdda2yNa2yiFgq44h4a4MePqeghOHri8XJAWCVEwUq6Ki/BNWArWTE67Vs3nj7dV
ctUiZEuNhhgkATlQXzCxNbXJzeAqapufEYg9w8HP3bgW6LKzuIQSAYGeF874XrGFyqVf26zpaCfh
LDqTz7nvCb/398ryHlHpFYebZ18howrj+o8KXfGozTtvvcOAd/k3NQaNDX5LZYouGf7DSqEwJ35m
CXjwlZAZuvJVURCJjS8zHOMcMesEvVfXv1Oj/DtEur6pjS7AApCIyqjyTK4zqUXaCvowCg/EMk3x
1rzmWXklFOt1MMJe9pcudHYZFwmYzThP8iawyZf7ZPOLDQhLhG7wb3/0xWURjqfib9BpCs+HL2bQ
pxhKTBUvRXtwS0wYwecVgoMzFE/+vOHOCfJwYVIEl1RCtb3gb0c39Ka3h9Onor9WySEJkUqguZHP
uaDoMJVEQtlFYzvMGC1X/YKzDKLusc+d80Oky701mpkkbVpB+S4CtNOv9Gufm2ywTgF5Lr+9z3zG
foKRX7SzHUVsEEIQ7GcXm7aaJWgc72zOO1FEDm7LPoH96ED83rzrx3wJMkvKE4JKzPlUryqaw+cc
kP61dMW6B0PAb3Mppel4vH1tWyzZLQhRlY0FwvcjUEYy3kH0NN1DUH24c3V061eC+kp8dpeRyaiO
gdmqVb605s+HC4hYs7DkPd1dSbj+kcYHlg26bEmx7v6EOn+78xb0+iXYgy6AXg2Qmiz+yE4CbjqD
hy1huA7wrj/JG15W9OE4/aYWBGIUbESRofI2F9EyzSZ0ZqdS77zhSjrlP/YC6ylm3ljg8xwPaQVv
oT+kUl+FHoStulgxfLE4Jsqbvf7ICO0D5LLjekiclHQaua2zPRcWT2G6vpLuGJoFzintdAZCOeyG
Ja5XU7pmGY5hD1w7UQEKdvVjh7cN9KX3hX5EXetfLxQNrpy+1ck+eeF5NcADJEp2NrZasTZnzMYE
FcN3r2rWTlkpcKhQE03CoT1XqGtSkzy3gMsuxyoGAuYbwdy6ZRL95kErvZZIo49La/GQR/Sszco1
YHlJemdjUGmg8q5gfbmGQ1xWLMVLSMQRQg4X7/BgYLhR7U8Eg0/p1uSMwOOUyU3PUg8QhY6ipPas
XAE5drSkX0Oz/aygAVIfbjbFo3hxEothoWB4/ed/IzddKDCK37jtbCVIFGyDD/uJaZolFLHXdAr1
c3SK5mvFKMdgDbB9h2jBGjF2Szl9tiGffdNRPzpgYsvgGGLH17I9VIF3Cc5spdBhO9uSk3WrTAnL
KfXPf0d8dEsCaYM5Ryya1+KLJSPTjgCSeXT+j45Sfbd/7Mv8KdFx9AgKPDRGiEnVEbgJ69tHkcXd
9fAVriLWXAxBEDJT349BKs0SltW0S+VaeFmXHamOAzXNhj23s6wAFyA8gJcBViPdZVqqqQhPMAGF
YDxbTE20E8BZSr6HEIg9VzBZd4OriiiijtwvWVtjBE5hp+hA4rslTrgHlpjMUpWzCsQbsgg/pMHO
Bnp69yPFxnCupV213c7fsrKX/T+HncD9a9DvFoViobYV6WXnaUN2MNUI+K8w01Zfj74+Cut32iNy
/teFD+y4HaDtynM6wOjXCUHHMxLH3Dwpid6IZT/FQLqIaNZ/eSneEEuIGOhp0ZRzEJseQ5xU66nl
T6cx4sPbJQT/DKRBAhg4eaEaZa4BgOG1TBQBYF20EEk9Thvhb+Uq6uC/iqa7ngxFd1uubvR2GeyZ
402eIuSPaspwf5+7ctX5LC1DelAow9H6tG3Ei0V8ZtjIskubfWAEIUp0VTWQV1IzFtRcr91wFlMz
bCYZWDY7ilUHJ8+EnQgn3JPEsU2At7wJDX/DdmnbyZNIUL2uP5TjdqT5SNdoAVceVLZqF26z6hPH
2VHhCesFqBH54IpfznSjBNX873zDC80djaGDxU9gyHD0hLSBnWX3DQrV78o2moiirj06BZEg9eXw
qEdX0IVG+pzBm9AK3KysqIJkFKYV+tluv/l+iU20OZ+beQUQ4FViM/3EKixqjHWL3/er3cZlRaPq
92Q1+dRpTYWqxyIEi4hscD3wJn9Cmx0Xkw0ALN0eiaRoatHO95LPWHi6SPPHy/vxDRJAg/f3Vc8S
SAo7aXKGuJ4PjPu0t33GRfDIG1PDnWg0UTzCHNSPxAthqwlBN74AyJWdpzJmTKKe8QlCeHxqJQ6U
nZWn91Wyz074sdAgMZW6eB3deupbbGs0IDoSlt5HAhJyn9EANQ2Bi73GvJEXLX9CniNFKsGxp+so
vvj9+ZpSZMTixooOzLDF9X9GQ+D7IAQlykjMfdVKg4lud1uVLrVodxy3rwan1EDEH+4KlhHtP7NF
rve5iRTsBmfeAY0zVhcpOyTZGNSn0XHacw7sQtXbi1pYFUyaKGLXqwx5tC+Z5BzXUFYYcyRgM/b1
XZ+EmpfEGNIZMfm2u4UxWEH8AFEinX85LtB3/ikMyalzuvPZO6wu3Z/Mk+zk1+R1JJwSTq38aQyC
lwpa+FbC/Fdc44EgvJKBte73S2YNIakOM7GDGsyR5Tmum5x1/P+cGvbu4Z6ZD9euS1YvvO8HBCYC
6fE+AYrTHyOWGIMLQC13nujcYv50wITYBmZXJG0Pwd8hwmbghhDHYk9RpMmDXQHWEi7EZBzql3mb
6q/RcAZzt81rQbFfXBd5HNeK53dgpWn3INyHZdMO6WzhSmRO3YRI8AJABN2RpXUzV9xzjP9v4bWk
5u2oAIepF51T87KSg4W/ZpdRHQLfkP3Joryy7arGL+HAmE8RhI9niEV5HYa0gIoTzjEMkCXqOOwN
QOyngp6T3sThIf/oTaQhfZlN0xY6B1wPP6Mt8wGXzwEhqQqGcuQ5enm278THopilfVGPDMQN60P3
2eEcUHitm8YSqBjHjC/sRA5adyl6RNPCTvPQr4T5rYMRhElwqzkhWQ8e+JShJlr+bjd22uDnyLWG
7AOgEwys2YZMNhp+90D0buVFc+OSbL+MCr3uOCt5bvSbFvGEJRVtrixwuFyhVPrxGd9bvtjViNO8
NsM6k0pua0+CUwfdo4O5YUhSOOv1uqcjKdmPci54M4glYnvJcrJpf9qqyKBrDDUOJqTD/2Q01c1k
dmPhW+2AQqE3QHOBYYy5EAO6FgPqJusJi+HDMezkD9Sl03r+ml6aesRuBQ9MkyhLugiNS6Ba4zOW
0Z9NN0mIv2Utin9l8yXFrLG1TFRW9i6xoBmCOe+nnl0trX9QPW/yQe8k4pRuh92iFdcYwgxpXZR5
KGPuBMhLvAzFN4uyr5u+kwJkRO4fseVn+9PwC8Ndm05K3Knxw79K1f7Owlw1aFMRQq3sYLcpsJfs
2tvDDCXS4mXsZBIVY6+2OI7mDcdSwNaKNRoTRTnnoCBB7iOofh8EZuBLW2w7T/fyKD1Y5MMGTX2r
hXjFJrjVkJSSm1KCpaDxd8V/Ml7HX8OAq+AYkBpD7sQLRCijdKrljiRBCisyt8e3XF/wx1Y5boPJ
7bALco7akvDpyKunrrnFNDXbEHgqq/bovo7J51pcuWkBLv/1kV+Law3rtrHQF7NAO9f2iNFdwnEM
R2DMkVlB8BG7cL91ks23Npn2o/NDIbkBJJ1ph9JfZuiKq+cWy4sTotnty6joTxwHjNwrWeBHMhVU
2xALi6V5r/2RSakxVVZQNy2XOUmRoME5xa64I73JyXybkSNUEVMurg+OBekBR75D3VY5pj/JUu3s
ok98RLk8pWxsG5xX9V3CEHLu8JFt+n40uuWeply7m0tkSyeZMaX/o6ljdw73rd2HBXBRS2iad5Mq
oe3F3fbTeBJJsZYql4mpeADEOPz/Pb4HaRA2nvLFwx7oKodysr3lXJWmRB8NC32cydwNX/zQG/yL
E6QfBQ/9D9eLkzF5xJbBoiBsWV9/+44gLNP5nv3AaDHMA7+ayJIIEKP0oyR/tvzVCfs5x61XPA66
0Hiwo/awFjOzG9UjFqOK4e6cTRMGN93g9aWnz6i3WO3OZYS12cmjOgXZSp9LqnszD3gHcit8K2Jn
ovQT0YalI6MRFAqOD+mdvxWUYeUhyore4g0FDVRz1RUa3XFoWPOv24aeMHBn/YuZrEoK29Zpxh3h
WLOFbba5ea27SquGQHxk7I4Z3VH9dQ6Fk54h7xYT4HzT+XgO5T9qsbBfQL7XNTuJpc2fZxevU+jR
4l5ioffArE05oyHgsPcaScTcpr19rVZCQFSmHEEZoI9N4ybfcTgYklV0eognEtip75oQmIwv5nNJ
a+fwLh0oMNdbdujU5SYaaOZi5s485SddGlvCfRFk8Cho7dP4XHT7wonVjJ0o34VoZgFMRFfgo041
Cki36ZPhceA/HUk643T8+BSC0sWqV/EatRubfvhi4ooX4rAndGVw0a3N9U6fpfotAj1OscHoG3jk
o7HmGUO2qtbNE8FLJHO0q44bqZXcKeVTdFyzH/gA92QgniB311YwrrrO4VhKdDiF6W3zSEiswvm3
FSoditFd5PlfrQDXsmaOrX/GJiw1mcko0poZ6OPhLxIhMA0oYTyM1e1GLzwA3KkZ7W080pf2r2NI
5W/Qu3f6BPoZzebT2U7kbF6di8pLfZi9yFIl110/aPDh8u8kFhjZFKQ0soEv/DUIxGm3vzMvS9AF
r1IlhXzGPz9m80gydx8A2i0Q93asnvCRANlMKUzy/9jWEOlWfyjuCcc47XrEvGbRxqvmYez9HZUk
zLD7FizJUx5dqZntjpcLcZcKMqtnOzFTR1OYOtVO7FKQWlOHxSw8kwmNTHQS9AGaUtmcmPOCJ+xV
IvIpBDZCNG/Np2eZrmPKmjPbGWLObdO+4gM9uz9HT8u4t9IuEQxAggLsX0tSheM5WZ6oo4xFlw7t
UBuIJiN5e+UU7pkfDQmmyrqylvqUpmD29Iy8IYLum8bnWyH7JAQZvuBPGY2jXFRgdQkGg2/9hf9l
axb4yrTIHlUeJRSQtVFyHvuDXr5uzg0dBDbnhBCziKM2ETMUWWfUP83Bu+kjI4r5AXvR8PeIviLI
tJqaEKtcK+Zqw68V87eqx7Sw9R0A6vzXjUdpPO3t33OPsfimNgVlNIukkNBKIRZPDgp7Ga10sjkb
72/dqKdw3x2WZ6vf7NFPM6k22zMOZ5MqsCWFc/J5MxdeWBvyF9/FXrQyoNGuD/240ykMoDbWvGmV
tfs8cdhjpLr6qlzIUTbjl3A96kLdVoDFwNvJHplduG9lS70KQEUqP1p0PK9wjaut0LKdF+nnlPXy
9+QR6DWvg4GVKJ1g3/QTLeHv2R0ctXBhOJw4oTtkrP+dT6WEI8ecKs5WbB7fZd69l3ajWc43QxTy
N6Sp+w93WaUIAG6YUf4Q3lhBMzN5tX2hfAPDFnkeB9tFPh4c3ANFnAbJIE5ibr7V2HMJUPtErayW
9rL/I3dQdO/X174g+5iUDEW4YGxqyAlcE+Vyh17RB2sYOEUCGin75QhoTApygvUOvGrOeJorcmVE
ko82d73XHnGOXtgWYuQOYxSzytYt6n3HJvmzqu2udxz/jYwQiV0zkOmTrm8pgs/95pmEhJMrQ13N
ivpGfKl9kza6t/MDWK0L/82kBCoGeeyTVrpTMIcfsSesINRpOo1d8IQySYb2WT/zRb9tufkeFI/u
KY13yof0FganORNMNvpCbBci1iHdJSGra7YVMYSuhfAPn3OL/HOK9fPVS2bkN3BMRPpFJwy1Bd1H
0OjDAZnPbhOpn2/MBDBp5u/flah1dEsHNtp28N4mfH3tKniWIFjlR6M0DyY7um7wwe/UODrOQfm0
kAiO0kk6l8ugLr1H9h6Aiez+QuqL4vioFgw2yoepRspJ62blgVP3E/qiolVQ00JtHsZeKc50/AzQ
A8GC1k0s3QGjRTUW/Hgqv+Ve3Vlxwwoo3wrNIb5OlKfeqmOd7c8c6pTrq6sgKUvcCAFnQ2+opx/+
A7qvp+h56ucJXCD2kzg8aFoBT0F25NHH/EWTae7AdpcJG+f2QdEwENboATdPBsi22ZA37sr3BB10
vDMulmxwIBFU4e8u9Kucg6UOVS0yNMhPHPDuQ1L6T4WIgLgNT0TGa4WKA7prx1wIsaxQRBodP/c5
Mbqnd3OyWqvz31OYn30o7nKRisRBmD8fsiJG4C5DHEWKpQfTgw+UMlnawnT4BstL2CihCmZBxsYl
hluKT4GiT6rjSJsSaTBbqDOggG7JwyCswH31kLBu99DtqniI/5tYv+9nzbMI5KpDOcl3+x8sXC5i
TMcIRitB5t8Av/NPK3+xCbcFHfLehiZlSD6x0Iq5h+9fvW3N6GJEA0A4qjPOR6j6iZo8A15fjc+X
gqqyawj7XJQXFvAoLWufMdW+1JLfzwFrmRThGF4ye/ZEfKNoRBUKZuCZB8Tjak0hSK3VXxTRMeft
rbZge9l4ABhV+SW+wWNZod9Wn3hOD9qcGNwN50ggn+nCKCyMigi14uPxcS1tTTBwNmSQc8N7AYJ8
KLCBJ8cyRrV0yDMmpzM/IpIibmD1jMsgUrpsrQtLKwltNLoulmd/XG/t6SAr+eyNtWC/NhbQKHKb
xuxaNUecyajsXtwDWY2QZhkoSkbC6nCKoZhc8FaLuSGr75KXb7hZ5GEa754QZoK+E+Me+26t7rRF
ULRY7V4wwUA4PKWJU/f1uAAI6ayK2+u6d9ry1phCzTeFup6RhI5bOXqziAa+hYNMSTEN/qvWh35w
le3UdKQCl+gsXdtGxg2ZyUgAX7LSMBzNWsdwwVv5s3Y2c9F+76MoXWxecIRURbwY/cbOZkLiqEGn
nWitgbBAwik75tdGNUM9Re8TrDttD7ruck6z/T/7oOL+WieV4Q3aZg9iKeswWvTFMEn4Fp9zajaA
6rbayJVeI67naSADuZUsh01PDi9yP05hPZNR5aW0LRRPwu99l85VXxcz6hkVE7PuD3SCY0DUZdcE
skLbN+QBjM3jx0cJhO83A3zcJXVcrE+7wpT6TwSc+qCB5QkguyE9aB5WdNS6iXAtSozZXLbMdQgk
lTJ/7tKjZ3BEFDsU+l2lnbguYq9FNFXdTX//YeyopgM4/rPUN00HL+7BzPu6T3Xj82+QR1S5aDh4
j77BV+4nAMxXXmkOY8KBb48rrca3kKVS0TinyqhvT5UUF31EYfHCbfNZdkIYK3+iwgZVCtNqSAVy
0oQzshSqpksieyrHGde6JXz4RSTBJEf4dfkky4fNyIeu2dtJwZQhsCqoBgveeu3UP3xGi3NLQGKf
c5yiw8vWjNK52mrR2bgKKe0bXORS1eYH4euQbv1+/cF70mk1YNJEOUAWxlZOZlmtKrcTiRiwiriP
iqVR+//tH8OO4cDwFt40Ewu70EppRGmMZrqQ1PxlBTUuAGg9DDPEn4l1WAH+4FXMN9VCoWqRIqTE
yTjM50OsayQQoQ/36q7yOejx+ziZq6YfrBgpWv/wojQFTN6WFa8e2uu4R9xiJBpJM/s2NdVbvhBv
Saioj38xCa+WsCCoM5QAdpBum7b9ATxZ8AgZG+rA7V04JX7SKGYJDszlHCUoW9l+UAnPzyrRlmzb
bFe+9fyufjZNoHFe3i/mztSrSytwUDsSuOrjeJwp9J4/dYTu5cipFauDi2knTbUxUMtx1PvIZAe6
oUcNzaT6j/xQouYTm+9uWGpf3SBqfVdZ8RyuyVhDSdMQx25E43rYzq8G5XPVL/930ig8Abcufg3L
xUSB1LugdYTKIP88FmJWVFzndtQLBSN+SqW/Wporgr+wHW2S5pUO1hoYmRLh/KbPxoOWB27luNyy
iYEe8iOjHRxlbeJIYjEMh8nB1eI+O8F5/q4coZbvUVqj7bvyY7DbywDua+xVGkEnYSbBwWC18fJ8
7kAbCGNZ9fVeZQhTRdyshBMeXTbQ6rdKlzuYjn0JZYrCSLbsYFYRnsFcDAZilPtK6MeTkU5tCyyP
G1FSzQ4JciZa/5yULNIvMcFNcnI+Y7za033xc4qLvGneWezO5UOoLmt3H90AgdrW4vPjlTRsr2iE
xzgzTWFO8voP/tSkl7ImQy2BaBMepeVu6DFmlQND7DRvh25y5zVmFUPRI0pTQlVDotbWVS6y6GPE
i4Bxxp/yR7r0tLEIqKy/nV3JXwvYz33iX4IZYBpHMoy5/2NVyRfIO4VpE/ibV71ZcPABFCCJk50U
i4808P3N3Vyh6tfZ3My+pvmx6SVOD8NLuMQPYoiv7ivgLvkM6QwaiK5PrnY0/TRcdjaznng+7zZS
f1LF3iIC9o/Os42WVH+S+aaPR62CB5mJ6fQiEKDNNNPcsbVCpv8CMVuxcx+16/vxnBOjrjsU8mw1
HzMyFOZGIQRPqk8Wm/PC38/ulpUzzrakzRYitacoRMQDt5c4LhGB1gS/N9I7w01AhPlblQzeGMvi
zz4jFzTotQG4vVqelQUNuoGrFsJ4m9VS13aeyJBYEWh4HJnCsrJmcWsiJf9nhA0WW1pgo88kcicX
rcP8C/LI30FihywNfyyMYZZPS8I7ZhB+1IVrCbrVshbQj8gGVkt+Xreibww2fFLxkiAXEwhgGEpJ
aD0pwyVy07yz30dHOviclxn/TmJoM1ZOZJOBkxiuEJlI02+MWu5f/dfZLVIP2hMGfLUiLgDw8pVm
573+jnFj3j5tY8d9U53usSJIO6qk0L0SkUSiQyv2jYLlXPXXopmuPRmkBBMxPGopVQ/kFemDeMiS
ja7wSRH43RjzaBWcApI8X4PMJ8vVIG1jEu4Li8s18NHGoiDJrk9RGJmKu91L6/JOFeSWQAt0MkYm
yNTASbOZLEYKeTG5/lP/BH6L3ph87T52JT+DprYJeGFa6MPS/HEVU/NrXDD+LR1Kfg8Li9FEpOBd
I3gRztvNxE4O+TE3GDNxcFQJSwu29N8vP8mX83i3j3Yk9sCyacSAB1T8Gb37FbbBzMjNgmhnMi02
Kkf7Ly2cUoek2WDCyU57uX641AlXytq+8gX8xvNpko4qYHCfz+kSoEBKq+K/AzYb7Ell57o0rzS2
I6pVGVnpBZGPoMCm6kMCvHr0pjXifrnMHBjr7HYq4XAO+IGut+AEQPOuwIfj+H5CI3nTSrmNauOE
u9EFGI4qTv96gAQ1VvkW72tRaaNfD8AiuTpUZsNOfkcQgUaPyMCrx2CKrtVDpyGNwsYZpEel+8GT
9N1NiJACMlCg1lY5um70nChwgxVeO5SgVFaTdzGDMSlQxi/WEzjbZb7rnwvxDDCsKOA6j0V0LENu
kmgxAFkhkpNpBLCE3ohUrLOhqQK4GSP9c3GuzOq02QpKhExjsHjtTHuLk9OXqnBQPLl1dLXXIFMA
w4cwF1eZaCx2oc1GgUMY7ymeSoVdELFrRrxifo60mEHuUQopYt4lP673mdlx3W1PloHn9IE1xdBD
FpXq+kM7GGdawp5x7tEigL0bDw7DHPvo0jiZSoH5FGCXLFaonzAAV998OxR6Cy6JrWNgrQ1Uo9tg
QOl0o9DzjhLSvcvjGBhE3L3DEjjLY5D7Hn7u8Mz22v0QeBZnkkYcezHsudUGRMVlUII7dngMDMo4
MgfRByEPW+WJ3C/bU+FHLVkj73PYsktYz76rExlYLgC4nVOuhY8uSTP6L042zDymD3UcafuXuszz
Si3WjA86ZdShWL5Eu2VX5nJd48I/24ICDhwDkWtpZav3ZtrH2AnC67677KyRX5f8/Z3lfICt4LNF
eEXod0x5r03mF8HgnKVl4uxSxpsMdoNeUr8xVhKyrDVSSQiYx6TlpQzhn00FiZktc3PhDMYXAPGH
Dx6WnmEhc4Jg6mnA2FYkr2kE8Vi8VyMz8zCJoQEUKJaVNqIjeI/zaj8fmXHt4P9acBu2iEV7Veyp
diZgqmtqXLo+UZlukK/s2SXEdbwrU8yDtf37oEKZFPPQaKmJ1nP5l5EY8k0aPNT/Xv55fk30r5bO
sgsRfp8SdARZa/ovTdm/UIlL5tTk06Op3IMQGLQauVna7rn2yAXAvkcHPIAEdJQibbdEULLtld28
zGEaLpWUQDeik4y25CfUN5Roy2WRtlMqYRuvIw9EnDB6ERsQaMWBSjmC8NNvKOTqOv9g69JI55/E
uU1u6hdkUZe/r6Qzvk/37ZLAOWegPZshUKLHJTBShuNWKVxKycaP9h/tXsXft6KFbhGz06PvgTqE
UBmFvyRy9IT5OPC12u1XGsF3CmZWu9qLW2YWmvNSaHRKGmt58/8Hf1DcBJFhOBkoZ5UED/QBxmN7
TesckBhgGYKspSysuVPzqMKzYo2qrAvnCB7DtKFLpMe/dhLPeaIkAAz/v9G9LE4wZIcjrWJBhbSj
j7XYfsWKHd/GkvqQQDPC2X1IFR3hA36EQlgeDJHYMfSwertVqOynDO1++rZGyjtGQBFy1xtdGRwR
MP7DR6+0DSYQEjYZF4K3iPtI8K26E7zyBljAAO1hnm/D5SH7W6Hq9KHM6CVmif0g1gRH4Gi4Z4On
OKC2+i9in/yVgZ2Ndu6gA7QmfB64JUZdtdOeQgB2LMveCyZWTrOTtsGz63Mth2GIeYknFccKbPwn
pxDTXifExZ03hJ/0U4Xg4z2OU68fld4HsPMRr7ADcyC5VDg6GA7s0M9l8coNWGx2OlhbHJ3T1Bvb
wjWf7iaYsPQt5t9DEOOyEvv1Oe5V/3h7b8HnPbg2U5dSUnkBjgotve+JHBOhLiK3ypG5ykxwr9MY
CSDeCD0tmJ0cisSVxGNaEi1laLh4K1u+C/WuiwNehtLAzU5ZLbnd5DjxKpj8p0xWOIm7nl/5+WdY
+aGKRUrdVrAdsHhSTbipNobuEK9fVY1CAUhsXTU38YpPMOUkvoc/Fc0fMs8kkW4DnUNDVcPfleUw
vzJ1eO6ol6mA8N22UaLwbYFcvNW32hoMzf0dyDyCYdDxsLhlDYtKpfGuqy2ovgYW3O0wLQt+T4Ki
2yRG84iZdT3PBosgpZT9uM1cEDpGqK0HJungcj7qDk8xdcDlDaWLZVjE0Klv2DodqTwHcNpSP6NP
upct8m7/Xc/rjhqoM42YxV41ORegmknXcYRgxxdwpPD7Ne9dyEIBK5fdKBqay+4ABYE154xfoUjw
D5o9M1rOAvxSz0RyLlB1xK6x750SLrnVVN48zgiIqHSaCYuYe6loePfgHwRHjedhC5sWh3CRWdsE
Fin3SW32OaPutGeB2v9QDJqb6lPTuRVL3+yO5OXE7I/1O6FPt3IT3bM8U2RoXntNowSHDjWnlrWU
llLAGo+GKV3JR9sOht3lJEhqqHHPb5DGmanXy5FRtTQUZx7aEKQ+xD6K4czv3Mf1Vx+8lFdveGR3
6oYe4xAlXF6AW3xsbk8SYf3f6C9cocsbQ3P7p6AHehwp42bpJZMeb2o3XZCwYHQYZ+cpSJEQ74Sz
72LvSNzP7JWQdf+JMz1I46JJWnjr3hVk8murRhWAmarcutNVt36WtXZ5RttIuxG0Sp00ad5HykDt
EFRLl9j8ARKr4DvI14JS1O7anODcNjEdh4OSF687LLm25RkYruWugSqtOWVEvd3IJrJw/zCr+9DL
MdiAWTnPIqVXzEQZ9PTcriKhFp+IIKIjCF9mjni/0gsO/xTtHfmtnMeeW8O7hHz3609gAaSPXLMj
Tac07hUrmNplCAxu9kZI2imk8C50agbF/MwsUUBwUR2XOGMc/HCGjhNcvStP46M2YnBGgcYit0NU
sWNP38C69hhwm96mvnXH5AxoBtZBQ4hIgT4X6ZVWX+qdCm7stNfBzNedkVOCEWRRwBokaKzuHnPW
zBMwKYVxGYL0uBvQ9C1V5XXL3WymaTrq2r9Wh4YUm/DG8ilAWITpGkOCW6DD+wNa6G3TBDzxWCyR
1zTpJUd98zWYb/tIV1ibx3ZDx6vzBAe4vDIBqymF7313zv/y2mor/8NNk2/PWmUQv1uad/AEyDpN
S6PpqVfAGvlmpD6JTXOZS9k8VOdjcmjRJGi41KyGwL2w3Og9fGqAd3dHqrFyVnKS/MXZ0pC1jGsX
xhW7nANtqHHEt8hD/27MVwePCksr1iQJ0BUFBBYVUKHaKWitSe22e/XbKwvORxK8+ToVRnTQbm2H
PrEpe5iiYB8DMDiQ198FWLFbgw9YmAkNWhQQ0JpMUfJBDFZ/r4inCHaTKBtSGXK9bPKS73NG4haL
twl7SaA+lo0YZ0MOBhSRtRbs9se26HuT1QVIdWkysCygv/8o8gtj11HOHfHgyZh3fAyEcbAXjKgb
JbKTDSDC3n7wM8zgvQCqbxJ7AVSNOIi1k7Vmd0OWEsrZ/AqnK0O2jnojkptkRjaDkiEqk6q3EX51
97U39SdyjQ686iavkWHQOqVpbKCzCXmYhjKmGANbazHRn70GW0kmBaYHO4vCiXrrZzh2Dovpmj0h
AN52FfWJl7a3vF3Ll6MWAMvrHSQ5RjwOj0HldQNPE/2VzN8TOTU/r+Ex7p1sDdfoUfaspg7rJbR9
yR9BUURgIO7d7aKiJcBQu6t82ANEuqjwNPwEfYepDLfFpx3/NFJEcYdPQgZH3nFVFx+T9ssPheMM
M59FGoG8mtQeFlR/X1vw5tnjswDzYsnxhPjsj24krcXc5LvVcE5fhNuJXqEshdzsD95v4mrbVzRM
3iSdj/RqYePoLkW9oeM0yeQ7ayByFrp1MVmgfeZZp/RDfK8eDaiuj3syRjyCj5LC3lckZCtL1k+K
kH6+eNl+BEKghYtKT07msQmMa+3v8UBvyQo+7xxlBwBFuO5S4HZXkhjJtxQIg5Bn/Me2goCcHQhE
64NqTXjfZBcVwCluBkB+/MPoi1ouqXm8qUq0VzrTVpacslrkefxdA43qiA4IxCee1Ez5jSaFNau4
685J7+zwlbffqyHi9uyJnj8HVDcxL/u0cWBhGiG4mkB6CmXXvrBq5SLKQTURNrqqZsA9EZ21SK21
x8jpmsX7rgOJwRzrzw0Wny9yUbWsMgx+oUT8AFTM2dtnTZ39+EYDRVioci0vK71hQOULhYahMwxQ
vhLVLTFYy7FVaormYeEf8N3VJqvcg6Uutv1tiXZkkhINDDvy8ZZNZiVJnFUcUOUwI2hYMaIoThZt
37XVWbmw3bmAztMD4GlXqRZsMrnBup6CmvIrbjXKY0g+J+XnPRfAQwtTIChXLRWeJOx1zJGMQjix
oJgJfC0Z6Yy2D7TuTLSUW0n2GkQxosXQiPm1qLjeVeP3re5ItTM8Hg8rE1A2djN73FZwCguhZswU
rCvVWrA98UVBxQvg2ttVK3fiCdAhuzuXtCqGkh4F4F0lJF2nHYl/H1t4Q8KuwnRmXixF5YOBFEPq
V7sNjyxB7GLxd+JoNhnSIQoqA+2JkuhGtWXKhMqXg5iw5NlhgqmxOdg7WVKBWK1oAV0j6JJFtGg3
tz0GcJ4JmyYl0b+/FAivFxnlzmsqWmZGdyzROgSegIvJe42Id+eXC+Mzq4QrRAlQT5ACqYoSAbXe
0aeR7cneuLlDWPeZuVnBAiA2Ln8nYKCBGZd7NsLuUcXb/nn8cmsJ93PZ6/TqWg5MCNR/cOXfkrFC
JNtVaXom7V6fg2HmzQzXWPSL/UinaFnnbVTBAGEWgbLx/00Xp5sVo2KsLdjxGlyIbZiHRzBgL8xm
XweFAe617MpISmaTYeSeiUgMXTWQ2A6/rS84q7/kp2tAEWixDApDqS1qWyqQlxTu/96yrPNhBbaC
wjOUhPga9OKBy1g9fMWATBEnA5viuaUBFeUavXRt/FP/zth6kjAh3QePRnU8KvobrIxyQJX1sR8K
xwpMNwgzC+k0T/FzF5ktkSxSbfqMBF46NHp8y2b8b/uZ2xLage7bQP8sRAPKKchWZxSBcPxLh9kJ
eo0nL6q4xnQxXTSzbwm1hjIGr8B8MoLgFhW5cNP2mYljhgUkPLQC9wiQEGv081U77HrJoG3WR/Nf
JLjHYQ/JA/MHoyoTauoTJy6kHIf/BZYbQsgUDOatmk8m0fQoUW3K7pU8OlyA29LC7ss58JkW/Tms
pMqUx3YA5HzbkKwWrIs5Id7kmEriQOj546oV2wjdQBfvGBdDBab8wKLwaVbKmBwdrpZCenSdHr3x
9lHCfxzAAjdXXj7+Vo42vAJSc60H82jYehXrvLUm/7Lr0BsB2Q1Hz0axVRudQQ3k/zcsMp19Sl+2
lgvby6g3T0r+sgZ+GG6Z3/dbA3DKxgo5z41GCsNtav/x1fgiQ8d4d/Rj5QC1Im0yU8hrBZoZbA8W
rfacAKiculdPpOC1gIQyAm1D+mwZH689P6zqZLnQznWzcGg15aI8RlKAWnvofcGvi2oqvj4IvLGG
KW0fYyqWItXT8qj9wwox6JzLtm6Ct8MdRs5E2u/+AcgdADG9OqAA6KqWkT/htkpIg5gxr7DjoUR3
g3+z5WIygSWAZgQyR06IbyNwRLx9Ik1rJ5+tiAb7oDmKP0FC29EUQqWWQkHDRYnEbrsHgi/63l8B
tkbYSP0SPGSBeyZYz9rS0y/vJEnYC08KQARWmUylrPNs1AAa42jovMRJa14hJaioshlZSMvyxDwD
EoT71dInXw9tlT/LGsq/lxVryf97AZUnIDXPLElgPjb2ZCl9NwNTzZE32VC5xzPNukV/vemRsCWs
gwTuqp963mh6tYYF6GINrV+/ZgRSZqG+hNkCpvpb/WQr1q3tmYE2UkWknL/nMhLZQCklXHV5u+18
QW/QRmiShojQuELZkf3yPANMjLtbA1hQqMSLwxOXfdG59QyeH+PP3/BXkPcgezY3bIsy+Jky81Cm
yrQqLIuut/2z1oIthaXWh8TOQrJDMbfj2bQDZOlKMPkd+q9Q0ipT4Dzu5iDGg+2H5nt00iMtxKTP
iphwIdUk20V0HDyz0jswTsJNPnjO0QvORS7RaOKo87pGI/QbHiFH8Mb89wKcEacqyUjQh01VDj0o
2CKCXm1EsEkNxQSEed6Zh+Ki310e8NnVUBddi/bNQfyVq/FjCvNpEH6D70lzYGkIl40tZv/bPj+Y
EN5AkxpoF8w/HG0SRU2v5RlNX+jW/c1FztHnJry0uP/iPEY9ZNRDdllTrrzXf1ncJLCevB81VImY
QXPeAUW+7QcXniozXehxKx18sUV4AEOZaD+Ir1rcE1RkEE1Gna1TXiXljqpAGBhD4sdZ2tXV/2Xu
Zro1QH/dxladSqV6pkrQ/vzjuK51q8PaQt3j95kvPgIRMbH+lDAvMq9xQU3RR0LL9B/HM3SnFsO2
M/LGI7VRXvB52IayDajYwJlNBZkx+T7Bmx9RoBsb0rXAszaOYBNUg7tLdvDVA+Q7xEI9GwcUf//1
6111Qjv64XgogiN2SHewUAAhVmqv4QsZwlXl0KmhEXTAe0HBcBIkXvQjSkob5ljjmre0zk/7GQpX
LItCEGKqITlPkL2/xrH/GmPcMHiHS95QHt5cWJV7pivIGmxMq7ak6hy3tcJ7zo4ZwDUIIRTrGxK5
77e4WyWv4X8pX0dMyZJ48BOd4iZEOHVKvQY7X+H4N1PTc1Hmixyaz7WLl9XAGu4LZ9uo0FpWvWKP
D7+vQ8sCDl/UwCaVadh2J1j511c2f1BWkgDOQUW4a/pd+dX+t8JxJMEpm5N2rZl5P6qE4catrNXc
4J+lJ2msuqVVoqhm1RLAHvAFpfe4ZCdVy7qDKTECUQKU3HspW8+9aXJleFf1Uf/L/Xkrco43mDfR
hFNBfXloTSTKLRzuEhSUTiLLMkImqlf0ApKuK9lcgq08s3YnUEIipoH/XjsXyWJRD54N+5n/ae3h
Y5voXfEicSCvTBlkwCbkwYCoA3UVF800PVimi7PeyLM7Aeg4s5FmvnBaA4nkiWTFepQ2jPC3kQcL
wv9FRsec3qLzUhUNXX7hLUZYNTy6l8vFZY6K7igzGDff7Qi9DbzY5V/aayVPS16uXRIu9yY1jf2A
QTo4v4sJj99VoIAKDu8wSFr4LyZEkFDV4cMHBcgk9eu9BT5E9EGKayUjTp64gdgG3hV5Fm+5WSmy
fj+7Ggto5JmNEKDlc1fcDcJqV/cVPYCFE3a6i0cho0dIYjZZPwCXX/1Od1Js2ka2KFWJGd94Pgxc
49nG1eBcXz6qFVT0DnVMZuPaCbuIIY9xJbzwiEhDUPAsFwPIRVaGoHUyuDrcVrh0+jC0f/5c0r2e
HV3gL4QXvfjHZrD46FyqJRk8Th+dC/IwQkNgkyl8gMwzmUJ8vKSpemum6DvKdl/AkMkdcKxsDEOE
kSsJBHC2hVnhfAIAWo7bZEW6OlWF7LOrhlQR6feaB/4lrF1rcGNRvwQ8Rva6qK0tm1loj91nIMnT
s8w9Pca8Df9Jih+CC8mFZ/zq4UM+jKeSgHPUSQ03jVrSgT8UXAo/5ko/PvCEjjZkl5hbgN/miU0T
2GGfsRExh6h9paGUKxeIFRkkQvZBD7DS/U2L2oBRWYy0yLMLUrt5qXX9OdSZpJuhy30YJsqYrIfu
egbmIEHKGah4gg3KhJ4Vv7RI3SJ8X9gT4Q3FqeSO2imrc/GLp50hSVItY/0E1XZ2ZgUcFcbOmM1M
M6y5o9Qa72rkXUN0op2vP5Z4+xSedpwKwSqbzpQmp1QwhmnfeyLAowYjARjybwqdK9uySpVcKpSD
nOgyD6E6qubPytSPPc7vc2O6yg/aMzI/cmh3586yvsVkknUkRa2a5secCY+ouK9w5n7YwgdzCtFc
h3losTVWSZE7YTXOOfLyLOSo1mRKLOTTnGmknh7QP7Z0Au+V1YTaAbMrm9HBLz13hOOzzuLvNLis
G6rgY6/sDwBkRlDbthyoNRRJr/ohaK/gKl32IRco+9b3m+t9gBwQnFDKqAEHSgSKGBJmaBo7BD6V
oU1HEzIUU7ANGw3xhNIV3JOkO0aJ2kq5NH0CL5j+95BJ6bvKrMCUmGOkQMxIX5ZzphW5qIbaz+VX
dwWo5oi7nBfZgh7ZjkaNtPh6CFgeJfIsTJmf/gna8dVR0TZe65zVGAg5ZDhset8GNNVadLd6XYew
Hcvkudz04zj3gf+CnzjXFNBfnL0E0DyjfTNUeZ7SDRMC7wuxkhyVyCkHT4ZFvecggKvP8FrZUtOc
c8bHaWAZ7LdyI0yaTipHvD6PkKOi1zkR8nyn4Z98SUZ9YAgSUlOm4ijAHpeTThpzFI1j0YCLWiVj
ZQ/Ip/156PPmgt0/FSQNbCT6pkDI5ZkDYRZ/oTyVw55raDEif4ffG7CVY8XVleKzf6LGCvrEdT7G
OIjggB/O4lJgnaMemoIMcW1vJoPvsXIWq0Vz9e8bBhwyU36Sp8Ga0Yr7oKyflqfjk8kgCwXaWS8a
zF/H/CCFjEa5R3AwmQyaRwtsyq7/Ef0OVjPvXBYXsVhROfHb68o+27is5R/SznJLKDPWVhGuMQ1A
scKodCCJknkSqtjTmln2tJlaPFmU2Im+kfKOiAnyCFyUvIBoywx8Q4HzKBQjk17X1tbj2+k64k1t
VyVfB5woAdLusOZElJVNBpLZGP+g2VrGvVvewuw4kU99kw9z+CSriU6x4RLbsfJy6qdcppPDdFFK
1qKbItEwQbHFT2Zu5Awz+gSBHx64SlXoCAxP/cO651ovcPz52sSP2HF+YQRitm2HPL3mPvTa4nFQ
TEKxKEXSA2qfOJAuBFCkwF7AsIB7bY4ZgTSDPjB+8MwDMUmKeYcbEyBizKWQhVT7hrSb9szQKyGE
gQXRLAJMhpljILdXevwIIQ5XaFMf1OJgwbhNz2Jcgp8FhPOYbq5WIdhiBithXHLVEkrvSvIimEB3
1k2IKwiZtsNdAkrzaZxi0hVMRfgqcoPSYjDmoZfnVNrc+WnIgr/n0EPKMGBqW9cPS7ywvZjUNRpl
0pwFOEOJoPtYXPxrrAyiss/R8sVMmj2z5KagGwPcj71o+Op7mwf9o78oJLjJ4j2FkozeCd8PG9o6
Gysr4Zl9AfbBhY7+eq9Hnd6XcZVa3MEhDTBjIO9ymq4oeZ6otnIhdmNjKiN7JHObvGeZC7D7TnUK
0XIZwZlHql3ZMfTrC6NQ4w1U09iQHITHQhN0XpY0UCmRtWWmGNsjX6JlNPXnkZARFnWoxfK0ObmI
YzaZLzPbvpHxSa6CAdP0ygY73gjuViEoyDLI5xQG4Bc/NEMUYFHFNm43usxKPsKmYTSdiek2SByE
2IERceekdzBCLCpQP7Oox/G7GCvxWmAGSmptWdyw7wXbSZJEqgMHKnzbnSdy/K4Y7h7jG+f5LcH4
RuaeVEb0QDMTRoVQBEnHvkWC7ZFsZ7AW8CxWVQ+ig6K9gE866T9GTdpdqMUJmMdmffj6ZjbNzl9H
gsJ7uyykc8yONtFVoEDSichUkaTvV0+mnVAU3e2rZeVIRbTqysVcueIqyYBOirLhLYlv1S6Fc2uS
42TIdGZiPqB1++hOdkwhO2PiRluroI4COdoe1cq4WL6j+oytPyTcF/LCyJ9Y4YIrDkePB8Z8VfgG
jhBMnP1570kZVVVyrGe3rtD0broP+E7K7Wsdt0sJQCN+xeK0oQLf3s9Ds7Y+/JaJG6a379Ie4yjS
tdDYBBewDxOKDAyzjDgWgiYqwidCpZRjOt4OMmqKP1w0ka0FdgqHa7VG4K2OEjgsiyNd1LP3g9Zj
+jLL/iQ963lacSpk4fwMpAad4yGiWjFmyp/8seRs/FisR2nW45jIjo2GFQzmjbU/FF3H76+eyTdx
fGvhXKdkKl+BS6Xye9YkIFvOJa+6oqBimiMDIBKHpnBBD1sLjNw1cR9MMQw4FSlZmJqN/faZunjc
ebf6/m5e4sXpg9XoxfE5X7yhaCBU35wGXtJx9fXV9QVfyFD5fcPWmZaUtoR9KaoRSNDaBvQPTcsg
phZHLk6ESDGvrkoC+oxRHZjgGSVR9HJz0sbTcJyYJ0jc7DBZJYvgRKlXtH8nQMHhAS8b6frsCilx
BRIJmiS96eyh025ltzdpzy5DRjynXzqI66HukONlhvhNA4cKxYU/pQ9o6uqaFwKDds5/7pxAiZw2
y3r1LURCG1CvD8D9vVdAY8sCwYZLTcPly8CNL4gwZvyag9UuM7oTgdKT1KR4Ls11Amv2ER1sLBeX
+phcP8RSYobWWFVagL89Hk59mKOUEv0p4jtZqEcXNoj0l3tuV27E0mJqBQ8s5nSDaEMdkJXx4UeB
93O3OjjwAvONqLE+j2XAjQ3yfsCFHcnrXiXNsM2xdtZGdD0Oq0ooG1/oQLGBN7v07C0ter6UXYav
1EYYFaWSRdYxwphJM08A7NEW7VC0SOTvUdkIqM372EmmtsQrSaPjgjwpQp8fTHL7OZIFOy4nutEf
nSI9y8lQM0F/uC+a2iUZ0BMWXbkYOac+LNeay9CtIcX6H0M9otPUZ7/h8M0qT+pLyRLGe97SNGQa
0pZfWUR6sBeIB/qGxyj4xvVo+xZB//WK4Gvekl/hm2/7VrpJdDewoTctn5Jrl6xkV6GTav199A5k
6SGPHuYkbS0yZaSjD1ppQ1G7vZcCMe9yZD0nGyAqX8WfS2zUzQN7TG37zZzQWCq0qVtvcQZSqhjX
FszGkuqDpnKlepIpJcVOS60Vn0kqe6iADpluF6xJMCOvWZ8iyRmVD3ZzGACnPV0AW7a6RlNMxsLq
eCFjE2s5ptibi0vjitTml/5q1SypbuGdAALm+b8qvDFNmSQwwRE1dtyooc9W3bxpvafR+rM1sSKZ
HQOmZ8GbF1WBEZUhnKfxDjH9awuOUu/khTa1fFUdAPDdzKut560qO7eoZaUwGhhB1G0MR3fTO4qV
pJGdhfz+j7c25sLI8ZcsKTa0K+ICoZ2gpqF+D2G4H4Q8VcB7FzruT+sZRWUoD1IiORJmozycXYBh
1sL38exvgnxmqMlM4yxdKEMCABb2sw8Sdc4nW3jdtuDOds3XH7surgsQOg+buiQ2PvcKYFv+VN/m
VgpJuAcwrvvZrexTBcZfQbDEHQht6tRoO951FzDbulcPHEnZIXUMRqP27cGFnHlkGossiDq8vNF8
cCXts9NynOA+7s81MVtwvQ/YuBLy7HiH2hrvIeyHU98d6oVNjfR4u+FiXTdRYOgShvmIU4Mcqa9x
MdHIFxnmbOVefSBrSAbyiWoaRf5VWjc68xtHmSj3ZJ7KbPFSDDK7Ydl6BdRbqrq0fKQ3SHjDj2XO
4nAXEzMyJN87aRFic7UXlWgFEm3ZHWdofn69VnsTUC3fW0wFrcUtFdPUzsk/Y/htiQcEADE56d/v
O3yDjz8xzuf4OSKi+qx8RnnbMAj0ymNLinjWKrNeriC36RCjH+d++DHzUh7vrGn0RIKU3DcLVCr+
5kqLfZJLgwlACzjrVR0fatl4F7XVzdMcZgjPOfbAuhXnNJWAoqDrRP2hFO8nAaIgVLTe10pKHpOa
axME9abbT/2bPuvRsZS6cLRCI7GZk1VwhNK3JZxOTAUV7QgRtilXKmDYeMG30o+eo6jkEC2NEUKg
7vDn0vw3uP3p05ovOx/G+bqYhqwkYHkq7pQoyVzjq/SUkSVqG7Kn4vGWjpTeBLvm+AyppoldDzcB
ys3i7ps+//aDFfflZmrXa79mM079w32XkAatlGtNGDHHE8UW5JdPvXFKJnEuaX496UbjyGcGYvEP
T/uBOA2kdDxm1xOaxN5nEsJeJ5H5sac4ujcDlGLzuIoqqhUhEGlVBgiJZBpRJ3e/zRMYH1l7XHGA
PPc9hFlE9N1wOsteXvZmIx+aHRkbMSMhQZhmA1tqRkwyic4qOD1DHjLbAUjIr5ipMyeu5PHargsf
xw9oC3NwaovW4ZQIyBR8bK1WArHSVzMbyr+fouPL9ekaTxILEdLCq/zysU+BVSfeqAgx/MbcbM0h
6OSdBX4EB2Bc9CQpbcfGJr7m2GEz58NJkQlMiWnHMV14tohv3UIAunxwHfvxXdUiKlH8GPiQUjLF
YA5nt1xHtrXcFfpmZoGF/hGwnxvV7MxbsPDDWXkfsPZg5nMW3aIQFvXTL5taAiVzh/F8/197XpL3
BXV4bKBNkuOMmLXD68d7dLggvSjuNqsr3wKnGD0r6EXpAYHx9HJXRyzqD+k1hb6MNy+kegNomizE
d4ZcYvMhyntIHMkjQ0g5eiTIu2J/L3lJkpuMLNCUw2xzgwDnBCjqSBAqO1dRaBXy9OjZu3pQzSwP
HuYJEeJa9R+vezq4CyAziIgPQWiJy1JS5WT3ZY7/rktMdO+ZvQVYDHk7pPHQ6QlewvJszTCEAX5+
uxyGC301/ztWbKqkqhl6+F/6c2UHV0BZVVsNMJzoJ3c9t2z3qV2pw7hfHqRcUw7bjAkWtbNzNzSz
6t9ybuyjkHvMlIGzcZylBKw3GdIf/GR/q5HQLyZUiBXfyJ01RgJf+y+a8jf315rIQArKy6dib4vj
7fXI91siyqrmh8vObUKAwYcL9P478L+nAgYiJhyMDexeg3BsaXrcMUyeJP7pBZNOnqt/UUh8x7a2
n5gIrvOrfRk7Z2kNSz4DCqvdLsOFVxTu0qKkmGfvey7WwBcbLbDuR0ysknRvCsEIx7SzK8YZ08Bf
k8gFD6CbFWxeyu2keLWHRRPHA74xAk7OqU7HZOVhEpi27ZCqUT5/z16/N8rzUfo7iQHU3s6ePrI9
2JyYx5InF+LwhLx5kVL5M2e+LETM4FuOrBJYEToPO1PoiBU/6kuOHjJbpB0wwaMhYEyO8oC9xUbC
YxmEqoC/ND1qi11CzlKfdG/TL6nbf2rcd15ZTfMhU0A9GBo9OWyKKmG0KdGtrE26MpjRi/UMPR6V
FGu3lGz3gp77jQFgYggWeln9L5z6kA8eaCECoUQv/snMWH6tlCNmwB5+Jbb1QpEjdYEzosM03agW
H3Xr/Xr4nZi1pZNO6wHdFfR5eCHltlXTtm2ihn6h3dDai/Q2MsEnKfBJHv8ThKwv+aeEty5CkJTD
QTGWQ4XKMQUGr4nLaaOuGCwdRqg8DLA+uHQ86SDeG+djZNjKdRtyPMCu2xOcNM1WtI4fnnkSBipE
oGD36eaJUPc5DCcQKH7hl0wGDV4YprL7g20TBCF8UVoclsQ62/e3vDcYGSTycDAiLCukPp6cllbA
Z96QUkkC45aaWXKD4gLoNyxC/A/zxvkZK7fHev9nKPxMaKc0zNX/RSwaNHaYumFosJNkL+o6i5nq
nwT0iIu/jLqCcbdMO+IAIKCgwWIzUWVEPZGCmX8HbVIbbj/e4ecmHwbNx+EJJJ7CYuM9Dze2VP1j
D9bXrn/xsh1jcHzk34gmSMHUQ9zDYtgI6gEhuGM6yS3vqYw+q8biHPDMOcm5+4JjrlzUc/UdzUhb
lTuEDyYJG0G0sx9cklTQNuf/zjJZrGZcqcSCWYVeStmGO3Z8VkXLLBL3rQ+GZyMboQPfombY9U4B
sNCcx9Y95WLD6XIYOLNakJJXPLHJIte2ZcOnuJ/VsFxT7cFjhyTR9lJ2kQ5QThVYiPnlAIwdn4+a
hrGXhV2jLYnbAEWqOHpWSaBbDdtIEYdHMPUFtjzxvvSAodpNLDM/pxvrhGXNFYFXa/1kCIu9uf9Y
XPLc20PqyC+XKQTRxfG4gMP8hF2Eu0qUloH4wf1dKLQArii1QnxQeU1N4FD0cCzk/M20BfqmSeM3
seaZj1yhV8EPaEXEVJGR4ZqTz/k7AV9V4KXjb3w1rVLxzuJAvP9aAOQOU3ZWPT6AIPh+RXsA4lMO
EMEGe9Z9XsKEneRNHiinFV8q4r+Lf69mVtHR2eu7TloTEWZkzu0UCeO+MlB1TXgjbe17wPpe8E1j
Bv5eNmpYWFgPstTVaYlQz8qHMtNVPYq2HG0MGLK+A+1mRZ0wIIl/u0PguDrNCKpBisHvGKFubUI+
voZj7W9p1V2+kxeSC0mj6T1tBEw0hmn/bJ4YZ2tmmHUC+toSEJT8G6ijliJyM5hERLe/HDuSbyGs
cR0vWhwcb9wrp4fpRxtk02VsfWmIknVjntXgBx7rNF2zjuvZQi4/aE7plOtqQk+M6jqIZP5lkbUB
pyiX29J3tEQgVJSvDInKlpUYboxlOrw8ElBu/6gEc6xUeZCkgKN7Y1XC7UrCB6XkdClbFd6erBBN
l0NZOZiiud0Nl8Gy4lCyBR5p9X7UFfSw2oz4iGhRa05v7O2t2dpbI0yNgbMgkn+f0zmcmEgv33oy
HAaLHZKr4QGLEyonV4BhiOe34s8m6btCdYshvFvxuVLklfp0OtPhlfM8ZY8fOI/sDhOUd4FG2AAz
YgSkua7lB3y2AhRLqGIGQHkLSj9ibBDLAviH5GX0zYlk8hwcDNIgqSEL9iUmwBPPTz4FYzaPNiG+
Q9bhWbQ4G/DPboyANaRMSN6QHLSQqwvCYwDsc3h1TOXhmCjR3RunIjXmhr1S2vlQ7a9cMSlsOx3+
LHzRf+135goPeUGrHdfqu+zLKWExk795Rrq6baxmJhSFTNAOJ/XXPM3WEiOaKF2yAEkh8fgqUPt9
Zr4XPfXtoFurAAEYpmGunU9eGlA8r809ZGetFqCsEGxdAyz6RHAceX86weMTL3lbGCArSFFsWAz0
o0YxIzAN96XgYasEBp9F7qcUIdvO1IH6ICuIcUIBuRMGnIpGcxJL+oVmYTOsYRFu+nhETub0HBMD
qXVDeLhpyYRrOlelM6Mt783IvA3faJLQm7BRmMMnNFu5o4exS5fDxwabv23ycT/jDMNQtV7AOhv7
AfI76LuTgMvzixNqt1GVr3BfIYVwiaAmqn4mRGCFppRmwvuG99MS1zhBGaqFpK0XgdxFJznDXg9/
ZUQrFH+K4mKc3GOasJkAhks3/yLJP5oZNuyt7/hYCwt0nR3LZbfisiCleky20ws4GNnJedaTWp/j
/MPT9N7iUu903LgFyh+KKgH1BJSp3uRiNjXNZyF5QMgfeuYs8AOi9afGJY+xKUAyfxYk5rHhW+CQ
i10EMldJGrjH//3aB6jKB4OKJuRIa2WlikVAtIeHhSrHrzgfVKiyrSFwinaDSvVqD1y0w2RQR2+h
2v7V+EUh0EWosFPzirOZuXu2vlTcH423H263IXnyBunyqoIAxl8HVb/T+WGb0OzEEbxs0rz75Fa7
yyMiOEJ5NUQTLolSveykch70mUDz10fQKJS3C1206yU51SuFIud/HHI6Fm3nE3kRCXeYQ3Mhdy/v
tHXBK52R08GPvFmhP57gd2ilYs8X2HB6/NJISdhRtS2yUpLusLk77mCu7LnH7xzW5iHhSeaYVukJ
rYv9xXw8XGKG3IdirrVdgW6JJrht4bXSN1Si/BqS6JQjODBw8+DHh9EoOIdrn6BW3pvgS+rFdQ2k
lzcBoLEDshnLOBrr+649xanLxhcMR69YGV7uvbiX9UyTWZiYiuH1apRbhuNnX8tS62eIYJamHrK0
tXvPwNgMuKkgXIfgyBSEr/DbmtTOhISNKr6bk0aHcqOczotYZuDpXxK7Jnz7PaQSrimb9KrAdczd
uxIfZcXm8NlJOzeo6iae8LLb2ROBY6AFsyjIKsXf5XYafLSQHIsNaOP2qThqS4ra383N3KS3ZKNp
8BuZPuxW/zAqqJTQqjSJT4O9z9SLFDspp3HaZtvd49vIxrAfcFKv3Tn3dx3WPaRU/hqbaeVRUmB2
uYSU11dCSYpEijefVhAiPrmA/kfOfyhTE09ETN+i8b6mOfFjfEkpwi9bxTA3oOeekkV7ZK+7n+kR
xe0aS8wuQ41cd2Bov91OLGLyBpJnm4rwIh3vo/5sFiK3jfZNSEeVXLhln4A6mnQNBRCgOAktnGoI
xmOHZz8qNBd4o9UNL8Vf1StycAITK9bRfxXSo+CBSTNspcAKj58asiuA6Wb1DMY43W0F0aPgHGJx
VG/YwYDASwMqkIJWj1MJ91ek8oif16pVr0vCs57oxKwsSsSD/w3PyLzPSCDkBtDVAUK++vb24isX
W+zZGM5TIeOu2+IhgMamUUw4HE8N0TjT0TRVoMlnBzmKSJ2GldP7TYzGSfEK20KIK8C/ryyK/gKz
a/rCP160GdLItHbw1GdAiYQgs3ft7Mafvvvl60eM/RRZTKLXcakD7lyj31TTdwlTq/Eqwh0zHOLz
wOBhR4wPq5G+p36z/RWQ7jD7tqYYkmBrpFphX+xpw5v+qarzJHbg8Bwn6L82GuhYk+C0YYHvKUOq
RLtBhWQpZMy4+xibTaXt5VXYv2KUDRGxumXIlJ5bQ+wt0kW2sM3NTScRwe6DrlahfPEEcyPBN+dM
3pOrTr1NmUIiolPg7AIoWBaKOFVznWkahd3UDyUnmthu+AZyn3Qp/qRQy/L/FthK/N8Dl92zIdSH
KkI0366lLuKBLA2oDZZYTc0tHjoyrNBBwG31DhRRvvSJ4w/LevC946r8plI+2HWdZChbuZaPqfgD
uQGX5G6/dQn/kQR/L8ygflfIJBmIOphpZGl6qBimBoc2grW9dq1603IMCtJKZoYVvlWYUFDF/DFD
LU+HUk7s9GNpNv37yTj91up1ORNDdycXdkp/BXa2jOMR1KnkeIArpAVX7g3XarcZBgXJcYJqvkhD
ibU/qZ7Vspl2INYUpk1WntK924W4ymCATTxMIfP+obllcQU5LorUG1beJI3zW2sGYsir5kehy4fd
YMyCESkEG0QTfLb+aDGjtf+veIZgc7jQtNr854TN4zUmkTYI/kT0PSewRBLSIXy7SuBqUTq8mnf5
tQNxV8x4FFsLciR3PK/HBaWiFh8RtLpt66z/96SPtCVbyb0tfgdmRT46bi8k8kLxkSnmvzMqLcmM
maL9W40RkgP7qB3V8oUToYYOm4HdQd9pAfS5yBeLrLVfsR0d9wui5oVJsCZsP3AO7b2RYXcL2PJ7
WYKFSlxL5ferBzaiFHQ2J1GWV9oin2YfuBnFqXG6yelNVT+fFIsFXudJWYOl5xu4OgVJB1t0XaE8
uQ4i+RC7W8P5rjQId/Z7J8s/YV5axlXwUhhUF0NaZffqjM0Y0CKuU/JvtJQABYwFobPX1jDgoeGn
LOtBcQTuwOaTj6qfkBiyWFU9qnEsW5DPOf54BhXunjO53M6GzdEpb060IOOTAg01SzfMeQhC/9zs
T40zugKZC8FMQPhoXVeRmFQTMSxhS6BBwI2fhzAy0zTqoTGyvB5qLypACkQGmqYFeeDBuGGHKgx7
GLgGqIH4j2nnFdQFmp3cTxqC/bHa/ZrKncUDexYMzaeh5TT9Bz/hwY8iQVxVnamOL3Uxm0cAjIYt
I5wFBWz4Aw1+8jhwCzTMBYvYV8aoGbC6bvwA3xOekklV/QO6FcZUkRpAsTDWEOhvu0MCL7/IjBQa
yeepcOCLBEAehqaTl/GcroNmhFFK1viaKZPqOAIwA4VP3iFm5deQCA+6ggHdDkjOM7uhXoChJizZ
ndLpGugjzORZfFxigYp/+Vad2Gr7fPEloJwPnQnXGSXDp1dxkJGSI9DnOan2tFv4Uuj0mHk0Jgzh
IWPtp1hkdKNJ0r4X/x8ZaGhWruQTdjI/5RRyWvoE3RmqMUmgYMDYwAQFKFGeBqS0TVM0dAwjfsIn
/V37hkudBS2e6nWRZN5Bku5K3VDMTSuMVkREHuQC6yNBU96k42w96btp4dSSir+6P4IGwdh7GiH3
7TalsHgyxKN2Wso0pHe17QmznoBmJpuyLjyxtXMrT/Quh74QCH8DAB2xG6fEtv7TN0p88E8HPKpR
lfVgdYW9SWBY05wWZx4UGc6EuNGAY/XGxEQbE53wrF/NYgaNoQ7U64STWb7/kUH4b40jukUFfWiO
cPqrXdxiAX59NhmSO6KNJ70n8BooUXH7cUaRiV3JHX6w4a3HwI3EmNvepE8wEnHJgN6QM9C5r6cU
q9r1YBZJToZrwQ605OxcaEsyEZCAAIfzuvlV9uPlC0MnylalgT1lEoLhFr++earhN8wfmC5Lv8Ea
SKBpIYsQBTwGI4bIBeIvm7a3p+oR8WRBsmvQ7qfhJL4z/8ouPRsWAhirw94KDXHurdw7ZFoQNQfA
KECPqLoQiaqaHaVD02MgPdT6HIVjoeFhPHqRg1PsRlFQAS4RGw1Y95+bS5v2clyUcwiQD5ozTxIC
fIP+tlxmJkY0UXw2fT0RX01D6WKU1ANv/LviQO2kn9ATHKX3W/COO8gV9oztScqzIC76YUVcCLHQ
BlY8iOK+0hI3zY50/akr89t+U8utvAMH5QkwGLBEV4jPHQCYGy1d+dflcpF9Wi9HZRrEiP1nHvbG
ArZcCEi3R3ozNnV837fFFWV4QY5Q7cv3Gtz/3nnBK87kFc/mjd0pOba3lg2TyxvQjczrZn+aq2JN
URGO9IpCp9bohk4B5wfqfRTYTcb/8Jrk2odggnLqZtu4pvj6A5VfijPA/tQaDpkIw6jR+JC99fdb
gDfTabEvS/9Nm/atSaAlNfrTUflAicCe4ziqnpn+MdBGlTF0g8oC3kqLt4No9Xu7FCRTkN+KIO/H
aDR8nKy0YZuGztX+3nnYkfOHOabjJSIOTFQepfbF5z7F/6mAQ+Ly083Y30KjvG0ycmDYmOfsMLeq
j+G1cGs+gD4xgMRKQZYqim1bz5DUMHGzTfj97o+uPeUI8W9g1akaXKWRD2pQNS2T8o8IwTi40ZzD
rHRgpoARU6LID6xhUUS+t1hFz62nw461WA+lkhl+HDulJRHJz9r/RBqidzCEp9phljVmUkRYyjer
yvJC2BZ//BNVHG68zJYQBX2gGxqE9VPAH0RYaKKaSh0S9SWQpwdbGAErQ+46W1YqEE2MTbdsU+Ru
KR5o4T9tPd3tcBDtJxsJL/dxUyICzF+gLU2qqOlYHjgQKNPcBKC3xlhniDnIh9V4A6NNLcKxYm7j
lGm8GLy/oo0gKFufIfjG23ULnkx39jdnRS4k1vMzBagnTD1ASybQjcQm15ZoEqIwOC3n3MARQupS
IanuXioIU22tU0Srrb0KOAEApl0meFigj9tQZNLrfEXBtYFE+beRo/UqwgU2pdYn1FjUsS5V/87A
wvnEwoCuxO9d/Nu3gxhupYkl46vPfvs/P7q24BBzPZg1UlQNgMQ9QNcTR7iprIdZu8a76KrrosOK
6NLfB5TSqN4D/Vi8TfOz3vi7ZlGsSactthX0JZxzrZE6WyIbb3QXlKhmmLKRyIS9HN32UhX/aQSa
WgY0yaneQZCW3CoAk2h+Oj4RYpJU7GXkTFpvZmPMn7exPkeUu6BE7ICgAJ92nKssSFEq9reItb9L
2XCClmlncCoMl14TAclYakix2qFp2sSlzxgBIomJkMRWoAnRHm1CGRYq+clSEOmBO1ANneITUjve
6qTf5Pqv8Y5totpgFO2H2ZF/kCmkcNqYuq/CL0BY0jnaTi0uQRJqmrphBi5OVEy9gvCqftbe2rXK
q/ppbyChhFS4WuHSl+NeTNdAFZSm0nBCWnXUboEj22BSbjOOQWCefjPOqIqGY8qKfzZOf776u4EY
463Drxmc3YSV2TieWPgOTaeztilmL7iBJYhH8qMFCo3yuii9YsYyGX0lFVBa61autPYGAJq6Qe35
lUA3CqHkaE1WVIXDm9EbIjFpR0BGB/MM4HkUkxy4d6y65lbZtW0hDO7cMU06EySFzuT/uXkCN+Zo
LwCFP5sI9gGMsd/yfVZyuohiKpsqyhNNVYGUWFO8/RERb5vkioIDCbfaKDqS7TPjedqBYofTK/eR
vyynNdBlSU+PDyIN8rFEAdViBcGY1oJ+Al2GT4Y6WzA3eRy2vrrP+YvmZ6jJlT3nZ552lPXAGq2b
sFNOpjosMLka0yYtIIi2J+JCxih+0X/Oz4hPXts3YNPUyjYbTQ1ogWu3bR/O6BpSn7nmI3+L2Gkk
cbr4O+Gld3dOYyWRjRc2Qfe40/D7BgI8dUSJBjIpqtIlYEVpky3mk/C/tzyAaHWK/BCiVG1LSH8q
j4dwubL2EaHfm3NQUIfPhmAnjQ6p6TRplgnBWZQnOklE+Wmnxuu13k9tV8TV/52MTCsn79lJg7XX
Ud318n/TGgRMzdqsh+m55tf+l6mltiW7JZ/4CaVPcccT2ODpKT+WZZuSqfz5BpzwJ5F7cjidIMAK
wtQDZp7YJ/DWSC7H9HvLGEA5nIpdOctYOcx65rlmk3HJqEHRsHahPvp3ii3eFHYiCkJT/q5nOgDr
tSVACLqzrsMUTC6SgMfsG+qeMDEr2AGPBwFIavrzr6lIQZnUN2oN30x5MTceKVSqp8Zi1cI1g3Xp
gsBbn7MKzxEtQaQSIMF4USBEaqPO/LMnX98YXym0RvR0AHW9m+fUe87yFZouuBIwQXCBzwRizdp/
3GE+R2cmxHlD8LMGvAMrChSdOYPMbeSjpA60Tru7sxzbWYlYFfIXl3aDiN1H6yo2zp5/dsMgZxYY
V8PInvMRxTxEGDgcU5wtH2bF7H5R95NEgZ24XIRs1WBseVBXyvJOV0hsWXF10JpAq34JrvvkNF7R
Aa4q09DLJ9/nzBRb5a8bYItI4MHMgmnf4u2kSy+hHnkbelXmA2KOmCZcGdezrxsMVQoGwt8VFepM
HHfcSjuGZK4Oeg86QrY9IDISO/dJ/jQGw5M9qVLW2oIuhrbx/GDnuyFCWnrwfKOSxVXCOZmESL/K
XzvX+A82Rsn4SV+9j47ocGMsZSBwMlXVR8UCtJZTTU1b51t4psaaX8nH/AtlyzpfC6hKDOE3Bjrx
xGToYT+0Ldha6h4106IaDTawHAwmbH8wRwGnNQ4NEJY0dHkG5NdgV3pJpMdb3H3A0jSBV2+dCd6x
h9s5JeraiRUeSPRQarMZG/00aVkcOqJRNQoaIkXP6Ez2N0jFCmWpC+N2RgM/BQ9K2FyrriwJU1QQ
i37yT6wUfDms3GEekRphcR3q+sGk8MRmxHLbFxUOxMOaiPbU8VtjB0KEt0sCLFuPp9HFZGYKeuhg
tGYd3XfioKlO+7W92LPbz27ZQdJ3Met8W7VgeOS4PyKXQh/HSSSV/Q1766YUdEbdq4yYyg0S1aAx
er7a+d4W7HJ0LsRh3UOTpEnLkVSIAyEcwctaC77OKD3oFUSYuR0q/8+TvnsX+zY1U4Eu8RCuShov
breH26H5d3gcIuSqrCqdiF6s6gCoNUcdeVYSWQIhtzdpEmB5BsYi8EMgUvc7W+lp/Jf1i/9aeld6
aBsmowYamjvexdn8lpu6K548PpsM8ACvhV1rmGK6m/LGX9MoMZbzqAkwGRdZnVOOsEApiNRfw/fa
B+sC2gDmDX9Bptp8wh5AEOUIzKuWAQl7knPyztnoAUoEh1daHeKCABk6fb1NNVEmxnNbkxr53qDA
hw4SWTZ+MqnxOPlJTHOLV007SidCeCmpUa+vx3JEZyXi4/f2oaYqT/GpP31Qp4eXNff+//Uzy3Kw
Jd4e2ETQMglLOvy99yCtqbIttEH2MPprbV+JhfOWYVIymuQz+Lh9UHaGr1j3PWf6qOKTwLuKd0el
V827RPxKOtpfiS8j9pGELxs88WbGgB4Y3/QH84JXoWLGiy7sKBrp568ageCr69wyZ+JUMrVPF++A
LzfCJrf9J29PWJiulHJ5XqZCRha5r4LqpkEp1AC7hHtlltTaPZ1DhCjpD6n9C/DEq7JINzwxeTfN
0Zfm5As+PnL4If1FFZ4rmuKcfTkyr9QHNbIPZ01xHJ2eRz+KoUKNGNxMYxWx7gYUfMcJaV6sQTZa
XU6EfQvN3qfA5HNdfPWpCkr9TFD6jGV6/yoL9iqP7aMlPpWYYyA4R6QW8utVszHVhd2FYoGra+u7
yA5o0AHj1YFQbvpkJ4L3DmHQUa/iJ07oz5V9dFaie/VwTBesoDV7sQz8DlZ8rmpmQ8V4In3c7HHi
HG8MvXBC1+v4Rq2vBJfhM8o0UW3tRiYk1dg931aBrXJpov/RBVz+oVsC0XU9ftfCupeW+xcyFL0v
eah68u2xwVNmcgxXigHOPy7Orv51RYURARCgSm1D9G5wXY6nYHhSIqdJPDeC93aFSNEv/atHcyB9
zCLOK/+9fRw7Sv2/Hz4Mw8ynUX14DwHl+uTwcsYi2neVzq9AhoojUB+IGPui8d7A74vTXzJkf69a
BJbOgUzrs3WuDlc8rCYyfFrFLchjJB7HsGEyNgqF8/zqmE6z6YBb9vn5yix0a/TgfMXQ6x5rOVSZ
y0Popf+KCgAhfVWsJss0ENQD2yJMjXGDUypMO3UK3yccnXs3o79i650CYrL1LrPUDu+eB14Fd8WH
jZ+zAWtSHJbtTu7F8g6jqnKZaOC0JEPRMasgm7hOSUvGy/SNp5BEcXuTxcHFGRMV0u2xHOrsKob+
vzdlpV3vYjT/1Eh2xxj7DjSsg5Y64nSygKMkk/hhWd44EWB1sAKMgqiVeysylFKAQEsea+1LbKnd
IsZMIFpM6VpRYLUpS0RB4BX+yYJg2sefIaum3cdEqlE2Uh0kV9VpFOaXRIpnP777MRql0QAr+Uj9
K2U2eScvwfKd5j/ORGz4zeoBG2EDI4ojRSI02WRSVJxVuHs/fUv/ZTWlKLtvUpZgAptwEIGPri9f
vCqvRVXi1zYRCoa7FtWR87eWId5NhxZB6VuRqEsxbU7H3Hr07rY5rzEBzfhzNg1/aBhr+8ex0a0d
qu6WXP2ezywUB7eTrFpDk3lpOa3LrSuXYxgHERYjSdrUJdg1sGLNBe0Fys5sIgGZya7WYyuv86Th
vfkrcrtm2rWcwTCyiErNpxSBL/M4ld8AKirR1XfTUu3QwUlR0gkiRG55mJi2LmJ0WvfJiodKzD4l
WQteBSiRiLu5O9nq6BYO93dG4cdz81C0GYpI8eTfg4i4ik3IcKJSNpaoXKEzTOuDAO9cBnsZ1dry
01ZM0RV1Vk5Eq+j+SRV71vcU/zdLeZR5Z9QvPJ86u0Uj/3pATsS3U7uNfCCi/iiwUfwxVRwDEut2
9cweU+oRHRDUp/r8xhejzGf/KckHUVjkToqmqb7Z227I0tUYhTWj2lGrV3SbDEa/D+6/k4oGYzG5
7A6djgNIdeu1BpDpYqCDoV5L5xs1A5N+4/mFxzWeiZKgrUdHzUzRCfVeO2lBkNLrndh/upqjIEIv
su65b0XYTZcmvzBAjEw7GkbDGRryAaJkLZxoJ1RJg07j91hmzaAdpvv5nhFYZxXUiDF+r6EFfSq9
NI21fljuPOvaesXbmZFWIdVigs61+dymZ6uDFOLbBgmd+LdI7MJizBle7RecjXHQukWBxNdrzQfQ
wa/IsxZJNeW/RPiW/QAjIeimH9pJvZrgm9h9EtOQU6XOgOUVKOr26/so6BX9sHnBCmNx/jWyxmjN
xy1PI8bswzbln66YaaZ3VgaECU6g3RZKJrblYCS3PxpSgFdP9uKPu1msWe3O5cQgnT/0gr6jyHi3
5x1ve4+FtOYPBxZ0oVfWq51R1G/zZZKu7UqzLGYT5TEtdUYY0nEEDTlmpx4mlXz1vFFmvpHjrr9V
+kWEiEakYfu6y2Lil2i6OJC9VpMynw5MJzURW9C08nAi8rCC0NWCRwTguFrVF3E5jIK6zseYukPR
5vMkqiV25bc61UCDBMeAzfmD3UmPm4zeG9YcOFsaVhQXS5UMjgpKHsblsmQJqP4RCuObFEsb2ngT
xKTPfsqe6PrzmlIa9OOsxntAY9ZK8d9kPZXH+gqlW+A58ZTAL+gIwEkc8Y6TOw1zMGVrGStaVRUJ
NDZUe1mnYPZ1D/feCYn1GNumBH4U8EJ94W5h4qeGzRNHqDMWyEfnG5qfL3F74rkyhnDgz4/QDk1Q
HwyOgFsyuLH9JBTNivc2ynCA63mUg6j546jz13vuFR5MhMssHY4eSC2GIeV1xy+F39uGMbBV73eB
kt282whs6wxCICvVMI4zwVC2bVrd4xq/bTQKdsKnFy/+dkiM2ZNKxfMuvv9eJt+xQIhRiD6B8v45
YXn0XX2DxEB71MKThhFfxBaRseMpFJIiUk7CkZLoehXF0+Ru81IewbEBjmOoKPQXrJmS+0bQ6DJ2
4SADaRohEoVjeSMb3y6BIN5yL1m9n2IKRmM2JHNkQoCoqlrpRhXvLOlwFT9pNf4Rr9Q92t79Hexc
fgfb6yyok3+4rrbPvrFrKH3J2vX7TUNTimB3BmY584DbDVWrSfuOMJ5k5M52vK0c9SGmDddg14Ca
9cOZYNcTyLP+5HYdkkqZwJPDEzhe/G2mLkEOARJgL088zs+bEwAgPSu7wy+uGPmEUKKAR/cGAW9n
ASHbQanLffa2R1rqwJjgT2JB9pVTUgU/BSlWtcUr/6uF4i4sOCZ+vFCZmdt/2WtztnmFbc2tinee
HXVKzEwrmJKxrVeY1qmtzH1RRNrf2nOVq1VTJ7QhGO3Rtskbx/45P5lVtih4QduuOcvfCTnqLbwa
kHciQ88qsOyGfUkDrnZwTf63Npc3QrIKX8GZAFksAQTVD5csxw07uiSQkeLVWVelkaX2C6psGp7Q
54szp/s05cKfi5EqKcz5i2UBG1rJToZsyXWj9pGd1TQPa0Trj7hmt6J1xMKhayqphs7PfzW0Eh/x
B39JiEFLgrYlo2Yet8z7aLLTQvPIzPDuBNk20PYG9Vgj/nn4U7JC3JzzlYWgkBHR8o5rg2T7bDRZ
lR5acyA3lH7ikHmWrnGZ76XpsVs2xQC/QiuveI7IOy5wN+Oq/U6UwES3pgZQchq9ObwWk5+7SqgY
7o6QMCWv29fFmQsb9UyxyHGXn2DtKZljCbFeWTHQiZWtww+ADar54SoN5w6ZCQFflnVuCMWGVuJo
b//NEfGTIDfT2mv7n01xwCeNqfsh96qU627imeaCPvkB50x8ncG0Y2LbpLt1U95l1swmcTG6vPNp
2y3siePAetnTIxrzH7UK+KuBekXr1X/ldN4VqktZlODV4rJh5oY/kzexCPhmGVUZj+lRecOFip/o
P9ISOG97Wc6dnL+KZCkPrrrwRpXPMmCvEXBIJ2H1bwVMJWIGbjXAKHZhhrtvjFL35XWdlSdqS18+
HqIO46FqejWmplPu7W2pOu46FjvnrN7EbYLzgMbmKttBLV1p5iJEhnWpqPBnR4RXx9DU/M8jjTDV
DZmT2BP89byPCHZVfI709rmemP33z00QZksou76o5HlrhM/oUtmZwGnG5JmTDjFkMHfkTnK0yGRZ
hIRhf8EBPYIkkDACBQEXyH6tVY1PwzgHkofpVo8791CuOFN6BdyvKQmDIj/AdaLvAXurBfN/rMDc
jIjXWuRUI62HdgZI/M9R81DYG5HwUdBuCIOYRc+odkYOyZiS4fUA6RMhOmq8bog0b7ezhhfqC9aY
S7xo/rjUmukUwACAp5hb34/O6cQ6+W/I3buf5WPBJmdexJVCWUP3/MnZf78YqWZpSJRIintOrRbz
l6gU1PtEzpcIdH6epWQiw6Ww5YPCzmD8RwBjojJBKIwVUIrqdxz6WJrWs4t28I1yVo2MQRMRLd4o
gh8y0/8xl3/rx1SYHSwE36bk1RZ4jE+GW+E2HtytxHCyGg8x5UHJVE7HbVbbSVOGQUqceczJFIuw
MUtfTu/+3M6+pV2+OZD0vl/p7oczOr+ed8FqH7MsyxvPKwdhv4tbue+q9Lc1lqfrDVeho4gW1Yor
YUs3TyYTfIy35sKHcuUW4bFIA0QTCKqllDLy0IRaYMwGo8LiGJMF7YFvOQRl7e466cZR2hNVCS7h
rmeut53tA41rqWidsp6klo3UNDSrfwopF6S8ad8de/lBhALKux/n6hlBmSV6YOP0sYzIc3nPq6Sw
pokCmqsIEI0HfzNldtwYbzKZRKrzzH+K3CcxG4Nrlw+yjF9H8Qe83khYcHEzUQVtKkBb90SLk5To
OLEnkV2TZNt1B6MLYjwnPD2Zhw/Gd3XFBXWk0NT3wVwUxyzj2ab42hyn8g27bLmmjdB7kpKjU3be
vLrnCmoW4ohUw6d2MrK4/uJ0iM6Fbt3htRiypaPwdvhOtwyxyZtpajfxrVwiYPAIN/s+DQyLXn7g
oU1qYLRfd+HmRCSHf82e2r0o1jmBi+oN1xGqd2MvanlntD7DETO9qrYodk0LwTOGocMfzxCNwfUp
VOPntgmFkQIxgGViA0DyJWPIJSEW6fwgIboTf0SZd3Ti0+6Biulj2IGccGwQHrZRJRwobDqSPw9z
pV8TIE9RnHfMxfni6/vXcG1Yn19HDVWKWmrXtGx3ryW5BQSaD3BLGKDCKCKnwiPXeM1p1zyY/CDg
BNxN0emJQ3pdDaqeGBkDhdmt2nlMHDiFWPAJL2ljHkgeFV+YgngLKNuyLSyNxQ610JFErDUqZPqJ
NY7HNqXyjbxZgRQnH2by1zoyoPRXMSfTXiHU9FQVh/JLrJCCGHBuglfv65YS/QK79AYLGM6SIhpO
1TxznOZNaXJk/mDh/awRsNwWpOYvHgR/T7qeJoQOHMm1qYUZg4ZyPTQ7NUNrQmlXBxI7EFxoDzQq
BheQqj/254U/Ffr/IXjdmV9n+myd+FDYNCta21DRvscKMYJHreZOHfJuwYoKmwOsZ72bIqoG0q39
cWiN0E4Z84iTmis7Qd27kLaLf2Zu4dyRL/PopxV6rU5OD9aO9eCW9PGh9FHf/p36X6o3Syf/8K4m
xa/4C+PM3hPBAq9ufDK7PIP5FFb93unp7iUkVYg9RywypkmZELKxLZPVISBe4cTGXHZ297B9nHPS
s43OQnWzi1x+BBdV0/hg5ApEw11OX+XZla27olXPUA6WsYIC1CyhfhbKdJZ7pJjWhRU+qN+zgGPU
jYupdHpTFehHqpDQzuUJ1XkhcC3iFV1edlkarEHx5kp1BAuhHbig7ZQJJ7a/nD1f/Swnv+nbIjbP
cehrbkRmtc6/2TWi2UGLJuuV8FNsjuzPyWpXp3Fwjk6Dx1aEV0JT8a/6Zcm82lB9O0qycDoBeydl
DT6xip9b3/Bz4GqHACWRofRlXHYB5+pdrlzBMoTLR2tN/RJFtcDMR+8HwW/2m1aULHWd7k3rXBsz
KV6Tu2lIePSCbSRW72bQrgLXZSeiLifkTRf02w1WpsDaKMo0fBWEMMMfFV1k6EhUAwRw9XLuapSs
IR+QN8llqX71HGzNNJu3X261O37WptIL/8lJfbYw8cQPSNWdSrXQBstsTW6ye4o4Pks86Sqxe1co
0quri+wXj7vZVORErIb9AJUq3MyMjENVuy29ysQ0TBFsEqFkdjyh7arG4lJN1G6e9P8X9ifq9/Qq
WVt+wq9s5DpqqiuECxJB7r2e224WdENigeSvjk7NV7VADS2nIBS1A2u6x26qwCKZtCPdI1TPsLax
GeYHnc/KemdXMl3dPrwJXNC96XGz+fwG//SJmF+/T7ijHnHZyLEN+24pjvXyDRWqH9jRzmTxLqZf
uEiBfLZhMD00RAbWgjZxJpbQ1I0q0fX+KBpGRkRnpkdGTiemEnwQ8HLkL84nlXnCHcCEdWlIs8vZ
Xt83bsvm9zUcbwEKBq0evWcr9+x2XX8946crqTZ1ysjS1xiaHeg1qa2E+aQb3AcJHmQKAUYWJVf5
sTja/Z+/n4yHUwg151mMEfB91yTu0PhwsenURCcKJk8QP1uH+kZ3aQLkuc+s994D6K6H9bo+7OX2
JqcT6PcgMfaYC1EzGajTZ3cAfkQwRscQMFFO17Y3p/4Tlp4gGR1F9Cf7A0wer1aXHs4VNAQlrh3V
ss8GiDpJuQYOILrOOlptBH3ZI/9VlDHFnnLChjvYCrFTKAsZc2qxuihUISMkGBGgwZytmKcJzVmM
Bn3pl/E/yD8XpuFZ5g0K99kKNjdE5msO32x7EhjqST21+bTMK6oEGmziVHksGomOLoqa7tXvqoo/
YoRS/Kg7KOENOoYIZPkb0oNp0YBTZAzmHepESWwLUQDvZuAIwUxJuNYscf/GtY499RpKQH5EtLAr
Xg+GsS1K1VpOIlrNKHf1ZRNzFOIlW9oK6WDcECnu1FcozYVTjOEYPqe9n1E8kYoS44uU8yL/J1Rg
fJ8+TrODfSqEzrbshfYBoNkt2WqsDbXYO4aInZeYagQmsEh9H7CEYcidR4no2n7H4OlSiKve7dCR
JB2HeoYnWEuwX7E8aCtpj8ug77z2JH7WbjTnFGnOJjjC6CGsEJioYD8FW+7wUveikb/bM9LaMdP5
R3iJRAMO59pkiCjFXEYgIEDDIfXMKBihDdKcBhMT8UIasCfIZCq5bCHbgXBvtfzegZS7cW/xHLmE
KDl0YChqVZmiAgOWrBBBWEHw1Hax1HrncXQLp0ROnTQJj0Cf1G/ABqIhywIFTNW6ELNqQY+l3dtt
7WHp+acZEOYW0UlyfpiEhq506n3ps+UWafKmMa5stBKRo2NvKtUveZ7ACMQ19TTY9bpk1H39GTQN
Tix9cp/M83SrU0NP1n4jdnyY3Zw61Ex5jMe3H7vmyFn7N0CRLXHfUGSgNlHblzllGaTcykmXeHs8
s7+C9qvmOvnbgIv2bDvrSTPHdhAwO6g1DBOyM2HWAAIya/+nBXQcK5oS5EVmrpbQY6guxJLSDEeu
YohiYe3QB6i4b8pWMVBR6ViQv6CYJtT3eZ3ZZQhvPgHS7trGRSO0M9lOqOLxJbeK7mznvBTJ30pz
GOmu6TphKOKgWJXBcAjYcB97sxX3G2cxCIkMo1DyLho8uadkbovqsVnX+WqTsFLyCvj4AnjOtK2G
TaCKMml3NGmUBluNqAxKYgiaG6JwKW+c2zj+rdmc4AdHUuDT4xpfx4C763zXz44JodQ0u2+sMchM
LdqbhjIW3p4DxYIHOLI7PEvtCzx2a+QS1nqpeEBqGLr4RLjZ8Fn43YPeAaEka8zHut0bA1pD6t5b
gIzjsbovSkonvLHGleQHFK28pIB4Wl6kxnoE43HRrPTgYzsrAb02YoDnqoXDvOnpCZnMbJ9rcjGf
f7KIjsG57FGSvGgCglRsVHfsxAySxRMwBqr2k8Qyl1c7XUFFEdy5nSCdrLY95f0aOSciQaoDnPA7
wRHVG8vwirgOVRRsxoNUvRQjq5viBXslHvOQfo6VCZvOZ4ER/l7+E1IWk1Y5wJ1ujcV6wT6+3zQU
6dfZiFaHnQb8YaYO1/obUDZwhGlQVbn/7/SRmfSGvl+omsjNqOXoj11/+aQyL4a2Z34jmu42cnl2
H+3pY+JVPiCE8FwKDZGn+iSZ4txYW+A7RUz/HmLXeoVDXzQw+harTCMvC8W+19J7sB6b9mORdWEv
XgyiGNh8WopcYUiNp3F9fNfcEUtp7Ir3lMfkqCSIyVQYpk7dM6BsHuQy5PVcagYpNgzd22CfEAk9
wz2PktlWhObTKbTZCF669IetsKoSw966kyB2BLwv3e/wLpHJrKs/GSx8TZNIyHilJPCvOqcz9Kab
csEZKwE1EI6vMvpL+M515UuC+ad0K3z8kQuA602zlYreNz8YHF5SdngDTXvMyPa9/3/QeC5A+0Uq
oMOI38S1/010oFIzjh8aQ0wxdBZLAZIAi4Hxk/VsEM2ljbMxSNrq0ZrjDS/XePEs5gjad+EEhL9z
N2ubZ7N7j/bTWX3OYm4LGsc6bQRBcBGhC2MwFG2+ZujiqzERmaOQ/nb0G5KA7sND/Kpni9xXCos5
wOudxCGoykPhZZ7l3VNgB7AR6sbXTvgsOaiwNj+4MX89pmQbolbN8gJq40pJ0vlwJpGK4+vWazZT
mB1d4Oz/Ahg8jl8EFAuCSBJww3fp63WB0LI7X2Msr5hZ9Im5etlEkd5+uSPVxa8FwC7yT6IsR1tk
2ARBF2WNTOQd9K9Yq8GJNagYnfs7NUUeDUayNSiAll5KPP4NTvGiKfN33axGGstQlKyY7NFe6da6
EtVj3DIolA2h3R1KIEwcg4LCtczAyzNK87w/m7YSgpj8zkKvdidlbvQwE0/Iu9Sl4AsthslJ08M5
LJf015W8KP1E9C6aJtOjBpxYHQ20RIKJihUVMAC6gbEbMHUudXRpjLMGoLFlJXlfYAcQYgxqM1P9
nMMOMYhaDry0p+NN1T+wmWRf/zjKlzg9degtL5GyylWEaaLUzbY1Tvs+vSlRpgVmeHaKIKf/qMAt
MGWsb3BQ4qpXRBKyp/ZlUYp+MID4SkpGX7ws6bswkBwLSuDrLzFfskHnuvNPFQgK+KbBVqCi12SV
8diPi8hXE64eX3v9eFiyxQkuTnRy40cMC5ptdsOuMK4ZZq61CKATOOVV7qJrxixQn5WDSeqKqkso
0sSpjmmbNZybmvn8mnNGZzNBOfE4RdXoanE03K046ukMhGYtkJ9nNXfCZtWmVL69qbkW3KT/WLw2
3DUKqKb99lzVnFNn4c1NI4qvpbTE3dLQUwZG7PHdPaZ85yxn/yABkStwCKrKTqMAmIblmgj4CfrD
a+kxHs6bv6VvN2G1p/kz9P/ZNdL2Ph2fvyiFhCki+2Uobbn+a5FZ3FhDGPUlx+fq6Rd1UIkUkGVx
lmjRq0kboeibUFc0Renz9u2Xd8ITpVDkNZ0bKYQfDs3ydR/9SOPda62kDKh6FwDaeyO9s9+jFQdp
H9SWz7E+Sqmxhm3JTQKkaDQEctG6Um0EIvx4ikcfr8aO2R7iFGjduTlSpyt1xWGmpfUwF1NRIXEA
2gdxmKy3/MPfNHOC7HIrhLPUXcGQDGNQxBbeMPsvEahb9APQJXXUZEpVp99gZuvz9hknLKUExjIv
KeMBZl1UDPs/ZupHXDFrbSkHwgTJZe2Tc1lwBnDcfwBH0KCrX8JTp5Fb/BnlDoNsFOyu+sIsVMIA
99YggpY4B4n/ewcRS2RpZi4l+8QlZvvQLeYDCtkoxrhFc0sUlYfqx9tuzJpDxhh6Niu2FXUF/1y1
sGTo8q2XXxKriNDvXgqI/t3PoWTiXs/QFDmgHSq2HHhmPKXxjI7MA9RJHuTsoLzZJCEo2j5fRgn4
E2gay1JCNALssPpEO7DROQpSWFPGIy6CMo2GBUtdQQTvN7RMIRZ8NXsCQycvkJ+20iSNOUMHD+sQ
09zd+5SH71KeZqLj60v46uh7A/uU9QJ6AYkWLDiQOgUIXNb6NXPoLyPlAkJ0VzXPa7z13GSGfazM
QKSPD1DQDhhUGhcJTSJGx2LjuAbN4m27SENOXRwl+88fKcFuomVpNKMPtFN7BRwM6uxhYnaDu8vk
YjaFKRbxIlbo0xq9SJMK5G8OirjiqON384Xirm8Da65FZDsiyYmNGOZJoUW/scaSWhkml7hECTZY
5JB5y+IoTc736OvfQUJ63UaYO6/eX/OQTdC4AwNVTerTiizbcgfMHPJBeNDWD11atHzUZGUOThpX
Fh6jIp1jK+XrVPIY2PDgXE7ZMPmHR5Xbfp3gTBZNYH4m6s+6HfT7yqAJ+9WGmj2E1uWuvgdK5VwY
eOeFXDvNFnrxQVZDhoPWOyqKtb6Ol/cIpBGZiR7V33cxtKGS/a4ydVwoDt0u8fxQ/SKJgFYZP+fh
b+V+SPNfupJLpub8Z5VKg1ZxBO65nLpOh3jKS0Zquy5+45XfyTfWkPLVwX3IJOImqnmC9GDT6xbc
cRNWAbcK25QiA0wzHjIH5uI6KcwLV/D3MwGT/ZsS/b07yGSVKr6Di8rAYUzngf+MNaRaOXL1XiJ4
BavL3nTTa7DgGo+SkkvY1T8oOg1NyWvHH9M3GnQ/1CWiGMchWAny5/svYfLq2QogrxHfakDepFwb
G0HfvpqYzF5ke871OZ4Pnr/Cm0WQQ7vO1OM8UJH/JMWHceZGgIwTn4wyCeqSHR/eNvmPV/bo6twL
Mt8wKJcW5Jx99WmBnIeufB0N9vVGyaKGA8Iyvo8yc8ytfotYIzJQN8pmrhdlouxqolM/9CPqriLf
CxoJLNPLzOA6iv/+3CvTVm/krm+stK+dxIcTAVt1ZsLnw1UC0AdT1ioakN8H3UZ1OdBRrmyVg/El
KAYh6gjSTvu0jDAL0KgpihiTP+kmLg9eYufQRDmCMQJDdJczotXNchAhy1naejx0HO/gD5O+Uuri
ymuyZl/RPQLoHcRIKu+LcMLISlGtls/ZqQT5j9rXDpGGUE9kzrxNAZQrqX3maq3ca8NikmkeLYYx
NHKuwwjvA+SDj3C4c5i/NnqIgDHfIPjBGEkM6YSWSOZyENunxoPEi+bLugKnqWIcue53N2vPApSB
uudTpYqPjpbg1JAOWUfX2n0ebfNvIAUn1UT9ferTb+NQliYI8TJ5Ifh+r4EuSeUdH3Z9bi+9isVw
IcpqWtcnD/Pxh+14qUOie0bBoQVsuZs0h8N9rxUcZD5yLM49rV4I7jEr8X9GiWvzULuTu7x5yceR
VXIXCT6fngYJ3hYGCeetBkLsWTdTN+uEUFcMP74FzuOJvns6Hsnn24HUPOmdtixFVjrLAmnQwaiF
80md1fvu9mk1F7kxsR/ev9cUuL6RXYwtNtAyOai6YOnnu/yjQgtFy/XERHdcmXOoe+quwpzJEQDz
2Gkimc7n7ns+iyBPggo0wdKNlZniBC9Osw8d/oCVwzNqdqCVyfZ5XTskSKmtPBCIdq3ReRdLx1iw
jA0KrZtM/O68j3FW+p84VYBK7MWEB6yx8tjSMZoyLKu3wCGeLim3u7UCXCwzFvqMuxKQOYcGApi7
UpYk4RlPfTDNTYAUFpmwQgrGrPjK2qxu4mo0JXaSR/Vabjf48cR5gzGPHw+oqy4QT9Vm6PO6W/W/
umsgDIdqxqWyzY2KORYLqA1aGJ9fRsx5ZPvXCqDZg8h9VwMvzU3Fx2xU1fYQ1P1ZCCoPJKbLujxo
YkCM159lUXRO/J1UjMYrcxrB3rUhOAl3BndSIRZDJDObj+zg3y3EDayYVRfvAcdlPUm8/8BiYCOM
Hb1wNT35vaKaxf36XdANBTf7MyOWAeG63W5tQPoi/W6keKV4mTvygqG3CEyu9zFiiI5CaQy0EAxN
2TwM+A3YQc0mzAtEQnrJJKuYuLtp4gclovWcQ/8/Z8ZIx3A1wql/Fn9zZJ6Tr9sU9SFdIuOrXvaX
D4d47gP1Ztm86s7zCOMxsPrSDw8HlcREWgrqZkSRo0cdbqR/LqLpAFaVA2DW/mcsGtWG07yzl/YQ
WktORvegfu5LwlEaK2HuAmgcA6jxeiPqGNxm4Sa6U5ETfEtRTSTsiWRN57Sl25ufMxMvHf4N0odw
E/3qmxinEeeJYf4sIB6gH2jflK7RwAxMXKmpM4ukXg7SVu1juqPoB2AehFfMMuubuNMkzrpAd4j8
OQnQwPXEoh4xNzE/qBAxB+A3sRtOGa4eOux2m5W1misE89qjnqRkX4ItdoRx+TW0LC+pW7hCoLTr
/a/H6b8z/kZXf4NdEIhWDVJf+5dEG4BRJWtOEnog47IbpgjCdUMlaNHkaJ3mVoVplp/ScUJoJBE0
8Fpqy77+D0wOXvQiA7BoyprkvpTeB8/ZC5cRLVU69Gfu/lla1UpOaA1dZbdIAIe6iz5YFdNibo7Q
HIUNAyXGbjhYxXkhrpTrEwlCvXQrlumd9IFrAyRNUbY9iVqdeCz4PORLFPpapjh0oxwJ9DzvpQSZ
grn5tktapsO6OUzb/8ySSdg83l/09IhYIaY+83oSvBjEacCM9OIDqlWApcDS3wFRlZxsrudpk14H
WVObbBzoq6weaa2TJtCRlS2w6dYrSNuGUBdo59OrvITSAuYtucYXFl0M5x/Y/0pLDyfMJZx2GxWH
fn61eeAlxgWtmrTz/V8EplQAf1C6gS6GK/+rid0+RBq6ycG5NvG6+jkp4aDNNKFdKW37VQ6mZPEh
/uTcQvrs3GWHg4LNn35czZqTZBbNSTxqPgaQGyweqkPEDCUTyBuQFkxexhPxT8Ka2KyPLnSj1S2D
M+rwcYN7zZGqVpXUzbS46e1DJdBsZNwH/klxpvno2TPCyCNv43f4eC8NntSQXL2V5RfVKz/q8xk8
+VfoiZv9V5MAlZ5QKF+sZTGDiqpfCpZCTys7xYSnJu8alI/PzKb8xrRQj7U/GqMTOA9KgrtV58Gf
zwg6iCNph54P4Bi+RhrmRJoWHuEhM5y0N5rEWbitpSWg6DMv/fn1QqCDA7G2DEaZvtq24rKbI3KW
bg8SZnm+jg5ImRn0/8Qr57iaZD0EG5ewWdB+KVS/RE8ERtGFeJHFhUF1+jS85ri8E0Pd0dfDN10x
GBz07RyjDuaCIy+MNBtaYeWcpjys+6VT5snA5Dg0DtcJHiiG1BtnPVUd5/UhjZ0EjzPlbcP8cA0U
Ni7FsVEctKEhbcpTz2PT/seieVjAO7gGvZnj+i5OfJMet+DEdCbYFcFiYW7dFYvgSs3nr8iac34k
GD5veiO0AaX6v5cyCpjfQWyCK44w/2g32qUMPvP5MqGtzfn0L+AEMkwtODWLXfQAUrYNKdWxx2+k
SK2za+gELWrtmE/ez1R27rZ8n1WozHlyKhICGu7SZZ0JFUNCP06GXzpZYLHIQlFSjd8I5MeeaG/S
adLOu1EeKTO72j5NEhxVm2Am0j+ONzVpwJItaoCJTFqzks4fPy/51C0lIcdI2KK5tqOTMRSsUXcQ
8ngebziM2o8VdzP/c0nAIOlZ7KdCJx2Ngcg0rZco+JecRGE6pYW4YUquOGQQ6USf8IuvkYdQWamq
zJNLqnOJ7+Io1VWXAuqRNjhwh4GQtiz1nAMOF81D4oMqzHbuWgpNl6F58FMgiACM3+ScVEJtl5N6
Laii+jYD1H2PokKXHYJFOFASqopa3qb0izN1CdKgkIvpYFX1tmXzA1TRX73IJzUJUnWV5lYENl4m
QzlV55rssKBV4LuYZ++OXK4lkNQbEM/VNGmIAQoHW4kh/tMVoSivJ9qHVXXvKEi5kGSQqDyH037n
n0EW7ALF87WKhAhOISbiILrwmqLTALrQnq6SUQqkum9VgTbBRVBmji8PrVy1Z3uQoyljYTkjACLr
PBan/GOUHY38hM53BKb7Z5VFhCDFhwcaLfkrZXcsH12SU9+rCA/xDxX1gew2qReyTAd1iKt+UIFD
Q10hS9J7UXbHh9VZ6+B27a4ExAVgU8CQRE4dhATvAh7uPy7e8BZzGRRXTclEJGuc6YxFdM+Hxo+S
FFPr5RElde19E3BY6v2aD0rt5p/HuIp7KKBvnVOMo8QTTqBm2i/nYPjtU1mtF/5qJ3q0qKLJvAEN
WlFxaZrJ2xkVF+3TZTDicvGX3rJo0/kHEd3YLN8tXtzNoyZxUA2zr9aQlYfpFlRWddef15cDs1e1
JkZN+GBl3XyTI1mdwajQfCXFotiIiKPPAoShtnjug8iz+Glz8HrSSLILrfAJ8bd7NgeGZsBz45yf
crsSWLzmA01dlPDyME4+u/ZvwgBy7twSl1WOzY65U1dtnvSRxMpYUiLK8Zu/ohgxqtVlEzOPTlCZ
TB2YURKHoYB3IjB9XSXm/uTS5Wm+WoZlmHy0J9ZYZclMkKTnFx3PhY0IbaE5XoZsygFgvd2eNKAO
qlXE3ohBtdRRozMWGTv00F0om3291q7Fe66ylEB+lGreD6U3jbHUgEKTY+Kdh8+RspQxFYLiYs69
zyi6KVRfpE4KXuuiToV6tEbhv7NgW6LktBe9fPfFuKrY8S9w30X5LQSy1+UkliwF3OPeYoFkymEq
5v/fkFivxb1gA4zS7Xll3xSujk9AxOI972yLZB4EEs/Wr6IVBsyaTXrAABCdzsFvdX5z8Tvnp2/l
6ywhtSA6kAaa5l+rCs5T/CKczHGo2ezjnqMKaz7YpZKhv9/DlTfEUsez5a35RfHaw2W7vN/c/s/E
8h5XuWyB/d8Y/NU/W5dCzZH3hzCd2HKb/IVUlYTRMj63Vwbdlw4a/wxhmoxxZXE8NEPeHDHb824k
R0V3snpJT8iTipttjzYknp//a2PdlLEPtFapbAaAa1T6rzau3Pch7uAJehtBy8/D+iDL7RcVFgFI
xpfHAVnCTdHASXjWusbzJtAl/BofQrAOz96lnSFjpmSmq2E/mIkUy/qiezS12AHI3+PZfaqVl/wz
+Z1h5FUXkfokRW1tcZTgGqYXmbHcJuV/6vUjC5otMUUlaap0+qGxhKRSX3yICoVe+9+pW4A17BBe
/mMoI9qrVe/DqpfXvAXifKs7F7OvSfRpb7hvy9nLpx3dg+euTLetp/CG6+6jzP/NKllfw4T4gM3E
1NaqxV9cVpr8PDuO9SxYMZl0I7Ue6Cbe48FxuIF9gVoCNuzHykTJtj4EP6q6hjoTDybNA7rOgakx
WgcSEjcb2/RUBhGVxDBt/4gK7X0IZRjkpANsLKntc4wzug+2s6iPTAY50TfsqCTatVAcC80mYncz
PlnJlE/ljqr9KQxeJJKTr1MQDIlvd0kNSDv/dl8+BxyYftcqB8HuNuBjwb+gQEI1thPPFI/zQA3k
+qoPxSvxy9rS6ckf48pRdMs+3J21+XmbGEThO85jGTpmQ30xK6vT+mD7x/+KK+QlTWCnsj71vY//
rGI6aV5XXnuo2xjxlXW+HSNfmksqCn9Ngq0wyYLcqSBt2MbJVzPDRcIZbP2u2EV9tdHX/2CBvxlp
BjEbEI1SSWAuTBgaESK7BzSE8KW8+cY/IypTOn23sxMayCd7sf6LziHoQK3fpzM9GB9qGkmuv5+T
fuKkK3N56ZWhLOo+jGr67snSgfs9xtBo8ZuFmOVwca51alSdmcluAnUNWOiNzo6l0+gFGL7/6A/B
2fCgAlj8CR6Sf+10R7mAIox0Tjdvb4iaD4xBX7eOinwA9lMZPWzHY4743uhcjZDXqgOWBbp1oHFP
EXwS7Vctga8IWKckieU7ULEd7GAR3/PWeIP6uqaiL0tVE7x7YyKYBSBYVZsFAJGNnWQsOQc+A+bz
xZoPuHbjKsfIIp2NYetUtIIHV7w7hKNN+poLmf9nC+3giRFsicOcK/nO4G/37PoITtIu0prytXt9
sZq/hVCWvrvPS6AtdZNTTJWrzzolUU/TsH9fWKtQgX0WN6x5f1CkaGjn1Ucs+cXHt46n1lKJk70j
HOsWcUE76YkjEHWHwNXWYiYN9H7eK3qV0BKCPzTz8zI4JpfqyzijFFkgl/93OWXQ+EUY/pVS+4ef
t2QoN52GqjC4EHlkxVyHo3PIjxKvKfwH2pBOeWWYsACuQw10qhyNBoqoIx5uvIQ814FsP7dAZ8g5
b2oTjSKXchcdtdlq7zmUwFpldazh+KA9xTwgX6fC0uyQTTJ918RPpOTlbOHj36ITuNqEVnbQ+iyE
6Gd7vRIJFUCuQagpUEmBCS00LjbOYBvBv7zR4dYZ6nJp7CZzdJIgLQ9Zf4LRgcIuUoBBbVeinbqn
X59fknRoYlD+uNa+UrCALTB2KmvU6CHy+ikccKTGm1CSa8WO82m0pqeKsEMsSHHQnfdyk6QnjiSj
MIDQIZDPCVkxGGdW6vtInt/GT+LPvQ5lS5vhlVcuUnYKujaUepe2rrYMIXT3WnVP3PIjKGukmFj4
VEmMgvaD3UerA8khGDsoylLzntkkrLMgZL6JTfgxP1L/HBkYGXw6hDJ8IHkgNyph6eWOu9VXCYSf
tyN/j8xPKRFyInhdptRWq8cPlGOiRLu8bEGAXiYfOnmeEZWnIKPONuXzhep1Kh1RDt2c02w2e3H2
7dQ1FygwP226qT0c4EFO0baKPb7rys5K9SnA7yQD8zwTHxVdoRP7unkoac95oPPeTnySKRonaS+X
l8ttHiZdZdtfQO+SMt6B/cnfMjHT1woIeKsGs8FS8nzKQT8Lzm4qQKLBcOj3mCbOL0wQU3+uAILM
c3Op9gJdmIKs2UStFmkcFJkiQV4TYcso0qtHKvVQV9h9n5LaAS18Hdi0RzeRTPNlkjYI/BjlNVFt
IpxTBJXCs9JcALw8M/W1XE2aDs4kNCM/cglvzOQ2+YHdUIKBGL4FET/sPpGbjvugmtkYuRRfCjJf
jff6zQurypiD7O47kXVnSKvE+2b1CEimLOjOW1lFMs4CiP4Y8+dLgb3/sQvUgW3iX3GgeAGeJVnx
YCh+7LQ7QD2qXLcYb7X1uxw/hK1lOAFl+3qK2Bua/vsyb4wNH2skZX7GrTyXi1R67F/07C1YV26S
+pPuCDX0feLtaw6oxDquNaL0EkX3vY6PE73CAt8oHLTk69Gp82Jhbzwqewk2CrXA3zjMJTtWmO4v
o17MzIZO1aDr1nA/lFraAs99i9rOEjNlykHBoyPG0uxf7uBEcQjso3RIgGyW9c2i5B31Jc/mk9VR
S+vjktGcIJxD3l0N9rt9fi20Dxmsum/6cpsmIROk43AMoPORqbMO58NRfZpmpEhkx5BFzQfnqNw5
o4bEbFp+3HKC/eks1kqqsa9P03P7HRl+Rjn6sbk7ajmKwWxP/gAveDG9Jbz+ToM18njGMBOp+P9t
912BcYfKCAJQQTxHtOaUIjVQG32ao1Nf7cP4wavhhQJC325jVpluAWTO0D31gglwZNtW/em4CJYQ
AxTp93O2blO4hqzpY1XgHK/NYyakHRU+3+wwx7g4u2Y2Cc+COh2qK22pPLKSUUHVZ/9ur+SZ4JqU
D06fvXqSlh+zUtNJwtSBXTs6SKCO5LcFLzx3fR82k4J8vWODV/Tn/fYwGg22Z77kNLzjc2AD/Woi
ThkXxJRT9EPO/XYatmbBQG0sdrXEvabhF3h/usuSr1/AyQnehBov9tKmRQBPXn6f+YVnbswpHIEj
1ttWXgrItAPuUQVJPeRws56pY8fOtMgvfMBGrHueGczxG6bCmEUJzgUDfUB+UFwFDruo4T7NCnjc
iFrFHdy5OXzIoFiG6yeeubhzxJxcZGB5CrphfVDwWEXo+gQExDudjf3rEPj9/mCpw3VggthA64us
O4akRdVbIiC9QWTETOhI2YWO6r+lN3O2EdD8cv8YcJhakGJLhuDKuP36VkrtOE4JNKgl3WsrpAux
O1fWd4LpPxd1Jvd2cn3KWIECiVn4pFFMfquXkzc+w2HZfSP4d2H0LkXVSIX5QlNqA2w4nnjdYk+/
H/Auk4CElv6aKj83Pde3vYgz3DjnRF4Q+iOKWeRsMLxoYlwmU1FKRB/x6302TRTyxBBxw2/e4h+n
ajWnJjpSn8CcJBecxW0cTFYAq3/qpLEdVxI+BB5OIMjMoOv61HuN1i8CubocmAxpkSsl2LzQ11cS
MP5/FGSCa+0zKkbgHXQCO0B/84NA0GXu+7/kAB7Ybhm+BvD7kjlf0kFlV2rxZvVyp5tFDSxcvsCh
cDz65Snt4zHWD/ybOVBB8wbGp8N/06IM8mzuHLQxBYgCVKisGV+5UQJ/FzqVWGVVKcO4tU5Hk3kn
hZRgpF+QGY3WRQhP0+wcCBbub23r0jbX81rqEu9MBVAe22K6cSBsKbZDoDuKmWj+QOSdjf+EGfjU
w7RYNYud77acQlxVgCUR/qlrvtK/QC5R8JHhRDmz5v8T1BVBqr47iYrNl0Qhu4rNMyzOY2C7eEGi
ctTrCpAVBQEt0/x7FRmZty11wxL8P9qlfS8MYxlwTALu88IgVohO2iTR0cSPeTOGdGucjP3jxTjK
Do2AiySvJyBFPBdxLC3XHSlCIT8JYa/Whe/+qYgpMi9c8AtysqXXGlpNS7mjs3QOvStjkE7v+fvt
zB+nLPwewPSAYI/bqkRxWQReHX3GORWNjk8LxCfscfiEeI+7HvqkZBja3wgeBVvmgMqE0RgJL2Ec
DLYjenJ7/Zh425NlwrmRDSvcP1cPSXRYy9ylX0KgU3UPftJif4cErm+UKu9hViYLHfo3SWo4LxFv
fNsNohJsO4CBJMWVvatrr4GuvO2U0fKlGBhENHw1zRxmDsCtkLRnRjaA0TfaAH6LQuQjVcSVTcSp
nYenJLvZS9Ge9wbjd773b/cJURKycDxk6640H1LuPgpepxiERipGX2O9DZ1+6fSIuzxFLc/AmofH
fg2Jp0qD3RiH8eryV35o15g7Sf7aftoY5f9fcbA4J+rJfOEKuHSLk6ijYhrwU+Hq3fZo1ODFXsKE
zFksFv5qD+zYOgXCE3CxmRV7kgnp/n8sCBfO8qd0pU5FXnxGWpCnmH2A+ISPAs+UNcmXfiFmWc9N
0mWfiff2Yj0kwyZGByxWjHpoovHSmJq+WOcfaAX2KiY758hKQJce+/VI2IV6Jy2qvGdC3TGuNT0e
X3G9yDV4r31TOyFKBxCuUkKQKICIGW629qw/inW1PiiPRrhuayK9WLTF7LW8QQ1CN6uFSHNAC1F6
MP3usKWq8CS9p5O2h+KBpon2IfWf1bTagu2Z4LuoVjBVLZoEpteZ7nNz2pKn7T0AW18fiUjbY8sq
Lcms6+VxA4JnXjYSsr9lKfZvdHmCn/jFn2Sq4L3rvQWVx1om3cu6AKneKHfDoKzm0wdYDK6CqsOn
YZVib7ufZXAFVi3ocHINCq8sI0OWHKpCtlydlqHd4vjrfSDhlWOjEs9LEUBqtE5y/vjFEBJd7Ddm
R7kgv1UGj8txDtrQGOlJ0tV7dAzPwD/jhQIEgVvXFtop9yBD7pfWX/sfava8/Bl3h0tdvMX5TLX+
i0NHZ8B+0IKQCcETGbqeBkC3DBQLuDCAALgyzwUxXMPkowmv7EYSdxK03zpccXUUpxZfs9vJ15d7
aDuAUmdZKKjEgrhYpMC2PAJVNcnU4suc28zztSgFFfg8IVihhZm0XujsHaLSy4560AAPdjszeE41
Q0zJiwfNmF0j68iG8yEAu1DNMhR4mC8PjoXULOyzuscC0KlsjuO8VeONKpPwHgUA3cjikV4Txplm
7Waiu0q8YVv/iuFQe8zWZDBnqzByAyNo4hLMYlYRQx/G0VMV+B5px0kZxe3MSSBeroREbRXKI+m9
bogHh5e3GXyseItTT5jNFxQf0CAW+I+IzBD7zIUYZTPcX26rvcgpGmYC899BG29kvmvVRan1OaTE
VKIJhqMUVnrlnK131CRjMUjXeQOSx6ODJA0kVE6EhYucyWLYiE1HPhaFbg0wRkRt9wqOwSaI+bKM
1yRiR7p5+SFGfSfrUjG0epel1ElP24fQYyJwCsnS9ySZEvlvP7Ser3YBBLUt8hPELMPIxXI3vkdV
nWkQ74cqbqkKApNah/cnOWo2ZDg0XKhVUJ6Os2XHp3x4MQoI2zz5/mLBckdUa3B3Y28BgHQn/tP5
AmV5iBivqhnS9eRCt1AyhNOs/RQO2+4YhQ6fJb+/+0yIr+cqdfJNZSZtOAtYT0llw3QIu6WD0iSl
YNyKObPlQnfWS0Q+SbLueCyuAokvCY4D7zhqqoBfbEAxYfO3Nb02REsqqbv/aasOwiV1lEmU3vgA
X0jQnAMhpbtIEau8Xvutr7QxaIWQ0xpY0wjauMmfPpY0DKTWUEAZljWrKkPVhgfB569blm5OpvtX
m/D8W10H/a6Y4XtYVhAT1+8C26lY6WC3VkDe+5+rvT2mP9TilUdcbr+BpEqqZ3x4Nd5AZr9swbZX
yv8vzJjCcIbn0p7zoa9jrJkXfob4rYWfeAlZs4csRKd3FldrF7wcOalw3VI5t3eP4QtEyql/FIEE
wsCBLSpd4wwgEyJcf2q2W/a6MB1NAqKc7aU/PceYdM4fvl8cILD6KkGB3z6qx6Y/3cgVilcoff09
tyJQXVf0JelD7EDhCYsuNR0X5qk3oaHN8+a3wf0j0IsS+K1DC+dFrnLBIMXvfqc1QJgujDpGFFL0
5/wu8FV0v+TJR4UuisG8D9EcpWmzqUJu6L0EY8HHIpZU9hunbCurT9BWEE+LQvVwRLwNntJxNv1f
I7bptwpC3+XBDCzlZhzHEqAithIT25sTYFjptlf3642XyOwcjgATqdRUQ+RVmQPDqzf0MifNVwoD
2mJ71wIFM27O+U5jHpBHm4Pjx18G90uvkxVTwrom2ASBepAC4qyzxs/V+ul96b+Uh+YePXFIZ1qN
c8b/LqEIxW9utHQJU5LBdXOwFNGifWzaXPL+eqtbwydnTDZuNBp4bBKWPP1poQ2WE8mk3iff4heB
v59tyO8VYGjEMsONu8+EgtnqiT2KYYs4MG10IMtq9DeYOvzvG+wv+G9pW9r8jbcRfklyCeN3Xif9
vaC9PwqbaKqbxlabUfnMuyAivfSydpR8EeGAKogZrL8aJhVT/YKTszQt4amXEQxdgsWKdAkgCIRw
tYDuSQVXTV0VsCZLrzUOJVWXCexemFN0hIYU5r2Cl2qd2U2+qW+9654NoIEtkuQX+9zalFEEzL6L
wKtKo5uZnsVpBJML5e82EjE8PDjbJYGoIxj8AfmrzcXled/QjpYVkrcBoW1Plrw4nqDdYAIQ7MN8
q4DyH63dDnBmU2flKxfHdBM9mBk1Cy3Dgzk0PpfeN/YROq9TDm/Hnru0xTO9mtmbRwHfq49oBw21
iAzbuRzQkXmMG7qFjRad0P0mY2t7jNxDyJPiFKUUinm++BD/PpVBoGA70J8RV5qkQZM8J3vXkLJj
0fNyTgk8eOQTdGM9VpTO5a2DFFn7EBTGSRp8/VMw5M7Zo7tnTzGYVYndmx47te9Jxfi0qS16MpgB
knzbn9NjOZUjlWDK5dCjtOrykHAlEstsc03HSOdaIPMjcxQ3PbTZ1bZ82ecoGFYJIqEf9Ys1+H+u
Rdd2VjBcP2D7nZZbZs5Z1w7o1OzJ1K8P4PwlJmqiNZHOI0d4Pk3hDmV5S/s5IQCiAHulIkZaEYUT
/5dxuDZfmEVoCQIZsO4bmiZN6ZiGJSkXQiCiJqNvZ87M3eqa68wqZLIX4KrkLvtOy2EswwshZ8lk
CrUsN7Z3SyeE9WDOn/u1qAdHW/0Z41Gn/7Shl/EyE3yQKB4YH5E6ywQKRiZWj2L9qOwRmRtcw3of
X+gxfVyoYRNPtxsXjfuJ+le6uGi0LZ0l4eR06FXoSdSDcXazPLqcoGM3UyqVdRrMS690l0mapoHb
dUomaqmVzX5gXYKdkAvWnKR0DBE6fboo5RXncuth91RVz8BE1D0eETkmREul37LUkah0iLBytN7t
GdZLh8v9/CYZG0SBm3LIzuNk0be5UdXwMmMM+z2n9ZZn96gXK+gqXacxcF0xQiJldK90x18CHsJD
11R+83CGzNCGwyqxqLQCL+1L/KfYJHhG6V34gRILpxRo5XPwd3L+8XBWUWGNw6opqLOc6dHlTwAG
BwfZ+QrWDcOgOLGEZIzAKCLEqbC7oNkv07aaUlGu9rVPOetgZ2zUpgU50006FSEp5XkDfRFHbKFH
O654YVe09MQqWXiqbtlNzzUvDV2Z+mIS051lvGuPAYeEt5QqIMUtNYR/VbkLhsrlmbDrzN4eK3sY
MiAiRNVnG3fvrnkmN1m/QOvVLDlXS5umvc0mnzCqUUBmyi5MOwJ9CtAMqLlERNzE92VpgmavwMB6
wbfbLDfe7RqxHPYIEnTeH1E5wvGi/0P3f2tEgiy53/LSFkUQIkv0QBlFCJNhPszoDH/xhoEQt7Tt
ZMHsn3t6c1Bb0umta8rNYtG/tQn6Y5DOkvVkkrkdsiJRw5jBdCDLxcqM9SNlG1VWYuoYVSnna9GO
CxbBeiMNFUVVDZTuNR75d1rTGoBuuATr5jgzuNbGU73wqZlwbvvhMgQSy19rxoH0rClfdvdJk+Mi
OFIoXp+VcEb9EZ1IQIvfaoidCFlCWAUdXIflZpzntWNxXUkFNQLb1J6UFeyL6hvRfc6cL49p2Q0v
pR3gs1Br48i+5mOLLamVnddR23zOpUpVdRi6KyzWndSXrGkyviz+Wqwjy4eF75Qlv4YhcEpIO+pO
F9Is7E5GL6Mhfk3nCmIQddz7SvhujtZ8GOdplRvvUHKPEpusmv94M48+bJy8AEHFs4lU/77ihubz
YTKclQevtORbYf81pvA0k4zAHc2RcpAN+47nSz2oERVnxBBE/LmfU70EbxuKo8NV1WujNqsFDXxG
whSJGkXSpgZTxWcJ7pMhzw0iar/QODT27iCDHgj7AqrViYsFnHtJh/095jRPX5M2MNs+gxiTVVjF
XOmiKS54t7XxSD64ehTTpi70dYJcdSp0GARLyaUu7Ztx/SnE0NULFzYcRfOUqUYtbfk2k3Mtr37M
Q32an4tJAAoDq49fRl6ZxbA00woxQrTAxdhf16Q+jgks6g8GTzQxt/K7WpFN3vdQ1oPdRj4ORvAc
Acjf6LMvr0gKFRClX6an2IZQOvDFTdl+eBoFfqXoIpYaQvyUOlbz9UrYhkCnoHNTO0+XRZxcB4Yl
DdFp15SQ4yaU1CQqAVIk8M2G0Jzd0CtjYSFgoi9dVnoVjxaitzZV+DnH0z0LxNGzIzqUK+56LLvs
PGpXVhe8tbzNF+ewdOOVLRUUGGt+c5w4YVg79aWpAkDlEJ8IvA4rk4o6/u1cFFMLFT8FpPT+G20L
BGE/nlM7lN23QIHRfyIfODXkIMXp/Y9eGANyVrnX/88OmITMOsMvRYFiIcA4S8LdWXfUHbLrG8kX
mDdhS6ikz8SYf+KfA5b7AWFQLIPOGx4OdR5nTDQydPRdNTu3Q1hU137h4k5FpEXDaH9NGQ0uXZLN
cmBH6zofg7k0JPn5wypB1XZz3JOwZ9iDuFLQ/BnRq+d9mJpW/wHmhyXs1CxWOm3YHX5DMOoosg+F
gvxRQqkAkT0eYfqdaLL+hehiusIt21w7vMrS58qGBv3umldMgoJVxdQZRUuwvb122NtosrCehDKb
QBtv8FcqNAih/yyUHNtPRad/PQRdDJDcnF6O0SWP+DesyY/jxBLCUjyZ+JyUjg8qLb6hWVmRDdzE
cdG6pVL2B30EUFydETnD+zgBTY351QPcQFq+yWfPhu1u51PZxsLGfA6DkIFELZlZ+6f4+j+ts1XC
Ogk5F4VZ/nurk8P9m4+Dw4RqwreCyF5eM34hKIWRoUrD+0E9AKPJOtd4kpBbPCOLP93u9DXicOqt
khGwies8Oc7zjqidzJPyGPR/cG5dsxCImuo+tnS1H1XAVphXxtXUZW76XDLn0d1orjXA3nQbTf+V
zrOqRlVOpMnxo7sag1bY4h1Fe7RLG18l5dtUIXpH4nt94WTsiJhUS8tKgVEQ5ML8SiCOrOal/dLx
IEQQP4bMOw9GE4dC0j9E8bJWQiOx5VVBJ7Z6oGmUuTRqYD6VTYa51ON2YWJ/49zXpfvg9+TlKxuU
1Un+SLmlGugRq+rgx6cw3+VKq1GDrVKWSrfUJ3pRVXta0eQ+XknARcu6tuB2ZM0x0kxDN4jHmTaL
2Y/Lh283D9X82fI3vsnUPZi1RPl1aw0aPEJyinyCnJ2yYiRzz5uU0D/ZzBvqIAFpvhqZx1XaLiBO
VKWjFNMXMyMRbBEzU8miYIJaWjSqAQJwplX+2zPz7L8DvuA5SJgKgpopPMjk8ZcYoYhm5tnwWhc5
Esnwz7YqCZq1Ey1UYnLWG+aox7r5H9xMZgqHoaoqYCszTnCiaqtqU8SLkKvmUACXBjzBEtKDpdpH
JWApckc64HqcmgKfnaOWhVlSf7EfDjoBXYRGpor8rvdZFRwivrcKG3OwB/ZZDF8q6xYRLXkFvpSH
IcV3YPJIVLXuMBKrc/yBy1n8CGMLFAxBP2aOr83oBAGC0xgxSQdHglHwacFZmHtRzcjEVbG5Vj0S
g9Tn+Ko0jRQtqztu/2m/zCCuF4syxl//Zkynv54q1QL++CreDv6nFUzcLax7fWgk6w7N+e1gUWdb
xTPPC4zyCty5ZTqULOTBcHgoDrmdTGu4DWwqivoLWaQTv5+ghyIuaKDievl6Bpv8e3mSdmqmZzTO
B1FUsxjJSvDyyEFBWxdaw45bnsyYLVa31eOCMfdcF1OCWk8g8Y1Y1EQ3z+qNfg9EYaVMl+h69eE0
5lfPI+HN2haNCHlAxfhuV7FwhOEYF9AkQFx0ZHe1SFyK6wtlx3SAxKws70PizYpLK/7VTcX8B/Ot
Dvt2nfcgI6mHNmYOpNvAtNsA3TKUZzDjVcW7qQ78S+7k1bSd0ZvhQOtomoEaDvxt1hKu4nlBNrks
T9Q0/qR9ojig+qX/qPJYYnQkfIyxz5ZpeByIFE2++q47A/D5Qf+bWe36jawcV6E+MLoep67SX2Q6
+XVdT2+CD2O6j016MaJMUoH2f7+CVKojrECSK/r5inBI8Uqf53XCHUOj1KRZRT3wO3lBbhstCq/h
M/aIXITiUe3oXrusHfKzyIMCsBT6klNE7ccN/kSn9ivtyU2NFnJCeZ4as+CrzeQCfkAcyK8XEzbg
3FPnvKrJg9H5oEuQ0SiUfLESnpupQ/EgeSGWdXpHhR8J+3lZ33IrLuhdx+WEqeesXEuHX5kwB5kp
SMIr9qmPx10KwhENPFYQbxKATdd0gLipJeTiI3xgGcXuuCe08zRxodezUxEsdU9H+outswMmB2M8
EIQfBid3BCHtCQtDOnWmTNpAJgDEXleFMWU4LR4sSGQKWZTiosVnBIXE7PxD9m/iGT9J4RwQeSdW
BLZzc/E24xuB6wwhk00QhGJlQ61ViurROt9VMV5+4KbDCnsubL1o48N+15cPinF/4r9saQOCaebA
8EZQfEF805qKg4N+5neKyjOqPmw6ziSL9zMJuuR1aV8AhplaJYm1wAUTZ4UGkzYPvBdUAIykbBj6
9m1n3h3Dw3b1Kobo03bJVDBQiVn0gN8FBTLjrj9uKpjlABgDg8XO4LCrdwmy/NJ6Fkxemr4TYYQF
V2aCjMmUdQX3WaVtcqpekPaKi7Ln6vCGSykm77gzhAXid1aCBDolDT27901RDCw80V7buv/h8D0Z
2Jkg4VSaL+TUMlJXJvO4Bd2Nw+qlthjyguEoNJbuMn1CG+LrDMc+fAaLJMMAIevTaMo5eVeIcNh1
Jpuq/hnouApzW01o5D2Wi7WmST4ouSj//3G32b/7lQd+qeHBImoEq5UDbqmjN/VKlFXiaO3ZDKNF
gUU7cA8KOl1Ci8GD0pFB//MITU6IUgaCNMtUIz+2TjHaJgbyfz3oCoYfGSgZsXYFMedBRqVZjNRF
CS6F5IjiU1OosENAhO4l+ab5AKr+RaiTPfdOwRmOnF6Uwgie3IAIoe7wWEnsR0D5mb0gaYFimw3K
Qu5fj9dbwF46+6hEUi8A9TJKkRm1pkR+PdeYHrpogH65OCR0XoU/RkoLIWe0BHYh41KuGTc8To84
Eim7tsYri09uCbaCwt+k4XjW5pR/27qsRtXRNPRwiCuw7kQLsnqSYllogsmdDISSKy2JOpYrPMDO
sIEBAg9zR/QP3PeiyxmRO6iEGg6hKI4Xr8LHvC9m5VxYNUeV6kxCOZ01KsdCTx8Ql1AOvhX5mjbc
Wxhh7nU8SYWlCvTrvuKGMCyovgOlU6+BdmMKFw2VlheAhZQlU/x8lHa8IrfvHN2MMGoigLGGeQzJ
cQG9T+HcQ382XJh3L8SsTRtVihIzf9PWsWvCuQ7f5c8JSiC8axk4aUft4F8OfbXfHs56InzaOBVA
ypmWbhRYB49KIux/jalZU1NP/VkzANhvlolMKI4VBe1CmJgVAwt/sRxqsDEQVPgaeaWCPKQ/KRFA
8YBC2HgquOBv1sKsub4b5t8pgmqXgT/qMiO6SzudUmVqMLiLi7f6kUsso0ySJY+Dv4H+WofjxxK4
eVktwzVDrOd8MCMMIcvyjMbmY6+oP+vcGPO59iZVGwQA5U/qWK5IL8CX0N20zTN5eLSHYiySyBm4
pWi5F2MkBbLox2aAoM9EgjVEPS16mNkf6rNsKH5VqO0PmsUIuaQntiThRQusluZSchy8UOhyFfax
kSx7I2FrrfN0WlXoAxJp7iaCqKy8L+ehILlN+0u8on8f3hiehlwsn50+pKMla5GmVI93olKag4uX
vM8KblErbDoxK2IF8DQnVMqwA7jS0xFbNzXSFmTZ9tJ3X2VoK3d88AT+GeHd/nsV+gH9SJNzpeua
QSpkndJqBmCJHH7D1VdntIMfFsOcF1a3I+uHr0MuVewS4EC9GfimTCanG5zB1ROqKFnbuTY11Gp7
x2lPPTR9MWyCZgMt2NqKD4n6nSrCeP0eHO5O6oUX63LXMKQ+F8EpX0ehy3T/yIdb6QjBHFUn2EUk
P3h1B7Byf5XPQ5+X59zZ8ZGbXCfwGGOKsixixZGtjN9Xs+cf4Jv+yQGUQ7myliMYHupQTfPyV5xr
+8O6RS9vuPCh/A/IvCY6fHwKd30UqtS4ExPzHomimfNj7rbSOTQlVPJ7WYrOjL87VgcuyxflLD9Z
A0qj/PTht23Hql8OiXaDk7CcyATuN9JvHCq6JFiBCPo88vZS/2jNeb8uUf5ZTEAAG8XEm6vJgYL8
E8lMD1akaH6ybwurBfH5jKXUd5Csydb0OhF7pd1S0pZFtS3N/WaJaJHtRtWs7Vh8f9vxRktBzuqZ
UnbYa5GZnzjl3g0nEN4c/rkjg+/NNC+qSYgInqfql3C5VHwtOUfdTra8k7uUSjUddGUNXHyIcedC
2n2mCqx+SYG+CnCoJX8423gJP3D9AfksFE9wqnOGEu57XfnXn+58nvAYkvZIIgrznGIZ/3VfKK4G
2Az/nZcyGY5IJr/ltlWnQCdDtLhmsswBFukWfbm7bpiMSeOfgYrebYc3oCudG6dZH55+3neCFK2o
1//qM/AGmivU72Iv8pr2wWpPf62H9hbk5QQ//9/z8Un7jAbKV7lcz6oJijE1E4QLfkEqnZpBM7gu
0tYABOvzPUUWqQMZWrZZhCToZnniOOCXKtFBp821mhoFbvpVr1kE/6MPq3+MxAwPXgl4gOhjrVb2
5MqdgbLh6XJXhU7gx4GiVENp9XOv/GVLvmsbfD9+rbFzqY48XMWh0ymmgaAdiXmm6dY22B/O2+vA
kjzh24Egr58eEe0Q0D6Vmg8Jv0MdgpSKUC1a0+JU5x+uPFsp8WTRSUQjzKp7Fb19fHcyJ+sFWI6f
DAmOoL9Q/nSu6ldoMNKEVYvB7yAwCRg31IcnDaaAgQ4RPjUaZwJxH+cz9Zu4zwO0ViGOGnhGqcZq
3I7ugZGAiAk23ou2/a84+RVNUBDf5t1YlLOp9XXTk/n0LpbbRNpylZI5DVkuAiN5UfLTRnJckNwv
BqCPEYIFbgdaDM2WaXQifBJLeihj7p3yLs2Cbvf54u8cyRnbV9upjya+e7OVcAV0vlYo4Hklz650
5L/wpuAvRug3W7ahGzqOwWFyxklCwCI4jwcdVYDluy4EriRtUmdmullLStut8Ygszua3Jghf1DBj
E8gxVQGJrQhb1Vax1PmpTmqVAj1xveyduXcWxGpmPTmPRaDQWiboSoyc+bnsXnRH0O0PQO7hTB2v
y1WcOEDcjdH0NsHDmG3fJcqYfKjzMHJ1g1DW8jOcfDwz+WTZz+6AHc+uEyR9MSzeiR2cZS/Me7Uy
aJSgNa9het/zXDkdYnDnEmrQ/U+3FibqjA3IJDuhRGnpQaWXYdROGQQA+pNWsdm1tQqIcHQC/A7W
r1hofjd8NVW0ZfBOkZZEvjeaBY8EvLW1j8dzRFidGzof1V6iAEj0JeZBFAuGmd2V+DQDV+GGTnc9
agTzPxdmCP+rUh0qsyPivohRVdrvZpmbUSLoQv5HZukhV6I1Vgf4B22rC+hh16D0+x2xwEXqHFtD
YUAu1nIwc0w7d3h42/qYAOVJG4jqwmJ/7WWt9tCkuXlhinAQ48YEgIb7DAcoUb1opQ0KTOPaet9b
6QN1En8UiwyWwAc0ppZeeGE/QOVtwGegcM18irqQ+pfIu0lM40b4Xik1OJ/oLrdh5P1dT0RWWdlW
1YSwyfHpwNPLJGAtoZHC34ZN4U+Eq6gVFGE2zNthHDMU02rbM802D7rXcB57FoKcd/xBKSw76hFw
wgO01yxDu8eY9Nhbss+jXoofVxWok5GDF57Tf3P1KYDI7UxetJ5ltvt/cEMinxn271Xpi9rUWUVb
wUfvP07J7XOlqGgoYOWuKBMwMwd05Xwko2DCXgHtE34naXbSx9bd5khgPBTNWNaPZp9KHofEnTb8
BDXoSZ1JaKrfA1LPVTW/2Vc/IfksVVmD4NhF7fCtFepE4XjyQD+fFUWuLHoBEqjsW2dQ+1SkhZiO
9u51rEOZHk4vIq2VtUg/u3DV+U3M0BqA2BChKnFd2ZWZpUrEruIFI/eycHrDlL4G6tQuzm3aJkSQ
xVd6l4kBNeh+ghCevnUWYy/BUO9uQoC3Ztk6ncQG30jVo23Zq0sYZ3Ge5Mtbyv1zjNl6X9D/Ipx5
7segHLZfGJ32mOrpRquT/MA1lcHXbWhzzdxr85pgwvGSwyOZSD2B+S6VOa995G5ZgMCc0+IfU+8Z
QME1/10Rtz5m3aB0zLLfjZ4VD1N8vEnHrsULPqw79ZSL+88JjUO7rGO7R6RXdDu3yxhNb96rjWRX
CvVtwWwZ7ySaqxJDsT3Gd/Y6e7G3ZJk4Hd3t8/pIZLA30Zl06kyhGrsopDqVhdWj3Mbc2k231/JP
4RrydsrXEmQ9IoIEHQ9oIgiRpZlh9JZKHevFNvd8YKTAvNlfOWlaziNUgzFMyExJOBw7EhJ7LFjB
5QoxxCnYqn4Cp/LvnJUzHajxt+Wmda8cTRn7HuXQxLsfQAOVHMl09WpjuZBdAdP1Ir0nlLS/GoR0
UCahK4nxnbpEIOtXZwD7YEGPWg6wxZWOMwo9qFta+IR5bUo6+QZLXU8EfH/zNiMfb7gjMfH72Yuo
dI7eqG3ZJIKHW2kzAcME5GgRIaXPmfXqDmuf6gD8CsRi/hgzFtETNcjNkTFAYx27K64Xj/H+6oPr
22WbmxVW3sojyBG6/25r3OPmcJph629dUO/PZuYFvl7uKFV0+NQUcQFXsVA5KJj1WQv4XcArt4bp
sO+QhjqCVX1FMdEboEIdTsMXZoNB2vIdSfE3Km/JzjFAN9RIaRKaOldWkA58WbVsrQBERZ9NTMvs
N2ch+hbEaCDyDxWQXs7OhkGl/KwQVdVPuzn4BmVROibWKxHf2vIQnMbQUaH+cHM5xptlo99GCFVE
snlfiWyWljjkIyzpb9EeW5YonfkvKO/AT+hSQ7CSjTgpHC5umYwV2sdQ3EKpFL2YVFUaqfROxrL3
CFW3QZFRdOvCzn4TmLI1V1TIuXqr8la/KSoDqclye2lQ9Uh3055P1shao6lP+/6JRSp8YIS9bSVJ
gWHIW2Vt/iT165JiHkYIRAscZz55dC+VEvoHiiPFdA+zeCNAsjzTgTYCONwSaFhQPy+cOZ7w/SDY
8EYqhUBZtNZHAvfEoJsKsghimiWj3Z2FVqQ39tlbuKzoDpvhLkiiSs1/Znc9Pgieom8nztAJYdGg
ZJ95OSFPOUAaTZyYGWu0q9P+P5dWWl2riHSlfE643NxFmv26uSSpxvIgWRPlxkGWpHXFHGlDKSPW
SZ7m+59YVlheD2a/MB0622KxFqNpJ3ITTzxVS2ZQBU3L1GJ5QXLPQVaTgoqChohqnn4QkdLwZkP8
u76OkQBC3HA/pnNUu+K7SWUGuXAyhgg5c+VBi5KDLzm5Cv0k2ZZk0xziuxYpKs789azsXBit+ygb
uEGgGK1PHHK1s5O7L+Lq2LPKEEKkmdSXr3gCxGR6j8Mstg7IcLbnyyK8F/qizPFic2d2nLKFBmQh
+gE0Q1Dqmm5vTs0Fyo9QmQW8GkLiwuicG9dgtYQFU8+zWMcV7bMR876hZTMf18txCwKVd1BOwRfI
/wjbikAjvmuqPDRv+f/C8g9w7l4fBkQ05KFx54Ose4vbNeg/Z/L3pRa98KgZdIGXglC1nHEmIxnX
/q0FGLaZ55UWpZNrKJBVIPa0ofc9Yfl/eBa25VllRUOrQl1g49cDuvI4Rbz4IWgE4tct1eT96YJI
63YuF9CaAhJn0vnwry2eOzdKxbvyeo1w8cPNkUyiZ/awZLsplOLiiOLxucLDh3R/wwM0Fccr8+AZ
iKXgQQM/q951UUM+7PUJOaUgjVXshdryMx6ALZ7YPsGtqKAZLNxTISC2MJlRW4HuykmgTJVAJpXn
3nD6GkQHhQr/0iF74GjQXKNvFXWZh51xS+tT4/3I1PQT10Jyql1Pvo7jdvGg6U2oaWXOUCThpR87
I8RfquIWLmocRC6QEAyEZTnLzanH3tpaHC0fKet8/CcSQ+Watim0p8xRVEEwr5NyG8c2bGeB65kq
r8JrQTvwZ48zlD38mNxUid0ZXw7BKPTEn3b1tHzPWIecKDTBK1iiKvslIVTvm49ZTjtUINFAXzdl
NjzZSo6XS14mcyEZ5DxG+8GmxqJYudug8JgdOERK6pKDJppiSWUq8hK9bzxQMQpZg52iGeYaNJYq
uYKSwAzr9Bm0wvjwk+MnP2EdEt2FU0RA/sqdLLxVZaqaNuFRFF3aYhkxp7+12SRqsu9uXNsO+QQj
9qomVND8aY4UuanDrkp7qJUEhQKvWp8QqaoINpe+lvXv0Bqz/mypgHAYREvvCQwHtSdqai/x/VuV
DVCcoWPk994skZxxSD/vKS6Np3TYejVw6wEv5bqbMReNHyFv6tZB0l4VryS4M9spCiG6IKwphlUj
iuOWQ+PdYQdTWq8H6LfnPqTN42qoytFNZx59a6+AxlQE6ShXQavf3gkjTnuBlLIhZNp0WgYDroSn
GGHL5pHaX2Db45e6Gt5825LaVOxgnzF493yoyg0bxq2Wt/L7WS3FrxBJcZDnxIBxTzZDka9+eEz1
H9MCoJ9LVq/tHSZlTF0tyKjNa5sm8ANuiMYTf+I1i8vpFVjlQy1AM784cTVVLnnfpGctFa/FvvHK
A+ACpSZWHXaIJIABrsEFOYu5dMSzcVM/3kYGz8RlMMnFe/WN8/EwokRLaABwMqa2AMySXbhLyQ94
+PqlK88JTYBI5VsH6dFjSGQ+G1+07Z2vPEmGnY0C4cOtqr8RNlTzqGAtcMfKoK19vbcp/sEBYu02
io/DjTQNOzZdfDht3leuGrHodwL/RVWAgRNBuiuJNXDjN1hBV0cv6EAFXzmv6mkEzbq+u+gf4iGF
kblX6TeH4z/kUAhuOHI0Z9akXYpYaBwke7dh4Kq/IY7UFU5lESqRK057KpJymX6aPy42A2vKDQC+
htnFwRARGJ1Faf3oTNlS8rfhp1nj9olE2iA7VZVrcfBDSRqen5WCQhexf9aUIj3I82rdMt7lQL6m
65lhvfuFtiYkf/5iHKD6lT+pE66u0acdqOrTJ2saJC6P1Ov1uUeWEL+pDdk807587JvhHCcsOeOp
BAFVsV2TDaWKT1G0RNb6wtPVCx9/BEH0lR/Y/QRC517DGIu9revH7X+m1WmzAmibS8XclBJRKpwi
TpwJXRfD1R84oTednHkkgVknVgPCWyPkrSRdLoA2+Cr7fycG8JvKlmusXdo6XsjoS6ZDWPHEpVug
Rg+ufgg0N5DnMB/2Z/uowaC3cIQ1fC4iWwEc5CpqA9pCai0HyMRycqvpg2eKG6SU8B1QGhLUy5f/
UExALJov00ZszJFhrFnF9bcoLRfdXYScQSwX3WblnhbhXNWeh+wtSvSY/91vtn+nMvyyKJafX3sV
AajZflLfM8HJQqRx67hFRbCpFwYMvMrX6NLIU4DLnGZHB4ZAnbj9gplWLb/3ZQxlfGNAxD3MwsUg
IojXDc+m0t4LrropasiE8zoJAPbL4624os6G1lx0PHIS7bVoxj/kiaRd3vOJiG81Tk/9yJZure+A
v7OQAv/R2Gt5Qn8pR5bkOyJ/zMpV+4bKXWoEAbNB/zSsxVfXT0n2Yp83mMnb7DM/PMrMSiFPVcIY
TU4YbWw0PIo81X74Aj0PytSDnIGhT2waFMqw9a7tznY/BY+YZ4O4Ne6Zwbut5SRWCBV1kSJIFabJ
HQL6MfZD8jyycW3n7qJvnumfl/3iM/OlYYotPDvEzIDr4MWz+a24C/sBqnQW1ceiZg3/i4g1ibbY
/UzAzR6Ab9J1JkJfvq69LbNS6GmoH4jiE1eIsJQF8P0G+P/7/IPF+8rUKeS/h3xceZ/dqRDvpR9t
vBV9PQHLu/fSyHmPe9mtfdbEAosz3MFn2Fgc5aPWIns9JiEP0frBowfgQDvxjgH2c2iSTl7yjQKp
SLBtO3A4SnN10Mo/Kr2FB2JefXZm8vn86eTOmHZyWBAFsP3H/ybyVHKo4ahxYzazDOS1wuVkkhNb
pLLfDjVmA0nu3SSi3NL24QRstINl1Ju/D6s5FD2I04zJBpikwcyPNmHl9lDD/LvgzEwOFiR/vk36
4tJxrDsj7DP/TGY0ofos4H1CC+QoB4byuQfqO5JaVI2G3EAwRhjOdXG7UHnGf9GpuyvHQk55i55+
d0967aEqCRtqFMHgp+Jv+wpi/JZliVWRpVRtn61zboysZmVQrgE/EOX/u21e363LydR2UwmygxU3
Y9yx8sl2FZLcgMlIKz2Ygbi2PdJk3hMiOVKGc7+UGf2p7p0XAj/hHlNcBxs0EZJL3xfF4bRBC2kR
jJAwiKU+GUkDgoCUyWgUXWORRI3gfE3GMQwzPMSt83f2E2fSUAyt7fa0SC3jyKqks56JlwL3wmzH
hUqgGqjU2u9uHnd9yVrc7UY87nY45id26Km6pF/c0DNEk+O7cR81zfKYmyq2gz6F74s2UcCpMamv
DqiJdP3Xg1SfeZYnMcEgP8LK0ND7SsIQwip5NWVjrLe5j4HQfhnOD6v/IO8l6dDM5LC8y3Q727Hm
YwB/JwlID26hlVtg4GOHag8N+fsTCcqt/hZJ/In2Ylnar/C1Y1MFWMxAztwJwdadWoWjEFmuKA+x
1GtRkR95i2K0x6vP+QVn54v/tNKxexTEccY5WITq1S1L0wGF0/7JuLsHtaI4ZPCKYTWHy9QpwC6B
M3jSop0r8fjPdHTHOs5ODmHNGjX59UyU8a8Sf5/W8o6/xYU6K9uVmCXa6EuLS4yewvH+8Q37XGzb
CeU0H65k4TCBS7V9w2O3B8/WE0+sM0d4tXlg4svr4F57eOx0jUmsVQ43PwxMSEgNCstuy3g9o9RG
xwjQCVmSp7IHU6qvNNQBQX5aDLjv0/SZZeF89tCDxtGlRHHp7HDnxenYrULBUTA5nJV+hWb+mdgz
hBbnGrGjoDFmX6fJn9D1m+RUs1bXubddLBjWRci0NAibn9fn73UXQCfW9u0AIC615DthzbyEcghj
FtyIF8dHHHw0HWnTWP3IMHyqqdO7pMvFemjGxWgljGD0CUBKZ/0any3H2m+on5gAHXRYDxl6c20t
UfxpOzdEBYnbZY9PK/l/yO/NqWbRbmmDsTcfvjeMexSEN1q9+ieQwbeLhxy832s/NNqiNaXL6yHw
85OxlOKPumHfrPw183YNOZwoI8d+tCjwwNTI7TY+vQE9yQCCXLqyyb7QwHHBVc8MXAEEwaCKasJ3
dBhKDeyRzCS8pdsTiOIp0RJhw6bQC8XozLi83JEzoR21PwJXTQO97db8YcMDHvXht+07wysGJsUE
S1WQW6nJ4hccLPbfiTYOUJ4shpEXwtKOaeM3lVhHYd8gVwEgJ1JJHmsUKK2alHEvOCZM1VaLHK5z
Vudc0MY9WJ/zlXZnbsv/aY39cY3c5CVKO0VmNivFtwzMO407DfPi9on5hrCGtbHALk1tvY6k49yX
oZcqKQt3tBce+FnyrA25JI4eRUmZ6RLB9Q+BmCUVo+u1fAPzJPzFhVuh3D2lhT7vuol/RMW0Bm+i
42hOiRMwlgoYOyp7jz60TVUFm8SjHbDVkX+hPEZ2jSqv/qr5lkb6v6qknpCOKZx/jV67rFc4dUSe
52gkLpKpbk6aLIGBbOKYogHqqMV6+iy4EAzWa+z67V7lgj0ukst10edgvOhi7NTUms+YFFjxMSVk
APySrpM89bbSPm8gFjWVIF0X/mrG6f8aQgov6xjATu/RKByMlXJbpUXeI64kwBYg8uo/phSUqQwP
ma9sxiEGbHHQJFRG5PPDzPi4RDDCEROBQNTA2jPjRUzxQXwH8htqMjvBoniIzJH5cd2/LCdfqLDc
RnxImC0aVnpiQ9gzdi7K/T+gnR+tcUMJ+fSTuVsh4Nsuopdr9JA7ovFq8l/heRLxJEUutPLCDOqa
qXoQwlvsxC3x9vGR2DVcDnvnEAULELCdY8g1l6yVuVVfx41v3imAeX+guSmPp90Zr3rsFt7fLAcz
xoUG3jhbRu5WF79+qqmNogc58bFxlpKq08jmDmE+lBFvp1RTgzn0o07njAZuifGky+OT3cjF1xBA
syoW40psb6qGYry5RojGWPBl2WEiksjQPPxzwOQk/a1/SF2WmKBURqVVPspcKYRIjaF3iA+zrdpn
XLFAnib2o3CIq5l0vf4fFEUW0CQlHERIoEFBjRsDV2zGK3p8MUoUK191S8EDg2pqknuPGpE33Len
PNfeJGhQ/w3T2w6y8OUttk8DDx+j905ybg8GCL9EQqGQBPh+xeC/03WUFa97euDcENygEvq7y56b
1nUFvoqAsrN0N0lD/Vcus/I9hSURtrSAYzRRPvU50IEqzVm6UTzblWqpKVWkcbj0E4r62Ug8r+n2
wmMX13s/iEhmpfYxHqH3c8u1Vh9SGGd95tx7wu0KI1aFKCegk2Wc7uqrGo+7+fw3CzTEVvdn3pf2
MzhvaIjpAe0kLtrHeR8FpvqZBjHEcy0YYarcpCUCAM6mpPwoqN1f+rY+fECFZqswXoI6KOFP6n6S
4F/uTAxMLNPtrqWXZ2v9RC2YW07BK9qdyE6r3CGM/nt8dk7R3Y6wA5Kbr+7CqASNqTwSUKAS2/0b
S/p+25yFPqi6kDDpJlGNsXMGvRB5wBY+fiKVkwI2f1iN4EwXNL3ZHSpW2cZeV1gY/3551sKrPax0
FV7XfTi+drOGhSs+Zw1FO/ttgs4NWxAsiDQzKVw6MmPi7wdNKB2m9+5LGxg/tPZSwpoIyr2Ww0fF
w+9rx8J44/ALYsj/dkmo9sbfIOhTC/fHQDX4wdA8rK+fdLHtrzDY2UBKdUdivPbTJbY/ZwjSUJ6W
zgDNX7joI6jH5P6uVDs4KAX/IOShM4q2QR61r2W8ARwlIyw3ckxafxjkIjYpGpOhdxrlOHvbdWyQ
53oK8PjkscEFz4W1aEhK83vtYc27fhfIZb/XSB9ge7jes/BEsw+7z5uxv/OSFaq7pFn2+fRBc7pe
GXNU3su6rzQR3g0m0wx9qESIyu7/ws/druIlNQbL8EDT3kN5uJuGdof1FORhx02O78+DJ3A63XwB
JQ8jPojzVuuilaYhzEckAjFxf8JbTOzJWnw7U08YQ/J2MZNYqF+mhmj6CMb8Uc3MutWIfYBzLLwB
PFGm2yuB596yjKF3txEbgDb4lWWCw2J1xIehc7W4mbyP83Km0sBvP9IrcpgY1mRuL6RRjUyrVvxV
qZSumNGNJSOixNpWGLRYYC4xu468tFbh+/SYYRAN/Dg0x6DgMyIcEWIAIkdRCTEaKBHexXIvuw6/
eRvVcDhAlanoZ8lJfJHepxYDF48sGaiYSfK4hZoefEFydfrHcdVNWN9q8cjsm4BoeuQDrP9Yv2YI
kus61/SKLwLUyeN8izjhAQYbhX1dht/TXJ7Mjkjv1Mcbuocou9bsIaqd7M689Iqfzoj4buqz+gep
v3bRpfNGS1TOdvQKGIbfHaBYMFUGoh0uqA3WV8+r2frH8lXgcpO1nhaudxzePIDg4TINZPNgcMgp
mPh9HwOAKA+Ry4ZTVuWBk6U89bQvbIHbZ7fmAZJgjwa1MYlGY+sYQepfbnUnnxCfqdZZgpmOPZ2c
HPH4kMnGvbLzZeDQ+/sbwIreKL3DXSFc4btGvI4RkEvq+PhrfQ/3UDKx07E7tqH/QNyUukedEmjX
EjUVVqd0MP10NGLP49Law9DTJjz4EkSpmrrr4I/1HEANcnyAzbBfdkdHaGid1Pv4Rc6pC++q42Vx
I75wDAEQxcZQbn6TyYonxOmeIZ8hh3D8aPzHl7z125sha4zu3HcV/GrJ/0cTKzsvLgYOmOkrtGX6
aole2hV0tbPmUbQ///XoXg/eSurqo0k0UxqHdtdZi5F+/qiRal3turI9OnJaV3JoBQH70q/aqRWw
Z917o16svggfAY4OeC++g/9q7zKRRfs1/yYceatm0i3tUNp+jr/SPJsNNGox4LePM/AVfKEIfzcg
hVEEErGs6DFMjIDdXzb3iIMK8B0n4k2/JUSLncW5YN8elKOZeaglIkmWmqBlBIpa9Nk/6NMR4Msp
tRTPx7IrkmpSgKDPu/dEk5mb+xoQAYEWd7vyKoyKQkvpSyU5Il1Jl4Oyroakxc/WfQfLhmsrJzvk
eOalzv9BlBuWk3hNjBU0yqF3ummz9rnmip/2Fy8RZGJuQ9ZUiTao/LrADDcPs6LDdKkRcdnAUYu6
9umaWg/Szvpblxg4h3qpy5Hx01sNYZosetBsLYjaYVXcqUhbB8GHTOD+Xjqg1Rof4iUPWHvduXWa
GwOGxUrXTnswRPpglI+msOSwURjGI6A/iMyDFyc/C9ugRGFzhHqkhxTVwabzreEaJyxvjUBoUn9h
naOxK2gqXtRQcTe4eeCoJAwoQrEl8JATDH82CNwkK5V8aWdrs4zGL9INZyig1D6KUzIMxZZhl+Zs
pgY9podjDuW6lGUv78Wg3BmI060AndbAdD/javwknY7rwHA71aZ82O8ZHY9RGi7/rEE5wka4v49p
oWcOLwhaznxA8i3DADWC/6zWxlNgN5zHegFbeklTAQtt6/tt3ArgkJiXEFYtWiaQNlP81U8yqbxc
XCmt4LqMl9TQPTHhNjBsC93Go+Yb32tJ1ySij9OdnRFEzJ4Us6cgJXSgR+ocZBHj2D/B6/fzCwRA
x5x/zgTI6ZGxRh8zpZEwovIkA7tRyw/CqrlVdi0UTbOrbPXcTb6hmUwikL5NAeqDn52zemd+4rJg
iY7Pb5j3FxnXl7RiD+X40GhLXKmPfL1GFC6vM3pfxuzVb/LveMstnyILJBRpwRFhcNELYyszAv+7
JHPfiEMUzj+198IWKFgkPXmEeoe5ySdOJTCA+pM+dv0Lz6IvPM4/UlcPYKP5LoWluaUj7lKaz7Cw
tw+ZRl/MKeo6sZX2LimXBrKrdxplda9VALyVq7WTaXz9t+PorLiuymwaOF9u3B1aOjlzwqgj0Njq
sukbc/uXOJd+axuqYXuX+uc7tTTqKJkWMWhV7f8kKG95BeBsk4vVE1pDrCBYlPz1xbokoRryz2Ld
ZHAU7YbVyi81v178wqiAmLypDbBEwRpm3wKmhC2AEFNVZyHEimUdrPH2r4g2HGhqSqVV2NEgUxcl
ivuKasGkwVtNL0PytJQGVDuh4eN2+oORlzqSXGjDYvDsI8hXNoqLzmQKtbfa6U1HweTydR6F0bE7
wJh0gxiQIELnM/+vky8XnmY3nxuGOPJ8goz+yE6nYt42JDzw3yMDsRZP3N+1T+aqnIt0UEKD+LpP
CqGXqNFIi7PHW38rtugNmIbsdOQIOUtuQVN7dtKgf3uqof5+dqsvKrTH5TVckhBH1oUJV7XkK0Cv
oF4hMA9RMmiYMW6h24I7pWs/DUL5LpysSK8U+WtShDITNu4BrqgFR+AuNRFp5kEU6WdsiFZ22SFV
v0s7Xxm6bea7WYp6iMm8rfbH3t0Qfj2oJoShFhlRJUuvhsPxTH2AmgUjNxTXKFTfCXTZeJTcDcZ3
S0SIwSubaoH0rjn6Xr5R1b10pgEKyND5WjW1wyRbpUfDYNG7D+hHcKluuAfCX4NvgXStHCLasYL1
bfXuAoa5fZwiILrTt37Q0TJXBd7DjPNrPGPezfZPEMXaivjdyrLx4+wbZbHxZa7gIBPsS/HGhwDg
66muUJqDcWcKDEknDvbHDkx44vtjlpWNe9hc1CNEamWaBd7pzU0YKUqBBRGWuSkLY4jR4Uvyr85c
ty4B7aUwlGNx7VFr7pW45JnIR/dKlvOTJNPE6IcsFoR9IIXPk2nnOnk6OWwSW4xWXlh3dReFKypV
UuUA9ve+j0xHKh6dwDpfHWHYJ3Xsxjy3pyESFBmo+ibybe3sZxt45iOhGuvZNCuec7+Xm4FV/XHy
rV4B7675eSzZOGYjz4I8IzbEvtnjGOJ9phy0QnrCPqzM5S9IuDIf9kYdk+7jTqFdV3BUsHU9wqnx
DQi2uTVulgKcGL9FbmpdXA/5pto7b+MwaW1biOZFuKO25VUoxtnnt2fr2+Z8Yrlhe+aIMuAStyOy
/YlbWFcNymFryu065PBM2KGQ15t17h+2igJ1WQ+cgV927bKZJkUnfdNyTf32LhcHCywnGseLD9Fu
CoYwa3js40JzU27HlqOYkjgBkE06qb7aZOulZdgPkOefnYay/ylqxvW9eHoN7Hpy/3/6aYvPw0Eu
UYKALi/lrIjbEACcpB94NoFC7PU/6YM5Cwf4LzQZeLs2+7IXhbE+LClzNcImC7j92k/1+q182sFm
gbPaOVEJ3+dpOYGfFyZk2KkOErQ0BXoLTJDOPREfUbHOBXaXr4s2Fe7a3oG8BYjjF3QrrmLWRelg
oX/xfVntNCZt6ZIhWDjgj9ERigCOPKMMIf2hlVhsGr6IZcFlorj8R8PtGZSSsna1p6wJ53lVtm7J
pExRkUGqbZxB+T9/gKAOgHvWT8c4JCitH3IG2lSmj7NXGaU3gcYsN31EQtGTyTTVATmC6MmT4zr4
8dPHOJBWx99WX+weUghT/by9CXZblBY7zyhYXs1nEb6vRtfINe5AASrvmAJNQp0JwLH5dawDYe1s
yj5E6EyFtj89wa4JXEsKXx6z4UJQOil2fl1DSTJx9CtLhFpm7oV97ygGiQIEe46weHsCdx4/wpnk
2w2MuD5FLkgp6OOo6QK6keKNXV37C7hbCZps6bcTNeYMc6tpHNDvPZWoLFj3RZYovPLQs9JWnzIz
/OkOqScTLJRf8MPlqevo6gqcAkV2JGcZw1x3QC7FYqmm9Knxx06bq8B9WtoIHBezUwZNJDYfZ39u
z/DonvE/7W+Scz0DKYcVmtMNbR3SiwnwI/29MJwL9+2wOW2//taXI0n2NbYs7jT21qgiAjh3AauC
2PQTI7bF0WPlqwPBRRed7fP9hMT1IQHamiWZtbyKSz1iq+yZGE0X/HF0p1ii9L49PDTYVo4SWht8
OCVh7voL3Q5S7pUe4aXGEuHvCYUNmq+nv1kXODVPT/KcP6tIeWUkK+RFVmsZnJMH1LA7ON874hSb
NX7yUNKYO19fZdX5Bm1vVaeJcT1LqbZeMI+f3NWtivZy6XtSnQvob/71BXKFjaoFtDvRNMnQRqGB
LBIFZafRkJPTVO2ekvAz2t1+SBIwNfLIIJuzgIBAq1Tnho1JmaAPF7fMFZami/1v4IcRw9z5rO+Q
QfDh/byMai502uABO/aNulsWx6xK54bZEVPiin4rsQfAVWX1abaGmN/DTL6mumEuKM+NHRNvI9Sp
94o+zDF1Cya7qWkX/qFY/Gnl5VZAxSYdiaFXqCrkshEFlR1/0Ev5gVT/rcpHWYrNxxxhbyy+7jLB
7kuJKJYO14FjIQQ41rUkUCJ6D8Wn7etF5hpnpsg2/jZY2TfIRd0g0CdIp7NGwbgxioQaIJJgzYyv
E0+FNkxIO8nXjHZ2UH440N9FxM0caffX7qL5dhpRENlqeJG1f7gEjKCbxhNOD+3xPdGkhxfirfcT
RxLQQLI0UInUNqxqeddelGzWdxnNVPKQPWH5Qz5nZ1789MxBHUC6StUjAJ5D7ZLoUbM3iDaRRxac
OHWbt+Kec8DbmimmNJ3k4WgzHcq/ia1rqPLw9lIaHfXKlC8TU22mdcBZ0FfRx0gM1dLy11Cmhmpu
mrWstPK5kkCtfjCq2nNXe2ZjZDzFxtP0ceovN2TcKctZXw8p6UEja+PbSPZWqc9D5I+M+ZC6ulWr
nX6fNXuW3p5zA8Lqw60Gcw4Wpb9NDWNPBIwHhqUZVqLsUohQqquW8IxVxee1hnIWwrkt7b6OKtFu
uS2KQtRdtMKwJLG0SQH5mncKj8hfvvt7gUV9FjvYRRB2fFgTp2++/o7doE9RrTpCLRX3OJ6XUeJb
WD9R+OeULgdgSliS+l/RAhbDSj9ZPVGHiJGtJ14sYbNSJnvAfsPbHgn/sLUh345QKdK9lbAGLxN6
FqoDYjrfCoFnvtj5NmwEwCtFxzRzWSKApHNdInwL1+npU19RLG1LjHA7YRzgdUA/JfrunXUG51Jj
M84F+Zgi8TvFLYfaUpLBOu8rvwGChprdiE1dtl+muZwntkPmo3dXmljWo+fTrG8DbHOkgvm7VJm/
Cywqe1LnIvDYlykKfip/3PcDNfrTCxrWl9ykj8WqLDxlTHBq7NIOyZmUY6mDuGrev0Lp3zw9dYKl
JMfiOapuiqWgEW5b64S3UTJZ1Qpuhfq6mJOIACaFki7FI+9/83UZL9VdTPI1h7ZPkwzaccCaq7Au
25WlIjtFXVIGry7qiG1q9WU4uvFRMPon8txlDTk624VEz14IPKGE34yuuzV6zWoj4Mpgt39wVmx9
YN0uMynyiGrAS6+MGmAw+L8gWAHTT0t9yPlnqJbXjtyu3+IW908Ao4vzf1pCkAEVsRs3qNUT8J2u
K0vn42xvmERuJI9G5vgMqK6Fdb4a4fcsrolo8vl/lxph7DVuHFEEM4NIEKmcUGb+kLFH9UkckNi1
VBGErXxl/OUesdEGbp988qHh4COf8qXV5+ssAUWsYw1a5RErJI7CzosQV8cKNlpCrCaMcYMedL8Z
A5ZNXxqwVLEfg4HsWQNx7y/k6fFYt92FHOA0SQcStTWHlcGBtm+yit4C+Dz/JL1rg+0pGtuzPdv7
Omyf89yzvXEY83BgsuInDu6RlROPAcQfc61ALe0qFAOrtrR/N91HrmW7Xy4UxzKIDsVeTjRTL+ul
O5o9M7HXVqe8vbPs0mK8Et/vKxs3FwHOvIrcJdgA0TCGAD+8OsvHw2OymqrduQa0XTTnQXU4xw5c
+hYAzA/fUnn9o8HD/pv80aP+N7qNueSL8LOtO8K0x3A0+7LplE4I+Xi21yeSVE9mJ5ol8NPmyYXz
aU1UH5TU6w8JbkLroq1qzkcbmRJUV42U5+2zKDrHY7IxYDiZ8UUs8UbdnFYx8LNeSn/ROo8Rm6xJ
r31cCzErb5NpbTQh1gOz5yhI8kD24xG5BBFHSGVodVCXD76fI2iPf3zRz8DktGJq+BcF3WNI+kt8
BGQ6NjSGRQI3J8qU3wL4cSSyc/Wl3Uc3CSkwlf66Kkz+2DaEvUGJLkI+E6cvgC/Qa0lwM+uDr7nv
nvLKZBAVRbdEfD0F6igpXXfPxvNcAK4OWOXxEGh6/hUUvb3Ww8tjAT263BYw2XQzJsrXPcrx8bM+
bNVrXHXvT70KX4PxWsWCaHElCpLZj4KFt3RRDcMYmVIaKIjhKuvdkKHQamRUslA0pe1vPyYjZBlz
KbOaW26eLrp0C8/1GmioUHYHHZK5L98MtsCv24AnfD9pmXHx2YX2o6clJSXmx6expUKtKc8Wn+z3
Ad/u3vmxBkYgzlLsKtBFxgNyLEgP3QWBL6rV1W9d2Dl3pH6fThIWwRkJJh3I0o/Wu2y+D9Yx8jp7
grUNpj52Xilzgps8Xsb6XWoTbP3WvJIO3v2WyD7f/E4ObLs3dJN7/vZlh4TzsW2A5r1IXna2d6tq
rlXPrAbvL5FZZHHcahavtreiDSOwPEpIv1xymjgzZphAX1Af6ysrtWkOP6753dp8S9HdDzJQonu4
4c8RYn5VLAwO3OD1Y3w+sWUuw2hOu+WfGaBmqKHL2AoSg8cwYELxhOXQmEiKjIQmNi8GoqeT4TeV
A7UTbtcY43mbm+djzUZ1kNkBdRo2Wa5sIBZHW+P4yU1Jo3PMzfBDl6d6YXKgIl3NrSg5Ogvlk5WG
6LRFlgjf9yDd4ZfHoPXiTfeu7m4mu0OtWdu1pu8VTxG7zYjFlvLGsctJoFaiB/Q/BypuESNXPT2y
NhnLNFiTiKP19VdSShXcz4PyHn3kFWNx6ACC2BYDOgzD/frtu9aOyMs0dUmpFNGNwEmnmlltL6mf
L8sF1r+ACIBErAMu/H4b/rDsrGf1XD+3XGD7d78wJc8d2bLp6mz8GmdF8l0Pn8XqNl5BxrHauq8R
CBuvHkIqZTMRpS6oIg8w5IIWhSG6zODGjKfBDrrRP03G9Cv/4iQ9HSsBxngAqYp1BoUKVVG2/bWA
+OfQQO72iB3ZeLTaiN3N7RIa05z8TqW6sr/4YqbPdFOx1fEFJBvqNGeecoOKbooow+entDWDNkc4
3c7Z7WMcbH0IcYju0ykxB1/dh0dQmw6btUkBHijyW+9PrCO6J3bdVREWBAxkOU1A60mRhZsKt/XG
vJQxFCZ7UvaHlhww3R2L4CuuOiMPFVW7ptMndfrpzny1KuLBfz5xIQOOTREkfHO/hLgQRMCC7RAX
4SlvsC4zriGNB/uNUU/SzqpIqZ6jh6EJu9IRnq1ju0hsJpfftmh9TtPUHkxoyv9NOuleK00Nl90b
nudoKzE0AVJ9nC2npcUksiCn/niVWKSMDXzeT3O0j/K+kw9TXKwHO3XalEUcz+gM1LQWOHJ7qIsC
bXpTMtiWihM4q0kJsU8LIPZR5oBK+NrknTSL8T+JFotSBj4HCr2B+ztX4swdNgS6h9Ixx+HmLhrJ
uN6TveHOFIpd+kOuwNZqqyl6RfViyc14lUSxZaVkWpHMBF8cH8WYy6/ndnjgmHZPW59i9vu1Ek2X
aT+gIYpnmkeJKt5I56oMQ8A28XfZwk26COQao/QWj+EjbNj8XvFENQ4931EzfAB9PXphdVzJaQbv
wCiWvylBpiDVFW685iPQPC595nwPov4ev9h+70pC7bxi7N2u+3I7t6R3387b3IhhcwG0EZ1Z0gFh
eJx3h3ptk3gdTbSevy95Y7W959L/KfUAIQUOEccfSvOyyoFLsEyfgyqBlQtEvGl3Dvvpue324zQ1
LOh5PDyhq0GsRUir4Yo5SUmTlkGMoDnA4ZWjgUAEA637cxtdzA2HNubW8VuvSY7fquFG1lv3w8q1
GqoM8DB42pLNnALkWpbINV/gvZlgSnC7b0rswbLuxy86i7Ys9i422GbRFbfZ+4OW2RTetaYGZ8L2
ZGYHGVfGeVl5QFKYU6eMpOlD3Vpdr6yjW2foSULQYomoifFAXG1K/cpB9i7E5Nza7KYKSq/lStR1
XHpw9Aw0ATgev13Fa2A+/9kMyRlokqdNpuEEJfgpPGBvJHsq8JGvhFC13eIljpl7RDBSQTwGSR7p
w2dwY5+QjBwKMtXJxM/Ve23bJV+qQH4ciFSTT4mQS+dSm6yoAopPVS9/4TP8r1PjxoYRo4qs5T01
NGIxypjdUBwNTEWeJe3WHAIOWUIwy8OojZGGE1b2UFLjxuALronuu+MU9QkVa7Kjf86GhMWjRhMq
YjW5DvOpH7rMWWXqrArfJxnPIACgoxXukPO81YwMeT/kCcJyCU7sMgk+52YLYDrs1p92avTqSDJR
2a28ZSxR984ZZAbH6OwT8JpPKhdXXQrxWOjuU91GfZzD/ynlFYcFXAIA0+Q+ASWzgdmtJlSqNecw
CEkMCm2v1A8IDVDG2SYspXI+1HBsjE2PepzkvJ9HUxOI4WPjn3z2d13mg7zPqBzic8f5QMHyqioo
A3/OhyA+xU9BDwZfB/vl7WcIHXlMp2NAuW7R6KtN0xf9Wi/D9/QsIruhbJxBnZO0mhqzDi//HqLt
t3AZUghcEUPspsKL26yXUSNHnkYOGERHc+jr2J9to7kQfC0geoE3ihy3GiooDwhbGM9ApLdQosQR
u4Kita/agJO9LkYAfVRkjBZ+Z/U/5uNlVw+D+nzRDtrrRXf37hsbv7BBhLvc81ijf/uAVIp+XKxj
+0eGgpvxMcymPCj7/rY7Tzhj1MwE5A+4UNZrvIpknRkFqFq1CU7yQoGle9W2D6N3+5oy3fvZS0Ze
G1w9N2znh7rgITLkPtc+trRbdrR7UdI+JeeKeD4/k3RHHuzRpORUI+V0GfO0425vOihWUKwo6lYr
Mo8GhDzYa+9Q4Kns7STqs8w57ssw8QUIGydvgiN7japzGqAy91B6CTeXCa+eEL9STzyftGSt9ouB
x82AUlT2imqU7YdRTvYHSf8A0Tcn6sDLbGwOQhyGGTbsSBJJ3NZKBYUbe8fCWpBEaYyb8Unelm2I
T/IXDKYg4MFAmZ9y9oJ4Y7pj6tiAmq0AnEJUKGHyIbIA8PIZU0bw1HocdqulG03q34+HMXgx3z2n
j29lBCJ6VJMFEZ03dBofU+9GNxoaOns1s8g4QWTNPFLAerHbFxu572APUcYlLm94+6UAB1jYEuBF
knyIFuNwi43rO6sEhSTKCEz1ZiaG7ccxlf+LBZNr+ZfSUNtqHezFu9m+dBDG+BUSGz8g+giboeHN
Vy5puZyvT8otPrp/TLEpRcLavWE8I9C0GnY+XT5JRjV8I5LsV0eVQ+5SQMRIuo7W/L/Z8nadfyQW
/UfGauVFowdBFMO5qWjqL7J8DAlDDpnfmdYI7eO6z7CIGYb/0KlDZOcyAzaIVoWzJf8DWQLMr3AA
UIKnvFUySc1JAg+J0LOo02lUSQZsDIyLHUN9Plt/ui6lpZWpPm25fPBnxwCNJVHJocx+U5rTH38/
yY+SshL4D+9ybp1ncoOREQbg2mdY70YhwsOHH3JHTEOCWZSZgD4CdLl8Xh1h7daOoEHXhMJnxfiR
E2vo7QWYJhhAV1vpfcuprHsVSdeFqKi+TJaqxFw0BQkro8pfPpvXY34jKdC9t0hJ+8tmWRRW+fbe
sci1B1qnjguwAbVPobeA+/NP+3x4wksZiWQ7oMvHv2TqMAFsdeT66iLTb6slBfFRo5zHxz36TmCg
BsP2XZ9Nyos0aevJ8QUzBW81kHKH0WybN17AUL10AuV7knne3199ypEgPvjtZkk/eh2YnWsNPvdQ
gIW6wGmtQiZmt1Kb3Un0elbCzrk1tqKA0W9XLdNhWMHDli7Lj06NbE4hKpo99jQpAMy6nd3HZudf
qEwnYMFwUWIlynoDlVR53nf2hKyIgdLp+bg9O7U9yfVn0hZQreX0+OnTTyowTgdAZI+lDuTmIndN
oeJo3usR13UaKu1ceygnWEDO2TzoEvukKI0ss/h3dM0Q2xCs3953FzvCS5HKXom1XCvNJ8UXHzk3
50ThKnpXgHRQx6ha5MbicfL7J+T3w1yTq63evLv71+60/fFUc1Qkkc2ZuEng5I2U9+qPTE4bxs1O
ACyynGttPX1MZ+W8WLljf4MmztfFg/PvIO4mKQdpQN3dBYs0tRelC/rR8Du4mzHdCPQ3moLB8SX0
vOCllGNrYiuPD+StFjyAq/haKcLzu07c6BcwjfCc+GtUoZzq6JiJubpGgdXy7T0kT8OUeWhjs6Wn
h/sJ7S363I/ow0tXk0LEIw0w4ybN922jkQ8e2RWRUFl6TQ3wAnNHBWEKXjhRLyjiCyCQO33WGmYi
7nVO2nTfbNPHHn7uiSBGFrytwqooa6SvQWEjKjUK8jVSkElNgoF8W0oxMwtY7oG9GmAxUKWhhghl
mZYqTYuIXU69eATH2in5Zdq+FLikIin4V8AN/pUWmnpgHExft5nq3q10g3gFFYlx5OuI9v+eZgIu
MebTlVT4asW3dHa2Ze3BnzhQpZhmSEj8OomtyRvyODyqhrUgQ7LUU/TWWRmE32fPzd1jrVwQHOQf
dgFaHfd+cFSmVeyC9DKTBw7lMoKG8LbNfw5rPkAGVmxsXwOXe6j2ddTu7rzGczucJ4VLRTd/Pop9
kkMgXP0PdsetMsiUx15DnCopgamiWyc7jS3oEHKVVxv9ijsCdS309/1rjhtoJg7WrJgIarK1pA1M
+leZ6sXr4qFfHk0pGReOrGZe5iansAJM3DgljkiYsCLSc9QYka2PfJxB/Nw9VZX2FwbIPVDq2o/9
yQzfFKtCUNn5yL+uZgDNaBVFLTHVt3QPCE+LcOrSXZheliVRhdR6VagpFL0Z7BZcdMwa5I1igYgG
5f0KG/0CjiT8svSda67EKcJPJ3n2R9WbcnJexP1g2roLt2hOormNqalALO3Xmy1+s01a3ohWdkR5
KCI+7CtDbfO9oNFLl9PKZIM0E2ZxOrfZ41yVL/CJAPe97kwND2CJwezsi5mW2zttsRNpRjHiEDYI
kmrO1eRrPDW55ArO4wwBgWu8ZPKU9JwMQSfzSbWR5p027j2mibs9jR1DR4Hx3xsq4UqKRHQR6iOM
ifABqUjPN9zMWqEuZ34IdV4+d2EhzUVRcQJirDjQgaD9D5yuaL76gFJqPuL4KD7Dt0obmg/dTftL
/0Ez73Lm4iTWy4Rtjtx0C/qg1sPChshmp9/PbC+T5Pd8oXPjQKhuOybJbjEBdDouPPbNYuSzop3s
bn9c8Izx6Dp7+ekhMuEXzPcQiV2TFMX9WUjMI2PIV4uW5ZyBkCOwLa+ihnraz+saMNb85cLvkX5N
kFGZhBSEkDdhjFnBoLStWawSAdbTOv8OCg7zoE73RwrNoahwX9YxrAeKsQfXu3tlPY8bzDnVWE5x
R54+O7NQGawY3kFXcfkhl/DCLnZ8y2XGaPiGKkRG46dZC5oxvuxPLtCMblBtWfbfk8W7EXV4r6Cm
B7TrSNJlIsmSKBnevy4Swc/k8T0RnZpkEfSnlCuXbB4X/IMablNaOjc/1sySN5FTpF5njbT5eW4T
Zn4EHQMTFAzpXdRA8vR0cn5JXEUj81882qRglVUc+WWlr3NpdNAC1CslgKJu/BROqZbGCDGP5eSx
+4w50FJ5n4TLJ9nhzKwj3Chvtjc8P3MC+IgNGA3hMCFwOXE00vtJiBEmVTKZIjCCxdWgtoRqSSOW
08w8jeYV3tccp3QMcUvux/9vv9wGc1c1frrem49ttxvdNv0aTPPKFUBN0Wa4vACPgfXwkACPc6vz
K5CQOfPczCIH9WM0CPboyLJjnHsdZkgnwC4YBJ0f6qDkLy6YEtDqMvxG3BH6D6SRsmB7zf45MjnH
g+1dPVPz/gMW+a7aU28umkbfhyUWBAsc20ku+lBMIVQNyZ4wbm0Jk4ByaaQLdz080mjSa2V7qsMV
DeaMo2pWupqm6JeBbsof9Cd5birKj57Elb9gG9TTP1KKYIGegrRUVKZ+IeaqhxzwAR4+ws5CBTpI
79DySWrhk6h1qV9YcbmZtOXPWe0m2TJQriUPB/Sn+nYzn4htsyxLUOZC1BDFnJnSH1DsE23hg2ov
AXM5F1WfYfA34NHg+9azvj3UYRQdD8aIgDBgvow8NVg6mmUBwVJpfqCo5hMJJuJnBAW6fsL7bj4e
6tVXdmPo6WI5YZ0QorLoo1F/kqkblaLa1I6NhoobzjBAh4LU9pZC7BJzEU7cJXEhDsd/TejbO6J0
VNTWOsXtqa7+mM9Q6ClS0+cMXrvN+495ddbdzl+B+u5kbkmYZYNwuW0Usvprpu5H3CA3tUng8CFn
EcKbbmECZCAbqJXqnX1yS1HGqDVzHjJFoFkrfuu+h2loPkv+gsMgfj2CbtMVRFNs/MnbE5O3EMeU
lkRDBn/D9H4NbBUG2R0grjO4zt1dVpJ2kF+z8qiAxyRO3tXwb8VEiZAZ47aKvim2wO54651L8ybW
Ppe9iHpAi5SmjTV2vtI8U0sxHImphSlJ39uykBMYcEPgqFHvgja4DGlwDW1COBtg+lGI8K4zfiUn
TFV8hDrQooulx3RpVrU5rh2aWNfAZ686ATvtGR9SYshDrYbNkEuL7AIH+JGE3L11fSI0hlNrq+DJ
qIxQ2SrsQuY5lsifrjTYCj2l/dwdEyeWmMzxp5Go2RFwI+yATmUC6nbl2j1YRcCL6aJS8go+NmWB
XWfEsTN4AgVLJj2gclQYnQTz4mHyJkRyO+7ynysGFwRx6zB+YvBg8KS3QLuTk+RZD+nVGBt1Pa+S
675+6xFiqpxcbTC394YaBl5oQJjSs4oNxQMar6QygzFn2Me2QqQBxgU3QTTaS6rbC6nzfM4/oUG6
EtYOvSNnKp4M+ErW65WVeuI0IrjiNe8GamTZvf64/US8jUzMRlVeZy86PzQJ4j4Snoh9iAU1lVNm
DlTNDoMSOpeAL8q4au/XYFt2p5jfH/pW3xqVTAdu5RdW+ihTGWKByeLunrlSN9jsISku8JPrS+zZ
UL15BWS23gdyNS5LKwubVMCqhP7Ld9jn81GCy6MOa18RVCVkO0VId3xaWJYQY6R6+1uNqqiS8kWv
c6ctrXKvH56G4ScQO/7UhOzspPSja9SII4em5+Za7KAONXejGmFxWFrZqW5xiPfDFJ2fPnIAclBg
kxJ5n0j8pQ65Nf3wKKMDi/miUWCE8RWhlmKH+ATjYxNtols1i5GNgv7M5/kno1P4RR66Mc0QwLGo
mjPD8pxQ82BX3CRLYm91t8TRXIQM+PVC+Htf60L3304lxfVI9sQmbaasohBJAyw5fkqZBKDZEuXW
r7Q/o74bLsG9ckpBGuhVnG4WFSZ43ufWEmHE9RZCEkQF4R00Gqcy3RiVoANu1IUFocYyjGkmvOn2
6lasGpFkR5UpgykL5c0mS/7xJdqnF5rBMk5wp/PI+/Ctyp2NRWy468SMjy2H0KSnM2ubPfBvtHM4
5JqkEKgab2GOtMdFibqgEHLPsHMfLXy6Z6/YzUzoKh+VqMXaD1ZnRf2N9p9rK5U6+IC5yIjKy8Ry
7V8HVKzttH4kLkbK3qG4hkzSBF+A3dBfJxfqJDZdexJRk7JKK3cSCZ7X/301kLfAkdv8ZeavLMTK
nxlaUtCvMCtUaLhmJQ+vJjDUB/2W04mR6ero5Mvgl6f45sJAMu0kQSWG84GO2hwrknsIOftj9qnC
qzizHBJXfiq1X4yOK3RkDXeTKKQCovPzqwI25T3jVE4Yc5nj4skCHsz1AmSkA4X9b27q6TLlpYG+
yz5g0mH+0HZNyWxarePXldkz/LDmAlnV+6KOhRbL/Mqn45Gxw9l3oPjuR1IoNM+VvtcAMWoz57yt
RrOFPJbQwbeAzpFjCH179UutbpFwuGva6APRBQVpwS4rlhzDruNwv/eWsHLiLaMpw/FHVN9LYIVw
phH7Wp932j41EWWmzTuhqm4PIWF1q9RZo3g8p4ylCByHxj1GDqHVhq1BLjibqBTIQtnBvqJ9wdBC
2Om31dVn6eQPUOzu5HlP5AJiB4pA1LEt9s8s+PkSYN59WGBklQRCKXS8AB2gO+bm5FLxFcMDwJ8N
FKaplvwB2hXZENaFlplQwNHOeWb/FMUi1l0X5remKCC7kEbwDZNxmW9cn7uLu2ijXpmeB+0VRsKt
yINaZUqCfV5R+ETr99I1+WMu0VGCh1It7gjn/rpSo/qAYs1GDuVg70MVi5cqhz3RvwiUjqetFiIV
QLdRs9kXWZb3ozN5dKWBHNfuVyF28C7UwKNZX02A41LXIQ3P1ndkgBDxUgpV/aApBoyiax6Ke9BA
+ytB2N+psgaT5BhQIJ1AGOZgQFWGgp1qoMtTOiun0XBoXdeA4mmlipUYViFFScMLT6/XWKT2MOip
NGJFsq7X+zuuKWOOkjYWB0ULT6gVkjwLljvYkIf/psCR+hFjt5PZEgEJVNvLa0llI96drrVbDqIi
HewTI7LqNaSGQMPMNZxq0RtH524kmkQELYqmiskZA9u9vYVJZC3LpPJJ7hTGzoluigynAYRi/9uV
kLdVn55imUXYv4ew5CTwX8VLY3wHhlJuq47u+44O0xWaB+A0kAfUjYtivgOFO0IKVj85M+dqOw8p
bXbz8zsaDMyV6HJWqtfBAAXm6CPPeGAcppSunD6AT18B1ffPX4knyzDD0JXTxpu8yXKuRBir0CMx
4oMOU1JTBydYTcRrdFCSGBKLgx7K0xPs1Pc2oOr/o7ovD/cMlfGp1KNBL8VHYdf1EnPvKsgca/PZ
Oxk/qllHkIxMTU/RkedzvUIj2215tEcIA2lpu9fT3oAPrUwE+F0zoyxMMb9/pg2EQ3oOhWCWos9K
hgsZ0LuSWYXMbmJyscPIB1TXekP70V7FR8Huxz5OpHG1jZLRYyLHnvMFLuwce2l0MDklQ3ADzITM
j1YMnU3mG/l4HVDyZzUKXruSY2yajCM4JJlj8HDWhcaET6L6PiwO5W0N/ZqIECNinUaKxJdgiw5V
MLXb3hsSLVKiy0zo7X5JX+YYL14lzvJN6AD4qgaUc61ZcCUqi1/gX+h7ehl7OQiGSeECmL9/kMpM
H2kMELyCWau0/XHOVkQ4f7kBsCZOvxmtS8MteyHvNkMnS1upqK0OVBPf7Pqpwe5+CxZ8oevvgDVl
YKF+AFw3Re5lLg+ylzo7FSWziXP7SL8fvsMCRG93wYPj2oZsRpwV4PoWfbYlxowFpEtnzH3F6OPM
xD4S5sVr3mWM9EzM91BHx+FeWTpC9W8RT3DZ//ll6YYOcwzblYVGWNpNwUkHrG43qviwbLfJSsHw
L6ABt326B92Z7DpGQLcTIAvBXOGvU1T7pjYnMOqX9sJ7oVcsoiW54bPvSr0+VkOrSvF1DGTZ3q5j
x+s69wI5SRNoL6BktUv5tykedg0IVuw/qOdeqzZU62ijtTx9qvVdMBDAKnAfsdttcQBpll0CqFok
1wTiG497uoxJxTo2EUTpSPo4FX5G1zsXVsa50PWkoOBQFvJHMQkLMIFGgWTMUxeqPN6y0r9zDUh4
M3GJehAMFo8xSEdxc8l8S6LiFhj7YxDad1WD4om+qubB92QFO957fHJHdgPnf3aCJLj1XdNDNxgZ
xBudJyhfW5MDyRnuwzZC+Fm6Y4dE58Qy142o4H44+Isfdun9EFPzOD/wDFVQWiDXi7We0gvIo/cy
Gg1gX1KJtX245ku03So30IqjEshL/gA4hQolIDv+aBTwNZhv7UKg1ItoALQ+TZ4CiEB6c1X4J/BF
53aR5wJIX9c+HJnLu1JcQ1foUfnhUY2xR5pnJQrJyQH20MZRbA41a9N1+6djBFJcJ/cjteqHw/cF
91s4jiUzD7fIt3EGfOseWIrcC4HJS3LKc4KZQuBa8xWZcTH6qMmj3kuGiHStHLz8uf8vCUQDd88R
5CTnyoJlJHM3RhT2kWdkJrlrU7zU6CQj4wrkI3+ccsm8z5+X9TqWIt8oXlSZ38qF8wlLi3I8Cfd8
SpfkvPKiCni+O1zzgOZmver5evs5rkA7yU4GsJw5DUfIfwd6Ooekyr1K5sWKbVeUbK4waOujQU3m
8oLYXQeNaJAuJdYqlD9XtLD/Pwr7TVJ/L3G977y0rPma6AAUVzSlAZMSX7TA/BfX0gNVE8EcdIeJ
Opif70RXPklNrasr8T3odZRCWpNuWeC2vgQ5xkt6M39jjB1ctFP7+wERfek++2dL50L09wwSckMj
vKzlaRQIghJ0aPxJmRUNM9o6lJ6Gwm1BWgXRBufiNlh1AtoehQfNBkcOmH1YdbUsML1Sgf6WCe7g
KOgwADacAgARqEGlM0babSigA+H37D6OlrMF1hm4JPR1RiZ1vlU0XuHoRIKXGHmsq7Z2nRK+wyN9
XSGCMaHqrolDmzNnXOLyuxJxz+Axxr/LipyW+EDTQ179kU/XvqpplZJx31/cQNhKWq+bZa/W7IOM
Rbus0cxGvKAGx5DRMXGK2ELGaFBKhvbhTeDeH/Jq4WpFS3//BIUa/S1ce5noPW9WM2/RhLg+wjm2
bM8BxgnH3+G1X+J1gGHZsqCmCWpFDyCRvzG11UsfMBnq1lbLVqX9LQQuOZbl/MQaTyo6+yKGFlAl
gr20jr4eD9NgsIr/eQIjTtTXrj/RBetA1mqxQAX0XyDneRhXYsYajzPFlTXVRZZvSEeu+y5lklpm
MqrKIef3TaU6GAM7Mz2MKtcDqp82bbDEtS+LfDbuXDe3Q7V9UKdSw6OQglj1RKEYm6l+CVK4oXfg
bCzTYGPCGVq+HU22wixVpgoc/JLUqvlwHAORjs0u5ePwiu255pmpwKkIII0lWiiHIgeBgixcbuji
zQ4FF9pES8ddoF3gYHgwLRCCW6e/ugjw2oAoPaf9Z1pCqzAMKzQNHnZeuUqezvGkLZ1wuFf7R/zx
SlMs5uTLCLHaj4SRdZJSjOy3jP7htTr6f2EJj/32oMhhstv7Pk+rEPtliWMewzancLI9tVseS4xT
vQf2wonhrEv+Z1OawXebXGlSXMAI7sAdCUNfopcGdGSo3+aryzId/QINv8ghxhIPW/FCWxUA8U9n
XV9fVXgPsH+ZlJHHqLVf9xFP2WwZSTxsC/AyVaaSmHd2xQ4FVJ+VQE7YH1CmEMLousllku0qzfXz
gODGy24a4X8qv8rljFDMmNw3AJXQWDLYxfFqUIHoqGG/NJK8RvmfJcx2eVnXomt9Bt0MxWYgLWaP
UfXRi7nSK76DI9HsCCNKiFsKUN2EbxHWoYVMELYQ0wbLDA5A9oS/DKPcL5L2Ucs5eJ56USxxg2zL
Xde7PzfMkzzVMWJGCIsrwFEiFIZhRbYYscPa8Kc7Xjl0zQRaOwvztFlMB5q+nmXaS+gI2UUqltZV
ZtOsct8wKEkuuY+tGiv74EjUQK6YEpRyx4P+oK05EGP9HSCwWDVGn9JoOp7BFbWXvjTOCsTZsHMB
tquuc4/5SR8dLl76TMXQqNalxpLXe/5gdWL77JH/gaRjwWvu/AoEQpa69u0MAu6Ce8pSWaiEU8Tq
nDQ82x01nY6kDEtOnnfKPYMvHu+cCdFp0MyChnGambHaah6RYJM0cgjJI4QWQC/K5Q6ZtmUvKPZc
r+ruGzoyHNC8pDUaqOBaZ6toB2rE7fbJfq7VZW2m0zuOwl7IHlFqpA5g948s6NtL/xeqPrAZv42T
iXGRuI0G07TfNICyrVjt3RW2mFlhtY2lWbQWQlbjUL+RzvO5J6r4l6RdM8W/ZYwyfxKYME9w2n22
GZ7m88KgcvAvmzoHXRcWhDs9QA0uFJoRllQ/K18b/yQ/+vDSMwDWbC7KGP2Z+Sr1ihF8CZddl7kq
LP0oUkhzw7Zwb2EEyc1xzi4707HyvBhCtxTIaKeyasMm6lrGG4VK0wdZ/hY4P0j1toIDqHgWoJm2
zsMwG8xal02W7HL7aDnxKA1tNudjMPzNTHahUsaJvG3S6eojxNEn1vwDZBxxk0d3VZhsArAeZeEg
kd/SWTqalk/ppSEhZ1I/F/La6voFqDegFozHC/tSKc2+bn5cM9UWUJX0LRP/CcUOQhjnLTv2JM9G
RpotS8GJgbQ64QbJsWkPx5vYClweCV4f+1K8G8MFhqhxWiENgE7W4p2E6xCzqe/5vU8Nm6nOnmj/
60tqYFw4LdV38gzwSYypgyt4W3LK78mEB/GKd+k9gFLKSWGjQSt3DqWHaK25kZl7phlAjfUdWjGa
eNrfYapGFHDcRwYc36hBwXeSuumC9F8/g7DMcdWRZTbmznRpEyQ7zGDwoN8Cx0Dpzc0MMbLo8b41
xicu11FgGf6GOw2Qm5duus1wvCB6Q1Pxmgx/cxCf5faJ2wWLoJinD98+x5z9aJYSaK0nIMXn4lTv
Re7Rf9VP6XAWGduprJKTi6gQsbhxc+gxHlDvnRDCmEX/1x38s5nfjIM/m1zWfM6NJRldDLMe2aZR
W6hWzrj1wZG/Xt1vA72FT/f7iZBQ7BOXTOqcYvbRPz1rITOOeZswYUakJ2gyR3TgMrUhRWBPLJz+
g4aQh7j9ak5uWuhIRroLKA/T3tyZYZo0nGwEOSSp4gc5AZrNxga2ar1/eFyjgpWyh5LO3k6rGpHw
Fh2SSlSLku1pBkuAzE7CIpn94qkT4nhlcPwZ/tRzbeXsaqCwcHf6vwUGMDHdAWy2wMfCmcsv8GdO
daHa3dqWYncsP0Yrc6xct5JtUMGMPlzhptUfXB5z7y6a8i48Nu7Ik5fMZGw3TB1rd2eVs3WsM0WK
nF5xr/UOC2ky5TcLiHjp7A8hOCCWfcDjn08Zt+t4PHA1ClBPvYTe0nm+sNvlK8Q9MWUBoHGJLKXz
+hxisgcGbM/AqlY+Bn9ikj0jA/3goyCU1QvjGoz2ryFNapg/3I7ES720MGGTkzLkEjt/u3rp9CRB
gGgMq+QOHHbTYWU/REva5nRwPGrFv9KWOhfqD3ItI5Ngk7HXlgOXff6CMhyoF2J3bPNke2G2vSS1
xghWYbx37jt6rst3mmdAOf92yNWyI0y4pXni1KBHs4MsLiNgR6wuz67KJ+FLFUkkW/lMtbmsvWze
Fd4mGD2dTiwYGnZhNzC1vtXNjIrDN9xK5EbdZN/I161dk+Y6Kjz522XpieHGJ33fTRGx1HGyai6X
Bj+0TlusHjH1GEhWQT5ymKj5DQqyDi+RNbki9eSkrhnfjNODJuE8ZVRGS1JzczMzhelJwW0KwcLK
TcM0yQNnw8T5WeQdU8jEmTnP6d67/uYD/eK2sX5kKQ+JYuE73ZGKedWz86JNY+Sc39leK+5JaPLO
nWYTKfXCXPjzIa87D7xYYhmCFqG3yKdhrpLO6maUwRyNz4RnebRMA2Sx2jrpz3aq3/DWCWHCyXUy
QMYkVKtaW6vrIAwJSfLCNQDGrPbF6yfo8bZTENGUGqyJ4r3SQI0JMphdihA7QTtw7GbNsOM3a9Ej
KRF5UtSKmK5mC0QgUNN+u2KfPKuwhjgTmWWXIJSeYQYCVT4O5gTuUdJzDRqTuX7N6MMbDO8txwWa
Q1ZCImR7enlTaPph43AVsaTVF0XGzUX03y92fqSSK88vN0p30Koue8DFFzMxG/wVK1HvzQMgqXPT
NmIIUXZwHtqQoheiYmaFgWtHDqLKDyJDFdMKV7iRLml7ko5xOHSOJr5Rv5V9UGcC0mc6Pkc9MVH7
tKvgH4x9t8+OPH8+kTLJp0pMzzXq+lztnEs5/FHAdxCJnBtAp0Dbtao0i4lSp/+S4iOHXLLS27p9
cZnLbHXjfKt6cn905zNK0fRQHEm39069bdBXL0w/OP/N0Ayd2V7cGfOTXZ+lr13LnGdM1LMV0bEO
p22/+dqzuUzFM3k/zKGgZ0HDffluvmeha7cHQ3dL5XfT8fPNf0aa/ZVBx+33F8CKks6Dkz9kxjCa
lcEBIXExSXjqo++JtbqfyKVaijgYqBEiQbB/0NyovDHlWUqCNVGQTJsTnJQWjTU9nV6B1OocPHDu
9Dlmpgh2cSuBBb6zffo2BPdLRXptcFxWm8LfOq7GfSN8wOLQttz8Z6rLyp0rgl6UZi5KM50cH92/
xb0eIrNM1DF39eyHcsHfvGYcBs1Omt1/0ADBLSLf6Hq9JdUIOVWn1wEk6zGkmE6CZ9YkbkCGo5NJ
yBFjrAOVlvJsU9PYhHP5e/DsRmYwIwoPczeXkfA7Kxkhr14QQiC+9iIHNCkVS5SKbVsY7j0csWBu
ayQ7IhEP36eb0lXi9G4E/5ak3ZAW1HDPHcawWYUaTBhCGQsoEoTk1lrO+jdNa6ckWq6HlkIAIHLE
yeezPDXIkCadGZgleQ/Sgp+gvZ/a0CeRKjvMgh79R8pvz83wkEvAjli18dWh1F5IyrDwqN6pMOBz
ikgYyA9V84g7xDp7PfYDLvLfXgWqdgPEyYbdND57vSrUBIQBC0pApP22xChMxRpOnUp3tGNhy+2O
38Gf+hgpSJh7ql0ahdIFgZuai0IJ7t9Ld56I5xVOyEgqbY5jhmxIjnHYLaYqlI9paOd27zE9QL7L
guV2SF+nSJ6Hva+1az7aLS3yfRUZShuTUvVqPcYtk/cD4sSHbNMkRFToWjeJfXV8wPDMkQ1epIbF
Y3MoJ0w5Oc1XKo3Rv1EBJTHN8DkNA9oVR1Rx1kz25zJc/AKCql2Xk4V8D8R6cz0t9K/bw2eyJOVN
osP+DU3JY1YO4zKfrsh264sRTHdfrAjtNcRAsOT6QVjo4tK/aoe5Klhq6hQtw1ckdDwaBt1vpmav
lqusS6vsozYXWmKUES2RT/lOJttZon/Ba+hUB8bjuQgNcBF4F9PsDiGvzxveRIQ60g9/0HNW9khl
eWhvCYuidWRsp45hBZpUoCuyOp6yF8Ie3V/KifiPqhpARYcD5Ld+p9QGrOgXDbkvl65XJDcxrWuV
yDyT+qj3SC/5+5wewgQedISk35b1ZRMRi3f5D+LafCjXKzQPURIbsQDcmbER/fpXePGpRb1Tf+k9
Fm9Z8LqRkTl0YPLYXdvn3ia4vWyS8SAp0nXoSiAMiLnYuE0/eHP11YGJyh5HZuDFff+8MaZRQWXT
r5ZUz0sezJtCsHtCIN9M7IfWWVQ8n3hhMPp9VkjQaEXbci1drdZ47fYvmRIVGe5+k8QOv/GXD32k
ASQGSgadTKz9Lh3G/Dd/OYu5wiB0axryfbCvDcV0Lfb0X4rjqMYVnMHBscGkcnyHn+CyscTPSXgX
x8r9632F/OLXA+ffgQjXpmHdwK3YhU4LRDQlLs3jvYMM6PEnyMC3vctDBKONZsybXhRQJeGYpNHg
lyn80l9MWWORIur2ZXeKdmfGGu/OUqXt56vwxHxVLy52MZumi83kYc4vG5baHO6BKQmlBM4hFIum
2ez6hPDSBpNlsoaDVoamg7dzXmv528JvO9bvNfMW7DVwaDXxJwR6AfCIoGdAqeRh3kT7/OYT5aej
btLXWIUiNlIZAhm9QkheBMef/eOdyyJqSBq2cXrDKubm/sg0oyUOqgB82FxMPWIOcuQEfnfScI7J
I4QmCD70MNcp3jZB0UHy5G7YXV7mzu1rHrzgKv0ZJMaaXcAHeGtsvDjksMBNiokrB0rnswN77UR9
128QEe1Dt7upQ0VOjUCLVJ5EyNnLbG91JIiI889ma/hUWpP81x5RLUL+FX6/SslnYK2PWx4nMhOM
zDirCG+Nk5jirwJV5LwWZVIUfVUdQFcU0sUEAs6bmWMTeEy6TGHdr3ip5Zz2MiQxyv49l73urgpc
lx8U9jtC8GQYFFVt8u+QTiiNFkkbmj9MyVb7CqKQFM6ny+vwyMY6EKXgXTYkdhD3jH1AZUj6biZN
vll8tSkoVNBP7l+fLYXGtscWur/dNsMQbFZb0QBwY4iT4DbVfeZukdj1hrW2Emle6mOI3oGZBkC0
G4b+NDiBsJGfSTJw6IFrw/VQPYFmHw5F5kdH98caib7gy3xn5UsijvoDkFL7uJsuU1phNaZkvBMU
DcAdKuVVXsF3O7rG/zgif2CPGahLfh88hEKv9MavepAyMslKnwMofH9h2wUuAYuPNndxSehakKTG
U8N7EpPx6yMbpEU/wS9UmhRQVqY+He3E+FREJu2KFC8bBnEOBYQmcEJ+7eEmV+wyV5WzeMv+SIil
U07m4Ndv0Y6pHVwq3/rw7NOHZUU0QnN2WkdEcBp9eZRq4Ud7iWqdRxh/TN6F/xmFVZHR+Llw0cE9
Jh7qTLoEj2VLNDCMq003F8cVhcswIb5L0av+sBZUL+aJD9gUdIKO7w2/lZ37bz3r1DyJnxuVndio
OXL5nxkBJ7GUnaC5+ek320Jcs/sAXX32zs60cmv4JnjDytQnKTljb3zZ5eLHYFAHbKoeGUHy1KdA
KPkFzvtt/xZgf225haY2cGfmjPlRoURM7iFaYTaj0j50XhBQ7XvTkTlra/gte9PPeZSHG2Q/IeY9
89Fq//sR9psQPYwoeOLmFV9DwHthcQvbo0wRsJSnnKuRR/pRVBaQenVfWiUYLszInNZ3/LxsapgE
RKvpsdv2SMwBLLqot6/jeRvBCS9s6QON11J7Bf+1ul294/yTHePOmD1BT+P+vtv40NubNWItaypL
AuJpgyyNuvEqI8Pga4ZObE/mF2ffPfO9jrW4+NEwCId8CUila6ktWwCJMg15Le4QpbkrHeTCmgxW
nozjR1AF444RewVJkpKb7wVshQCdOfMrgoGTG4ZqWQg+1lLess5M0d/AS4YMLlS0HW1GOKx8kKh6
gT0iWaa8CTCslpeOkTonXHZUO9yAzufQDTEtmK1WWJjt8NuRO4EmehJK+IawA0209vvq/BP3bObM
TbRTphQB7AgkzgZjx9F4Xbhp085h4MkZs2sjhZgjY4P1WyJTyBpZj7yevfQRXkh/fyIjKSbQZLUG
vC0KFEVZaEfocH64TqU6uxHBtfbO33VQsL9OgXX8Ps6UIGwOYhLEeTfFlL5tTxyqekVWY3Uzj95t
P/Z3O8GCg02Qls2K4iTPCNbmt2MTXgFmeaSBg8dx8Cu5333l1kzB8rux0pCxzjBu0xdrVHOlZttu
lMlNbU46ZtRFgNRfeM9uIFRbT8OOipaLqj9soX06zFMurDCtykiX9aW7dOQMc7EIcX43gA9vJOGU
8G2qp6yN+XjdnOHL1t3O8B7VbHVoe4nQfWTNZedAT3oD0fdvyFQDVuzJWYYtaa8Jtsv0Fgck1etm
vPylzVCNRZcWC/C8XKRWwCI/8BWX9vCwYMxcT3fu2W47nch0wkJYDEARrc/x06TzD5TwRuYRQoP8
MAVI+v5914B+uFGdC+ysu2fmm6Bl7nz2Z9BrEME+VSRSXXf6UCxVD2GnbbneN4MuTCLBeW01iPtD
SbtkTlKrEoUfvzK7OrQlmTeTymBSyq1ZmtqyEYzHLXdREgY6002yTvhxY3xfTcsx1WD/RBg5BhEB
ddI29Yhz/XcT01EIYcSmnsCkH4SZvf8b3sSsWOMajqBiP+qcuYtaToloZK9m9TAw5tBySnwdIpld
7kBm3Ayo69nf4HYORMCjNlmy1+EUDogLotb3fXHNyr53YmFvJhLJPM4Fq/OnwH914Otenf27wpEI
JdLDvVvmgUv21ZslEJejLpZ7jbeP2CGb4XD6/Ej3IJ2VMrswjowjRzqhaVoibsIIcBX0d9UStkij
ut7S0xGhJsW+iDarlaD9xE3/lq17BU66mFSG4H3mD0HFKBWNWZUiIBkDB2N8t+sCTlEb7cNGNxsl
wZuIETCojdkqnF7pZIma8XSAQg4JK5Ri3SSkOQB2TgaHvvepoP9CglDZrsNZRPq3kHH0EZ18Tk2E
3i8MaORz9N1MDaCzyqU+6s/1EWe512J7RK0hCzkGvQMHwUTBDAaWjPMdI77nbq2kqPQbRVBfmkxN
LXZr87sRDRZ8sSTaK+lrvFvGABiDbZ76SbraQymNOc59vC6/p2d64dfHLld1Zx3yJod8DQh3O7Ys
/LPS97fKeVqn775bpuNQ5t7xpQGYbUiXmvR4V/wKJk4BkBJpuPOxoXlTQXkqp652lguvJV+qnF00
ztACnZPv0TlDs3tYAoX8ltb9A4M9zneo0gNGwnSF0Qy/LSYtHg4WrD507bFkoSCeKMHg/xi1WsIH
UGcj4VBNZg6em6ul49e0hp2DvN3qNYj7lZUDJs9w291/JaXQc+81LilXOf7EDOItJv24bqM8KIqx
kPHAHeHS/1Jfveg8jRTGmLwN5ZW186blztPUMNE1HjDqLHin/BSZR6xF/4H/UrLj8UGEIB5KH2q0
XBYllLD27P/ti6JxWmbEPjrMrwqHFPYKhYMc6vO/rFh5TfMmYJnQU6sQntcCJKHy9eng5tK7xPJw
eOEYssg4wF6KUhQaZvY7vxXKlv6nBUKPoxT9hHasRip0bAtngUzKcSb8vx+P/+MmDBh802NXSmZP
m48cL3SHXe/CFwdr1PaZlt9ibdhxk+kgK3NQEkpxjgMyXYntSd2OgcyumbnUkLNGk/O5CB7p5vtO
3F6zVFS+1CS1TCdI8NdsiMMwwEJ4pk5p7pkltGfhv1vzlYpdeNWhx3q1FCzxD9WG0ivgMgu0Y3q4
h3dQvQoGBJbasm8mGp2MCZuFyOgSXFP6GWvWfn+euD2/pGPLDKHh6U7sG7vYwCLvagQuEV9hrEll
Q+W9NP0LCuWpn1RGakSM7ZXikk0RxQ/+R+gHf30MyqTrBZI0KOk7Rbo0X9P5b9xWfJYGZoAbudhs
Z6dApJPnFnAKDQhNkky5Br2mkVQu3g0Z4Nvn9NOCaIaRUWq5iLoDWaYRPiXkD3lcOa9kiwrabnUE
+S9Parw4uvwjYxGrorgz4xINzfgzCY0dOjDX7yVsTXQ+ivOQTRrStwMsmHfcDtWwOMkxHPZIjg5v
g/yZtbm33jG9z8IeWqM5M6i3OCTXOS6LupPFfeJJDJ61lZdureYyK+f4ew4GlehjRv0Q/PYncx/v
ruWw2eWsYHUWYjxQrI0u2hOvMtHey4nLH5MbvcQXYn7CrUCxtk6iesZ1pK3yhDqvLASL+4eEVAEM
CRTRa4j5m3R5/NqMwpE/15N0qMAreipzkmDVJ0PR13Enw0lUEe0ZNEpgsW5gNCTM9g1YgY30jNaC
ttcVzAEyQssM/7fHabGmRaavy9+ETcs9m66qbIL8fWTQbSsJKFNZLqSV48WV+dYPXZTE0oMLD+wi
+o7zh9Np2W9Y+CiIfbFffxd1nABMyX8y+MjIvZUAioebLvFeXs9Wb8hmjw4t1DWlJIQjOP8KdnVj
xAi9DaVg6kHfR99VrxIKnkH0XEFFDwoI3g4lw5AfYbluB2qfMGvz7QEhHd/51SEJ63RGyejxAO9z
anxNoIV/0CA8KSV27kESorKeWHfZn79/mzdSfoe9EZr5mm4Fj/gZTTbDKwBSnJ8UpKkidSSNVi4k
775XQu7XdoQP5bb2vVXDdaxQ/6CGES0XpK73SwCCzmWdKHBmF1SmXHLO9/juR+CCZUuYnuxd9oP+
hFoPxpK6bGpsZBkZuP6TewvO0RY3MleV5PkLt0wuGk5XuUcOMsBMP61fU75yWvcVeOPFDNXL0BMT
+QAZ0bFWh6cviJL2NHfj6LyaKuKzY7ATiYSZ5i60XQiBNKYPtAT27w3kd6zpHcNkcpcD+kIfgVMW
Gqo6UMdIUsmTXQihMU5GnPowb5/VHQkzYnBUY73UxG0JK59b7WVi8NjArX3wxY2IRUsKyV+C5wjr
+KblSQH2qWmGxkXrXRt/Deo8lElb7nWmhxSaI3k1OI7tbNs92JMDDjvjCgzXukYwyYqVbttlXpA4
YNVAOsgdmmYO33gVnPOORPB+T/Fos0TNC8rdqytgMC/I43HyzHSpipt2DcwB/U/epLp8MbUdwlkt
AykXX9dtiopG/SH1JafyTYfgQe3GOYfGTChRLdZGG73tC2YCC/UMm3miumUr+Iwdi1pKF552fZ/S
qtk61JWSz4rHaA8p/dhFkaBSrK5v3DmbSf9KnGzReBaXsQ+oqqKFNwiIqkhVnRfECNOx7zPPx78D
HI0DuuSzwObMP1fth/tsz00hQxmiMMVb6SHn8nOjfXrYH38r7SjvrmuEf4pAhoZNudl2kKThJ149
DLsdZYA0BYPa4FU+Nfpfgr9U50oaMN8pRHnQu5Bf9hJbmg0mk+3Jfg1QTeQd5+j9QgrcApReZ3Ij
piiAWbtvPVmsTqqQRt6NsolFkaoQtvBsXTAtGi7pIaVa6OyGDsMUA+jNVN7diBHPuGz3BNGOINY4
08nXodzFeMNzGAw6UprOvogFQ28zkDyyMVvCEqAwf5xBX6/ZPXlv3kXSodsq0+ZLNPXH43MgEBe6
fPMSnEVVj/+ROeWFC90AGS2+JqPW0uDnvfu+861B48rAbmoN4oXHKr6eDrIt+unNEB5CYB+5NmQv
L7TtpyG5v4MR3eZZAnE8OwSAwOkjM+zMvM2BP8U6oz3r1+CMhe5q8hmVNNKKKfUn1S4kGrednhgx
kmD+I29b8bSebHp+WKTjIl/LNmbV2Emhlq2U0EHYxJpAEcl015Z3xSuimtP6Jg8vNv6VBQIsKnE0
lnh832f41dEwJxwW8Q5Yp73ap+UQ0INtnbqJze2GDYG9Wmfxng8l0zx7QCG546mfGp/q7EchJTiC
Vn4yBidLgh6aBYhGIili3285oTALaBoP3p9EwmG8pAtOekj+VfjC9gCMX54Fq8b2T974FT67+lfy
uXvxWHmsLqgF2GEpQLhdE2p5HpbQcInHzYcIzUra/6up1i1kAMzjNBx3Hggm2r/5p03qt6MJlCgi
1C1SeBySjRpTHSIu6up1b7QIZyv2bnT/G3zh3x4DEVfSLtY1EZh2haSKrzjPvhGPnsZYJgJR3lwr
wbbbOAFqswnpew4JqCMB4hyH/v/xtanunyV6rq0OvEEJyTBXzEQkIrk2JhflfFngI68RtI/tr7nd
djv0kf2XcznA8QpGPcCiSwEx4VjCPzwCD6/lz/Yd9/XA1EvfNXm2i4T2BxRwmYay+v5rgY/zebK6
7N2xeNxW8jXbWSRmPBg2Ib64uZlssOVXbH5HIgpi0IbQmPxrLXuOd6JfcasUACKK3yzY9TrIxfc9
RPHpjt7iwL8kli59MW0poUiE/S/DQEdbUUPHuvLH3ot7CiqJX6FzZjFg+UhOvQWtwdCZtIoXxg2B
YyhoOdeGzXw03MLPThAj0OHntkEPv3yLxz/pqcjd81ikiZkV4ndLkysr2V/GpOOTvJStllF7Wthn
YWoutJX5NJ4JoRhha5iw+w3+9/HT+CzVuUv+phZkT+fM5dy3Neay1RXTuhouRPYWCmxjKgJW31dg
63rL4tHbBTXlXndxlqg2GnQRPQpdbbmoWLij+H4NWWNCjD2GfQQKDJBER7YBp4A7Ndemj2IrZize
aR5hN+bYGiso2OfMQevdluYeHlmWbriTf2EUfnqm5he2RNXLQ42dTJ2ZyZt6YVevItPn3AU95il6
nvmWQz76itcoAAy9sDcrxI9cKBlkZSwFiFGs7EJdE7U/tvhpTxZxOzDmTU85u9wnmCkrs+BJKCCq
VdQZgj6FjY8BYbg2GG9KoOtBHXYyDttcs1iUl4TOAI2b2PHZvn28uKciUx8Pk8QoSkBNHRCo7Iph
SH9mnmEHMFOrVk5QK2g9f2i9+HdNj9f7RgSCinVOyxCIggO7w8FjJ8kBJCBorGaNu2vZCeAJw5yp
s/n9VwntVml8XQcbHDrutfOQiPjp8SSCVEbOMVilDaf08ONAHjjPAnzBYUJoL+S4l+TWGQY4g1vE
r+T0bJUbY4QFp7ESIJ4vMzMAhCHwWN0s3EG+ciMlyCUiPhip6tJ305h3bsMlAg77F7+zucWXpE2i
LjwuCYXl08JztBjcxPrefi31wD7wdVojCXnc9+UAK6lH3PXxXPjY8ZspFGOFakY3R+Y3axsaVzlg
TT4LS2LvGC6kWjmhyctxjgbmmGXxr9QqpA39Pt2VuxW12HcInmDsPT/Izyw858ZKpP4CKjTZzMiS
nHt8Vfo/rtmjksTe5IxgmjxIBeLTtWBLrYBBntXCrwKqe8hX0EJItDihgzlQVQxpycE/QB+I9S1m
2njW7mBIBGOEso13hJW5Y6kogL+6XJW1AMp9tuD7jRh10/u8RZj917ggTHQSvicsfLMUYJKbA/Cy
lnrlf+o4R4y6lmB6TFwDRC0ppnouusegyqjKmVs3bFjC1WJ4hrZKCSVIivQoWYFEkLMZiEqt6ayG
/jqdLeJUXHhOkx7YSY+h1Czsjnzvgkj9n6p9iXe4q4djoclakpWqcH68EWeKckPhL+XPL1QPGrFc
x5NZPb0GZw0lPiXzshtkhBdspNCZT6QMofPE2hdloS1/JMGoc8uApJcpZ34si9pSbm5LQocBVxfM
Za24LnGIcNB+G/uvJ3/ZftVvQoESQkV8E9eRHIe47KYkOAHXFfRpJCU2N31rgkjifI2ALBunUGMw
5g7luhYKgbc3ZOZHYceh3/REeB5Wj9FKySuYAb0cxABQyF2zRC+QlVqcCpoMcHI1/bsa/4sQcMsQ
eGxZk8Y2WKxC0IzzXv9LnfiFElS4TMJgbi2LK7x+owYDGQlBocfuuuQaUuEeNShDx6Rfvzs9wjFC
smZy3/3NZzh7qz72VuN/OvWfa2gQeH2pB/q7jRp2WTeL3cCmCmHKMXcDHucMwyw7Bcfh8jfMhohD
js/rlxT+w1NpEOMzJ0r4+vNrp61LTkR82vGGUD2axSCh0kNv/wVbaZsTH5xAW1iUyUOQxkjFU6en
980Xfr6aqm/gMr3bqePj3b9fIUAC44bSe39YzcJZ+UqnzAPcjfZ4GQbOPRJgbSvqwhSOy4A+FVtZ
3zIvb1vijmni74Q/6ed9R+foAHqTi/sndQLKT+pS0nVBL7jjfkB8IWv0f7+a+a6NmfwOkAIorDLB
q7f6VHYTGMGAmNZZ4Ew4D872ceNg2/dWVYL66zeEa665dQd64/OT0QoC/8d/lmRnDWjMpLtKnfH7
YS+DMd5q2CSXFVo4EOH2kw1tj2B4+runFhgaQvfScOm0jMca2KdpArV5PL00M0qaHpQXLhaaArzO
p6N7/Q7NccOgMJkgRxJq+O9PAvN+/SYzq5O6r2uYEr1tii50+4IeCIiYL9K/rdgOs+J2OTfktTlD
d2whdbiILJcbG+p/M6xc2MUlOW8xrItko84NsWvXKSb9D7fksy3fKjXmX4W2V72gSNGpZDv6exus
cx8IEx5SSnl016XRtQnQcn63DeLLx4IJsSesa9/uxndxTWjedjzsTNKJktWDB3bRdHMP3D+rjKyG
GGis4ykg9GY5oavhCpde2kNGP8SFks6hYt949P6a9+JicuvPaHOJsLeBInY3GMJ+mdZdEVLDqRER
xNqJMKt0vwGocqqzscVdEalXwWQN+Rp1hZ434Ln7UK4NHtrRV6t11C4+whyU8ILUYzApwRUa0Uk6
G4dUbeBBC5VkrYrwENNlXJXu0EO92g8xz3xpzSgW2HTAINQGG7zIrHNXFOBViCkbsrVKYt8WxsHQ
A6G/oJI7D9juezab1aeikAqnsRHQIEfVbLj4C1Wb2Mu7cW7yzODDn5EtZXjwdhMl+EyLzq46YIgg
JIUQ7gHiGqcLH+WrSse9YCCxHOhF6R++zPv2hMm2/6pmOHbHPdilf8gLdLbyGbG1XDnOB0uwF9yL
TiD7C+Q+3qKU/VmSGJP4MlfQyEIvaPipGKoe0Di7KWSWGYFVk3GdfQR3S7bcPp7yP88lG816Zojy
pZg3rEb8+8KOzymO1HmX5m7GIWVzargM5iOm9jhUUpJzIwJDKhvV78bRNCAW4eFc65t54yloLmtB
b74Lo52ARVabwZI67UPrghsiwj6rMzqgMolhPgyGa3j8PdkGEcYxFhxrSS1ZWlkFYaZHAsis9jZX
MK0BevNafemjEXmkhNhD60iNVEdKP9egplnL5ESzV/79Fkp2Or2EHrlnm9jnSZKfmwKTazTxA0O6
JOZXiriE/XPvZjjca9ZZOiGcQyDDbSWwWwz/veO25HpyK3jlwPXKOuDEkn3vmGHv2r2YFW5pHqkv
ce+2nRFVnLxNfngyZco0PxG8B4XphNybIhb0/aGtlJHZImWBL08D8Sl+wYHUQI6Fhgfn5QlMJ2UV
OMJL73NZ2izh3SCCX2RjCE4xj1n89USbaqmtf37rxDzO7lEVze2utgTFhkdHnq/X1KRbvkm0XV+T
8LV8ULGyoRDjUD+/8XxmhJTTjQWT2HpzZIPEIGP0+BpqSH4YjLqTk2tiPSpptCDQsr/s9Oa02a3p
xPhfwaIGjeCuDYBgsZ3hlnqomOIdiljSf8S8A/LjKfhB3NdP/cnC4i3G8Y0vHVxXWT3qYsNZiUUk
S60VFIk9AKhwaLkyTUXtU0e4QoGloS+Coel4miXYhVLLj2ufFRoduYUgf8iqpl/yaDR4GXm91yon
dRJQKzMXyvBjeaEbUOBBDIkrytpZo9RP30CgtYb+GR8ihLm2cXe64pBx1402BQOvfWkv/n5b7IpG
rXKbrEKlnqHSNayMA0AmB9lr4hXHuPVjveqZJGhiZ3DqCji8URNDl0skVCm30NuKapoZ/OJ41HcU
zhaH1VUfW0QDjRbyyWXiwGcN0UElqSS0mnEws8pZcXSv7qGmDHR1UVmYI49EFz5/4cFhG+InVjBM
faJo3GBM7WKBjsUFIT85ku2E1Dto6gWxXBNaDYwHCPRn3Z4uCSEIjZGzQBDQQYKCSm0pDMGkuDNE
FD9DDZyaxrlRZNmYKZI1lyK015kIW8lPVd3USWcoY1XMb3x2iV0mn9AfTyTfFEV0Cplse4u4Pxd6
XOrdruldT1RTYsta/w0DG2Iq7Qv/nl/D4RnpSDkhlEmrRf6/RR3CuGsdd/8ST9QVllorSiGfX7zn
bwQFIXpnjSM4y8+LnSRd1Wqq5nUOwHm9wD9iiPtj+VThIK2pc2jpxzxZwnsqN9IV/7U739JxwTZP
Jce9oNARS5xMT5xYoHQGN3MzNou9YZ9XlG1LXgPzh+pKOLTmjHoS6a9GHgZL7dXwpsPb0B/TXjhT
9N9dQn8fhRtCWYu45hGJuaEaCqP11PrZFgusy0tq9NZZ72gdEYPXtOoXjI3d6Z1MHuoYRIQt4yHU
bmrP+OHm4q8SGIbRjp8u8BJa38VnqMTctSBlQOlIcyrZhEcX2RloAomMJljEA+FtdWH7m5hrZkjp
Axevtk8yulLFbQsWEc/chfRaf1NbOTv/iDsN0RkD42DClsxnTGVvjv+1MuhBeb9XHE4CkimBIa7y
Lic0dJ5sXxw0DQqKZBtaxn1rtTPw9rryxJwzH88jo2MnM0oduzTiGeW6fQjvMSwYC2NfToBTb0dq
Upuvg//a5h6CgpqBsPfbI8qcOmLYTvGOaRn2mjDOx0pp+8bNlf3NQ01cxi1bg4T2IJUDzLiRsGhr
WXpKazP0TuW4JUGYUP3VxIajELilMxaw4q9/pr2LWZmp/dmvRYRupQGScX/2INmqW5vIa0B42thu
T5GcI31HBoywcLF3T2gItFJhH4AlSi5qGZTamk5VfWN5otb6NQHwvMsenXYjV6GMeaGlYYvk3swL
4o6ryl/g5v6clS7TBHb7vdY0NPuFHa6qLD+bbwr9/O1k5u8wPZ3BLR/U9e6kxonYL8jrREzkY2s/
CPZJX6WIGBaE2PuDCogpSzp3/cy0P513YXzRRXuG/1LrAtO76rojaYJAkGFbgntkaVCUJVXfUWrM
IxuTJPh8uCl0V5NAb3xaYYm0vn3e/VwkbcvtE4C5em1++7/6gYdqUcC4lb6ybYHnzzs9L8a7jfcQ
a5QzSXvbxbc9qt/se+b18p+NQO11e96R+6vJaraNUIKCr0xHz190nL4mLaKvY+fceEuePeJpcn28
RplxZTwpD1Dl4nytIpO8clF2nNbU6Q1ZC1VMf5LFJyBjOo0+LhEISNicqEKdm5VpWwhTU4GGco23
GymkhAPPreNlCTGpAZIhxt57yosCNutc9iULa4Vv37HBq6tK0vnMOpS8Vno1WbVmexVejbQOqVsb
SVPGP2qQKUOqyxzzI+WnSaSSjljQIWdaR8RnnC1E2XLA3wyEhnHi+cHCOikAzABQr6OvNBqBXfAz
Bk9K2G6mexxEteKC6wtBUslQMx8FbWC8MaXZOgmZtApM8KdxnBaHpFyCitId4s/A6xTKG+SiWlUi
vKhLSdWJvnOAFm0R+hrKcvX+xGZaL+8CCm6/ANlPLP/pnwFV0zCd9ow9kaMb9po7gvZEJ45HvvMt
tVuA6yiartjUPpm3R3k+clHDb/4ZgmIwBbowCIblHeILq0QFS9u9augrQxq24QUluz4S/xJmtSzC
i2Orz2jVI7Pgm+BXfuXUzyk4czsegWNLsQmrzCJnxrFZNN6lzY0Kh0WBSoUKwxWjAg2mnw4CHf8W
zS8cLQ9Au7XTXf1Or995/oqcdHHH3SWFIZLCOM6iqPXFAqNwlpS74AdKcU12IJXp55OIzlhA/Jvl
an4xHaz8nMiOYMYyvEwWjTcFh1knH+Kn9OYgYFKQBPEDi1uHjYPemQW42nDJp599hZAVillv9d+c
h7eA+lpD5UYHkYrl0kHA0HnQ9Vq4iTAe69iIEGNjSVY3GqCDl7Qpbz4biWkm8KeLDwHO0jFKr407
9m2IMSgc7E0mN5ExPXV8aPy1O7iyxYv0Fo9uHEImS8DLiaRESAjSQrBtMsgN/uKXvupo4CBEEWA7
KiW5647KHaWccRI6GjwXSM1zX1n+pJvtDxiWoxCYYGWnPIKRoTgkF2t98MPjmYDVItokoVB1WTf1
m/oGGO+7Lj8Aa3MBYOTxUZ/c/Z+VaBO/gggaUaVrWNftMUGVI1ld+Q8st6ZqAlutnj8coeN3OG2V
R+ccVLgJYR3x81Bw5I2udSQ5eCh5vsFsNIpr5mpi6klwTu+VrhaBj6CKDdfnAlpbVFLFQxheKCnF
yfZDLYpsLYY9VxP7Pq4s1/54j8T3IohzaEO0QTNFDSXRU+yNztUmaMecgRSrfHlUa8zFVKgjcA3T
LmlE6OEOUS/BevgMJAhTPGJfy+mDacJPyccX2+WpeSMuwMHxh9QlrBMC1ek1W1413CBJSz3uDqfW
JECKWeVDQY3sd3RT9cBveQiTlsGI408CAaC2R+on8uwqLi2fu3IJg/OJWsYvedfMl/PvPfcX/swv
tDEkaxEZPBmYBtZjyX8nLU+SX3zwcP+rkamibTV4zMBdLyzRJpC0Lv1czdI/LzqZtM5R24fKPGld
ERa+MXu/MyiSZiUCm29PKfKvOb4aV7MSLWh3tEOQB3KGxqPO5kh2IbLEe80gxHWFFArJmgn50Rm5
7P+JcIwmNLEupxLdCCMyzKOucEkiYYtXdOLTK6+mJKmcFMzX8NBdcts+kJ8ej7F0uFN5x6Ywcbw7
jseHnpbuveD1jVZTVJq2qMq6Z1LpsV3mcTdv5tU4wW5KgUtXTEn4fb1/W/S1h9Q2dxzjA/xwupOU
vpvmP6amqXQ0MwBGDZsDR4ETx6pKfOicr9UGQ36kRDqPG4si/5Oq9oetBUZ5PYfKm1W5EsBHmGcE
Zsk9/IhM0M0N9vDjjA0r6lFutYM31fxepPfD7WFgQ04ja3pv12dzJdgrrPELWa5+Mr7bxAm4h715
eCNTM7cHcy76z6PnxMwxsosmNtGqJV3IDjjAA/fKkETwBKWYl4EkTBHD/08d2XdfYOOoevExCk0j
s46aFiXifGA79LGxvPY/K4/1jiFohxKrgb4iHGcKjwFqOedSHeOw6Jqbyg/xYR6q9WdIOTMEUV70
HQ8RgRbiOBk1xD+YZwQtdU0NT5LOiDp0tEPLd2NHZb8kjMbzb2RtcPVBjFg2joH4rjYtlLOT+3LL
FyN9442lPv16QYfV6xdqHATu8SKKD3Ilrx4bUsNBZqaRfu2oCD3LmgxxKl5ycakTayWIQ5pFjvaS
a+Edo0jAFsex2r2TN0s+UNHV5zWJyYGwwcpbbfxSyZQXpqQIkxA5l6n3pO0TkHQClEOb8GFIgQwB
Df5gHj9daTtjpGuTs+MWjoo5c/iya+Vtg/A9Z4oMQCP65/6lLr6N41pVC0okoMfObqu1E0D9vb8d
Pk2NBdyZ2ZZQhmLi3PeaXz4Y58fruVeJAA/G9jsJGtsHEXMXEUUX35eMqbl0/7KMZkJcmReLHIQE
ubIQomHD4FaS7cYHUteEnyKfQ0iRVUUvD5kZB8VoqbWcVsc27XsGPhcPqQqqWK78Iyz+RtbSn2F0
xRHdZrhgO99mkP5Th86N0CMPAMtgIrPzxhoUbgZbRPC3QEYcwWyYXdBfi81RGfy9Ry/9LvjOmjaz
31EyKogVx3PBSA456rVr4Q/2vNXJfd+UpxTHaWvKyvhJUgq/sKX/ty7jUNDHggMd+ATG+EG9dSc5
4boT5ZXR/jnYTRDdCCkhFECN9WB52oFxOcCRPhaqlFHuvhbl+vAkEpuy4PGTi0jNGqjQnk8P0GSx
li3l3RSXJvBZgBIZhKCZTbFXG3DdkTJ3yLhMxCLmjiLQBfFxBk9wWer+OeX41yMfiAfbhIUl7b9M
lCzkfjpQXSc4KaphI69rznefoSLqbNLAv/PI5ygyFl8/uzFnnUSTgVy+tmQWFyTjQpRbi+BZOWLP
JNL5K/Z9/NZ1yghrehREIldqCuWHuys1njkJ39To+RhnT21pm9QEOPdcGuxqMeFSpYcvrI6P1K3J
Yqrvq5aH6y46k1abKjAWyKXCM+E8k7XY4xxgsnBde/6cI1znLkzWuifb9mA9/x+88WKkFbD7D6RE
3G6ky3w7fELzu9Nd3aVoQmIJyKCFQfb1Q90OPrzQ4BM5KArDvVg42kXQEKrwM5E0D+0A2XObR1AK
zvbAT5Nw+J2EcjBkFK7w7t7XvCvUyyE/35YiuVlpNej/c7t/mSxFuKNqhbs1E5ch57U6DNpWFrT8
wDrfBWp9DQPRjvV+JaBXnQYDOqgx8qhb14O1UXu5f6TfB8q9AY8uLX+Bj1OJt7mDsDY5TTOosP0r
t9g3SzHX6rkBkJBbvcKnzTN32lPkClaCAaxP9lt+B+fmHr1gaPYDwAnJWh864ubr/zKFbsHT0DUe
aBGXUxV/fMWlH8taA1bVGRF3lkd/TsitbDN99irVx5VSARbE/2l0IXU89lUXZfa5uxiLk8BypEyQ
b16HlXHkoftDdyn4rfF/Dh+J8i3tPidlhI9GiaQEKzDvEyhFiO80wc4rjiISY9kwTHhdq+YiJ2QU
Rn3hhKpoe+qIEnJoR36ptIhvStV8iQqmDDe0LCR98Yv4MMM5rVfwna2FSXSu1CjTIKzuUsjntQ1N
b47z0+7oQuMGQ/Rek0VCxMysrWuV9MAlCMDdT1HgXrFiRey+SpHiO4e63O/lQzRPOg6DlA+d9kD0
HuPak5vD5DijHIHdKTv0ZhY6y8GNZ7DKV8jgnCGOmZepLGVgtUMOcO3xIzgaaNxm6pCFzpbPfrKZ
OZVf9qhJfZmS3Tx7jwjh9hrK4EXG6v5f2hZlJDFJCkCPMEQlFRQoUvBUUz1pl+iV+nJE8cMA/Uvx
Usk+ohtObo+8JN1qypQ+AK0SqUxW61zKsz9mmMddzITmUuCTTEVHPugnAzgWcFlEDEWg1KZMz1o5
k5WX2MxWT95bc7Oe0uPOthrQzbm6vQhhRrxCjZ40nlhldeDi473vRIWv6TXurt1hs9MSXLJ8bRwX
aTdAIXSe8I5BmU80TE8Nd8g21AzByWEmVvBGBO4wp2d65KDNS2KsP1CXyg128qlqRd/FeJwF1eEF
+XaVAjOHkwbBvydfhEc7IWWcnvvMz8HpAL1vnrFQGIb/CMqGp45BGNHskz4enjqC9VIoLHuQ8Ih9
UlfeXop45l/Oc3C0HGR+bV9EG0Ubav8TZCNw7WENssIGTwGiBCtFHIdVJlCfr+VF8gRM5o6yJUnA
alVD1BtGyL27Ta7YIycwbLyOHiDin1uvnvw7189PeKvqLT+fSnEoeD81kXeW606bPwiCu+Kk7lUB
gTSeSStn940XsoNycuutG3rVIOgwbsaX1h1czLKGa9ajPkIvBpRyJ093b9Wg1z1z8glcm2JEBwI4
yHqjkpbrcXAFytqLx4zQKfDKrd78yIwC1fynRUz6Qn6avJKV8xb4e/kn3cV7Vycl2Ru6Jo+GY80R
VX+p3IMR0BxRGlGRlGMKf4tBO9FykJjHY53d9NlDz4f7smQb2PqH7TCoJB2g686rVrNf9Byr+7X3
cFCl/R7x+fDew5/m+TLYCrA+ziEgg9AmVRiMeFGRO+LPd1WfRk5FHU95ZEOePZ3jz6vgQEeS+XlP
p84HMtqtgAMPp3xqgA6nL/xMMIs9XN32c7DXeDXyyDnnaJZ36eucN5YZAz3MjK7QRQ8c2v9awQwR
Y8/g+qbyaplqekaWn3SWUsx7ioIP8pFZB05Fu9P2uN6PWP6mWNjUIxjS5O1VX6if1Gl97amL8aie
MRAE+g3yeb3XZ5SoxLIaCBdqf37Wo7KzzJg/3UfEnQRSSbtf3kXic5c1V8HbC+ou+G225f2Wnk4F
jo9CwBwNv2r31+NmC+wi8chpZC134J0hNyExABV87VO3pdxzXWaPp6b9n8vqwIG9ok5yYqBPtxZT
qkUOPkf0ASzFX09cOhfS1+xMedz731wjCeu1xKk4ORFAEVYwCZi/+9Ai1zLxwqn2MneRBx3VS7XY
So5EUIoJ94EU3OgNFt0uVdWSh0mZ0d9zwBLYFkyy6c/HtFgyRAcIwhsp59EV3wubAa4Ii/YOTCkq
0RUkwHS2koiYrQu3py5LlXv2af29y2GFzCz8YC+V6f6sdFNDwy0JY2eU6vzFU+63fOK+RCrw+8TF
R3CruaiRB61PLXFT+4PyBtAtQqwn6Q49XPAZcf6Cn8sW9pGl4QpjzXbBiudZ4EHY6/qCA3qSD3IL
4MhF/vlPbUnt6hyQehCBzFflMjRP4dkw1eYZ9eVuATkWxHqk3kllCAqWXhjhKMwflfBVWpaKGTDM
7mak3aGOAOw6LGk9n0VYJagfr/+MdOqg42mNe7KgA2eNA8muqniQZqAwFlKYHmyp1LR6jILu+Xgz
iykK428MpK0ZUhZLitgjnrSUaJor2GENNrkhxlzA9B1GSFwaclOcWU6uINtbQkyg4BWTaNDFyZEB
8x2SLIXEVqefm2Ny9//IvsmDPTrWcvfY62NaaycUioDbb3perCN8Nt2Ki72qmXJx/X6AqR/JEfyI
o86b0S4MGnOa0XZZ0BG2G3G3I9QF4/5OQYRk8HMpL7OxkLlikz/e1Vi7QSmY/gpU0sy5RAH74oH2
vrFaXkDjghTL6skw5enxwd/NkuT2fiuqab8wcyjOPT1k2RWwwdlWY+Y2PZXfJi7bJQ40/lr55oia
hPpncOlRe+NwvrWt71I/5YAbsbz7vOJVPu3xcTjxIHwd1Hy5iPSoS8KIvJM7yd/yfA37LlSjCAsI
ur7cNvKUKk10JVSidEf4H0m6p/gy+pCd5Xkkb820UaX6RR+qeR2HUUxoG+Bi1a3NzfJu8kFUdjfk
skwj8rD8qnvuSMFSPD9In9lWuUDdFbfMyxLqGQJOLajVKVDeDyMaanj7OVLdhmO/lXJlzN+UIzVT
h5cCg11Ix9bj9V0y+xxBdsfBqEdGFjOx/kryWUqkhKLllfJDXfFuldDpcCO/ECyKayoq/tgsgygo
tjaPFJpahkhYG1fg9INl4DvRrv0Xmp7Uszjn14HrhLiA07ycztdGXAF1T5rXGDS13/u8juMW+02q
x/oaBFk0ZH+FuPjZ1O7cH3s5GK2r9q8lrqhQYmfPFrN/GqYO4EafoWyvcan/7Tyc5ZNFWrdJFBwE
vyLqKdzg3lGksrYJ+Qr0KPu5YK+2Dhj/rt8dX/kMlF3xlAuvX4CKZzPdNQF86FCZWey0roRLJe4Z
SIW0UGamVhUmX0TZ7Eg1516rQjnorBLoxdz6qWgZxfHMT9ApIHFnd0vW0SpKdrWJ6xl5/WdpPtRR
6MoEo4Ug5JX9EAQZvWp/JRPn3ntN/qxtJcCkWQJpPco+5FucF3hDC2u90bH+9IXjJNh3pg5x/4lq
mWosgcbp7JKOg93scUtbTzlYttdUvQMoKwe8Me2NntPgpwlAK6FJN2wF1sdW2fwd3rsPVsWpDutB
HA8ZZu6gXcM6RmfBEcCJ6jNzwqZJFVPVz+6CSQSUuztTbUdh7LJyXhA1RsxTQl6pnOLt1my49L7f
7dM+M7eTCgomwfJZv403TmHr8OQL5/T8GbQyvWvRPOfs6DFIAm+bZC+3U501lZlSIF4h9f+ZIz2T
H5tb9+YftUkdKiSHkIDLcsuKCgvMDKGsPqKLVs015wvIAfYMjY7FDvPSdFDCChinZuglEBz/yr05
vJBX3Nk57ZFKAoiaeDPtv6vNAxcXVXOKtA6YDTF3oov8Wt520KhEMSneu3lkrg+2/kfpAjYhD3WY
d0132mcblNUMeo4ouuX/S6iNosboH1SXF9wZG5TfYPOR/qDplH9R+En27JyjkFmt/XLOLyrMkQqM
7dRA1P9qqnbdqs36LPpZmjCh+g6ezm2Vzf6A3tOsjCSn1vLRouU/0rZE1Fl4yevWDja3yn3X8vrM
9So6fLkM37ZVKVBoh/YGWvY6ymMIF64/xHjnB/g7pKbGsAFzJSsmIAQFFsWXP7JYmoRnfP5VJPvU
s1FpSNjCbEBIoh2om6gpUqXSlPS+dkDITb9y6caw7cQsH3JbOE+xDfWWtBKqOng0XqZbtS1/nw/H
MFzH/W6TOh6nnLxM7ZipD0pa/eOGh97F24mRXpZszQM1srQhoz/hzfiU2yFVVRA+kt1xjxluk3/g
s5npH5xQDLLudXBlcQ82WEfl+jOJBNZVR/iCd2m61tPognjUoGlqcKP5wNTWIhBetROPDNgW+HQZ
h4E2fwNiu3MV7GapUJuXIYPSswZKMwPEU0exLLnn83iJroGWqNkUdtdbS/nS/xhaenGCbG7S6gcQ
U5peITiPU5gSwo53e3FlcIFNe19kklhcmZUxiujHPTKnZu7GHUzXdrnKoXnUvbnD6bsKWURBLQyi
1D5EAJgLIGOsEHxmfmAuR1K3zLz9gfQ0GQktUbSzYf3TCBN6IWehhnJRilxOJ2kzCRaPn/UA4eTC
T7qS2aEScZIf5gn251oLj7SA2yCgppth/qxfzWoWE5ANETLxRUizDu5zRuOQ1mUfNHtnQFQXyruG
5OvGcSWgFt26pKyRbeLFqutRv0b+8MsluFkqvW+U5MjciS/+hBJU2n+L3DAXWsDc+sHuxiK3k4IY
z9F0nhocI6uzOwO4TUBHTV+43NxwRnz3JfgbNu9uSqLUFaAZb+e78QlhTkj27DMFYFUru97OW5ri
EldOeOGD/xQM3IgNH0ABN7au966q6+NF9O1tXezwYASUabtxymIk2JMAXxsyh3Z25sDt2C96+2vw
P543AeYzEcaf6Sg/zK2vLVHQvRfygk6M/4BJZRUxXg5QVfu1TXJoWDxxUvwQhuIHpRh0HlWTdgPO
Dq+F5rtg5ZnDfM5HTqG7jKdCyK32h2/fIvmic1J4l0b/u86or5h5gh4Ga/vBpRgJn/83v4JIMtSs
QgYE5xmsame7fNnm90mOdqMRFiKLiXywPAUh4HOtB+tJU11r7g5942QbsBv6ypMUfVR3oYU3PvnM
I7Nkgwd8cJ08vc6n5VaNmN8FEFP1+qXUFZBTa7WygDsUla0JneHSQbAjZvhswB7tKWE+i5bdg9Xm
ZAHKUbLDOXI87daGOFvtTDC1dmuBOsckK3v46MVOEhs2RZ2fhne3f5SD2i1UdfffFtLFjGVQi2K5
whf2YylMrrsnFgD2/kOvFdUYUrZuXH70I9TC4XJBz4gtugv8lp9xKYaSeuD8au6rc3ZxV7tATjLc
MfOmeuiG+p9YRXtZgFOwSfl0TYybWJsHpXMo6r5xKccKsESTwDvxei8X4pEhzTpi9F4HTrQPUOXf
5UNJP21ZlF8NG/jo5UurBz6sah7DhlfwapYA1G+JsT1lWw7ZM9yp/TY+RZdMdniPl3uvKxVJDqVV
tT8sSH66YkYPNjXvg8tmZoQLwKmp0polP8S+PYvYqOyMHUAb+GuASqLMwXaoUB+QB/f/m2Kcmon0
DiJGnkDHb4840l++4FqolONbYqe/W9HSju2+xJpK3Vx37U084lSPFr3+iMjr1wPGxrWDP5ve4iHF
J1U+nLCp0qCfow0B2jupklMTvCFXN1qonHy2be+NS3kwwXtaN3PkTNjEdbqsK2O0nziL15FOyete
CcvAbsfI/rfDzrgNOf7Ndu5l3obf4idn97CKAfRNFVXmQHQFrKCwUv7xi+iHDTMWvZFBxuCb+wSL
cxiVsYgEbP1xjaWqw7lVQR9lLPLJe8vREGhrQUTDj+QZo6bIKotWUHbHGfhdTFQetUgtUWpSlxNf
Gl1mKRFcxT7Goxy7kV4xoAUbE/KsUBZ/yybM0UrF9IthbDkIpIcfdkv7pfvNLaKDtkuI7ZH4fWMC
cCf8UjmchqelOUYAOnJQtYAS7zgc+oYwb7MFj+MhrqlnOzXdNmIrNFMTmWAcCBpb2FvLSNZ4ehI2
HVz1LTSxkld64YKArnCJVMYfgWAj+xkt9Ou+y018DS+AM46uf9CvDh6H3zGT0pj1uhMA6kq5joEm
+JM6djLu18HBH1mypR0IlctznXxB3QcQMVfMEdGStdz6i8uxHRanOg4zU3c0CIIeJtqK9vgTdYdL
283LyAu4jpYVyEGTmFA8rAg+Ydp6JotROm8aU1eM0V96ru+heIhLs0df1hDqohgHVwGppONOrzxZ
IiNkstYqhVY5WmzYbxWOcrqcZf3Sdw4utca2puJ52vQJw8VRAX9KsH45cE3XnSCVn59w8CvTMsnt
5Mz3DOeHUJ3WMsjV55VVpR6g84CLTCw5G6Fm5zNkRPqzhMXU1S259fxnBfH3MKE6BizRph/CechE
aw5P8UFcNqdVVawjWVE44KBhzbn7UTJDTBOYyss/SfPwgQa15qt+RScqzLH4iG4Ou64szU26xHEv
+hXC0kubwCMkpVQhAq4/v6mMHh7u2RNnBbRync+oKDrz2UqcBz2GgKE7ZFa6CG94CBK1xx7HgCK9
M7v5US5EhOANeuYo15KFVZ9uou+IhWvzt3wTiuf5qklbNJZnSWo7R77XWofrd9soy/QVd4tsUQFe
5zyz27k1TlI9iUreNrjQCskIfET/BaesGQAY/iK/Zm6Kdjq/MPXfdWw9tXDf3I2IoCL0A1WOjHTs
nxWq1jlev9P6os33zQB+vL3yEfvZaaz0VUbpFWpHHLUOLHN3PFpXbxrfuAv05+TM5nFD7eqELWHx
5PZEh7k4cAhseg4oI94wcYITgULUj3SfYzOspGvo57wj0DaqXyDpdy125KAHE41RTRfHHRt3YCPy
TkMcR14kfLRNQ0Amr6UnoDRPS0tL7l3Wnwiz0o5NIimFa15FopC3J748jxsY0pgxbXmdsn8TRiBM
lNbbAi78VhPfeyOiGPQsG0NOip1QCUFE/pWYAr4X/M/pOi1FHkXd1owi65HoQtlhAKl3uEH1ePqc
4OngQEKP73w2G6/OaHnUdinOzFV8QY9bgpiqo1V2yduw8H2kMpO4nZrEhz6bjmG6/v6yWOwYH3Y5
8BgTVO/6D94MxarrygTmOTB9raT1TTky4ffkwXDWq5mL5q93g5/AgtAYZR8qwT+i19IEeq8Ec3oJ
bxvAHuawEFQGSfGXj8BB9WS0gXgJucpA2SJm1ERXFHSCRFRI9eX7htHQRsdOhrMuvX/hBV0L5qjI
k4hbN9Q/eMMdbm4dI9rKKaIO9YSSFw6GL5vMPCpfk/YCidOlrDmk5W2H8IIKtp9jVIhb27Sum+U2
s2/0on0KgRjOhuEOuYTFn64pxmAbMJzFLWZMSLNI3d38+g+3QKerGi5nsoUyIjlyOaxeqdQH9deW
2Hrik2Kxqk1Sh2uv89LxZMii2orK1jRaGDvGv0OMTeJAzRgkyi6uZX9Ii4pELF6qFGOEhE79ujp5
ASWij9azKAAhwtAt73MSG5I81saQbSS2gv+lPhEACkgKHVv+NM7JwQ8U982LxFUJ9qpjzECoA16Q
uF0JWuG0ZU6/zYD8R3H9FMw0HGVjtnDa5skhSVB6cVKwnmJhB/5Oq/T0XqzFkzTNMQfGoWLiheck
wzA3N+yYc0o01jZPrNlr+Pzt/PPseWSApftG+TTJ4Mzcjwz+YoM9on5iK7RsQL+XztUoa11a7wAM
wwmiLmCg0i/mQaZlJbEu9eLumQX3TYP1w64IbN/2hHlZWbwDbtbRu8LrZKbIqkrcMb6D5R787X5Y
viyfBFYNRxybu1H0/L3QBfggXpyfjraz89IKlA+PgBF00tF0LUnJZumXl3EHpVkIMBbUNnHTCVde
hd/manO7e92LbWewglIH6gKIElolECPY/npBgm4aw0/i1oRuOyvH0n9FYYHFfLRsRSuWFsrcWBgM
GivmiSwQtUMH/A/5xt5TW6+GKoFd3Cz7mUwvm0fj9CXlKWUqe52hEBPiJ/tvc0lmIbfQr0azq13j
mc03B0Gpl0QpC4UktmAKopcgzvRTOZ7ggvUjZpWQj8qvmb3hr+RTFopWCvaboyk0YI0Z/LpUj7O+
SHOskatpKTkNGEsm1ujkt/GUy1PfqafmX1Mtt29hmpbzuZuD3nlUvASt+R63MYG+ZUp1PvP30dTS
ZI6SmgUJd7MFANBPjS4j7LWMtTVpYhEtthCFQGaigUCghUDnDyRh0z51smw4gnaF6n8oReE58AV/
/9CHsPKk74w9Lk9IqEUPVJwyNZ1Sc8vQ+EKjNwsuHmmRJlHAfDTLfLOr6TP5C651Irv6H0KGNeQE
a3bYZD9v7nl7PExUGPrkKyb+WrDRG9/efXxpgT2QpACBRcEAcW+KB1mXY2px7bYUqUpYZOlffxIb
pSioyyDMvXKmMv3dmUgDVeaOvLjxEEaHW494qGmSX+e5u7wqyUVAig5hRZaLmjLwCOaSSlcNrAKF
WoLWCKKy206/HWUEG0/EGYuTlMRTVxZlUCgjGSM79OFdWI37TZg64p3rmsTPY6JtPwiPBC7Wkmvc
QSdrCPUvV4VDgDYQSg+0Rvmf69V3/mGfVmYcJ+fvQjJ6RZfAsKagogJpcsJZHxu4gXPaGvh4cEBr
iUeEoonktOmt5P1Ctc+xfVFUMD7FduK7wqdbK9VfEjR2W9s2gpJ7GnO5K+/G/RSi/CwEzt+sqzGH
CfbMLOvUFZ0Lb54WwIu+Md4ObDN/Ru5abzSt77wZf9ykBpjNzUXQYQz5i6p/YY8Haj6apC28yMw5
qp+fKp1YKJ3sQhS3mPLdydpwki7myWwHNfSgLra09EzjUcRpxUlAo3Qgo7McnLBeRjMtcHhL63nh
2r43DAPTNUO01pRczdG2lS28jymU8fVe2tYB8GVeRCpo3PN3oLr8Wxfi4PiJRwlaOTWV5FCuWGD4
xMAtYBK9ZTnVtoLA3K8E7kU3aH0Owuxa5N4by9tMmipyv4VLjwpZqK7Rxuw6qChc2E3efDry45J9
9CQQ+2C/7GRk0pj7Jq2HsT/5qorcHGvO6bpU9UMk9x3gMA9j98vxlTlDn/GLmIIG7MleQ2D/P7cX
2+CTbqjOZ2Tid1FarTMioV0iqKbw9NWYWOQKdDCsIaZU9+hsRYSxyrLSqV8zfRNAa3WT0cC/xUeW
7eBz5DvreC1BNjyNIhV41LEvPU+aUqa1HRTdCkirxRrE2rrTJMVuWRIFBNgcD1I7N4grTCBZF25R
6xOiwisM9taGy2VVG7/YKWcTUUwmQxoFXqWLSTdV6ftB1dvd/bMkuHCcyhDHarDRVmDNjGDmPmtS
6Dn8+zXsjxJL1exTtMxkPZlTqPd0fTsxI2FR4ZQJdD4gzi+P4folrV3GQU+Z3hqlDpG4F7KZvfrR
Tz/m9SWCIkBWyV5KPgMS4aGybBIWHA0tzNB+kwRzwHYhQWnTb6ag2HtL4gGX8+X08Fv/yQkbRtyI
luHniE9BiTrAcDYOrdUoLoWcgWDM5n8e3PBCgZ4i+/VGP9+eSg7BmtpL9A/i6rX6C5w7723VcWXX
hfmBKZ1+UvyhtNtk5543vAOsXE8ZKpliC17wa/05khR8fwUa7ABZQgCFydY2HLp3JGKXMYvCheh/
2+q5yVKqprYOMxoLpplytbWxfPoYS7LXmKmCcgLtmBLyKwR+jl73cxxJlTGPNKSEdIplkqmg4rWm
qYuLvLfLSMl7Ykg+Glai+CoqXrqeBIzST5KNMlRCe6hroCQGp5m5jCdOuzwAKaRUyx0c+KHnpQYc
dxLkh27h6h8refQIEG/f/0+HbIocYcG+hFOmcafvrnzXzJipvF3TgxC5umSFT42+ABQUlLfZtVdO
umiOC5UstIlgq1PyzY8KZlVnxOf1NcHpch0fhEHDYFjkeJXQyHjoNZ+9yZ166rYrQ6N0qN/AkhJy
q4dCllRwA1eWTr4WfB0f4eLhmT0KFAeuvOEnArAlusAjZj91AIGzyvPO5cpz1uagzIpbAjjhuUKU
A0oBV/nurPWkW9JNjrniNX6xkiRwmfgCv4xEcZ1u7KsbY61sq4fnMSU7sdrCaXmAHpU/Ss2OEMWa
qHpZTaUMHs0qOa3LwnBwMJq3u1esywuxS6b7NMtQUvlm8f/4wLHHAyorgAnxsgdb1ubS8iQ3bhmk
YgUAI6L3wgrhnA3HXZeu7khxwA5Qf5ON1xoEEs8tyfj2xIrQ7faDt4eVVnae3UOQMgxSdfjNt/LF
ky5Mq8CEJJ0TOchJZvX8iwTZY9utsPcO6ZzUS+LdstqSuihzKpCuDA756subcLV+azr8vm7KEIrA
Q7y63aJOQAcZbhdjSOb5q5atES1tTu+CmwysEujxXCm3ysvMCbhPtNMiG5JLbMjly/hGAfbPX1Pg
meanDxmJt8mxS2FvfpBC+cuUEuaI7jSUQNod4Mr2k4k8wMyFqzBdy+Pr6ouiD+JrZcVu13J/ENfB
2Lc4lF9T4b0nBoUGj6EK+M3OdpS14dKAO1n8932GPkF5PlV+b1sOJDZoQv+2zmPC704k2zNoLXDv
Y8foaanlyifXetULhj4nxsyKC7uwMp3aZprQtPn19j1LIXHVGtFtFoJgbfaG5FY4VnV4jg7bd04L
2460bBunDORMlYUE5Zd8or1M9asIvAA2WVm5RZYY6amsJzNX4xfaHOuprge7asiqt9zfvkNMdgmw
r+nassCpjXnf7K+uzK6w2cxn51uHKqaFGkd5UEXNfsaRj1QIOWl9eB637jmo6xo/r8uF5F1mTNa3
+cvC17YdyX+4aeLpHvniVq0AoYgOnp+DvDt/d/QPp3yANhMFtYbdQ5jocMvnJfQLn7A8pNeVa7vc
7eULhujwY0TZcn0IHuiBZrkqRBYu3wnAu1GeXNAX2psVUJkJJFq13CQVejQwP/7DhPdihsiAwJFv
6B4yBKzyALiGioguzvYbcNOEhkBzDkXY0aHChPrpBSsgQIeTRn5l66rBJC5+ChmoEugjLbIfjHu2
Rij6UlgiS+ba+2YJOgchj6TKtX8yT9yIC2FGtpQWpafCty42iH3JthM4+JEjZJDbK/oNHW32KSXX
ykOQ+RVxnxfQrYFXWSdQkb6imMtga7BSKr7JTMFuHaFqoAAxrSUiMO1hVQ7S95CcDPUqMHChsrgt
zbdiqH6e9gl2+/0Mtm+8/o0O8Edzj/Sz0j5mVVVpA7r+mcPiV1xZ/HtljEYv1wKLyi1mimmA0CNQ
HBJxgLFHq5nt8A9BKXMJOiYGxQ1RGPNCHpOYYb5/ZE1qOubTGHMVQv4KS3BP23km6oH5tDRM7joN
wc0V2dxC7bFOGph+G3QArTnyAM4AeHV9YmiqTG3HN17dfAsdKt0PWESnc8yzSm3kDVfEJDtTAHew
i8G/7fW9+p0S70FpjpOz1YxHs6dIsGnOpli+aSEKasXmkKefEHfbIypRkSFcIsKh1zmb46Mp5Fj0
XRQzcM+bBCKWeg4ig/yCwgaSdnCTS2ZiPWi5Q0LGRRho8HCIMmMUsku1VhoKT7INy+MUPkQx2cMZ
UJIc2kw3tiytxg1nq7NAXfr5bUUkQ5dvSSdlttOVf61yoMl0FKjq0gIisDYN/xKzdGqir68tAqEq
6aSy+hyhQna51yGX3hVy0JG+Qrn2J/tA2O3B7SRJPDTr88SU0RwdsAQIo46+kMzj1g4QAB6URXGx
XB5AA/hlXCgsvJAFGuWJBKAPhIsdPeDOiA2XXnr0iBVSIuUSenLKLsib0AbK/QZn3pfGE00/G/Vk
GUpVSXwATMPqPiW5rbnXR2LzL8sf/eW5hnNV74OqliP2jZmVLQ1pXLbHaDwj5HfyTSq8ZhBY6VW9
Q47fwyrB+5Zde/z8FYBh/agvvMWQ1OZ0gE4mNae+L8s5D7pn/e1mB/DH1lcd0fa8lWq/gLoygWEi
FKHmf7orxUqLre+nH3/DO2LCJ/BBNDWf7hWvE864MPF3UyVATZ4qo+dYg+cLYOFZXdE9hzR3o2zo
jFuUim1xEws4DzLHtj5FYBSGIQ9EHead/uAmiItIJSv80JbC2kfcATNsN3q0K6MwKqDZp3W/KBUF
tPINAE6cpZZSlB5mNTfubsyXepovOJOPzaBsasi7y1c0ixT7y/jA43zTIxEQH/TcmJyB5V+Q3ImZ
r04y1ZHvudC9pi+k+FruDV0T1fYXVxodlRrHKB3Lnh/PwJtiBiDvdwceKBOmY7ATXdg3ze5SxBpK
VSkjL078F2cCGQOvTOXDmOep4YWWUhQCXdjFVEBVJXA9oCvkEyeobuXjzGcgpuxj2mZE5wVKh+5U
LA/fzKLljt4lsXF/kMa0PApK5M9FtbtPioAEgSXTFa+4Ee0t40wayd5/xiiQsdws8R8HXAHUmQsT
N4yfn+DH2cX+hWqn8BRax+WWVgbx830bWOz07Kv418+UTDNSrBZvK2H7+molk92usx2rqpCONfkE
rEPB9iqCVZ96lI8hdaRr15JcDBiQp3JK2RSQFhB70KjTL4ttvqRkYOWCBZTIbFHx6Xfyql9HQx6S
huKdFNP/W2edjDlOQPpwubk/RpFTOOWnSrDAb4cowaPMuiZ5ZlXsFHfmxssF61NRmWVPAUH+zF56
q0fxYWU9Tbzptk1D8V/u2MUHUNP4w/zz6cTVhpVfkJ6oPNFecNhpbHbzkgPSWM1UmXDZKF0Ircxt
PX4aiPG0Hv8G9h/ZF+BD4cdh59Utc6Ajn1fZSnXuKrzd7ZOFjwKPNynp/DflaUmQ7QBivpaiqOIC
UkDYWcUmz5xNxwQGiaOmqcYq5Vho4eBj/v4/mUZa43hmQfXI0cJNLO9muyxtqotmwLSHTCBrQ22z
9CX/G6ej9onsB09Y9xVd0kLpDdXqBGuw27Do13b5pl6UrT0+0ifEwnDv0tkyXPmVOJHoSoha2O0S
QU4YdKBfEU/vyjrRmJwgHm9COzEHE/kUD8+AYjFd46k/IxeBSP096KkFsX2tXJM+YEcdCCRo01Wa
9UtikQk6mzApMIW/94TJ2v3JIayVoZBBtnYXb1VNMOC2rk1BZAL0G49lah1+DqvudXojvytF8J0m
a1iqPjF0yj1I8t9jVRpkRi3W7otZ4W73mv/merXauZV5wueVm5nYy/V4JDYoPvCX1MSXBDTbgoOJ
9HPLUYHMnIvWzXpMmR8yXAng1Qk5ppsMntIrfXRhrd0/UsK/98ooFYrsVfIuOvYn6GUr4OKsbx5A
o72wg27BQEq6pCLwIyPHMMA06/bxAK2rNp8EJcfu/i4vfmT5XX17DFU2huO/8afIUB8Nq4YxTgsp
poCOyqznijs05B2XbUu2kiypwBnuCuluSnrO/85m68VUe+2H+FqeKdzUHmIsse6nrABVu8lnTop1
2+z02OE6SZzUBwDvLqNPI8YPPMOjnRv+WcLR5EoP6JN8DR3bJ4wKrsXX+/9vn3K8Bki8B1z8Daq8
hXD8sTWvf5cSxtpmk8EwK+onzLbMCHb+w9u9XHuC/v+KjXOoP/AuowmaQjEqD/60jLAayiZZq1BE
XHdWFo2WWp43AZbhi0f/JacwSljdrOwKMbfYeBboHNW/mUAS3mcFjrVhdj4TMvqwMBbyyxkKFC42
3lqqwGdNG+Jawmxe0NCaVPx0cZ3NSvl06RUuXt0gArrKQFfmvKtieY+BaYj3VkIcnmGrry/kDFXr
8mM4brYa8L5kDCi++Aexb8EEwdwhkOM4KVqOHZ1+StfONSch6eL53A6JwO24tL0wnB8gJdkKQqhQ
RfeokVwcjTr/5CtdyWWfh5VSWgw4bS+uVJCc33LBH7iMEbtcLDFQCDhCzWrTCSEsp36k8SstmjJY
30FHDvnA3/QNwlODchT88qu5i/IZx5oMX1er+QTbmIOn/SIIb62ke87nsPsL6Zxjrirw3f6GnJvr
vvNnl2ey/bgIGht2pIZFXO4HaBwQ0zCC5T7gGWxUYGmO7i9HQxbLoLfLytN/3LY0FmJirB+rPejQ
QkYx64RwTnE82RjgRNuuTePEU3kqX83jYxsf2k275oT3jwdyNhFQ9At72c1NYJ6rrAEuOmOokumQ
rK8/30JMtwrtYTOBBcZhw/7BfQyHAV9aQzu0i7R9GlGuCVIrhPsRH9TYYgBtLQKx9V0VNTJsbCcU
RosQK1KuekqXLDw7PDrrUrScJ3FHMvVPfH0Zhepdw6P4Ts9x1jXDISxz63QXMn0tAeWrh0rdSXTu
7M2E80YrYpMVNVDkZ7Qi3Eb/CVsalOgxy6meDblRiB9YHcBH9CG7XGKjiGKt9G5K1RNwY7dFs+vc
Qnf06iZa1oG6w1xz+C7Ygez9zLnMgz9FPfkG4VpkxhN7rTjzIXrsReUuof4YiLO5WShgem17ulDZ
uuif22shLem07nOBSzhhvPGuDPA2cz5FFzGZBrZP9Nwcl4nUrRu/V2JXC+v1S1e8JRte70stkvhQ
AUZmFvryGw8CY4XiVcB9PbZcxdji3DdOsNQW/QnfYEopq1EpNWtw5nDxxcGIeTeXT2Sep1vEBRAR
oYlt3ZrnP5xdPR2KSqXFBZxC8kMi9lmCmsI6zXFpvkxgrQU2rk5LCdYr7S/psPldwQ/u/saAMerS
iMy6ZSIccJshpAVwgzoJieDJusH+TNVJI7Lq1s4VqHl7A1Zuh0y7ZAh6XFbUm1SKeuGPQIl6FyVB
MDWVgr3LWIqwJgmhU+v+n92yR5EM/BSf7P1HEXaiGyEz8QL8X4NNm4J34CKr4J7yykyqU+jHyHWf
U9YszpmUMgokRdMrgvV2qRWxoJvMxg8JNM9qwWFBw7qxHkMmJib4+G/KveiGB1W6EVvBGfcjDKyK
/OVYOA8cBS+okKAIhFbwkxTsaErx5okQtPQu1OprnIbMnZ9qkEj18V5rteFp554kVp245lXtTArT
qJ3XSok5vFvZ5icvfVgUYCC375J2C9uRZPBEc0unALoFmCZF9KJgBM9Rq5DXuXescf29nnUm1nAk
A2WJB9O4oTS/tDN61CCmPsNS1VM4DdrWrihggmB6ySDR/euTsnJEIgi4eTYKttDCKD1qb3apIvJe
apwKjMP9iJT1faq59gbFGkvMmObZgnGmkpTIorfryKU68/S+/3rDamA49xwPtckrBmT7mLLfCIrS
jQyvTfaX5uH+ModbsTdxZu9FqmD8uEEvltSZLk3ID+ujH5vJ3CYsONpjsaTi7Cg2z4q9NTYJyD60
XWgUgOTbh8BmDiXEImuxLu7OhEBIMCVv5Vw1lqdZGpPwI6LIb0n2OMH53kK+K6x3vWPmgahx9gy6
J5gcwi8tG2edTSPcrjwqhqQ5Xi6blE/6Mf/ID1gVnNJ9VFpKI0K2JjrNJh3S+REYJqTPCpW8az7O
tIQbN0oHUZ2jXOQG38M1g9izJYtfxohH/GGDYnKJ0ql919zLyveEeUL2S8A+gBpWqGkQsFgOVB0/
1QZo7jKEKSjtJcSpRn+M9irmlf9owH1g+NUEU6ONGckCRDnbFlC3t51wXFWqXf8czQqsm2k7JdkG
4oa268GMe/+lkyvgnRljGSQqEbbckF5fYHzXcN/ARiJhd7bKi9EcxJ2KOGNmmzYq4q0/3lU+AtSn
T4rVK6E6VTtchyQCpUWw+OMKwC0RtwQ7FMDXa65Zel9Qzm3x+rA1VOUw4cj1K6vu3tbKAREpd8iD
mdjcHDU2dVbkt8nVFxXuE5euHKjXFxweaQ3pDJW0eGPBv/1lGMbf5gXbVCAQJ4XxFH54cjf8743B
WwzgIydaYCyHKKXM4jSbgcwy0nU+QQft+2JSSmUHuWGVqamZXtc1BCgOJ2z3OO2maWn2x2KhGOJS
oQ0q3zlEqGR/e6RPi3h6VhGP48iX/K/7yQXX/+ac7N2RrhIIrUBKgKWEsPGTUtE+ZHEvjEJRFq5c
v76NYFnMrAo7hEzuZoDKcsmu5LGM5ZqZ0RPzNZQKvzg+RzqrXpgqh11Bw9HKQBR/YPlKsmXPiU5W
+kENYQwqz/gk0P4R8lWJ+ovA37wMRpW0YIDKEG4rbGnH1PSSDET140o0vjMDJfmXq+J4bxdjQGz2
HLeQ63AtWqZ7d8wCKBDzJjsNtBvIad3DzucuQMbvXTixV5qpFVDXM0v4PEv3RJm6TORZQPWSnwHY
C7XkTQTrE8WQcv9dvcZSn9DInky4tMfnpLb/CYZng3+AdtJmCaadyiBrlA54BjmUw5xueJEmqsCq
2lROfuaHSdfk/PxyHumkAxFd5HWM6XvYRpclu2mSnmxNuZf/gauNHwvYZnEiXhtzild0buVKSyj+
V25zn1YgMGOBmbs3hdtnY7D6AB00L7ggGETwrCqoXnq6DtNC5/jYHX7l4NYW9OXExoKMobGJp18A
HHD9ccGa4s7Sk+FE/JA0ZTkgspq/2y3PKCToWIRCjGmgd4rVFmslwtrXwsIbtbDSvp7uaf9g45EF
On2qTTGjofO2Z7ng/VrXaqV1YQLOJOawWKbmMEGFZulv774P6r6renhK9oOIjXZqLO0AQjnGQzAJ
pLgn94QlaBFPzo70mBQbWh+18A//4P9QSzVqv+4FBx/QqaUKOZTUe+P3ySPmPUyUMjq2DEdm96gq
IgxPzWg4ay5sf/kAojBbITfqV4ZoMSTkHCx3jBmgCNbIzhoQk991T+fbqmYFKwX/RShWXxociAzp
6U54TNxmIXXb8Sr4GLn2Uc/EQl0ImyvQw9GuhVr98Y8MjOdOZ5BhXLUM7G0nHQnpjlrubOn0RVT8
uQ/1AiCkjls4qKKejD7dmSeDhomf7qeI6MIS0CgvhecXfGZsK4vEZeqMfj9Nt4jMD9jO9Mzss4r+
LqnvNpE7wtt9NGhi9TIl414kwajXcJ+7Uy3WhEviy7QitNR8C4Obm4GWX1USKC7yT97f13oYa6bX
DeFXfxPObtrpFxkdE1Mt+5M6vZSHHt+x/3EHQyAysx76C+CrcLlNrrstSQBdWFVAqcP0kbJLWcfr
8MZgmmk4ArmuEBoeZ0Ts+Kip2/eo1QRrJG4FScHObirLyF40o97HBS5teLQKp+Ol3nmxnhgSEzbO
UIMwbLNV9kbO6FB00XqsZOjdlKOpI8B6P6u/kQDHJJKtNiKO5EhqTURo57fMAYQS6z6+3NBY1997
Cv+im9GTrQ5usTn1U33azd54o63E4iSzbBpckX0/Q2907AIcEqEdZk27gMfUijNVfObaOom3TQwt
nKlAI359otKKPW6nYGDzPr4TjLzT8JcYw21gld1VgqLboDOtHdxv83Az3vboyE+TLJgRsDqGCWNM
en/mr9LttzHsbCy4FuOqLI2ValPAwalfq8zQF0RWNFP1TgG2p1s5CvvZj0lKp8joYnoCGsZkxfq8
CdjnXsgLz0SMMDYx03H2EE0rqsFCGcGQWAClwN36P9X9NGWICEgNVpne8wZ25YD47cElVhDQW+Jn
vVP6wx84TnKPJ60IqoZlKaKCxRHP6hiUDl7ybTS5loZ02GwbQuiV6W4UgzByh2OZzGJs7TpWIJNo
Ms7e8jaDssglEBqrsN3uNL4z2Xf9MgN/1MppGAun49fVUVpnSRRjV6Ykhqq7ilhOai73nxpB5zfS
UoviO5b0Xfb/Lis2M9/5gM+tg4VnZ4dqC5/J3lrcCafh2yONV+o+ANC7mFKGCCa7Zm9tt6QqWSY5
bBkPx6Lw3A6O7riKPj09BDhEZpsT73k/FD/6XwTR4SvnGDthtsbc0x2PVun52lzoNGCiijCtkjZS
0SrRRF3uY2h7loJ06PskopA4wP1YcaEArRslzqg284YUPkgPsEBnvF9pVXwRrWOrfLs5N9en4h3u
ZE1+JVT8i4nT70m7K8eSzjkU+/SnbqmFecfy/EEgmHUKhwTabiayc6IoDouUtjYaSbrBlqDvCmcq
S+ko6TjZMBO04M2rqpETBrRb1K4e3Tl3olCkCMlF7ZUZFnG4mSrweA2DzXxOrOoR9k1zEk3NGP9H
M2oF3HiekCYV3VJz3QeoyurJEhma7FmWLM/v1vjb5fyYtqbnmlg7OsjhQtVwFQ415riihXxXbUdC
Nt9BDJwQZsbi7NFYiCz2OrxNwpnUVKt7ox6La3y8ySbyXWSp4Ehq2d7zu7ddJdeklWOiLXBkruI3
VtHgS0qCguxjmYCW3hQpCceI0HbVOdAHthiho8gpKG4p/rrPdLR09tDhLiOTQsi9iXBt/5XfTdHt
VGarrkj7+XkRbF7/qVX7WAdPv9XYlloVMwxildlHWcx+CcitiEZBb9jnyAc1YFPgM15amCIxUTAV
K8qByAQaExpBSldIWLPh/fy7ONhszE3Ci/eDL4pE4G3Gt/J1tjjdTinGdA7YXEmWHJmYoxLzdaqq
mXUXis+XUDAPlEQCb5Yyml7vS+TBrbHzMrrnuIJuXcC4bvGO0+nrZe/kPYatsc4XV5dS8eybzEYp
e/kYQQgSHQvWZn/PLx4vQq9mEgcLIwS/NQxt0UJDZBsq8ibeVPbP5oMS7DzJBkceRYfOiPPZklLo
uG8KVEErY1USHiJK+egCDZ/tZSJ388haJnum21q1FjWtJYBohLX4CEi6RVof6s7COgr8vfrzW3ef
/Dn9wEPoKsKyKgjZXu9AcR7D6iTrlojKUfAqr+KG3Iv1hTSZdJr8wHGmK09NRxwE5LvfJiaA95nn
WXjqaJnDPqArp0WIvbh7tFNwpe7nxyV6VzRsjqSGuZNnGV8TVvBN2usFNgtbgxDVzQeAQS0D//Hk
Gb0zEsTY6Fsko4n1c7LSqBkuKbnZkReF8w4YqMUgD+2XOpo2+W+v2oMdTkmaEydi4d6lrFBRPlmm
WLgmXK6xbCYaf4BafywCm5QyA4APAmVD3ZpJS6ao+QTXPPpkY93p2yRdMwIPMUd6xlaFLvyr5snz
NQDUxAYU0hht4yM5skxZLvmGkaZd/e99iiLb9Ju6YnqvclQKRGZgkGz6bRQkUJVzoHA1CLlLMFh0
IOjtGxyWscIt04nsJWitHcK1anEf05fvuobHcu0h1yr9B6cTYU4O8YJ37ys9/Ct18OPjv6vb5jaV
Cg0o7nVNzlzffv3J46ek235ZL8f1RD60MNkzVQRuwbdCSAt6N0gnQnuCtQUc3SRrChxAPjKW246u
IJ4sKLTVUUzbr5pcLfid6Ry5LrxQ5RFUlcKEml2EUiKf7W26i5uWsP1LNmkWc+svc25gk+LxWwh1
FRBERzyqTjKBMmv+qgrqBnucSTemraQ5v/csGbWhZSVzqmYXAYliQIC5pIWneNOuyT81D/yxi2QG
JQW89yn7l/J3w1bNNfS+loM5ObDhOUK7IrfiUur5L7vwRFvlOJlWj/REANZ3LL8bMNIxS2JaDDgJ
A+uD/aa3zUkb1alytQpCxzMxALz+Lvn+5m5BRCnlZfPYGRnlOyKEzwNJB8+3EZ1tE3iUJvFjN4ya
kuXDBe3NfHr2TpEXlZF40mOaKLqTyimilZuDEukc6UFH8Mh3LhCd0mJhreKYcwCVmkMsqMf07sc3
qMegPlSsEj3C0pZP3XdYbhBz+itgAs0rlEfc/a2YxG8bPwnjhLT/pny1oG0UI1HO68fSfsdL0u+C
2bbjrS4cIL1XbT/yVHiPj7bgWxW+/hWv9kl3hTnHYQ/ulj1OshqfNVKSpNpzkvDjkuHF3EHK8l6h
/UATHfx1AZepLkk/SELu+4LmxJmGzpuBzHsOG/3/miCdCPC9juYUpPl92GiYepEhkIR8DXR7YZTP
I0z558n/A6QYTINmKxbU/JMkmFuGeNBIMzSNkNKST82tk8KlZKEcTwHUmMO4udwgUhN4g/G5x4A3
x4NVZcYRkjRSyuljCITi1gGGII7q/qfNLr8bFxOcWgzCmyXZ5ApnXZTEy8GhGRpdK5Th4cLR+jo4
55xT2mmZgzmU14Thil1Qlk2ZX5Eekwz1+JXUYWfS7ej3IVoUrBht69gTIN8OfvARhF2QkBPUPfDW
MSADvwlu9UvWZ+bvjy21OtYDrGDqgqDrmY/rtVOsbLMZ4tBMxVU4nuq85iC9x5AGuSweARvpIM3F
zijjhAe4UrF1B6yHTaDOzRLJJRtw3NPSHXjp6Tk6ZvE5VRiwsAi1lGKH0x6/Ldjy8tbqXg0eccJj
oz6G+r51XOfUj+hd3VHDxDVQ1z2dQLTU9guwAdMYOgPHEX91YNMW0f/MdOehL9U31G6fgu4lwndk
WrOOFw8o9aTA+9siKys+BEdj43A9NS8ism+oKd6FSmoeYUl3icgcxGucA4O6z1kXom20Aoa2j4tr
b1akJj0TZpI9SACnE5DBblyw3RCxHbQf4BmEgoLtoyBosMVIVKrQv7MUtIAHGzVi/JS2awpXEDI6
OLNyrcF+oIeoCfn3dVrsbP97bip8DjfnndNI3fm8br8vOUdRcnEQlh1enyde9/qgaBmN1AFO5lVq
qYpeHLmdtl3w3GaTQ4tBi1vcB7jzVuRAI+8k6a8j5ZDjtYqjcAhyRyCKf2kaixzgG0Dcjeip7HY7
V2DL52Y5dHG8SyXfof84/YsgDRltYipZkdudnf7e9kVU/3zeXLBIp41qBM8fBdrdEtR+yjkG8cIe
o0boE4DeT+6Kw1T7uVXAXHT0/QCCRdHhzqFyTyFEXk/vs8csXwjRoRHKn2cOnGKMZnaWOGCg7oci
PHYYVMXofMfJ6CN7Kw1LAIYITL/tYlbirjP4zrWZk/aS4k/7kz3VTmBbj3JbMfU+1HIS141w28ij
/ccXulv2uJ/gXTis0uwvbOHdkEnom3gEgdV1AxufkqbcpvT8uvygtrNu2JAmd3rFJDWB/apPWUTx
wZHdw/cIuCkGPU9TsIOabt9JZnVz0hv5gx7osPstLsPGPrDb83T8/IkkfrKwLH6vWbtVcG1if0Wg
53iSFYLXqyrT9/0aYrpp58WLDi9C/HXm2GkHz1+BeWBG8T0R6EwAxDkh84hMUa4i4eN8Pe06bIC0
XZi9XxZcfAAcQstJwceQi2HBRnd3W1vGkvxAw1S3vyLy8KH91xCYSa7/bwSqSFmqc6lOQ6L5CDBP
8HR/4dZXUqUmqmvofMt7IeDgQI7JRAGB+D+7af+9qjC77iTTSwdchCaP5GMRZ00zKf7Ob2NLHPbm
btQ3JOSJwh11h83TlhWgXgwTh2p7VLILzHT0g+ghqStnr4Q1K88rONwUmLuuPdj5dKGzrl59gCUc
sU22N8oeT0sVozyI1hKmKyBhz4spNoPt4A2a/+75C5zah8yYJC2YnAzH6oZDeils2MEPS+guMvaN
63pXmz9Bcb4Ll2bJzIMcqVPn2Cvz5n4TPpNCJjkYMmkEQAJWHF20U54YILtyZIWc6bIh7GvmMGZR
xTDKz30PcRJr3P/oplldmvElW0ohEkdn2eF14aoRjGVXCD+Dm++UoEbWmvMtw/FwFktkmc4R+j1b
w47wcNxf6BIhzJ80kv7VE4uilezdkTFJmF6kb1AUHg+L6RX4PiVgoU0i3oqdyVgQwQ63yfNdWndc
v9SOokEr0enkyVNXPlJbldbEPWNwCJWhlYZyLRXiAKW1Aff8trC9C8VGBNBzdYxTDcCjiwwm6zEl
+2Z/J6MLdeKbvf+MVJ0FOKXOyOjLgNpaIEOB8MHSrTQO/qDvlxA1jm1c1b4l4GdmJmZhAJ9BpjKD
i4xUIJXGfIUnz5hg5BPYBcya2+nk0RuPPnXjTl6vK8oB8lpe5L4S8ybGxlVADuN4dZEhE6o9KPT+
h6XbjKj5R/xthVDN9SJmfr+8+zTK/sSRs9TnAoEiZArA5xRECNSGaESjExghl2E3eOKOUvXyvzri
+ix6o11n5Tlhn4+lf0pHI1E0zB+bgwry487KJAOIoohcjqNXfxmUTT3lk23So7zO+JPVt9CR4Uob
MtfmRo144fyX3B//42sMj8OIEzraswhy2lfDUob7C8I+ubVIJljswndXJiLqsIZrzPWLDzrcWXMU
eQUG2y2T/eqD3DvMu1uge1raA/eIqiWp2qcEOSt88JE9KUmWAOuBX8Dy9YbXcam/CCQOhRDL/8S7
MAnmZGahivQwhyG5VZIIKTiaNOC4SgaE4bufa+/UGj8joTzcbC4tHZjKYvkw3Ss9uptOTPJReepc
Z7g99D1g0E0ARtcFhq7uu8u58s2l5/cnMFyvYE4zv9PHaki1YkOwLMBN+mosaohVDLR60RzeDz8k
V3enKKYkLYpN76s7U+S6xXlEaGJT0NVwEATwOQ9ENmF6JvSdBYUfElXHAI/2zYKQ2HMiuJQyX0Jd
H7ffpc/p6iYfTlHqFyCmsEKSJg17wW+XcCCkYFCkbK/JWVRg3rS8C9mtrIA3dcxXjnuGP//NUW2Z
Y59zIHGfxigig/AB0U8Cd/4g7Tu/zw539sZ4/J8MICQW9EzpqoTDbcXYMwZd7CCWGD6tN+geTD+z
gxCpkhNIfvY1+f73GYVlHzxPH+Qn3B2vrWjQH7TQU/iySjLeUtmrGxEXMR2Vvijbe6+xfuHnzCpo
JPpRfMopG0dJLxPVwi9Rmma/ND+nMv85xYrDu13Efi4a7BJfujRj1FQONDL5J8gmSOV2eFdHb0XO
eMUjgzeEhNm+z6IFGpaWM8WdwIrqf6R5Mnz627UsErjDTR4YvITfsaVBt4azutLOKbWXl4eeLMur
12e1oZt1JDG3mPtZ0itqkGJ+8mj4ref5XTMSswGtRniwUhYbVTERrN7pN2qw442RiXoVZkgOzCNa
XsldHFvrs6k9EKYWd19XAHujGdhk0bdfBWnQrmiB3Y7FSX2dGrTazoAc6gK+4ElmA0EL9TEwyY99
Jw/Q6p5kpgvd7MobKs8hXv9uAXy6+J/aO4Hvbar8eJzzgmkMB9+y5Yf/H7YenYaELgTQq3S8zhQR
HhU2SUzqq/AiA98ySPP4Vnsm49eTtabq+3kZUuOHQZIdV4+dPXdMyQVDLYwakiwULJwXtY58RTVw
keszPx3WHPduFf7CEvTN1+e4QekBTxvTRnDh17DbJBl8Pp0u9eyaUrtv1W7KoLx87XedcuMiSWwK
2b6PSr/y2Sh1xrsyMQoQtL5ElPwWMLkOge13zzCcHCQ3osKDbpjpj/ki2uP9+KPeUYIqpRtUgYSc
rUZhrk+PKjxLwYjKaRNU8HknzfJaXj5Nw17O2GsNeA8E8ArQlRJQ7hZxXClXVUJW+3kKBfROTZ6i
KYFKPXP/2CMRcbxhYEU/YTE/8/OZqaw54SkRR0DmouryWDPANzMY0UXCJrgiPO2rv3S8c9uhQG8A
dxnrN79YLxJmNAqMp73BSIekW9qSnnrRp+YEAkDo4pc+MhpVbODsFyzlO7N3gT4Ld/V7pMgbs+Wd
nuA+gpO71FNSPoKKmnEZfR4Oaakx3zYa/ulKNTsQBOV3PfFwIhPqV54L9NX+7aYpNm0P9aZW0esX
8IrwgeR3U1sbrpq4lBuwWutwlp4pmJh7/zbS5tcmzBJO472gsO/PV5ITxgBWR20SuO0UH5pKuNk+
mU+XdOheB10QHUZaQONR5hRG+UmtJ4hsLioxvvCjSUTz+6At2+rAAxx7zu4RXgPvJHfDZoXlYjkI
JK2okPXlT0+VGBvafFbilIynYd7/WDB3odFYJN0Tx9AQpUHDAqt7NdSycRn0ngyc6pxR0IOvMv3b
8i4fSlQPggZSX/Aslyc2hfrLrtGJ7Nva4N8jfOHdQjihCpfFhxhkPoM6Gr4VvtfdM6siyz2hmLhz
mrWzLmn6sl7O1p3ea1SlpWggRC63y4gaFWEoCj4C9ki3YhCOSrBsw/4YRv8qquJ4+BF6oS9CpUId
oZfBfHAnQiRtHEneMnPMVAuyHp/ynuZxVfOU8uzhPNwAR3EHPvdrSY1cg/qAKNEd0PhimCfBH34x
j+L44vqOCXHOj88tDP3tlcpkVD22iEfvMWTxoEu4EUQckz976XulVAP6tEwayfVHhNudy1ejO9Sk
0amnzoRGeL+FkoKQKyarpG97zVW5niCN4O5KxxKje8vkk4wxLHqK9jgTAnJ5oAMEXtAbU6zh9BlF
201nGkh2y/w3VkYOK7exKAX6zr0r6+kfZ+dyjOJKMo76f1uUmlQXFYduaZIPCeJyF+WRe/FWISBz
dgOpi7Nu+67G1Mw1e5REv+jCODNI0fiwpmDp/QWYLStFefweJsYfbH5Os9MdVaRC9clojVK6EZVX
QaGnbS18ybmWX7xJz80seZYUPtBUw3jHkG+o3n628c8Oa7jGK5bJAJ/Lsw2/v0byky54c/mQllOb
DQQpW1IgsO2AfGYd08lCirprviDPPYfKVzcF2s8eI2Hg0lsJ4pxmtAEX8z7F/zeCe60MwLDkQ8R5
Z/K2B9mPZh9ALz8dGG1efu8toDdV9A+PEu5UZ+7C9VS6T5K44GBolSEhvGuuxu9dtCKu/v8eU3/d
8xDGJxpoRDU7oIR2BQdmi9sn4BrXrFGDjNA2pODe0rWosVcNRBFBdIBbPKOpy9UBvQvZJldah6fQ
U5RkMvh7hQgGAxbTFxNwsa9R8lCicuqcJDWAyNTFUw1ZV8rNKFVJ/3ChBSevWxhN03s4X/8MpZSb
39Jl3oh2RXx1gN++q6z1QBzYvGLAB3FeCTa2N5yV+WMstAF15t+RoJ9PxGPyrEAC/vZWQlPFxLZi
cP+7s21qQ9G2NtGix5wKNmC7s0aYdDowB3NeenRDyxKzXlbnHlB9aDKFRa1RQtSVxA66ZX8aNbKJ
iBOkbdnxt/rp1zLhcxgxLnlndoIDDP0fpgFeWAzmhy2wIF65rVQtKxZg01XoGLTLlmVM+9cDFMPV
mwFW4rbZMNREMm7lMpZk2Y5mjZbDJUoLrI8IHgsjxw7NMhBGQvdhXeWRjtlx9lZYwLaB2uOBY7k8
CEcx7vqMgkWmXjDam34AO/s4+DwhISbeRSLDCWoKa6ePddeDomY5PtBxnYZgn2j7Ej8r8+wOjjJh
+g0zjxFL0qN6D4w7WFs+4tHi29fzKGyy4fKTTO5ZdlpSv5YqIHz0+bnQG7C4Hji8SWcBvocEUmXc
NvcQVJC6rZiql6DhVI90m63npH9l7Uv74e01SyNJcZl+Zy+y6xp+AYN6qxkyypQ14emzBnddVRL/
v7xauHxZUPjkILNaAnVOLVIrVEqUsOINqojlw0hJ5bFY+W0lqSQKHbiLR9DieDHgo1R2qao6v2/N
B2POWVg+iZd2KJDwqDVWKwhx2nldNsdsXcqAEUtm2+6yB/dpJhvVUhp3Y2Ybe34kIby8sS+310KB
BppMBEvrHljj4DZWQ3v1SNZ+3HQew0FEnuO+vCZrDuM3eWNLjjyBi1bFEF9Kaet3CM70Il/KeRc+
iV3c92NQ7qcHDvC4UaE/ejQwpb9MDu/ZH6Zcyxq4Irfd7iTWnd5oLMjBqsMCG2O3yzuEitX7hHD3
3euFDfqcXbvYQqWYJ8l8xuZBCT1y37KGSTwbAIK67vduD9vw0a5Jsd+EBjjiF+lkDKrKszqDcn1n
+oTcbm65anx6wjDCxiknkfk7Q3uvIWx/f77qCtMHv1gptr4ZLVpwJ3jk4CcwJ5GOjE7DKS9ETLEh
fmqZcCaTT4IDi3XSoj9ZLmizTlj0kdVFQvMLCWI36vIgJlebGKn3bKa/2ezgQtC9qXkv4mDiFzJ1
2M18VrZwDlDnMWWDKpXp/lwOmaRSYRXcoV9Pg1D11M3Qu22pXaPLnajzW9KPtgXy0SVvX7OggGZu
jGDRWScAu9VePkWk4yzF/4x0lqnC+Tye/PH50mwlM9JwS50oNUxJTGbMwnxSL+l7daI9LyPtmj8x
D7bH58tuIMc0kq4N19G9kXESPq2N+AszsKK3WqZMeu6sUNxW7GzEyTpIhtMQRJda4u9jltkvLe0c
d2UTAg3Q9Pi6p6RUsXYoZ13K/f63Y0m9YUyCb5PauJlAg+rfC2u1mCZ7a526kesIUcD6pWig/1uE
yPQU8ix0thH78hvCalSfPmu/Dwx0U82vJaiSkJT4D8IF/AFjlzezIUL5ohveoWs3fZLD3t37aOL0
kNGIyGGhzlFiSTREM/uWPlLk1PopcuzGdBiSTqPLEiEMwYnBKXhC6Sv52QYTXZZjQlWbZTJuemX2
YzGX4yUBF6YwXULFDKBOegF/HTyay3oWyxaNuK7AKAnyPbkkupjTT4bwxQEtIGVaV9N7GrcU4itk
BJv5mvwPTqx+IQCMUnvzoUwJhw07mHPiZYhXNcXjOvgjUxdmXMgiUX6jdC2odsa3qtQmSm8Gdzor
XjkMz3lgtR+27FXJEhuP++8qoIBr6iqtR6FoNmlWx94kdsgdkNAtCrcUDqHbRD1ZPvp/5aPFDxq+
y8fw4vk2TGtZgYLdN1CwuiJH/DO7rZqqN2nPlBS9+makOVN8tPMAVAxa1coMOf4y3s2rAYM4x3/J
EE+LTlYD0WSXXN1zoudh3igSUaFZ6uWfEal3VVZnCn1CupfBTa0zSaLu37mKUK6Qtk0xa/Q2j+QJ
/oJPVXzNwTGJAzNGiUXfmkjA1dxpd3FChgrdLgV1CamcA94ZX6rHsHuEyRGF+XEVpI6NjfPrYesE
/+8ttGpaVGU6VpvmR1wy6J+NKZ/2MO4146HYl/s1P+VpH0qCPx97XM+Oarr3DpFYAKr2qyJWBz3L
XHne85VvD4DGhK9xr/0YtllJ4DHpL15GS5QzXhr30KVup8y63PDI06Jlxdehqx6dkoH3Z/OkHMfB
V6XpgEbVAWo0J3mVpbeRk57eFdWgkOXyROudmpo3w+MNF+UuwV90SYkWvUW6N/GkZV0+94V6o7bQ
/HeYVtVCDAbwpO4hX3ZmLcZRJVRSCFIgC9GsQRvqD5kmXeZpTASOuJGwS8Sj8TvmMHVa3PRCDpu/
eGxGZsV/qGK7kVtY2J+a8Q+I0yCMY5mQFPPlUAuZTClaxnF8T2oAAuvWVGs/RZ9taGqB9CkbuUGr
rEC4AaSOWfDm0B//yCOZ82eS7gDeZV4hByUCRDpfRiOjv2tBYkZ2uV1Zor817qrefT45PCbugYmY
usOlSHeIX+QQCaKY54lVMXa6a9143AJxITuXerrF2yZeehYJvrMJjHVvaCjQOeSHail+RjHImWS8
Aht14QvzTPBkAUzJQGP4yiK6tXFM0EGVb8RaXeWqlKmWglv18fVdR8gO/Eu9YhBvnoR70y8iDVPa
a7FJpL1hqbXNoOz+ORStEiaLCCqirL26OMVeRPNU82RELN/P7ca0U2BzP0wB7bgH5DNxhXxq+Hmh
JxNastK7UJgwylUSQt9yfkQmBbuqKusKcxmMcCIPUJwQHnZluB0tG01LsYJQSMf+ibA+/eVGrEEU
zoUNk3qJL+rRobsnJwRXfAuVg3X3YwpXVXbVx2hvF1PIB/9UqGrCYFfclJatIhj1cWr/jiimiNUw
5+h4hXqsjPArJa9xf+9+vppBbPAhVvai2f/HZe0yhI/fBM/gBwDHKnHX8DcEin+gYoC1EEx0Bfuk
/hgQW8zKM6YZeO/rcYMvheUqdnx87OsEoHONYnFbFE5QpuQ9buX9/ykQoUv965s6U0zvE3cDRT83
wFviB3ru3MutjfXhOuu4sZP0TEnLv2iTaCaVvzYVmx5hJxPdWG88b6DQuWAHnElOyKOBiYr33UVE
bypD6H4bW5EdxD/aOQWqtHVTbFzvSKwFboqfbPmIBjuSIVe8grVmATYImlqfTibWVO0JXlXdxiYD
9YdLLKnPtkvnKEXZY2tuBzUstSmtzsYtsDJtWPVAPciletZtwUvXY96/a5/GYvqdVLkeHSBDDhT5
Sf1y/CraYRgqoGAVh/SYI+q7/+cMl23SA9OnJyNxuy89UyMEt6a/1Nf/asVaYZAPoknAKE8qRlO+
CFluC2+ooaDz8CArEFJFcru2RoIkBDZ7bNmj89QSISoo4Lr1CCVnHVVWMgW45McN6c4tkbdijHxh
edrhEOj7VWCRjTMfINOuQH+35PNdYqe297xzQjR6J+SHdrbkMnZNr7meU0vSMY1NuSEhApTg+LQK
vb5BbTu/SO/jr/uFuJjWlZx8zi30+H0vzg8dcrjrSpBHtfCuCdrb2j191A48F1OgZ08az38CcPoM
X21QwaDvf5HzFPLYmhF2qLbAVH34YeIIS/sH9O7Ca2wCh2b3SzXl0DW1b3h0PvYJL0aQ66o0s/d0
1UOJyCk/C3+SPtg56fxIx1CS4/shynPI03K6MOiPYJkTmNVBEPXdL6xNd6RtJwH0jnzwRrQd3EGy
iNNVvk99/Rg8XPb6+z182f4w7E/x32ZdsEzUklme6yxL3yEMaG4+9ZyYKNxdhmp4fw03tbOXCOb1
vrMf6dV0U4Bp5dheYaRaT56JZDR7LDG5rtkd7El+niR79klPuImWBoxF2pdQ6gE2N+jAuT9eDIMk
TJHQ1odSa/UgBJHmasJTH6X/Mh7W7wj0g3jOrLVSD2Av/CbFeDeTcAPiVk7ETPhwlOD26EJqsezZ
uMlwj960Zup/mwschZBOJ5Hv99so4d3uQUWvHVpnr1pj1f6vzfdzS3jrLzh8dT3jle81Dk3jWGoy
guDXd1e4F+r7PwzB/HGZtC09z5hqY3GDbF1C5ZKCXDeeQLzZXbLQwk0p9REDqIT267v2lHNoEzSK
mHtbCoPPyWdNCj8MiuINfrtQYg/M7f1mhDZIlgYJiREfUbhls51BiwJMqSQKy5vkExYzP4l6V/7h
0+t+dU3adENjAJOXuGROhrRYNmuJYh2Js/kd8d6IFLiUqI6MxI3VReiquhqkg18TyVYUpnD1rBBF
F0XF0JXsyolREy+3weLqvCN8BrpZ3BhP3WSUrJ6+lb9NozB/mzmjpocp+yZk+gwP95zZ/yb7m7G2
GbfDQhuNKz8htwgpY5+fth1s7Um/ofqxjpUEo0U428IxfEkpKYDquf2uvtSG9nsXbh4vsL7B9JjP
nY7iCMCRTMT499A4sLNJaTmRnBTePxGFB54NA3WzGzxd12jmb62WqyzbsilVWysA6o5iVwQ0y1I7
5vzJ01Sgw6fQFvYA23JCJylmzbEYWLowV1yOfmzCB6bfwYfy5FgKxGYtjB/q0C9ixSDphphxZDaj
RDfrY+4xlY0cN8krvd/oRflYPNDfHkOsrUXm0ZCjwWcx/CPMdTUvfluVO7ACUNNoOj1AIcGDxBGJ
eiwxZxzwCouoTTlRa2b8hZa6qc2rZXKCJWxNJp1eO9KLVrRti3aQjORjJPVsVBLk61VEPO8lKvH7
der1AXlhlV9X2lEccTPNTQHFOUhvrTCQKtYmMI7X0ZEVD8caEKGYmW3tpggDihKMDWLnF600Xsom
b7TXY1zhzJIyRRmcHxKtuAUVt5Rky6QTX7IlRty3BGOcPKpp25Z8u16eP0wS5RKGBtoBbdK7tKxI
c1ni/VQCwSNVBDh6+apG4bKgE4AWlV/3az4LPihOtI6Tn/75Ocgot9xRP5C1kEcNh0MJ6jMPHSrx
ssWtrTxkI+52V8l7I3bCbQH3P+VKG95VIlflStufvAthSaGK6k+iaG2GndmG/iHX13le6t3tHLMa
AyRhve9iKHUC8C6iXIqMoA4j8UjH1AMuleFrEkjPQ9no8lznEFQQ7IsyGequFgDVllYwLkzvjS23
AVTWVjOHwSerwhv8BX3226xHAa7Q63YPHpN8ev+7qnBfVpB6NdfeX75PbrS60R6UHKH+vcXfb1Zz
8wjoMgxJzfVoJL/SqyEvbf0to3FT+mX4wjRo71THC96j5JK28/Jy5U0o9QUp7ikuTkuo9Hn5T07O
JPsvOb29IKMVD42Y7j5v6Lp8VNk2Y5Li1W+N8KDl5Q6h4oaE3PEMxAjrzKAF5r1rcj/5B/jxbbN5
CD45sh/whPwqUxod3VPX/B+g/AqXUcGTYN04HIvWilKYcnYJuwx9sI1d6PsFp+/OkPd3J7Wqp/rs
ZQaWwR0MSdnNQWmfHbeCzpTLBZVWGZV9g6HLm1ylWdFGnHtPPYlB2KRaocV9t7O4iD3KpojG+K6U
HVxx5TzAiymO1nYMCelWPVuqjpAzalMeIVhzRiowUucLHWL1mlaHimvHaNEFlibtbtuuIZGXVj13
mt5WLr67QLZMTI7oh81GIYU/WwjZ+S/XAuBdxy8+muiR96eJWQ16bbKto/jlG8RWDQZi0cyS8yEd
iDGbJjuQ0iusjbM5FHAQ9SEOTaxuePrQJ/AZ9Q/ewVT7piHylUEThN4gTN24LiqQeT1n7sKQJBsD
k/4tIjczM5TfQT/FktliGjOuSIZtsYst6tJf0m3RuSL6kyc+CDdqxIcs8tPaebJufNST1YKtq3dN
LRRZiUklKyNecUYkV6cfLkrkvWD6F19wrsqudA92OBDQ4vz41/S/YqYFhHBrKIJmJbR5dJifrCfQ
Om0LYRrgyFMaJaU88SZevdbyXHu3KfwnG0YjH64k2D3iTNix5nr6GdzhMopEEq4X7Yc2yef6rU2f
i4ojtKRHPmlh3r/yAaTAIPMAv9ME5XNcK80lR8aj2PARma7t/7ub3CtJhQW+hGBvKeIcyz4Kd/Gp
5lGofh6cX5+i5qhpKbOAcJQIRa2PISXoATEr3ekxVos1VlAuLmCrh0gOUvjIZQJgVr8fT8YH56oH
P8+AL21Tn2pMQnSkiC8XxkQYxAtWCkPkKfA9LmWirOJ2BFcNk8p+/h0z1XWMhlDtaG59kEDEvTXP
TGl9hiMSAQx3Gj4qFM22NHAL3+KDDwJAbvAGNPvWphjOKalUfYMhMYuFDBJ6Fwi2eEB+r5YGb8Ul
pUhWkytY70b/MxFLJo0YyOJiRe/iP2VTBS//sFWf7XXFjJ3DOtTTZue0AphFrkWXuWOhWAJtnsdE
q/l6S2xVuCdoB/NiGz+hG0+KpUj2cwuvgO2Uw+mh1i/QpmOj3NHAVw0coTIGI/EIpNOZy8EKs58E
zHimCMyqDBEelOHL7vsGev/cr7sZz9Ui0LytCRG7Hw1gYMJ6JH3N1Rk+cZzhXHLNhSg66ixb/0kM
26hpHgd6TmTR6imJn6UAvgnwhWZAfChn8/1FsLnGpmr+cJWdlHl8SIQnvZ90z0DzgIIbul5myICd
aKbg9Bg4luC0Mb3WWQUhoyLjYQSMObZHSMJP13wJcVhlx3DZ5KXkw9zeaEgCdawb34HFEJ2d5voy
m+9GTICqvnZRPAx+P5FAi4ETkiILJA3b+pLN4vPkliPYFpboJeVdrs5rYixx7tqNUpGnNI1Y5U4I
7JTPoyN/0EMO3rNKjBNp/CIx5AZBA7ddsWY0FIxxkWuvxol/JI7HDkwlZHdSaFfmxGlbpx6LI/8D
CkQ3ubN+b89escG1lSBoST6/5XFbA2S+5ZjKifBFn2fVeRb1zZtSTli5OjaRaY8QywKXvi9iWh9P
sY8Phke7JoXdkBnhSark5rBvW7XSrp9iKGA21banqwq899jSH4I3DLXflnbJZ2Ah67AqD68hLovJ
20b629dNZdYkZZRAKznRCelw7EvSwf+MlUAXORy4mdfIr2yI1dOZIu2OoIhGoau1kbR0x9sLpODJ
/vqrN78aSz3j7UcerTyGXocbQy+JX9iABeeV/t+THqnC35SGe36DT9RNwOkaI4OfS2KLLmoyv1aP
NovFQiWhbhLAUidRBi56HL/Bk7sP97bFwYMu9862R1lYYOAziTw6NFoICM6Cj7nwX6NsLJ1XasTB
KqeDF5dcLFdJu9RT6pkkCkDGGYx19SSu0N9Mpexkq4xtOnC47uJ2G57zKkgBx4O0n3Wk/z7PvwQQ
ZwT5PoZIsjIGQ5ESV085DtFzdXDCZGyAFmqKqOka/CPQy1YnfZqw0AGyRfP1wZryxuG9sTwJx/XB
A+xSTPvUfQUCDfzwMxW9DUCecpQJ9dajCSO3eHSdt1T2S3aWjTpfzDcvg6s7n2dzOG+mz3qUqcfC
2hi29zeZBY7jBeywzMziYHSZU7R2PL5WY1muRKa/BGVSBLLVTxTAv4+i1x/quTUZUJQ0DgJDPF2F
rsX9xR3PxMzyqOpvNS4x0cvQrKYHV55B/dudhCvc/WF88Ne8Z1fWkkYApNiisul61pt6knrvtXS+
EhMAtDfoa8g1cSIhigzudhUAyotWR6KNW3wYM9uuc5zw/Dqg3SdUnzPFdTApnkaZmaOgzrQNUUdT
4gtpmzPobV2OGm04UWXEpa4izp7WrkHdgPkIAZm4XGPouN/jTFP5tqI4wnIAW8HVx1NCMSK4g8gY
1+iVbmZqO6q+0o9Eo6tcO50LI4JyPXKj62DEoTIluXx/YsQcxIQoPIJhYsxcpIDRfd0qkQU83EOh
CVbrrLh8/eCtltCy2Ce/mhaM5zAr6w5d91EKyiZmu2IxW+P+lhK4GbuQZD3yBD6rhoXrlP71jVUn
lztvasmqTbI/jKZm1zigz8Iuy5TBCBbC2g9lcqc6xgNAwNRoD7ZblY2/Kw9KULwAbSmp7aA/Ys5k
RYwn+q7fCM+UHw+ARU++3SiGYC9cSpSLc7xWD9s7zMtzByWVVlezfaIlUJi+vogmpU0OKPT7CXtk
sIvkbpGD6vLQjb93bXo162bOWwty3MsJat7g0fvcMvpqQWiOhkXRCIdyZMsCcrKzGcfSasXCwORA
VszQfPFSJ2Sy71Ggk9vmf1OtsbK+zrCIShkIruSayyzSwTQl76Rdk9ppsMMD8F4w8oQfSeLhLFwx
bRSaXgRvGcSsa58d0yLu3RIn8yU8w6XDkA3PQWPT5WWPydQ2Q8nIVT/bcPBR40rT5K0VRw9voMQ8
aT0JldMkOTGx4k+o8CcVCxsgUuvKb7DFcEeG9fpfFffO+MZNPRgEXK68V0DLE7u+fNALjOSAMBxv
35ZOzl+MWvoYX5sPRQ5NraOxN22TeyTULXNk8WZmFfXo0t9pZF6Qi9zudPlldowxlZ5YIkwUkw/l
U0iLI/6Jr2MaS1G4R5YqFsGyn+q3N4TzwQZMyDO+jPbdQPTKgiHr13iH4a/cMQkxZHyEWlpvl1NU
7heleABTDsc1VkOOoJXIIhj8D3WAUNHpfnOuCV9xefnQAV9MRTrcqtjwrqeGVyLC7lCA7d1bgNCE
OdYyesa+ptMnPHu8HAKqVN64Gofr3l+SZrKUYsBAv3ra6DaNABfjaiYO4FhuA5SlHv7qQLqzHwFq
7vASieiIXyyNwr0BafDWPsSADLYVNdgnl1jW+kCoQtUe/grgMiCf9VBjKoDt/U1XNzGyhT4Y0xAu
xeQeXxx8Iy+BrrxAxUZhqca2ZW202syOnSaNMlRMBcSNV1xGnmBcqY1mV86V21FD0ubDeKuOCLVn
bt6J2Pw8ntCMmC2Q+J/oydLUWDZRMXkmJ5pKYYYpYg/WAVHaohNgot97BeDCIAbzqcnT26QHaGTd
s8FWTiwy9jXQQ2euOscr4sulaYv8SPZ+/PSQWX3hpzJZD2pbyl8usbaRwpK7RQQ1FPAlGRbUQRn7
j+DgMDUapdAOAMX39+WLeGNtoyDyu2X9MHNztITJ75NErf+fTvOPCSV273HNZxmGB5xGznFiWJAB
iHQ79OGI13rdXEYi9ed8fJh4AmIabTrLBZfuPtcooQIAAgwYYSot51Q7JTkpY0v4RXn+reUDWPzT
+7Oo/J/hcKrWDHcKBBTNld6dCrg5EdmuK7XLgUQA+a5e/rwk42+wZ4Qam4sVYupSbNUbrYrONjEN
qMkOJ0yYHkbwkyYVrwyU83+KOBsCNsXLW6oKZ+3VFeTJ4Znq4lwkcrlWmqBI3kegyRDDBIGESUHA
tgimz862sM1iw0xEliu+h/z8yimBIbNWge9Ib8SOwV61Fk49xhUdKA97zy20DecClLVooIueEDn3
rqLGZ/jBHQIAscyhkMA8BUbCAwRX/WJ1uFzwBG0TCYo0GJA8BdGUuv5MtNtWLW3ALFE4KljO+s2/
f+WP6zP+jIDU9wrL+Cla3Ji43cYDevnDxydCWhZA4aMyciTZXlI4S8O0nVvEAx8EWxYss8B/CRHJ
Q+pVj4mu65VttV/ZrvqrfoyhDN/fqSv5nwcLL9BHt43qo6FdXOLHNjO1lMN6DlwCLZdDeuU9mlw3
aT2tsJT/MEjk2lG7nfEu//2VAXZvnyWRtBKQKQ/5XEzQJAHkOSHIcKbcwzYTPqbtuQNheq8x0mVa
An6zz1qvTeg8wBdfS3RgumFndNX/Nm6GH3Q2rIoD+IBwPLblIu3McP98DWkX1GeOQHDumbUkerhG
ZF28u6AuLd+Kfbbezapf/ZgcEpyBxVYXi/7zLNzRXviJ9RGSLZjViRJOcDrscU+Zetpt6siivIEX
zj1ASzVuqC+msoxa0bpxJ2MPfTTX5bpp77J2h2P7jySZ++mkRNLRCMKHzNhACP5k/m6IxSMcWqJ6
8gZ9LMkKjrBEqW81XEjQDa7KVNMAbuxti/1NvaNGyhnpOi7GasUWxjrUav1BbQQ1t/WGTF2Kd0SX
+bofZ6M6Tck1VvxcoWO4hAUslo0pbOGqs4rW1qXupZwx3Pa5mX6tdlJAkp0AkjDRC/X7/G76I3eK
4dVyt/vQucCBmUZnL7+XX1oD2GtXMjWt9cdbzd2hTtsKZ8aqy1LSMcDyQAWzyLBoYoPVrdSfDQjt
cFFYg85VLKf/j5vK59V4Yd0reJofFf5rr2mxVwxFAIAsccjSV1eyPBrhBKR/ulI7KOW1lYfkKzPw
VDEwl+wMiLvsqrY60hccgOTo1Ed8gjWli5kBBZ0I0Fw4hiTJjspBN7WPto5yRfb9pklmscIIb3Lk
667FDBoQaKtQhgXU+efokkT+pqQQNOqSuTDvoN/O56CBQ+AVZcsuWx9Xz4okc8BzeQfePqU0WFv4
1Io2Q2Bhuq3h6wFLhGh136RYy+Y4+PQSXQZmLwV4NfmXme8FQWoGvBpwRLNLXzi2SYED8FTnVASt
9XpFb0TdOZWtz99dh91Db/8BAcE0exiHnyHxg0kF345a9j3bZ+l8ZbwcEXOYnA8W17+VFK/gGMDp
8gL24hM96bGuH2xYQCyXqD7fbUPQmZhUeFC1pp/NAXEclFwpOObt9g/HUXp1+IPESyfKI5qIhBdE
4qStrVm+pY2IOFRLUe1CWvcR9Nd8HD5WGA/9jAfQxPWzBirxmSHreZ1gguV/Gviqs1adIBxxeN3S
/fOACLtjw0WfP/OJosNOef1rQXXPnVcHcwVCeeWVKspZaWrhPMU5BfuVJ1/UlW+s7XGqqJTR2Gc2
WGYnem6IKz2HfzI23OGRt/I5JGlW/yeyOg8xR9ccEHTdDYhqBxoPQsvMszIyw/P/m6NLq+EpkXBz
ZnUBd3l63gVP3gabXloVE9teG+aiZUsB/H+vqp2ZcexIMlCvD177uteGQKwF5uAcvlOSPhOOT4Tp
MSB3EX+obNLPVMtXx3m1G/Sw/HQr6y6vAcUyTDtyx0qpokaRnRJMtLQ+kOIL+7jbu8Q1KkaTTrUe
6C5D4hXhJkFdhSpewoJx/thvs8O1Ay/5kuSROdZl1+UQ52hx6zcyqi+sqvMQPOVYz6DCOzaxvRGy
3VWvrDOeG+s+E8Ly/CVV+12tIhpoku7dclVa8FXXugq8WeqlyfBAbFreJBfyCUZ1Y2IwA0wamR+S
Nxh0GdxDx/T8YVcpW9Pe6UNYY6I+th2x7oEtirLTlJiLoq4nn2fdR4f0fTLK6z09D75nfCBrSKf2
kptoSHOt7HqwU8fKOxLmWiwNcYNMHbli+lEMWmiW3rwDAYuzlXRNJo2kuDhuBydoYGwLx/w+tvGf
r9XXcogpULvucAkz80Fu92HHAYu95f9RtKAeR6b/lFgBQknN3KZh+QEI1n6+4lu6hZzpPTgXZcSD
6fEXea6VkneXGsmpYVrSjhy2D8HXzuwq0RurJ0gveL+VHdLWeoHks5JPYoqPlI13RdOQbXM3bj0u
B58RJ7BNnH16/ILUE9Z1OFNh+bK1BKDQf0f8G+ItivSPTs86MHsZtiu0B6w9oJ+FC0ta6Ha+E9Ga
5m1enw2bweRlqnrrNTD+Uhw8cTSb9RtelYYOZMi/3clluw4RmE7XAsY3GGSoMndXxVEX70fFtfoF
eXi8/V5AHTQ0MX5lWLwgnjKaPHY6Z96HUoYA/9OLCfbZjsH9ADRE/CXsWJYrPToFCO+OJSyuF3/2
5Dj/k551Nnn3RUJ/zUOW7UrOwsnP1cZ7PERCCWgbGPL3aCC+Y2pnYhkka7f9cCF/IV98t5Nz/eU3
ChRa6Q8V65JaEOfux/jZov6g6C36jYbCpleUDPHm1aV+YtiP8PEoZLtgzz+o4/k6RcAg3d3CHezG
oB//Q6Ov3is8k2szfhsr55bZuzBgS0boQMKZofYVKxzldVPIrdO18kNj42oiGGQFv/a6wZIc+phW
fH8uZfLbs21P7L/OYRiyI7Vtj94k+NfW3k0CfFv32u6qoxyYs7zqVjHPWz18nXEEa1XtIg5WcQd5
uO5BFcrH3MwhBQdvL8As5DRBcj23yjxeDdx4gkpku98rLNC8/WJ8KQUqYFrhdEyTDKV+3pYmtHY0
QKfLYLZ1J/7AArDq4s0jQtb9DIQLG5xVIqqptuFmOpFD8DIUwjRM4WmWf6nk0Xbx2ypXW7U/c5bL
ueD5wD4pl7uz4OpRRTeblZfuBy49NT5xnFICAoCI1F1BEWpdqGFaPluCKSgr3bSKV6QaObEPCAgF
Ibx5aGxW5xyx+d2lrZGiVjYrtM1KViHYKkTPjZytHUej9zU6edLEUiMBqkynIqPAi0+mRvlAcIkh
v7bGUubaHqLiEK0XwPLQYsgRVIGSrrNbo4RppiS8SzHBUYU3leeLBuXieCcN2uMPRRmmEY3baoLe
rCnXTICNtu3f1JMzkgqc82JHpU6h/qL5NnzuX1kSyV6sQZlcf6ecQ+iG4l6eQ7/Po8T/tPXGVsbF
1DIO+42KABgYPzYoPkp35VVwgkuEnx74O+pvj1zuwRUIUvQGMw32294McTxZHyn8l+P6kNBPaARs
cyseMftaIuB/x4DnUSjnYtPue6WYH1faagdlqd+M1PCL7QviXW+bSrpVtG8gdpeOj23/iBkyqVgt
PWX9+yCF07z5OaHO55FzIkPSEkMZyeB0i+SclOhsDJbhcXo/QB7DKZ1aieHRKS+8oFTj6csjv6cl
6Datc6+yv8khAgkPPtQA3JH0C3+1XvjwSucha1PkNpBqeFmtcG0bWYEq/wUzVVJlKDhTAnWje8iT
J3WNCHH2cwD8RARC64Vbs5yIBrpYKBxpxdP+04YRYS9M4HEiodhNshFR6mOpOEUtnMxFuOkfA9s7
fO2fhHryH8tpLY8DOXEwp6LVumT6esO94yCvMvmCC77e9IuDYyyF/1Xzz6o127KNIcvlZiPJQ5KC
asVVgHBTyWIz8y9Mfich5a7JTx5JBtcbXfuIxBofpU+tITOXDEi13uPht71bi8SKBAGNgtqy6Ukg
WFz2xCXQc+FWEyLDBfKFuLRyFErlzSF5FSnPvGnpEeAh+AGT9CHRZAlrJ+29fFqS2zgzjqfDJcS2
l5zgcdqicQKuSa96eo8DfE4mupubFT2N8jh8oRehlTNBjadBZqqxVJuTWGAcZ6f4Jw3V6mRIQU6F
au9zm9pQJGZH+oLFnqmxidYygfZOPXW5/TEKsMemZfjwwc0LzN7GZiEawYUrs1vASWASyPrMhN5n
kgYqCEx166luZlRvVkI5IvS90uJBHJuLohlGWCIhKEvzu50w5LOWAATKc5/R7sbtkuOk6PhSVinU
qhzhUIVDwe446rm/K+VwMLm0YkiY9omXtfgUjuRYupJ7XKFQdvhTueJCjDBy+dmzePyysqTx+d30
QJ0Ob+/lav2kcwjPewjiVkOz2SrR6u7PVZao5qT5WzjYKoBZLSw73DKVggIZ6/dn5gR+IuNztn17
fjapCMi+cKPBfVlNmMSEQmmYxsEvd74ddgnfC8d/Roymszo0mPFKUE5gDqNn4CLvuuK78hVypUxk
E1TcKgBH4Il/+bAHQcmcvGLDgS1NXkXZSlxvW8QsGRkEsUHEcLybtdsOWO5XoUf3iUknCcngssA4
/sEH5lngMWkNXzYm75o3FTKBiNfwonKy8mFu1w62HcjktobRL9G8qt7CFJ2MZM+JK0Byqdu6H7tA
lfn1qLfe1OHcemMpwmK4bF3ajfAC54wJsFZNPHGzknA0IrsflqrA3+aCtZEcIouu/+ZZ/soC4zHQ
ysrCEK1ZUFh0DdWED/cQxaEqcmJwmffS9j8ka1t4vTrq5dDhfeNJBADps/+/xbEn1Ll0WcTnb57T
RhNxgu4+2CZ6s8eQa6pNunX0c4NBwsDAhw8vTHyYzbGbQl5Ka3NcK9P8yXmI1IOkRdvIAa8TWKbB
ocE8OOyl9fTK/q/SLRttauWHgONqwLkZsfGTDmuEzg0fMpD8EgHhDWSSo9eIF5LXDZ2DLUo33R4D
rhpkT6CftIwH0FwQjyyZjBxX3F6vd8ntMXFMXud1hkmH8oKbdizfPasPHfV5/fKGmDz8xF5e1Gai
qZ5GDsz/+67VeJFo4G0frtpUVUw/z746afMN6kqQn5JTaNgVBj+O6PmbfZO1wFWOhAMeO4vS8YkN
p38S0wC/5ml0/JuQMRmb3GXiWBdlqurTKf7MN5Iph1aqocyqBEHRgNv1UvKefiCbCBU79OxZ4+eI
BFT6SasqsNzVwMjfg01Bg3P9OR26OObDyEU9h8ZzjhmCE9p7DTcSXbHpDb7m6GEQJR/eCc1fJJAz
744XBHzAZTsGT0DCeHtYv6pVAXvhSJn0K0cVud089bMyHJFPKZ5li9TIVMrNIdOzO+8JBjJI/xxM
/bT41wkyj1TiyayVMbZ1Zh1ycZyAPcEeG1ld6SZGfmS/iBtrJUYXg0mnJp58xpkPPhLf4JewBCwf
OW1DQPruA5rYxGwCEVodJr4dcm+9Abedfb5Le2pDxTR8xH31kSIjQRF7qULx8jSHL6ShTG3Iyp6v
3Yb/14eJBKuhtYo6pgs2IlPqHdjqY8zpF3x/s9iG+XoTKYWT7xF1ejGY0dI0RoIrbzVmZY1/0u9L
MohHeTsufVRmlLW+F6xdMzZPoE78WW31S45PkMUaGwftnkVrxgOw/FrhS9dGLVM5H4am87nUzM9x
Mmdqs6eJt9SNwOes9xDkL9hqFWSvugHXYU/fefXkvWpYMcpU33i9rAg/vHAz/jom4w6u2UVLzMk+
4vru8EC3EAAsUbYtC327nh/YU2ECTapyn43NXfZ8R2L6UDGYRqX5kLl4Evh0tPx1j6P+49WQY8As
U9k0wOLsL7wxDeU/Qklr4p7gyyd5BAAcbX1xdqD76KY+V/Is0VQIvZkLn8x8kf/d4TfTrtScGXOx
cX+O6nZUArwz0bR/qn2pdgA/3Ac7Ej4Sd71eRdwS5Sd0jdGFttYzYe47NvqVOLOi4VdA8CqY8YCx
YwO/O8CeR+yD3qTSkONvkSmA9kP38ymzSUM3CgccDnMRrsDHqZnonwxvKNF951v7Dbfi4uTFVRUW
hnulmVZ6+26A7M7a/XZa/ZgXRHFhZQtJuGKZIKeKz1H0dmeTdBYyWkybLRKcT55C6gyiwuxDvx1j
8jcKgehiTE7MMvA1ILk8BXFubkqdjA6EH8xdDaoCf6Xd5IBni/Ao/fZbkdzXaaNBOfEF78Nb40vo
zDDZ4f7+KE2FAt/LE0jkV+eU7L/MBvjAW60l3C352tH0rRbqj/L0slJJOWExgLQbUH1d4M6UMW/r
dih2eI+fbtPVZ5XnMB2ARUo0BrsLZhhR4jMtd8pqIA+n7mOAvxtHwI5I0eDaV4Qx7aesJ4hqz3IG
jC3Gu7V2mwiksW94FpS8PFfokyFG0TwKZey77ffZsJBfhfG0gakc/H3iDjMHam3DTSaQUwh5KqyO
EwnpBxvp1NmsFP+8ijm3nAbX4M8OEA9xklqzOrhYFQXALHg34Mh3pHTCopLrd7m1aR9NJ6TCp6ZJ
URyjO5N2e8b908TaVAC+Tvqs05yLTGobFg+s4XkoxiTLTbqyX1s8ccpbQlbZk7ZyTkavJSooe4Os
0IHbyD+glF5cAE5PYfu0YlF4NBjn3e5506hbFcHluqSIoEHHLpmBEUry+grFgujK30Q7vSxqWWPi
9gLa8v15cDo5es5ZCkAXjfGAaumAqIJVoB/4bvVoSr/K8/wXbd9bmUpreH0S3ZO2s7u0xyorqXme
CRjYuAdn51t4O1REdDN7dP/f5XjIBZg+sQaIzFrksQY9rFa1grPK6R3jxQ7gjN5Lb8icyUK6bU79
Un5XYVZnlYmkVRbmi6UnBkSKfoM72ROaEdTE5wECnt0gq9eRR7eFncqc3nnTFwIeb+cqLbRq/cda
si+d1TZPQ4gyBf7qbRa7jbQke9B8ynFmaWzUmBHMN6pkGwgg4eWPhI77v8jrlwGXKhoDzUsPb9NY
QbP+lj/ZNmsgYZhptpUCnD27edeCRBtWrIfopY5DCFllkMe+HXNLvsURKbCkfHbNO3j84INH+ZvT
5/pwv0XMtKq1oYRN9vJVsaoKxp1Cqe+9CKbYBADR5ImFTfG8sWudgPpiZuZ4s9cmbARjkMUYDZco
eGNSzKt9es4JGcoicVCZHHOq958elCRZC2xm34Q93kdprjmIQM1AlAXllze47kZGUiN9maZXc7sW
HT59IzdCxY+Zp8joDv+ubPpcpHJtrdpJ9uIydvju8v5wNk/BV68i+jXGMyXXFyGs/UorTT0bvmsV
7Rv4wlwrj01WwCd7e+puweD0UvYgUVMurl/Xb3H0sopw8QtfOHe6Au0fPeYP3Z/3JcOXreVIon/M
uA8UFtsJdQZU3h9ZAZVK0I37pE5VyR48hnBq3bu93ZXZv4GfDqQkvoHNvqSGxZGlHZP1FoK14dBY
sOKLrjWL45LnQIPP2sSNMWn6wG2XNSrleldgTDdr+q4i47eHo4DgOoupz59ert7tjdgGWYe3RsAj
JJiFYAXtLmZLytDO0cu5xfiYK5Nxr/1Nl48gHepE8uDLCoTcd5tx8O7qgSuMrlxTZ7yLQsPKu8Ki
npCg0XrUo9aqV++aMJdIXB1XjLJEFJ5hG/4rnlQkjrukJXmTq01h2TQlWBZ9iolDCWy9CzdtPOEy
waQ33QG8RZeBsbQuMQKnGhPMCpdvnc0AztEvZ1waKfZf3b/TuKV5nkK40OWoTdqIMYAG6gI8T0oe
W+0Qjmks+Gx2D5PPNPvph/ZgzXxw8z/FRzHx2QUFgTMQ5bP0R58XVrs9f+9rabITcJ+is6WYG3cu
N8wkrQuRB9J3Ibx+z8HplcgA9s8JnJMq5t2WhECg41i0bz8H8d5Jjbf8VwLgNLqted9B5l6iZKnD
i4+z/ph3haVVh2gDhPs0SppksIKc/ntuS4uWvSjoM5ZcsLSPRT42zVm2VCQZCG0LyP9yBbjOfady
Tiwt/yD+7ZNw2f/UFb8YYz02xnGu37CBjf1DJSooFhbPfaSiAxwEl01ZkjHYQhAZHQVmdW0A0hPH
JB8Qfy6ztXuMzt1Fk7qNqPfxVv2TwcLxDdx/ovwGRzp/h6LhstswQaitKF08GWZnzY9NQCtmxelX
T0AX9yRY6TIIX6z+ls7OwQPuwm4fw4ZsL9ZLfdA4eeBDC5lnNPxJ4LfnzmS6R0SAe4JlOducFh4M
wsqMha56X0cmrNdUko03N5f0dbEpHYN5DtURN9pIUjDnG153+hwItcH7uGvDaQVKtzc4gMB8uod+
iGCC4WfkEjD1C1z1qYtYiA4lZVpz2SNZ4ZWDRHXcLGWiMw/mnghDQkCczntafnWIQ5QaVqQMp8Kq
VC5dlkptYv8Rxqyc0iJTSa42TZfnPZEQjfHItIXMPKNj+RCvV+HD9RPJZWaDFN6OajBsbDrWhdqX
uTm3FgnP64QaK75fskXYaHQU7hl3EkwuYH3QmFinBSLuZeGG/B8ufOYtyh0vk8TjeQST0P2q5wbu
Nzu2UqMPu1omv2ZeGz5KJHmis0GmVcSVrkpjJv4fuidsgLEVSaDPibozK7VVMXe09kPjCbVxgg3/
6y7AtU8lfcQpwJXF2hFFuIOT3myKuGcTfLxrNL011gdaRhs2uAZB/ONWhbxwxOESWly4uQL8D742
lidJetegKwCkISSHk26bW0C2NlXzCMh1MmB1saPBp9MiWCcY+waHDMA2/FjgdMDfSKyK3IfBSzGS
c4uX8c490pHJpyz3UFTpdiOq5YZvAO0EE9GWGC0GBrNMw7HjqNRK4LHQXVeDZ6zMHHk6f6Eg65OG
7nUH56Gtww8U5XPKN7kQVh6wzIl43zMdpr4OdoVreOX6+EwWy9YVDsfmgyuCsXd7PNaJRRR5wtle
4BLk0Il9V/qPbU0Kvyf4jHQ0upl/hZHg1+HVXmY9Af0OqZcm8t8C4dK8pcAovscvWaUWz4QBgBMQ
rioH+pq5x5Wuf9H/S3lokExL/4aazvot3RnwXhNxhl9coplm2rLRhS2CPFwsrtAG6G1d4STrjfn+
9e1BouGIrQJknur/LV3rJ8kdHSza69vNwgj1EKq8t8oGzS42CyP5Nmoxg0GYa/hLztRLhe7xR4cs
rObTCe0DIkrdmmdHtO16vZWZDPD70b2l/H6y4has1XXwvK5oyTNs75iwaWubOiZVMTIS/fj/MqNF
X6YS26zka/myKy0V4zF8NehcE8jwZEEy+ZgdgDSx/6vyNHDwFg/4FbWSPdkkUU86dRCNwMlpRRvu
Gm9UmDdMBNr6XnDryUrY/aZiHIwdl2F6OIXd0VHknhLCZ7CkG1CN51H9dljcSNBgcfPZxSeCRGEH
ieYV1hjdlTKi20JCZXW1hLH/tuUysauszZ5w/Q46hm0mPnfNQr/bUeHY4YSTZhrjuBHyE0VqWnhm
sE3LG43JTyLJJJwCdq6RBefcBDgaaktsVy+s3jN6H7U8fhpvq8UBDzDiXAfq5KuLU2tNEy8RXG0D
91l1ZtAMv5G88L2JYg4eBB9U/gPW5sF56wbZj3s7sW2WEq0JkUs4llS/CXS2amWuwOZcO/2Dp7kA
zcTuySSzn3uNFIFbEQc6moxoowOd8haFSUEpEh5OWr0MIlzVlxdz7l20HaV0CF+L494+YxtjkR8L
uyR/SSAJNZekJLD71B/yk5Sktwnq4RAn0ZLUseoc5SfBl2H4/5jy3a1b9BJelDaAgI9fJoI/8JVU
QylNxflG1f0s8TF4Foxmf0FuZ5lyICcH1dbjnUV87g2C8Zpj+16Ka5JgYzc10QFyklvlRPrxxypF
miChIqKRcLLKaJ5KGjEXFSFNtC0J+GelZe8H64L8Iu5KDvq/0MBW94eks0F3GT/Xq8veqJDcqxeu
DVpNepSoW8KpeAVpEc31eHcvgEsHmK4YBoB7R9rB/XhPTqUrFtZJTCvDlp7uBIM1SWlwOpRjpwnJ
9Tkq3iNMygV1bQoCbKs5EhsjKOXtcKC6BkU0Q6oGqQAK91wNOJLwicqSxHvgwQTQkbsHLjyoK/7b
9XX1yqB4ueYoeqbtirMUtTMQXyOU3XLCPRAOT9cfKif54/8kOgqfW5ehBJtaz8LikTVgC42qPazk
SaBBReKL2df5hTPKppyzLjMnrrTx2OP2pD2gIkd5+ucxerYyZMNvVc0ahIlQw8+IpNzl/KHYJOuK
qgtEV032Zjy8/a0+iTIyIcv4i2RGTWP0NlPB6E2HdFxCxw4Aw4BUYMVD9hROtu8RWwGapl3BAral
6frlJN8Qp/WLYJABzNsWnI/8DQjWWaxpAVmtzntpfYLqW9VhFjc+62GlS5D/nd13aDrmzzCAIl/x
PimsgTrIB4aLts5tuq/wAGN95gsJem7/tDj36ff17rNLVefVd1VTv3hQ8znM4uc/1v34EXlzvxtn
HhRZrH+9+38k8uzVVEz2JTo6xCMOMKsI/rIp3tKprBBn/vy++AUhGjlOHvpdB7HMQbWcESWw+h3D
+1gfAhV/4DQfSyD60jUumhxteQfKXrMlYGgGH63g6EusTfLS80vWABpErXY0wEXfVzvr71/EfqE5
HiiQVglhv9xgvhNxCuVsZFmAVIQ4ByytIQKPNNNpNOM4GgGCJJ3XoDgBQQbLscE1csrkIipAN3LT
EVWxbhweZNDmrJLRpSQzg/mJwJiay+NmWCzK0qLTSrXnKEu6bVU1oof509ygG+CEz9NK654wtSM5
chWUwelxaSokyAcoZrO+HL7l06KGFYhlb5vxOPudm60e4tTL746n1nlFjGcdn356MDQ+sEQhTYdj
Qz9mKonURNM1iAdG9gcElZxyj6Nvkpnw6BOsKOF+5zrwSXnqBUbjgEFq8qmkRCzji8rgXqWSdtJa
oiDRpJjeFI+ntl2vcWEZ3TmFIlLMIDmH7Tj0Gw5pIA5Cwt3T2H/em/wOO4v4ChPvUF06WLVZr4cy
Jtk2kMh/9j4FSF+P6AZOTRLhOumiZxcFRb9NNAOlTYLethtHtoZNiFssDxDHxkTO45Dzw63PM8NT
ZCuSRZSM4GGR6TW6cZGquTeVQnNoY1h4rCL5eKpuUI1gTyW1Iz1glALi7LjzW3GmEKvI5LZYf2Mv
vvWPVHL6FJ6WzjIbdTHRGm9UujgTFCBRj3QYnTWDDpsSDPMGWaDVgUKQqAUfddPYWbY5H4VYFn0r
rDGD2K6C3561IwmMYqb1bJPBzSbXJdpIctoiItSKWVJNloSPN+IDnVRWEfwUgZQr3FrMJQqp9dUL
Hpun3JEubSKhCy3eUyWaj4dWig441eHRLXFcJeaPF+VS8SIfZ66KMNOdJhg7Fxx5pypkbOvc7Mco
9p+cUswIp6QTOGSzkXPq2yK4O+rCdd4nnAF8HmzDNLDnKT2BH4NiuY7gfFZLAFkCizNmYFeScSfP
1qC4wQfXNIaTbBdpFty6asNW5Xsn9EIwa0+Hhi2JMyAivq0Z5ozpG620HqD8rHuEqqRSjqn2NGg3
XbtTk+CGvvWnHBhfYs9mlHLIQg4DiZkFfZJAbbwHihwkjQzMBxgwbhy6CvVcki9dTcz1PbcQXwVv
YGTq1EWxujMKrKSzZoV54UW7TyzVDIagYBBOZx+9MPgEOA9KcumHpnH9LPLvUxnfNFE7y0BXs45V
4Ro0sVN3tzrPT6br1Xtk+1m1StR1Vh6zLsA0HjE1A23JFX6qxETKe7BMvazwP63eGTEhpsu0P5Wt
e9w5ObGBNjcKPpIQUdpA/tVP5h/GkVc2KIB0y/rHUX6gFRMOWWM4Xnb/vuObqftJBf9Z6tUSgS+A
NT0F75JDYbupYAgVj9gGuOmnk0uhJoBwUh2p/vklIGa3RQBVjEDWPGhhnzkMDxKL+5jy2Cg4NVTK
6eIiI4vA2X2AZNXzoF2v/GojnGSNVvR9Td030tWDrPdZTNnlUN8JZnSPwtkvfxztAe0Y3JbFMxrB
B/XZHw6HWi2CqFMTIKV9AaKmqZIpZg7ufpUr/C2wITW6ZlSytCGV+9maL6OHboVOJvzW3y6C6M/o
F+Hc+6gTr1+6tg5BMytvzDeC8DqFtUBxCfDPitzLPls9m1rCpIO4avR0F+hDH5FA29QPfZCa04vy
3cppWk1hWE6n/tKa4lFc4SbVqlswpG2Oe4VoojJRvbBlHdlqgaUCLP6WdA/u/gCLQyttxwMae66t
TdjZLkMZcW3Tt+UKIg9qu7Dcge/xgYO91ahnMzouHeZWqUXeYqlxK0WsWTtlBj8GT9SaXRvpTBCi
E8rNCM7CmNzrqPwHMehZ3+e3a4jqgJsLM/7WuD8dRjoHB6V1O7euHgmRgh+xGDHlmUPR06IqUo0a
SEzsVsgBdksftKMiM/6zf3gW0fLg2OAxqx/0QkEZCO5Wv72szNKau1MrfwwpDgqOzNx/F8pssq6a
88GzVQIM3jhcVplwRIqaSSFPYtzhkva6apBIGn0/dTyi9i9JynKT8edxgxVUMdX5r72Y9ULRSurn
o1xCfJvZe3T9UNMe0Z7x0FlGec++IJn1DCEJ9c79j8FVeg0GGolitHWDYu55iBRikfDqMozNUdlW
0zd3LwH9NHZXkq0fXoMw/0y4BOCyr02AtHmjNAIW/HpYRhoU1P5KM6m0RqiLZV5W8yB1SgRCrbn5
0twQ+qOKApssPS6p3tQ8ZtbW7QL427AuOo7Xk1nhoMtXuVorRSpu4zs+aWp/b1/wu+g0cGss2jYY
n8Bjlzq3CgGtRjqnjFYbApn6aQddeIeXadImFMmVwWq5vn2+bJg0r37Uc7do4VpNdEl/X9rnLTX5
XtfqkSKbMNFC3cVLRffVrvLCwZyED2nVXoxM6Pfc3+AOr+5JTCMo27VAQ7tIqMnFE3uIANkF0oqO
EgCjpdeTrMdcCJY94gbmf29coyHwnp6Z/QDPpHp4Z66sVVQg6FeqhB2Dx12oCS9pGERd6x4nINfd
zOqobdYk0P2oB7FKHjM+xyDJXE82u3CXjf4V1ge5S6u7xIBfMi3SBWedWviY0hOs2XC4kxt8fUsT
RNxmkFTrw/75cRF0z44wrTNSmVRzo00CeKg3ffxC+pl3hU1iRitm9jR9Qo2z7ZlmLuM5GuVtwHWd
jnu5iDBFXieoUi0kwa9vpV7V3eZAtXlD6tenD2D1yrkVV3fyMW2w8GE5FapY/G81npEpxEvweWtb
YbYU8ltD0TYwKXzsO64CFv2hmNb9279FweAW2iY05r6Z9mGLCm/bbb8qx8omiElBxQiMBl9YVPS+
GzWurHpraaIAjoXxbCMWm8jy2Os3i45If5VgKE/bMSDJrjMRFVIn5v6J7KTXz2ki8fCqnnDUi5dv
H8Jm8E+6f0nzk5kbDbgmSj4r3pFb7Cbxm0mh5c7gUx/laaQdiIoFO2rG8YgqpYRH8mg+TcYFtk3U
1TGGTzybSGzEeXZU7i4/TlJHqwIERZpz1L6czUY8ZYa0huGQJUmSGGlPjCtbfMuMVqbWY0hdB9b/
0AJTR6Ms7LXEsupTWVMRwMwtyn+xHVgRTo3GTYBTF8/ZocPLxu8OHVuoSM+ZCB6ReS9FLfOhntof
hlh/9wVBhK3naO84g5eY6X02XkuGJnu43nOe2SD8zHqTSGm6NsWa/5/FW74ak6SYM3actZhnusCk
+LA6kZfiK+Hdnh4m/WvX5xjgUJKGLjo+nB26MaA4ORr7a3/tRLQd+mJKPClOoHxHpeVgnWO3Je+c
tvI3RgTsLNQ/pH7k8ffx1oNAlwFU/rVmpWX3YDR0jkH7YBP6VRvAWRpEeY8mSpvR6b6HYP7bpLNm
4PB8reooCtvqf8GzUmYaGCKjwlPwhDsugyu/A7zKiYHS1dkeJpZzCsaRyEjvI2xDy4j3mr1HzLcO
eOOonqm3OcXD/Y9goRWCMb3XMytT+edaoNc62b4osHrtwYh9v4tC0ik1jVahZvu5rHhMMK5snG9a
mL6MhFeRV9cbTWElhVIugS4Q39PP/SG926lA/v55cYwCGS23u5ORDnHp/ldOPOC24k8QOi85a//U
6gGMvN48j2r7uSO45nt0V/nf322EaYMoPXMaJ6MlQh/0NwC4iqZDPOeTuJf8CXz5QUUhR7lnaquI
zQwz7PMs0l/khrb459b4scjObw9yI0ehJvEWzBWDwjXZZuQ8nlMSWjvnb/aPlqnWuhhsVJk1v2Ti
PqkG41tddUvhexF3ThowWfLIRO54dah8Y7aQt9rzZ5ra4BSCya4bQHLB6mT0zn7/wcYjOt1ng69q
ikCxSQm/TUnFvkh0BAgueqp7hkRF0Wo6aG3IFyUsALxulWumtqgw5J3HZcROv6AA25wtB7x61llv
6G0lmqkbKPUsDCS4rxnR7evnsmNZyn/XG5+ONJyaXpa8ALNDkvBXj0moJrnVA7rerpBAU05xZFv0
s403JVjHBgI+PyAzb7BxIOwdYWQanYvBsPcPBK5m636fO7XJQqJY+JJ+FmfVhLw3ubsyOneq1Lvc
Pou5p4F0362dZr6WBwow11Ml3VM9H2NVQn1nTQJmquaeGzbSmXaIvM8I557agFffMqUk/gLdbk7f
jUvBxRrcsAf+/x5vO7thmMhahcmUE4abl/Jw3pcNv5fCF68Yb01hZ9Kp1KghMmmQNtbWF36exFuN
viQR6OK1W44r2OtTxH6DV+MAwyGrKxV3FVJgpy/Qgir1VViIVKPd+vOSL65cDeA00veUgE1gsCBi
pnsOt/LzomQAbLC8Dx+aeJ6Vs9j2FJeQNm9J4qvmomSpzoYgOwHjyj7y3e0XJbMaG1ZJ7AX3kqJx
uLWsD9xACDVgNoB1OLI6kPKV7rmcR6OpnwQNd7WtLHBujlfTCu62Zs1C96MzGyba8qJkbGidcOUj
o8g+EYzTuWQzLDaIj/6T0prCgL6/QCCiFtAy4TqUOIhFmEjgixAKJlsrmAryJN1o+yXqiFzbtDAt
CkAiSKjmVgAklrd+cB8w1kndX3KvYMdBfd0Pk9IAR4y6zsTrG3a8myplrV+M7qVa+x9BlGCbtU20
1W58JPk7Y+q3zc/2FHSzLO2oZXB1BARYdTTQr6n+kGBL4IOG3PPKbiwXnBtuEiFHNofhXzRkL0sW
BHAJrv364vye5OXNZf11kDJ3ZgIH2mxo33cSbu1O6WgFbNFPCsltgKUijezg3qlHXnponka+VCxN
wkP2wCZ9PA57W95x2pq48Aj9+kOCh4W6Nl3QNahEpF8hNuUcXjJRutnTHiIv6dB9Tkv6NrgH4j0k
HQ+U+n7KuPkZrLkhSO1atOBcF6LqvoJX6nRoS//94L8UgMTrtN3IQsaFbYZCFbtFyrc2cIs40TyO
QKDm5HWBEm8qYU17JkNNOSJIJjloidnW4PQ4mnTfTQ/VAmYylfMfnFXy3nmRP6t3st/Mie3PjVLu
qEPoksaAaPvTa2uVjoUnEKfoOtwfysM5bR4B1ERKrixPtIvzL1UxMWLd3gaj1bnyMe9ba0f7TnN1
jNysd/yTsweSSpmSjukpJW4PF5OD4i37sX/prZjQ8LqxMZr9bnntYw9/s/aDBxixVdS7Lq/9kyP8
FIzZ4TNdnucGFKe4YugA1hnxyrY1gYm7xOzv3NK1ahv3BaDoRFAel8slSuH0eX6HMtmxmm6rJD4S
wx23ZbZQnt7/WHEXKfObQ8t7mkUetw3qMrAoleriEefMuRfoa8gBwng0LiC8w5e0ZwOeW6WYg/4o
3cD9enJDr86QjAolrSQxUisuFBGIrmixJO/DXg/TKQ3NehnWyywdiT4rRcD++yxdgww2W47K6pas
G8ACZtQh8G2LvfvxBIMm1WoI05sTdKl3f5rO0SVCQzQRME1prp4n85T86flZ88082NivtscFxvUR
r18yBotVOnasqZZewL1BjHKKkdqE0myYjtgbFkMu9LCplaGB+ztrAxnmaOliilZAmz1we4XFILzd
leZ9fONDD62FfoRtAYfgfi4vmyiblx3ono0jhl119Vw8BVtmqBZSOrgbRcBEnbFYBlnPrtQOnYVE
I8dLDK9cF37Wt5rZOUFnt9lFClCy+pE+H4TVpTXyl8Y9FSs+puJgO7x/7344dZhnd8rV2VJrghI9
MlaaJoGkceuqegKfkcaabMbUUVYi9bUJxWcI7v3bscxAdCjWzqjpeUKcwC9sdjD5H/j+e3t9oQh7
yu57ZT3Pd3Ej1lUKKjJrCoutfedhtGNMyLtHqhmWmTuybuAbJJHTvU14C5glj+eBv5HFJFa+kcS5
QPWzZJDf3TDZTk36qbI9xEciQWfnTb8fBu66ni6zjXMtVXqBnX5NUmWyL1QTaU4VS17WjeamOQ5S
reIfpx6DcrqHLdZ3fRiuBqgMI/YZjIVvlkqZ9yCIK8qaDk0yRTLlhPg981KC4PD0SkOLdq/4VRpy
vZx+aJCw4nB3iDnwUKI1yb3+0yb/KK8fqIhcw86Clh3fqeqw7xXb33/3M8oWE8JcfcWGk3Jk7brR
YQcis1KTIfRSjUP5W+89uXgKLVrakvW4Fyk1Zu3J3ELyqwwGkaWygFkmgGqZSthSbOW8zujU5HIS
BRVOQIDXcVVV3B0FwpQwvjlDUeiV/vQaYepVpng70NZdt1rEiDbKffKiehYz3FQDt/PYUvJ2zRFG
q77pJ4N1xzbu+W44F82A0oCZuWhndGAy4kRZLWEWj1StneQIuNiopqQbPRUzTz7Rt5wNrFl/iEWN
M+qayiHOIkbc1TP3odt4k76LJbgzvEn/Yb6D0ikzLJw5nPvATxmM365xJKoqbmN7UhR5sDYC3Xzz
FeqHuVceEG9ODrRU+AhQ+ouL0xREtUom+WiYmlw60mimqoctzJPkwx7nCzxiNWAKRDbkF0s2rwOq
0ZGOdYsWplchqwK9llkNHiQ7c+HqoG+7pbXSXc4EZQJhgjq6vy72C2F+rkNNe3zMgRoxKDs/GPVa
V/Wa4nqwWANnIwFLoXy+lVKBFrpOzddF/EeCoezNltqZbP3zi5cN3FebZZHqKIsuLgFx+vqz4Oea
JKnnY0kGeL9TQgtgmtsD1mNzyG6vtu61NsXGsJa6aJvNbnaz+seFz/wamPXO0jQ6pgCd7LFd/Nid
9yT2SKV63b+vEQmEnHfWcS8EZSgrEDHqN6Qc2Ig9HSQkwo+T7mWF441tyum5eFZt3kjwhaX5KQlV
Ibl6NioPXX0hkmxavt8iAnvWr9h1vbapAvLx+RzVM4zyjIh5Tvxk41ezTSnQJxzqUpzUBkoBZtee
5L/tlNLQ6y1Wc9IlnZKeYSquupNNdSLT/wahGW/Vg1WI6J1TqWGM3zFlXmRtIyT64hp7NuScc7Ky
ssE0vbvoq3tdQOLecLIbb3fPrWzbn9krNpB3VAlKYpHZxRDkW9zCZtzAEAtlq16JuJDnieVGT3ew
U/wErN/jYoPwkSdKIbxZIMHns/J0S9bPsM/+0M274PSeSx2bLnvclvZ++N5Prk0tiF3MRq//+pa4
IoIZ5QvPa9b/QndO5AReL+XejwDnzoAn5qDo6BpZibDTbIPZYvL5qUWMyLKsxe/HWLkEbeNk8m0x
Z8xo7EQlf/57efD701iqVEew5F5uboDOUECXFCxrHsJdNLgMHK/FL6Mas6YlD50o8W2Ic824L+sL
f2+nkDFqPbQ0IabiyALG6/lUil36+QK/g2ePs93inZpu0FDr4tDDCHLDiHEsbXLzNd6zQPWij2TE
5DzLESiKcdkdVR/Lw2HjnqnrV2kcuaoAfTaC1mGqCKiiQ8+h7I51ocL4xc34WDVFivnHocv4qfRk
2smK23eqNmAgSYBj8fR44ZFvneH6yM3peKwryzTIAYTB9qoc2Mttk2D0Ih7W/Q9/Id7DTP1uWqDX
HOR17Ty+o7hfDQTkZgS24N+ESElKJdgu7dPjvdCJg0u6/ofWn0I5M37F522NGBzNHK9PIf1mw9aS
jpofbiU1fsxgsqhKLsAspLo+u6FPooNWYGS9DHPISPGqDKf7oXcy9ZqxLXrY8gKdfKmw9RKgNKAo
0MXYTMKJRztL8iRS0/KFMpdqA9e/PgB72zWQZVmsLW4Vwx6fJ7N1a+ZYQw5evX9sy0x+QWasJwZB
+y98AaIGSzjKOWBxmGSRivGFSmvWz7BE7tDGyVNHdDLfZJ2HsIVnvCwziTwVlweSJ2r7tA1Ryadl
JGMs3+BQL/ZRlzyTBmGfKMTCAX7+q016NZdxeLxKr8ZCERsLlqhpVlJdkbuvjLdMslb3VkrbvzQj
YK2F0CzE2pSSKxlXxgiETjldTD+YMC6k7o3F4nDPSJDHWWuXYUIoY6kfTVh/fDSGD5F7PZr2e4GJ
u0ZYufaP2GkqCXnT84OQYdd5Om/n9zcvV8vkepo4VjIe/CpmX7htGXSYt3vJNbMgZZGNDxxORzFC
sBv8anLZ900aE/gh/ycxZAWSyK2JtZG7zUbiwn/D9TvUacW5SHlBoXt9ufgC1V+F452g+RO4q1MB
PN1HVejUoKJXOXW6ZGMhrJFeI6i8fUmTvXT49PnJu7ois7Lf1BtHzFC3HxuppVv8CpukykA3shef
LnaTPna8NTJDzkm1wsBSeb4RmHoLY4PBG16t1S7BPCOSPdZ57XiWRk+He6EhId5/K7suTKo/6o1h
mLYIVxLO/98q6SGWB97mh7CKTfVCEDQ9xsTFHNBvd14KRsgTIJj9Rof/islkkZdTR5GX9kaN5O6+
6grku6aTu7FfvuF3aH55UmbFhiF8NNE8oYxWxdWrXg3Z5agcbaRQ2QFMqoMttBVF3S9Zb0xbmMeL
EoPKyxhb/Q33tpd+V3gn2eDJRSuTJgXfdbyGxLaFODvpHe4skuqqQRIeMnvFkDmE+2EB5yl7tSo4
0u3rhZA8YPw+i++d0GuZGorHD76Mh+dtWf7YBA5Izv3wIcOO5hFsdH2uCF93tlUU1Paodb4sEnGR
uUcnhaBgcxQs8CeokO2Z/bMkw5MzJs2nCtcGnnvdwV4J4LxrI6MhK1xSnSdTybzGAR3Kx41VDrfk
xBB1R7P6KE9C5AjecJnLPtwWq62j5XP4DnfhUGOibi2/Xrf2Srll3H7Pnx9xttY7XwamykDEREpt
s2U9ZJL8FI89D5idxBDuHdtFU39HGJ4tuY00iWGkkFvbAJJ4ttRT8KjVWGC8kczOCO5iYC/EvHeP
lSQVC9OTccYBp+QBiTLBEGB8NwZfOvIjUM3rDxWkopzsMbCNLMzLCISQpgOOl64NhR8baLk0oHiR
mfERU5xlI+1z/9qk79geprvGDeoZGd4mDiAtCE79tZ+CPApxCr3jA6Vq5mHqmDIM8fb94hA84K8v
nI/znf0xgDtPkaGM7AUEqjQsmiqTPV2cJOOUCkYC5ZxVOIj5iqMavkd/pXGEmSoYAG92NYpHOXsF
qCcxRyNh17mrxo5hmv7viXzXmJsfXnXHiRcHmUaDZKQ1PQsFQJvcyAx4QEQ6OgElPv06jipeelEf
dm47wPSLGX0+1egdGUul6lyRkS/G6+lZLEGAP6SX1h7J/oZCjTUeOqs9xSreJ69EfsGKYHaBVRMT
O9IifRGUHPiR51aL3U58CzROQFNminUnlIeF2gw7wxbEKf8/4eYP/QLFHk+qZkgrbjUiKA5dFr+h
4BzFwHmxjp5LmwvT9OrNHJru7udEKYGvxNhNttC4Jif5SXQ0emDK+ZD5d7f4QmOmYdkpDHvZFLjg
97EOinNv9HhplkRafIAUc28PXzwUoutX1jpTYAAIWB1g91Bupln+DN6Ebl5nefATSyHamc1QXc9z
7CIHNwh+Tcd3nPEIojL4CKYcLvYXw0jyZBeN1HQysK/wKSJmnwEFNEsn4G199ONXkpI+ncrStT9M
dnCLpeKcR/gR5Tpl68ZTt3o8YkevOwpxTbTSCi5WzJbRzGJ5M517s9hHrXNrBHMcYO37798TIg5U
PBOD74TMxRfy7KD7s2ut5Q0HnS6bKFTsMLmLL/T/Q4woPahtadM4K/zyWiJU3+DZ37MCYPbYZDk2
P20c2vhge0Y2KtvApct3641IROKIh8uqWxv5aOC3FFbhajdAwhhVTqzBbx4yQGT95TLHfRpvW0hI
Fi9/YXuxfbTA137u7ydo4PApU28tAW2KSFmiWhNOSa2wOU7OULlOcteXg7afm0Ud6N7Quoo5Qljs
jVJ/U37/+To1yCbz/jSnzKFWELLsm5sJQPGLifmufxpjAMHvhirfWSORJpoT4UAhnkWNqZOyFoki
0fmaKtUHJkc5Y9340jAnA8ceuLlDDc0Xx2Xc5gkNLWAesAcU2pV+MoXK1FhT+VyPtmSz8k5VIa9D
roMcsSjHhIUGJ6z5FvkEk8+mEnZJD3HlIogMiUZLDplQBf81tvNN6BftITsBD080QNcJiT53IkA6
nAFvcD2RBkKlAzHtL4zjf68t0udV1+9gmprKdOmLzuNz1huookjBU/6JWKrQYJlJaoi9DpanIRfS
e7u2yI0SAX+4151QkrF3B/2JNFNeiXfFMFafSA9/6tTkK0qDYkHtKK/RFZetxKiawl2WbBHPo1V7
2nTH3R0fptOhk+alTftx5eFg40g+VFvTLC78ukt3KbY3+ehgDr8cm4j+Boy4R829UYbRpeM+GfrK
syTkn1I7lmg5G3jS7eAemKssEYqYQ/uRpRyrbtztEFO420uD0IuuO9SXXjqEvCH98SoQFJVU7rKD
Ik+TAHtsXd1ySj3mkLQ3wqPc12dPG5kDLeUb/NOCvQ4P3I3aQqQ1TFG9wuiUOWn7cjFCxn6f/Zp+
x3KSLkpnRXb/Y5RJLvMkifSBmz4NZaDaTmgOzdhBn5ZJjNlpfBGgebtkBXeSmqywljj7aix6cyXq
qPqfjnrWDLUnB/NAy36LOA5xK+64Y7ww5f6KRZdVSg57PwTiRuHb5M6UTAuFq7VrxE+rDlsvim/m
tyL7RNhgZ0eYog/ef9+A7yXIZnpLtxSQNJhq2jaJzf2lCMxTvqOX8mzbEhtdfxeQ7/2k2q47m8wH
saGV5ajiXEkCoVaCdgSGT0Em8scVTY0hKt+nMWnEze0O6f/KbXxdnkkWtDilpbAi39tXFZIn+pKZ
BfjYPdpqW/+iYpgOvsjIYOwLt56dPTE2z5H2g2navJ88n6lmwIqylnqTf77CohRsCZFQErh9qiIl
03Cz7mJVznKBytrjGExoHog67gemyMF6W/c8snZBHjY4Y4d3ENJtDM4Z9Ov8XO417YKPjnz+wZ6U
zX+iuTmJuXSuEZb0/qP4o6X1qvr/w2CtUiBHY2kNdVZ6UTHp4ZkYl1MJEgZWhbzN+fqXuIIdriMV
6NR1CATVpGnvi2w8ZfP6FyotPHbV7F1bu4WrmJbvGuFxzNKxf2iqDncxu4yXHeWY4txM9AoOR6v6
DEisoYczybyEd87W85eTkbALQ8+8gjs/Jwg+2pGJCRL+uVgi7J3EcipLeVuQ/ClxWW5tRZJivclf
4VykHpeiCDOdUWkZScA2/aP8LDkO7ILIH6XO0WGO3NDhKm09QNQno8j5yAsSVDPRcwwQ9/UaG6p5
3k0DoLp1/2NyEMbLUCA4reBGR9hJm+SKviACreIT4tJFJyyAFIKcVu6nz9rUt6d06Wr3yQlqVIA2
xHOqYBDUOgLrpP1o+xgEvdBZ4+LWFH8Co6t/GexazOgpQswYL/OXHH3sn7/k5cVaQ6W+cxrd47Y4
Kev3Y0XDwc9xhQ14lwRgv7W5iCF+ZgxMWtNhTzw8ltMwY/9mOCu4yA8gL0hliW2dpwwfNjcOvGnG
b7NdHoNgyRywDG1JOJq/Ca+/BaMEdWviSnDK4wPyayS2fnputVSpIvG17O9glF1t05MQHOXGe/cU
WOGE3IrWvfxwbyUHnQX8mHXdMgUfC/4oLR6Dd0XEMZnzfvBujezxVNNsu9ID1IhdSTu+y4WtPeXe
xnTsJrjhyabVaGoIWU87ok7BHXsixNUWCWJjx0geHttymBg97w6ea0XE4CWWhboZFxCpss2sxrZX
B4IbSmt7Xs//AeETwUlg3kNOg+vCapLy71fxHJiAyn2YR4ozwcJEl8v8E10qKogo14Bw85DzKRzG
Ns+bQfWclfpaPREll/lxdUSwSxaN+LLUdMIojkDegnvA0/Dp/eu4rWl7Tef6w7Wzz6/zvKPGgoF3
45ta6+WPAxgMfPZdqFOlIB5AY9rNztqjNF3pJRhVK48AuoH7bzT+z8fGIGOTsChBtIFSNG4QRHuk
kmtWnKSkjcq+kaXJZU1mpixqThqPZjtDPAX6Crol7Zf2swFWBMhsZT+9N8O+tcaAO6piWJYAws6j
bN/NyPUgBJBoJaKgP415dd/caOjECtf2MhUlXauPpXiY8slQZ/yg5exL45wTD8iQOai2gIHFoHK8
vV90xJZFFgzRDDo9vTeNFIk5RgATVeL8KOZ7uAkTOrirhxy3TX23qON3A1GPrVY+Rqb3rbL3wZwD
DuK1ftY01+KdjYRhlOPGcMFcCbGN3TKTweF5Ycxj4Me8QMiWajGNoaVHPbZgfLW0YYG5yBFbQTl5
+iypSmCJ5zF7kE/xncDJArZOecE7DBvHJan3oXrveVGgjvPMJH1fayJvejOeJ+kgY5r9Y3Kpf0qc
rpKqW7G4j3GCnusRTcDFv2RNQz7PTC2yaqa8vbhhJSQfUqcYmW9z7Z0SxBQn3SkrBPCp6AZS/w33
pzCukuxRNvTOnJXFuLF2jKoSqvi1GQAsqdpm6bWolFPL2lSoXFXTqMqGXE1LkWPreUe0sIdXSL8m
iT1o/4P6PwT+3pN0iYYr1LNAoJL0gcO38YeH0IpPHcC1XjXtKjiohnhArFzcEhEZSxtlV96bX0J5
/d3CRgIh9Vq9w3JRP73Dhm9mK/ihfj5+eK0TLFeeN/0Gew5wWsVhVAvTFh62OSuvR0/jW22MWLVp
IdZRhG6tKHfhpcdIpNI63/YJ2PtKLT1hP1wXSwsmUsNc2aX+87UP9VMiElMtHWKpcFEG9eTvO23A
Pb42kP1MZfhKQIo3dFTYGuGASTZdHE4haeQM1cmUkwD7MoaGcE+oyTNa1en9vVqNJj5e4oDyJfn1
Dxjx+ok/Gndjmj5VXUqhEBWP5I8smu+NO8wr3v5IXUMRqHTe0ANm5c/LR6I0HjNDcmO9NW1CoduX
Mf7qFfFTUed689Seqj/esSVXg574Qwdp3OsGdDCM3x8NZXYjSoyj+Wbs5hQo4fONGelUevp7c7Mm
7t9hGK336HSE9bJKZw5kRZgT3Sc3BZzHa72wC6aCls/uQLubFP3XmWbQO08Ip1aZ0OhPlDaKxGkl
FGdCyj5WcA3UkXnLXBK2V7bnWfRZtUDkwNCZH7lWu01VN3ruTW8n9QaAtBN+GorTowg+XUuisbAF
WXGG47sxltRLJhMSPOna760JefFz7B+2IR+AvmXLOWyV+Vz3Ry9BnbiV0pdjno51QvHHYeZHZRmZ
Z/a8yqt6BuVjT0b/CcZr08aiCachTNCvTWrBG0Qan2lTC4PPBOKFW2BjoulOxfoDovMVoSVobGNM
wbObzqh+k7vDFYMu2+CZyIjz6HFBFmEjg6+aYrIcTtcEgBP2njUcI9kC3T769AFvZzaDmModlAHf
ceJTW8GzAO0iRgeWi4GnX/5OheDtrzkm8eArK1M0lqk6z/9FRVyfQRFDUf1xKxyD5FdmZLzZKY2M
IXrpi2fawJt36NmGQdY6/maX4OlY5nxBocnXJW+Xt96PkKqrOVaYdK6HissekQFwxfs41bgHFAsE
QAM4NwjirJoc77BdssblX9bFFyVYQ1rGLwMgag5pPU7yp3t/CPCq3aiEgJ+k9SyYy0WCLJHwHAbj
FlDZ3CmSS3MMq2Q+4aXqkae7JNr/GMnWv+nf2CQP3+SZkFp0sDD02iTIc7flO+VVC4SKBBoPLz65
M2qHUbL6DoEPiteQnj+OgYv7hykm7yyPUY1iBmWkbTH0V3ZwxOwBh04mNehaXAElxDFkOb9d8IFk
KT6MQU0hiOXiH3k+6dDwETqa0a9vfOD1CplXeGeqYadbXErDtkrNXssEKnF+CeeWmrSPlRG+wA5x
rQyXaCiPOa4FKcm/V6uOADFhs1J8yWGqWgHI9VzbSJDTCioonrX2jHKvWOfEFfo6td7Xi669SSLl
1UF9QFLRgUyIGdvnmt5KaLIO/3XYqqmIdPhh5F3cKaCl5dVJfHau3JId2tfyk/P0HKDO/yohouJw
qBPOn5zIyA+Xlz7opUoAKkNA/8LHl68qW0r5cSu9y5uoIjSWcGdr/8XlNEfr+yI7x1Gtq18bRluK
Pk+7k+kM7S7OtT41ZNMYeA8+wTLs5N1W12tiP0zx4VAVPUckehbjZ9oPdlh+SOdJ4PpzS3VP6nt0
1q4I/y01KnRxDpd9dTCDa/L26ereQAUvBfpS+fqrhOHpsg/w8T/GmJPG7hWocd63PZWe9ziVxdmE
vzYZFgRJ8akanHcca7Dk1MWSOfmNkRiCkxQ8QWLNgId+VyuQHGA7dsla/0Qpy+NGT8H7EufiwGlP
xAETtyPCSZasDnbvVh9Duq8rG+F3xXK4r0TU+UfuAxzqLlvRkpzO52wseckvz1lm/LfepyvyTLkH
fNzFNHTfAAM7C2x3qbAL/aafaevE6DuWlhneRp/xChxQt5aW42aWWMf9CT3d0Y0k6cpRyQyDAa/B
oaHqLSGE4ml4Pj9UQuF9gbi1xIP4xhfZOWa/fBADubQnOxfEhVJ24HScBPwBgt+gru3bgQVbviGe
TYngJMdGAvPzHmbzjvDHuYj9SbiyhuCUlgt+GzwMuUcaKEbUPekmRpfyqEe0E/kCt3/w20CVi+jX
1Ky4MAlJ4jOVWx2ZbT+MH1qWeAn2WtBfcrLohctG4+uDLLzsYmqJs+RqcVmeyZm5Cj1OXcXvgJZS
zQDG7EoK5Mpb7nJmZD3O446UGw4dSiUNLRt0dRRCToXBVfheioi0EsyneWY6JuBusPACyFNW2mkw
uvPI5LEyROGvMPVQyZcMYq3CgNYMkaVbpHq1ibNo1u2bGhlz4+WA6xqZVwszFDLF003Wnuw7TuMh
0142VPo397n70ezorLuEGSPWKe9QfoDtsJbEd7nFkihQvx6t7rbabWHc7lYrzKjhm8cqZmNi60se
ypIODhGzlE3tTdmBBOOHXaZt3+uogvhfVXkzbeQTY03cYhBbFJaBYewwQT5VbZ8QDBxamh+6sDeY
VxNqfP6C3P849LalB0trURKhCWW+3WqdQFPOxtjjT8oU9E7H9HnK8HmDngYl/oFgpEBUl5Mul4lS
IwHxrKD5pueWGKo+psrd3r2qq/UcVExus0lvM8EC0ivJSyQG4F9KaF5svO/RHNjUBV9ciBJyr6+f
VvYbas5UNm2YF9PfcEiWXPRRmiBVjanIWzh0WeZE069GWToBT1h8tfAVw0MBlvp8G1LKTODVLJhW
6CBU1jC7rPw/JLHJipSWEzafJawtS6/amw34XNGPQCZSPFIF5WJ71+O6PTHMQ3E1UaB2rHlwUvQ1
1SdXKEBUer5UW5dZzHDf0edMw3XpVHWhwyBbPIatYCLZ6RauT1XcdrLRWkyEzEV8jX4INtTyvEB/
lPNTrS7ipW4E49Gx7b1yShyqFoNBaoastNyKsbYVtvdw1lRSCrjqkLBH088qr79lHfm3k7bwlYEH
nMR0vEj978YhSQESwE6Avo6Uh9PfN5AZrL+yF2xely/xB3I8DLXt2QNUYP+G9IEp8BbizP4LqhKX
H7GG/vyj3OdKYi4lNDeCwf6UZR1dAnuQxQaepW5rPHns8kUcSYAwGD9PAZc/l8d9ThHrj8CLhPeV
MUukgEjyasNPjuP4KoGjOVzuW1nCo2MPN6/GkfWHe3NejDlNU5lgZ/sWqHNshLwhjz6pyif1POKN
lY2LtVoSSWeKeArYSAWgvrGiBHUBvPxTRKHTi0I+arX3saYdq3WQYkSIajhY7WFgjQdarkyfdzoA
v3r9gX/sru4AwHS9jsqAUayWfsN7KScaNBj7+jsOqTvIGFqi+D26d0LGWWRbT5jL8H0/Xj7wGxJv
bFbzCp7b9nd80JTCBj7FKvumwcfCve+buttNh6KmYpMyTtU0m5JguSWKebdoSd3yrQh3Ji6Exjht
PYkFVelBa0Oz/zFU4lAn+gCUYIK+irKePs9QsmnVtrYL7HIFN90WkmMuR6c7iKHkwal1qX+z9Vur
uAcBKrlWpBvM2wpGhf3yV45pTcdPHsEJx+QBIpEsG+kypDtFiGvIXtEwD+F1OjDu/a6z9PvQNf6A
iDRG44HoRPxJ1yGNfes3dbLj1YKcQHeWrTLbxacFU2DZDsib0sLyK1UNCtYTazzQHWBmo4qWK6rQ
tHVBbuWo4I8JK8LyaO3HUlYRVrwNDXhKMIDHwCvNEO7sG5oSVrGz5zRqh0klZ1hcYKCJLhQGChzY
jW35oCO7pn8h0IG6Wm+UINb79mZjt5RzNv4fJNJrYQ8P2ULCsyHbgh6YTxtb55R7FT+KwmF520kR
1VFuVyT/tO/9jsCuLLvBWxSsy/gpQZpLPEVMi3RxSm+tsedz8xZAOsfC3cTcgMhs4f5zVXa/l8im
Q8HS2JsENiDSjUEzQw3y23doKadc4E22lebm8eNZDIVziCHMP2fTNY3yC6C4WSHsOnrjCpHaZwpy
KngiKRO8cuTgnD+pFPi57o53r/X0k+Pgo3srSTzMeqYier6SlXoxkFkS0E9qRNtSLlXI8D6VH4Ft
CztuiaemgeSEt05LDMO1dt4/kifdYcFqZYAjk+KcDxyaLsABJ5gMZC23lmfiwjfRf5EUe/oJ7yOS
ve8VDecZ7BBnoaNNlHEMTfOa4/lnaRQBxfCd47gqB5dq7/22Tra1CZgp7uSXPUks3Ug/SDaNsGok
9203iAuonKTAWz/TV/FIGru7/M0YFanM7jmCIsVUUiEXGHUIN1s+XO5v+AZXNpe3sBmboKVZzUVQ
yvqVT2DJw+tUb4maSu+MWmD4U3lblrhU7S+HzrU5EEreAhthAgoPqcSxEgVqP8X4MTG2bXdKfZx/
hKp/Hgk7q3cdQ+Ux9RGIvaDwsK+WCGdwvVL8SiBQCU2hdB70yp41/p3N3DzrwK4+MKbmFEqOuiAy
BROkji2JlZIXGiRgrR0KNHjGXMHTa9fJ2UoJfBBRQIpo2kOrb8xYz9JweBg6sEqFyAFzC5SZK9UD
KAU4dfbdSBfs3RKUudTdABAeCKtWsxkSye6PXozBKQhEfygU62l7QPUmlGhyd9e4ixgn3iCVuF4Z
mzVbF3E5clK6jY4FKPRWVL/IWrs7ntekTC03nPUjGtya6oOtSVYAqNpT6gVjC5zno32X7ZaQYMTE
+DZ0WooeY11Vg3DKSUGXwrrEXsM3feIi6mk8o9+vw41+CtbhUvIqIwoQaTDGXyAYcw21+cggqYxi
queEd4ZrqnoWSMOmkAH0r4+DpZ8U0IwAA57VyuwTEFrFSL4vPvB50OXFbU2ta1zQxwd1SUKRyZeH
OLVM+JvyXQS4ZLScL5Oc4RuhrclJp9qGXVZtTCQWOebvcU8N8r/IBmc9UNAxc9GIPi5xYPPEHV+2
+TMi8avgkKBX3TpNXl6ZubSOCMIVBz3gM+oq8mfeKy2Elkbs3AW+VhgSee3N6W8C+hvx/2W/2w48
TWjRaZY2WCj3UUvV7OrN5qFDwe0ctRHqNkVfeBPXdrKPQrGfxtKwh7Q2Dg/DW+Nymm/jazsTr117
W/SrJdUF9kF0GZ+ICM72Pw+dPhcHL3fB2ZODu3+AMrg6EhCAloQqeS1Iz70ugxxsGE4Sw1xu9NBY
mLPfwv+tT16e57EuD4tOcUMd5gyQ6U7yrM9NekDWdmfI0NU8BiyebOngtrF+CFJw92GiUeQ/JOup
g+RxNs9fBjOKa9QTXYNTq2gw/l0eJ/FWwrxTiFdaeIgUVsPH1KsSGd23wVtMwK6wsHGLhefyFSAy
8QEpvQOcgVCuvTNZvNxi/XIbKGicW/GYeFbZRklqArQjdCkbiLIX68bGnEZ+4osNN4Yn9OSS3ebZ
IbIch29XMZTGwRNVgfmc8i5q1XvtUCu/odDp23a5POtLgBSswAG5neeMoWhPVpS+juLAGgdcXkrk
MNycxbvgRNakZHx9FKSLsXAQFwy/EGw82WlGeBljlo+n4MX0KbbrgzBhDsS9B7DGPokQHY9DE1Ct
MGG88Cs3rQDgD74i8va2HM1lD2YvK9+oGj/suIBGuY8eTiatNJfPJpoB8G+m6cuAVV2EccAA0ekr
KKXV6Z0CUJuhfRrwqCnlsA581Pbu7o7xbFipToFcZmPi3QeGItPW4bgwEiV9tLC9V3dxwlvyIEN6
DW3j3f1CNYDrrxXkrMv0dqj1zHxE1vRirhpB23bqXD4A905QjGw8Ai1xGwFvnQuvEUHcDSArR+DB
s9yucJnaBGSUduWld5duEGwN9diyWS7N7GKugj/04cY0vMuI6wicLxWPsflMT93LV8a96utAez8U
chdVdUYgJx0TNQLOvH06WJ9ISi0UIgnNfVx/RoQ4kYD1l6qBxFHH5YqBv3IUummdvV96a1NpXdQi
Ha2GKAFDcKJtm3XsMtd1zv6h79e12Q8LNzc3XmRIfL37wPXHcEy4Ib8JRW3Y+DHDnAoq1ix0Lp8K
b/mc9OhwIhUTqhC9wfGYyGELJo+XAnJZpkmpmfUmswUmQFIHbC4WYfPV6XX52vz5kcQ0lgFlS6px
TEcw5md7eznVUmAkUZy6oFooxoaVrL+ek3sKir7Re/3FW9RgMQHjccbZR4zZF3q6o82g7M0NV59r
x1s/+7sBhvOOHhNo0tTlva46u/et++dleCHh6lU+8c2Z1wQyUOWyzq7fXDcxshEA5jTp/r2vVBrv
JTTqvVjMsnqtvshmttbkSHrehQmg3uR60WI5Ha5aImGDh5W6kazlCK2N2NHz5w6hw3nVp1adXPYD
YqdR2hqz9ePt26X2f1vL9XHGnztdL77kkMpLSzmHfNpZf85ZEOYM0LhCymURaxKSd7Ch8grpuj4/
bzaM+cVigIq4s4N81KcfUr6q9NBrjUXuIUyacf5wPWjREKzpBP+n6cOJya21RuibZaQM2PBRgQWH
fiwI0vqqhEqOwf1sRw/J3FsQtXwbM6xM8ZGrbDFNGlUgCWq6kEjtOfbXQH8szxShkZQMoDxBVAIx
jZsb813gSCs8RsgLbyI6jr7q++7qCJC2zJojoVqxQIiVziq31tyPoh4xwc0ePNj0RvGYIznk5uLo
gHryHjDtZIDA3sP7NxaFjRhhmJWfoHwFWKdGvNWDKzAz91ylfKLv8TNvIoID7cVMFScHi2N9R8VT
KSfij+8OoRLiN+DzAuFFDVuNCuxeGcW+VsTlSYOl6wilrktC1xFucWgKcjw5m/IBBKYI5LYEyH8x
iNjr4sfzjc/zJiKxlkeDmHu/RFwiyl2c7ZwHRrFeuUumI3WWTRDwHjrtrdCwPyBFuHsuBm3i52Zb
yENjOs2FAomt3lmR+URGyDcnqbVMILZ+O5dqhT2gtsMr7GJm0QyBERGuikt+ul5DaSRdP666+MJy
bjZQAB0fsJk87wsCfxjyygv07LK4iVcpLPFgMnKSwvejzFipdsz+T+mS09mXcdTMjH7m9q+S3eBm
0gROQomChBGwQv66sEb6d2cuJzTIhDYSL5W+rnBkDsJGpJGcpDyyZYZO5qa2zByPov3VAbovCm0d
INTMj6IBE1W2m2dX8wQD0AKjwPdhY8adhvAHwssrsbd1ZUgEpTZwVweQVI+9zO5RFSMc5R+RNCZa
83tDdpdsvTwT+i9kooxf60SclP3PJlNCCTBsWgqzc8GuufLrfoHNTeKs4TJPDgo/KSH7qmcOKI3N
SwxQim8tK0e73CGJdlD81Ws9aPzYo5LbmuZoNuNI6GXAoWibn7MG7twxXSKGHdnrAPS2+6sYK5K3
hu8TtZ6teOeR+nMvKEjYl30U5iPjRO9ZrQVdSA+YzPCwwADu6OUaz+bg2kc+BUtdbzc8l6f8VOrz
w5BUlEGOfy4IcJbe0+zL3KGRAHTjRZS+04AteSuAgaGu9YeDg4r14Pqbq5lwIc8RL86PZXVScNBa
FWxY2TCpFYolISEcVX1go3Pez7lIoRxY+c8YGthFrmrSXg5JAqQe+oD2DFvzMFI1PDucAbtZFI9E
RJUx+TRsWfDEEZTdOYiOM+H18BfLz05WxIszHYlRQe1UUDWaqAXbs+9OSs/7MLYxj/KDhlbYY+W9
O40ha7vY3WneJYU7rBodLefP5K/omhxkZXkOY6L4qQdfduVAF7WNd6rSSv+houlOPekzKqvscIrG
/eZMMnrICLf99Q1kOwfY2n1fhQ3cfZ/Qaypw1wc2c3y90FpYtR2dyWjsXSfPrDMrARPH/kjjPGsS
97rvZRZw2AqJyrIDpdV47f0vQY2aCn/Zbe/DlIjYX/w7TtMTFTYAaZcwh4QC16odN6C+kkaFjuhM
V5699PB9Lprkw4QKrwj0wuanarzKqIPCLJ9Po4wH+RQ2gnAoQenglRtY8bxhlVOsfkbqStQEnLXH
UxS0o1WG5b+0dAdSjR9JZwUnhVTUQIcyXDJbf5280+G07i6t8u5QcYpj1tpsJdzgGXmfjLI2OD3G
/pqdz87WXEtNQhVkDzYWWSpUk9BrwZqa8C92KgFo+E0NhTJNRFSWv2Og/hsJ13oNrWGcBjI5cvpA
7UJlYUjnGisE/xFIZS3jp/wnUve126TjtvHM+jH0LuXzFfuXCAtQTrww56L4qIaRhJUEGjHFRZqU
jOjUJZNMg9F80VpRZsmP4z/rUBGco/XbNgWYpwiojjzmSCswLGEcGzTKm69aSvVH81atsJh3yZ6U
Pvs3qaTP9w7kt8et8KJ6S6c4zD4myH7mf47m/6fo/b8KXnfQqLNmOTP5uGpciQSgn1H8ey5wB4gS
4/n6VU3LIkCHhUtj7peOrwrp1CPDZjCyX4XoM+96C3woEt7dDkkYIONP+iqPf8QBNJr2O5QrxR2d
DZnx+C7K6G4NmATe0WLRLV5mtuRrgBrC36sqbK+Lv4DMQ07zpkbqzsmRjxinOcxMtR2bBuK9ez1Z
wHaaVHwt6GPKHK7EjZeAKO4b36AdiE243p2vFBcbzcvwIlyMtfZ/8PcYLST4yNy4ha888PnPPN56
7yIcfoIN6opvpvCgn8OvHLooYaBsT4dsL/8Z7iZmkYqu6xmEo6dsFsWkJoxE5yk4rphZ5ZF+58FI
wpaImcNc06f0TLe0G1CMhUIcOD+H0/75Oc2q386TbawZPmUO5jzmYy1SuX7BLgK+b9/eZc38mc63
rHL6eZUBHb8C2bJ/D/HFOg38dzwITlClQ+d9Tsrafj3h4XVIyH0sxBcnvoRssm85+dnsRIiGDmIU
jHSd/coXzB8S0uhWhBV3APB1CogBmQyAxnAhQAC8suE7avOuWKKqRRbHwNjD7qn70puS1jj+eqim
R2lsKYpEw1EAQm93aVganKaki8CUMcRt+Ed7ArGAttSbIcbCJVgZzfQGcen2aiez2ruExbhB2Zg2
KtWQeVuN91ej9SGSssytwU6ah6VIBwE9mSq2zcXEu0yzHks71BthDegggZ+Be+PNywOIg1qbM7UX
2YFa5LiKpplYhO6cQZV+k+Wz4+F1Zi2Y21geqHXQ93oF26Q7mNFR6TKXDuZmDpymTLtTeUxeLcD8
pwP9t40oIjtJvP9cNtpdI9+qcG+kHp8w/9zHRtU9+AvNcsfnPvs0gUPS6ODt88Bo4QVijaVvChVx
dpVbWD3leRmHiClkPbIpalruASu4+nMHbae/O3zmSrMJLU/jToSW3d5UKEk9TU/NNnF/ComvXg5I
LghU+zRa+0jeHD4TKSFl02XBg6ZYJ4+o/WnPHuPNzZcFxvbspVgDPnVG0LMRGnndJ4rHTYeZ1JeK
kEyixa517kjZEzIGFmFKh8NGlFl9+SSiJSV5vTjGPpRnCHby/Mfv8LfzPiDFNTp8IMieEChrr/VT
zqUmoIYNVsqXQ8W2ko0r7sISboId+muq793axywiIM/Bobs/CcZsyeuTWM3boITZon+nRkSbsbTB
IdrnpDtY0qwiR2IDBILxsiVKzgSEcW4VoCbmZkGNCMbjiozEuXFYn6a2HUrO/hxmuRcWItps62XE
pCSKGrAqt63BLAvLhr6kuBE++QaGy4I8ECrtHs+viFrmr+sH61V6eyQX1HGARSXvRVKzX0OfN/FC
Csc16L8AxDVkoLEyUfgI/vSjb/4V4byLwSl8f0suCPsLQ/YnYcn2Crm2AzPL4IIEroKdEXeie5qz
RrpUk86abR62F26ctEkD8b+ERm/K53o0DOvFdBBZYyeaO297Rv2sWe8Jl4tXaEJleMi+lNwRaT+r
nW/6YwkM/UddPOX8wyruAPhx5RJoj28Co/o29z2lGChkSOsAo7L94kk9D6gFds0zCosJEgu0Vzqi
7DWN4iC81Dc3q4d5Fdb7SJ08U0dD86Jn/P3p3+IKyT77wAdLNqbxZwKuMnKzSKOqFiGiaG8+Twy7
MzAX439YVqGCjaSm+OoSn18c3VPQ2VUgSGPKaJLmw3NgNQYQn9TebO8jWfoQEvEdo/0uAJMN+F8Z
R+0tCTSoH8TAYYEDhQUqOMAtbbsyDxgxADOJbIkSznP9wmAx8JWFNGLPLpAbhrX3J9CIe9Hx/fNP
HModTyic0mHKwZkDZjq+6nOEgxK8OUjAVvCsLSStHT5mkXnDgr96rnH0Jl84PrboRtgOPnHaEPo8
Sa1txkZRdKIuwqkzqukjoUreu5rA6TMa9uFhjjEXm5TVI3TUsdqGbN7pwFtweYRGXrNgLCmV7RcL
i/DwCYd/e1/2F3owWO6tzHj+G7knyZE2vnraLB1Ac3J7Epd/WK/gwBzYTP+MCfZLE1eNGi6un8pW
y7FQT4V8+gYuZYkf2nRfv5IrdCJWnU+W8c9aV7c5XXYdeCI6PT0rJP5FmZG4d8VApKXLmq+UKoaP
AAMjNPqZJO4hgb7mD4MOT0QdRMrSp1Vc6TzjxKTaBotoJ4vT6Qqiy2gcEqhtLMM8KTySyT2nMuGJ
GYbphMdWUPGTH5JbZB/QMnty7EyUMrofE3+fAVucWREyaOxMaQyY7NbhD1G029qrE7cIgKkn6Y2Q
ph2RLq/F1mMhebfvKC6CLYy2/MF3HwMqE/ltQPGYr32EzMvb33/huFqbdvOJq0+hysx4cBeIOgXz
v4pmubbNurzkdt4BXhCjh95GG6rJTS7oJzvn/YxBVvWDrwnNAnW7zLEfiih/jZcSGLRu8Bv3Iuo7
j+W9hE3aP/NUPgvhpfClmNrl9aX4CklwXAWv/3qocmb396vbpnUZLNn/GUNoz2PkuXKfkcLMiV8D
iG+OEcpVNtzWO574vnP4USB6nwAAWIeEAhIClX/sdfPPDX+ih/NxxJkN35ZO5JgkJGJv1cinuT28
TG9+EZqrI+HbOEpOjh6qHtsc0nkacEj9pNy9OTrY8tR854AxGQDzmO32h7vkKEUB3RYNla0clxSW
yJ0rt8qCqYD2juQHKqVz010celmkf3d+FAvqx9opAp08a9xdScLF9Y5BBUkv5OMupUYPWINzAcsn
2ZJlJjFh+svCLkdwj7ivNBbVs59/KppGmtZJFZJxb89Ehg5OMhAlTHerABLSu+Yi8CefBS4ibQ+A
63ww806zbxQqIBAGrC+MyQ82vPbR1f1/OBFOfXR3v4xbEqGQ61zb91RVA6462Z4GMMePVhGPgoSr
qvixTm4REOdRN314ysLlcUK6Lu0Xo4rOcfw0CCVShAqrnbJ633W7jMg1BCzKQkvz/ZFzQCQxu1pd
LLKSjPHIF46QhNHPlxpiMJYWOfF170wwLB2aC6rgUbavjvUDURS7ZB7gmhuDuUOoOO0BlpYGgLdh
1CPTMx/AvoZfY2kS9rOf00BpubE/xqR93JpLVaq8LKIhlxwWCxHfW89jPEyaOs0jpTBYPVw1y5JZ
21gtWE+9oivtQsn94qeol44jUhEjpBEloioy8csXGZNu7Jt0VSaY/fco2i6m5lcntutz58SAPExf
1tKsgqUNldu3R0cspJCJW4FbwmpsprmMuTzx/6QJAl12UBgSF/26FXEq41wCgw085IbHy65i+bAL
TAtOnovJSyTG6afSHmuDrrA6btHFZCobqo5TfFFW/n0JHVCsV2cPzUNxR8SJhPE0A9tp+cN6zRFI
0VOBMj/JPYCBSGNvEMWuSh/w5zv+GnHJNNVW/Nf9HF0LuZTWMnx6E0CZ8R6kPYvsC5PHRwtv3gjM
y9x5rvTs59anIWDkvUAV47oq8d/tuoTPkW3dRMt00LTPjrtOuV2yCky1IJBpsI58tSY8q/dx2Xz0
hFNYc2judf3On/vhnPoxFYScBRUx2F7UBt7iYInYX/0wvDgQGAHSdBMucBKSqTob6IP85O5Wml11
Wrx3Wnddu86z6QuRrK/djiWx26T91MduCVkt82uFU6tmH0DtrHawth2oMir88dkqt8zv+EPNGM8n
niT52HRKX/Pj17rGPfBVxVyuP9jvRbBKs76Zb57DfaAwFftWyovTdqyjAV5M59ESvmjSMKoTGoo+
DyA/enWv3I03uPVzq/RlSNE1chHjK2ghQO2fXCscWlOU5F8TUM2HPxHKEAz1P24BMEfiVOPEL/xC
KuceRoyH3bDAyDSaXu4eJrpMm71kOOMyW/K5TC8QHCLZfd7CKno0fpmyV+AmQDUaUbWlZnw/VpTa
Tgz0PbI/LuqUbg1thg6xaSOJ1RHsqIDLhWGPKl0wFWJj26oMs45jGJNohRl3SSagd79JovuHtPrV
bVY8AXdOpi1dCl4XvxbOERY0N0vWiIi1JXl68u+q1BeTYrvzEF4VpiKHru7LAcO/ZGifPM9rGagq
Df/NA6z22xEMCc/IEsY9Pl11O/WnR/maGJRpzNAcqvDuhz1Co2/GhbgStR6YXYYlBvqtkG9ZTr0p
kTV2L+1RkBki2i6ORLzfwxGOXIeY7zEvmNlBfWvKx1YkBnaVeMsBIuJFYUsXFQBrh+Qb51fTExEQ
FKrtr0v0AzL+YuZuTCIz4ge+ubEzE83b1MoQGxJ49qXbE3UGfBSto5sBAw+spB8nmqnxhiaEFACT
myGT1AwljNe7CC4u4AX5N3Rxjk82A7tEwfFQdqCU4NzoWlQyAmdlffCJuuX1oj8OvpS2WycsTr+f
RhzYjEhHNUvhF0oNjZiU/FJpre1qQSBwTobxgKHgQ6dw8hcXhdER1BU133g4JEe2mU3jU4aKqk6l
mOL8r5z709ZtmrycKQH5wuTN4s3eWQZ5legYN+IKPD4GceTtlS3bksnuBRemGKfGYVOeAV5Rjf1G
1a0ExxTIIdE3S7cjGfWTEzEdK5hY23IOucgi0EpO3a/ZKZeZkmsh0g3Q9NnhlfgdjyIEy0CVXMhV
dvp/YcMcQuYbLziSq6Vn1nGrzBjYU1Ntazaav0GU4hynrFjDVETh2kjwLPHzdyX1LWCRqATFe1pa
Lke/lrFoeZnViRbWm1exhcAr/qPUj0WRaGxvKEeBeNOy/YbliO/GcuEYVg84zmcLSk5EjsN1EMXt
EWrEOtHuZFcjw4K1Fx08AH2de2xBOFsCkGpD+ViK0Q/8jzCiv5u8TrsjGMemZCcuMumnoYypWaYo
sXSW4VebytdinQgcN4AY/2SLSZeSVfei2yDOrUYN5VGp1BILDgrNLuD/EtA0gk1WaGS1vzHHqayE
Bf6ajgg9wNipMIaFMPCIhpD1/2QaeqPb8Veoz3NPJLgv2SPAu8zlX71SOW9Yp8mHslOlJaDA3jkA
LYXtoaRyNp4leL8J4YUoZSPNmbh+vPalTYyICzLBM9XUog0RXinShOkKLMNZ3dNCMmHV8nD4KAnb
wy9a69DoceR/wA2aby5xTCCzRMYtCXMQ5QWvkmYMCXSw1Z5AbqCcPT0Lk6Y7pBe8zTv1XXiDKZ1S
IkSlTj3l3HTaOROh3LAerdbD10VoWkkm2oZ/J/PP/B+YAFfjXvBPR4q8rRk87QIIfFQfpq67mSBU
zsQw4fV/mVm/f0mIV6VAeiNeK5GCMyvYRDhboEIQ/a21e5Nv8+SslUTNN4NPgS9lpB5uKEunlv5f
RM9DKmliDlZw65AXUTlqrLWLYASh0qbzlWIfrPHBuXPI7RHsfP8MMQkNH5161i4JGqqeXBo5J7Fg
tTqM+NR8nJDIJsRygqsrlJYRTGjzX/VXUGBusYl+y+9nS/zGd/nvBMG8X/9e/2KjuY/A9TMWJOXf
bWu4XxSC1xb9B+WQ2eTy5XlgSW+D+vjk/UTn552caqrcVSWKz23ozj0/oFcDZKsdUCiocUNBCR2h
qKAHvEGEj8/lAFyZAWflrJMp+BAH7h6grzLtNMZHUehCfBPdh5YrtNrjbsI+bV4HoA8Pn8sirx/F
OJZA3l/2z54IELJeqXVYgBWSklPhjl0voueqbHI0k41+QROi1xS1entBBN5w77duFjawta5alYTo
wcnH3ttKgylTUd3uf+puqJb6fRfpLDLwg+lV404HoqzasVOswyY4q7dcZW6TmN6CTl2CpkTi/A8E
VPrKQ9j0LpBP/2hZ73RwAzdKZAnP5tA8z9T1yaxALXBZf9+Y4G8czr5zWprZ3xhTHWGRo1Tu0Hr6
BqNoChJXBXMiqRublNBv6q7pScld6gUBTQE8CKlfKYQTFQT6VyyQpWKZwqQcw/I4f9X3l3WLsad0
pnB3Nde19xCPReKMR3VnQQTtZmrYMSJs8RNYrar4GdXeTqzpEY1rwqp9fzuYJ2mhUPUAaII7cac1
CVE2KJ3OWEggU6jOeLcSwborxC8zlUpSCgF9oTCpzB9l+WhdmpQ94UFykBD9V3XT0/kTkom5M2eS
f9/XGuLNXohfoXleDM6AZkpJef4OG3wMuJLpzSimgKZqpE+qzSdZDB0eQFR29A+r8BGcOcgdYuUb
gorEpaTsCffyR/EgPX9YS4wWmk/lLMbbm6dBJSrhZXB1OEeQjthgvqsfEu2cxdjXn7bEeHzg79LE
B6AO0A/RKh8Xfbzjx5T8uy3kGKS4fN/XI2tPo8JVYwriConrIvYdMPXroqnUo5RTt77ZoDhp1pwS
+5eM7zTgQg630vavAuNWbuDkisAqzMv5kNfOvT6Xk9D/bKXQcdIhfdCFSJkJYXB/oURQNzf+4u9r
130h3uI6VzRF0FUgTe4eqzPm4Q2fvw4abKvE6rXJZjJTDGCtlzg1dk+uSCt9e/RpkfstKMg2FLre
mZt+ZDf1MSwwjOGeJWfhrZBp8EtG3MTf2eG0MaKpT9cH2nfJ1B7qndNV78Ug6bLXGY7pOgrVHG12
7NzG8vkkB95Ooi+3V4gYNX3Vu9MRp9wF0ohCo+EWcvUju9G9eOp3Q6G4swt0vCNu0wujNYWevAuP
dlZ4ocqvCfcN4vtk0LPHcqg5uyqEugy2WnnNGMSzoTgD/Vitmt8eJeNBkdnw/i5SB2lMytLGGojD
qbFLNtWnWnmZreaeiUE+oqQSQk8wxOs9Kkvu49itF7qg32bobpZgYREfjOMF/pLhZgk5e36gG4FC
XHrue5zMvo1Ynlt/6hfq9cUmcB5be0faY0wCUIlSGf4VkNWJtxQ1YxPxqupNJGkxR0YW7SE3YuOk
y63KcPJLvrz2wf8g0QprE1FZCRaIkkY+nxQ6ep7tFg866yaWj3C0USd/VOgwVo+Gw2XM/EOu69pf
giGeiLFksl3iHJvLcG0ka1knk9nyNP+qBff5S5Qimn/AVylTClAVuQxW8gzyOdQGavY5K7QtFljY
HAK77bsxbLArXtR/SOvAe9PbxvFtLraxDex7jCP8yawN4gyPDT+DpXW3idZXxsE6H2kX+hHTh1MC
KkMigVwl6+alZEWaLFZqtoRUULAHcXTqo4zOVs4NBaBefgNcmIEC4dg0ts31wyqi72JXANVQCS5A
IYh2Vec0A9aeG+HW33VkWftli6pQzr0OCZpvYfVF/n5nTC/tPMjb6QucOhUFFdhrlCexFmpjk8zW
eqZXL7kDlrYRlTypAeHesk+RM8HbcSqf41R+BrpObMQj/xBK84SDSdAmyBJSf7o6BjT6V7T3PROr
jwScK1yBtgR87EpS4fPIzx9S/UU9f0cJcEKmpEwfwJKhZAiiWMvnItvA1yp2cWzoNU3T6Sz9Csau
Q4q7N5JHuITpvcITKQqL65Eok+N78vfqtt+ydhMPLkWhH3NG7iiVtfIihaZS8dyuvDdORvfzozU+
Uj5QYeZJx9s3X3nB61LOipCYDI+o/HdOZUVlbq+wWPUo4R7aQaK4u9w5xvJVds17WDB9GgibxiV9
DdfDq4gc8z93vEmVMeJjoJhSxumDa1BlWQ3wJE58/YZ6CN4TUD12dKx1BOkr/wlnJo/Cwcm3x+jT
KR5JznOrFcqYMpAp5VilQCOh58y+0uZqK1t+EbY71dLQHkWUrNG7JW/CvwQt40/LaUnhXhuhKFxP
UEesEs+7QQtA12zwpn1Cw/EChxFATkV/J5Wf9Bp9Sw4VDOrUrbcEth+AIrxOolbAV/FI4/w6Ccx9
EckynAullCiK0R4q06XeVotSYCAtf1eke++LDr31MAKH0tqBordNJGq08+Q9epuGe74k+bQhbmMb
Zw0eZpFkLtV5eqykfOyRZNBIHjhnqha5uPo03C+SVB2g9sl6szmyUbXuclv499Iqwy50Y88YWdiS
E/2x675ud8liJZsDaJNFw/jkVDh/ylmkzjek8Mw25JcjX2OiRukQY4tUqJaQ6vhrhNt3ion4BT0F
oA80//VWjZo/Cjovp5mbtAI9TimkEw30QZFX3UEDaN/KDlfM2DVQYA6sMDVHKhnK65960f433i89
txQSg5MMLbz+e6ZQ4YvMWmDhyFqJWEthc1DA5zk7kOgDjAVjs8nWhDDgjbp1v87YIjcAR3e9O43T
nYKwMXEATS9ANiXW9g7XzPr1oAzaAwbucVkDOE/+IKKoQIT6+6UNqVcgqUAPr00hVBDJKCBxI8YR
sNXi+dx1eRwTGoRHM7u1rOThys/en0FmUN8DBkJElfQx0VMUDKAhgAdDtrrBE0g9Y7NY7lr455E/
0zs5OR9li7d6nr2SBOYUlJko/py+tNHS2S2Yl6cmIIRLw5x2wtoL8/nwOYGVWS2ECEWH10KgV6wS
JrcNIdRYWe+syvPC8JF9cUDw6VI0D9ygJyiGaDi/axTGpE+LwGXirL2nkX+h+7Df/S66iJdjwAjE
YVXVTov8me9Xszsvi2KkuFfXUx/F7qEw8BcnmLf9PSl2jNWRTy/+3zcGasDr3xUEMPVNZJZLPS6Q
9KnrBfdfCZ34qjaeIEv+7J/yZJLl5RQmz5uwRgivygvl/9V6Z+bEBo1+PG05+kbb5qXgZLjdlMnq
/b9eXPzqnzeCvfFoOWQ8W6LUkAYzrp2eDb/+rlzLv1X6uxNvhk1hQLchn0B76wzEBpMY8eYsKsQW
njrKyPFHZd9q3T5+XPBqD/1UaGvLcEen4q7ug1/STP+RftW5IQXRp86lzOy6WQ3kyCW/F0aP+M10
DnR7o9TqQhnB7xN4FNEE/LDhHbvQawILPe2a9Oijb5KFjhIJImgPCKTNsxBK9Y+MnfmsHftrOyMu
PChh2GI3WEvucRv+/PwQ3X2v3lxinAnRp4BN1YoAVnW6f55RdoWQp+U8hn1gHD+i9qrBz68YIhC3
URQuqDK75NB3h6ze3PitqkCozJ5uB3tgVp0vvbbvERcgwbu2D1ks82XmvHAsDViV33SY/IdfBW+t
kcbc9a+F19FmGU46kIudLXAV1Pxa74/h5UUXRWwkYnfdSLHjDe+LkB4DZcD39gh5B8DJOolJmHLH
yzmhVeUrwEjXpKt+w5hDUgyCYukMM7eFHeFRmisSgd+TgtOlGgJAjRPwSJvAp08fHBfsM4k2bopu
7sfFMonPUWYrlVL+3D4yMftz79iShGsrSkByMty3DHiL/iTg78MoG1EoUAGdKPmv2rwQixW8P0GR
/5+yoFgBs0RLpV5f8uYtcLvzC9BBotxlcvb8R57fOu4wb8KeLzXRB4hzvhjgd13XjoPiDGKZ2p+E
eovklIr8wcxL49j4haEh4Z6l7vtqD22P3NqCNCRWHftd3Vm2xLFr1oHr4PGgospRw+iEK2aAvZlh
M2eGeIvGLkjIfG+taVa+7pslBNiOsJxAwc8aDbdQeTBRJMXflGz+GHNbrfF7tpkrSfqnATpXzDxt
zzKH0rfS7fRotVR3PtEIZDbdySC4mKhsXBuWFnN8Ug4ek7lGkJfDT6lo2pqHChkc1kWPjagBrH86
uaEgwM6jWABGLf75omDsA/4q55ph17oET7XhpC+qB5JRQBeT3xSv64t6aK0AtV+XXitBzLDqK3eT
3l+xNrrNLaZOmqU6uJeTF8HbfMFJY5ph2tJ970DbB2YDY0NpY8WeLOxKgJrMlbSiqcgPCJWL1zAT
FXbGtp9HuswalD/qpXPcWRPJg5NzTdTdSZk7T9P02pzh6wbcEm1vkws4lqnPN9ULmme9bFc5Be7P
vy2aVXZ61M/CfkxptxetTMyKWfkwlb1ejx481f73SU6HBOilLFV4vHZkABK0bxUw0ZRLa79MYCEi
soDvLtS8+uFtu4TTkThdpWcFEwPuaxZf3ICCpLC/Q1+UEstEcUrKcZDkhqrmOogCJCWW81EwE7A0
dORLkP8J2eA/AYPTwKp5djPRMu174OJeCdrgScKHnYc1jvoopq222YQIAUkE0zRGTPBos6YXcJNB
WGYjiJ0A6eGBcKPpkLUViY5ItL5kJiWBJ4um/D+pjtI0zcXmtdAk3xRh7XWQBRDQDVpOtnryt+zj
I4tQy5hxJtIlfBLYS0vihNEJrjalHMSGFV5LZ9wYS/WUEQOO1YU4MQeMWNEg8bBG99G36VJiomBB
nb9F+hq0I/4PlyWYN6qgnSN9HdfTl9AfrSceKS+xxSXbLOhxtXjyDJK3cvz2d26ZZth/tMnFHvu3
h6vaQIEmo8XSFBJNuMgoETAoSSLQjdkGrGTNJZt8J7x4mwZAOQKlD8gPapbEfZ6TwqeRYj+Lcxrl
0p65jALElMCfhmJ7VqOO8gsKOwim1jhVXw0OziXbRbon5h6yTIvaUFPU5/Mm+zkrv/9pZRDfC7Kt
F4nSyGkVxyJGxIsGx9H6F/8nqSbCsP6eLJHViiDUla38LxlABJBe0gy7xgFtxpIOcnsAUYPR4x7T
VlorIOEn1qGzOTFZohmIRpKQDRPaHP9riuNZRCJ6KOffftF47W6LiCY3aP5zBqWdDogcnOJwK2iI
EbnHD83KPNrsTkidJT4y47+R9QdHjrN7+y5GOqpe+/UJNcgHfPPcKm9OE0RjPsFg6cWpUZSzFqPr
sU+8PylL+65hupR1rVxYh6ysATYby1eHXJ34xq06sQ9iikC3E5ljIDiFcjvtQvgTFc29cmIMVavG
l1BEQ2kAUhkfTie5fTK+2c6FkHiRE8//ByL8wu4FHuaniqq7Ckh5wDdnY9NxfbqKsz6ZrKXEJqcD
iTGXr5hCC/3DjgLopoJxKLSrCRpf4KQsauOniwzYijacveWlsvk+UXpr40m5uBQzc/h29mUURn1j
7B9rhEx4UFbGgdZYNqHdPkW6jmf44zkP18ozzhx8MUkuuLp/DyCxDunKu/yJuqZMX3EaEwTdIcKq
mvN3c8F4+FVZdXlNyI7psZGaiHgGJhSiH6V3Q8EKEmle/UDecN9EXSaNVDs+AgiiZacz2VXTE7fE
Hjvt1f/7FY1STPH0jQOt7M03WjOP5gohFVTA8H9VozEhvwbYB9OCXWKsni22knUJ7pnfBCvkvYIS
8mFvaQa7O3kbMq1nVnxYvml5cjfBhZckrgpgM5oByGGfcPUrNlrMaKFHqjyu2vd6JsgjAu0dDhV9
zs6qWlph5gd9pG0B9c+42H8c2lhsBFb+VF/tkVgzl4+PQZikMXnSildVq+JJdy/y2A1dStEXlC11
KB/76F7L5z79os8G43k/r+KRs/2lTQuaqAmwWLNHjyDu6QoqboaGbCv+Z69xV/v/yEHR3Wj5YAW8
vHlGM+3BlPv6UJyqXmj+AIdAHrdcx9wkeGHm8pfEIy2ZTqkGGTdhbofHSjfWZCT7+Bxc8qR12Bdj
fEIaUjOwBKXOan1SCxU9hD5JAGnMIP3azAX1b0F5RFb+gMK00XZxyrAlvr7Pq9SWocGTd0J5K1Yy
qyTYbhVC5wMfTkPVCBLHV7/lDd+2K95b1YXixuvNwQ6rVccIXegMxsgGNO634bSaW3yV5EG/RFeF
PmfCqv8b+f71ZijwEu7H4gdbdn9CxKKiWSJR2n/TfVQc62p3wfRDkgeT4Eu3cRTSK+D7TlKQX8QI
hsSOxFv/4yC2fVDqRxPhCxw992KyPiYtBak+VGIQTcy8TGllKDJwEEY0tnCbIzvUlhk5m2gxLbhE
FtsJvacTi06gaywi+bo8vUWJxj+qq/SZNEKkFIiho9r/O0ZjMhJhM54KkysNXJankWuIGBLsszjM
YceleGw+vMMAcDpKN9gEacPL36h5XmzSGvxRUbfzf8Ue/NKuemg0rwE4r2wAYea9kC5EUgzOILp+
sLkhY1HXPgCprhnTAyhlA0MfYFnxqSa9fkdxtB4q3V4VFyWM40l1W3ZWB9R5XbdY2LcCuVIvdYJZ
YxXmAjlM4kPfKRXXHJChUjN7GgPsYohRiYIWAji22rcSxSCHT91sN8B0jFX2oEPDZ4hIkxAvcsLf
VSanaHph4UCXnANjdRCZCBGjLbViCooMjllFR3xtpDHzSyZ7MUzJOVJyqQGiNIuh1nFSWJvVIlhr
ACaLxD1tIOPyFj25voZNKBS+XT3W9COZpcL24Eu/S7ykOySFF2vP4aEEA7Aj4+EVVGumWBtRdgDK
96LSfDb9gFhR2tvsEMysxqLGtj5b1oS4aIEskvSo2jL2zjHelSk5DaZoy8diOr8fspleU9V7bd/3
ESPfwpkqf3RMyzNXdOVE9UtK5iZyt780V9YtGD+/K41rKfc0ef9tL+Og3QJHoQF6ip6dW4SNXMu9
GrK5oQerdWJo83ha0Jsg8PWy68KGh6/XNXsNKM8WA+5cthNvLGwcu6RgWreSYN3t1Cs9tat+xRkj
E4f9XSHoijCkkC6GyiTsSZ6InRhx/dBP+Ua96OyawrRWvqPbg+8mmhnLIvo2B9goISqIcwHkhkxi
ATBl+YYt4ijTLp7cLi4ysWCgDmDuZEZcyWxBWXwhG46etoxJNTCpfRx0peFzkgyMDHIHAcgslYPM
ZBqWaAelZCUyMb0ybESUF6tTJjPO3rrjW8JH9LXKmPFZ2C1L9W6SCVxFrA2OqVLbdOoyFUkYlaEY
unLff0gVuFKfHTIn8RBiMxOg5nyEF7wthAbKytO9JgFVKlkn8sHOFSg0B53nyyrl2+HL+Srf8wNS
p3DPpa/oY00PaQ5dfkjP44kD0Rya1XcVikzgQcow2xMcpMmTLsDMYbqshGa455jKEKICKov6dKsG
yPExOdqEwonn8d2G5giGC+aTnQDA6OOQXpAUMV+HMLoD7aqusqLZLscjbarGDU3J8uFhxTw12c3B
RXFAkLT9Uhi3Ph44QDCcM45IHZnLz8SmOvOs186ea+uNVyxbgeX0k/aC/MrAyZmPMqotW3gqRRvO
JduyCbt7qJW2RJoEFFiBkQYXYtTvP6Sp+gjGELV4VI+DJv8NzK8F9/UxdmhspGrtTm5P0PSNm7ey
NSilicYVVfpTMZLA/nt/hQdTctFoyPbv0svInEuSRj4VaaazifYNLLYvvD+lXVCHBR3dz95p9l5v
h4Oqi5aSu7UTUrCyowKlv6mS2FIAKy1DAUU2QdJEl2kRb95JfSNKg0iFecfvBd1EGM8qBRiLdQAT
hC25q7Ynz0LZ6wue/JMtWdhMZItsGh1vA7p8QS2/uQZ7fcJCBmSpo1c4tCP6/dD1sPb+MqevZOaB
AdbM5NSnEVphPGj73/Gg56rBZ+RgATcnNn9j762ZCTTy8tVhM/6BfZTR3sijqSmMN0uCzMam7CE9
t8vX/1eCKKFnqaewAsAaHRGMkDn5masKJ/tUCp3hVeOjKwiPg0H1IvvpJf9i4IAaT2ve9VZ98y9t
2gRNAtO49oe2KxDmzVAjeBK71ndSIIulcUnopuCRZRdOkNFa4HY+N0iZjntTmhDH/bM7mla90azy
HRJClmQ0hT5szv4b2LDHI/Qp9FltjnlGg9ywLxTgH3GBSaRR8uzMzOFA/+6UDqsfPqaLqPkchguP
IdDurXq+3Zxr71y3RF2xDrlJKOZyoTOxaprIy6m/NkMiKTYtfUFRyhVYaGejUgW0YjmzC0K45Tff
8PVVd0/X0HktHqDioZnvU3LRuf1PGEzuuLO3unjkFaRvvFu1JYgxluSygdEmArhYKrVM4GSBaHIx
ieXds6QAMVnjyA2YZEHcLd3hIePZ0uGBKTemsORO5Ciq9VUgGT1XmVcJZGWtB9isVh6h91Tf5Cbh
vmZvDy6oYia4aCIh0ehGPxYPyG7JP+xJJX08otytBNbjxGKgQ6jbZ7ODZhhlKBzqhIdtQSvreyaq
XqkE5tV+Y89IC1Hub6atUxtIcRZ30VGalHSryztruF9mdn3gakAKubF0C/x9yrOrHbAfyUlCRP8q
UabPipVN1qp6/4kdUPlFd0NhA6HmECPBZVjOhpbIIXqGJeUjxEWRG3FX2+1BcK1dkiykDgiZn4Ja
BODYmd3UGibD9xV9vkeIqZK4ItA64gbB+6DhwMdPQOZcaUNmPjJMLxpIUIHGDI7ch41BEHAM4Fqh
TPSUdOlzOL5CFy2j6O5YDtu1UCsSRv+X5Jw7Yer7v9hPW4ZoR2p//hal9NHFOCNSd7D/tPQc3bsQ
cxzoO2F3nMjRuBee9lM+8/jYvSZRcBstq872Pp4q4Ypn61GFp/88jktX344fLscdd5tIZZ4lF+Mz
PuQqePmTpvHFNZDbjB89S/3VCgFAGPBxyufd4SeDjwraIGAk0lMq9QdkNxu1d6LbWsySgQbE8+ga
b8N4xTfnvXgud/8JJbchOYcQPo3eGFPN7g0TyaXCsDYB8TOtq/2Iuxorh+/edzisI+/7UpZk2Sdw
IRXjOLpgO0meKBazgRK4vdUR4VzOv772YgVq0PnBS4YyjDncjyqsHv99QTsJeKa7BZFKv5xf0hea
LbBeMkG5dsUrPICvBsoQbOGZMNz4uIt1D2NaZ2JkJIK+It+fpkRtcGr0ySxJTms/TW4i0QIWgDAq
O2+cwanypDdmSImeKvyxOmFCL9q8GUSFtfZ7yxOT5b6fmsLMZNSlfmZeh59qwJxlogpNh7Z0VXBp
HgQrqOx/kcURvd+UNl/xBbcsYoFI9adren/Y2F+AUQwOrkoiEcmRjvH+EgmAlK4s5BFXtxQv6p/X
yr8xuvkn2YKEynUmvwpipz/atdVL+GfOnPZa8+TixVh0S4CmUsZhQ6ZvPrNpXZdgG2mWK5oOmGSt
BaVz7DLKcTwAkXQfAjhOsid7+sOy5IjNTUGD/LHH8t8VD7MMXysbjp6Fy9WesNJUXzQ8yU1EyAAZ
8Oy2b/zFnGW3n0/D/LMlTMLY5FqQb3QyDJmrPtf7K1rM7j2C00dp+Cz5+Oj+jnmHyuep4jdoEPRZ
3S7GFK6xbPu77nOEW3XVzc7HLdEd90mGt9NHkUqd2K2swwRSP/Ahe4AKAz+KNGC+1etP59cUDGSt
XNrAlBD11d5aGBN2FaMZrf7JmJJ2OaQCW44NQ/zGDEY7cYIxa1WVS+ym5isbxenv7C7Pjxt3fvfO
IzImLWuRk07Eoip8VustBkW2Uat7alkTLGV+/wIQOA1LxcRbET5ihq6Fe6Duozanw/SMlYTvbEMe
z+cIqDRxfVNrYi5YYkye0r+qERb4QM0S7OXkc5+yf7Gc3cOTcavdXlBBu3R1M7tUqDYtVeArEHZQ
eQe+mK8F0hm8x3djIC2451eIWB7o5zAO26IdbPpro242U+KXcmmSqzYX+EQXYc33/iaxbm+jSQwJ
GHDocxQCXAtwyM1zzprgyxwL56WWc3g3GN91cRjMFVJESaG2GWtxVSFCUEdkGX6rAkPP9gBfAfoj
IZxhUPDPfnAREzrxGxSq/oFBXfVQ0DiMZw4JmthlGKeTdbSsqKNXdllrMPAcs4WmBg7ibl9KxKe8
QKGxZAmoOshd7OutR5ItisUVp/Y0KjkBWLeQRcxDPLSejNtKIXJPindBnpB+yV1lHVe5sBz0wDTW
kBQmW2BlXLYHWnkkwI2l+t7WyNTjlvJPRsl1sDZHfHWo3vDO+lABQuZolLl50kzKv694jLXaRC5H
BNAO52RsqZsSpFUn7nJd+685xjhhMMqPoLr0FzGuV7VlxsqR2jKRkkYKKIUh/lWeYiW+84p6Q45f
VYUWrRr489A9X66ttEoNnBEnbNsxwXQrFEb/Havx87ZEMfbkbrp8LvVeCgLO0asPECAX3ksJTa32
tEchNEHdgwOcPmldNvQCdQRLl6vpNn/yc/vaJfiSkekikIKQlhMiG8pfH2wBH8w4lLNEDo9kzP7d
2PkkxxetS2TU77PGaBEHg72d1ltNV+oU8zOXo4mNPCa79uNQrTHFTtihvTUbKLQlWqhOLVWt+cJi
0mL5CaxEiJeffhHQLuACrm64vIRtK1fQOZfTM7fUZGO4PQAritbvwsl+gIzaMSQ5ReSC5HGK28OY
RRgC2Caju0VUea/od/y4jbMnV2/rzppnI8AdqY4ScTnMCzGtXkQuMPW0HwGrWeDfoRSPBy32U3AC
LefgUMEtZ+K/7bSJsovFOJJcVrWJ/dbsl4QmEvuEkid21sxARkVedlVgaycYWQwlU9YS4JS0oiGC
JdgqdfSbBTxc6X9eJu+2WWSJNqNYC6UD7tPbnHapc3j4Sb9Xj9XcsAo3A0R4wDbkVLfc3XztJtwe
COC+mOoLyaO+dgzm/1xgDsm0g9azaiCrDxjJQNDQLuI6U/eY29LVt85myhvsd9bn2DQjfJTy7f6x
/2Wr+q5WcqrrEfwbbod2Y/ShyeifPlBMoYY0IOk3l+ln80YEkk3nEiRPxP1TCwpN07cU8twcSIEB
cIYOrljhQBQphxB0G7nalzf/vy4h5xUjvDpepCNsfrMaDMJWCr+ESZampJq0bcBIbQXVM8FVXjjE
RinTKerbksXE9xGljpKl5fLHUjC25RNnp28uGFYatrANdG0lxnsie88YtUA+j3a4a2N/GiwIUw6M
5IQeW2UMFZ0VkqpBG9GRtMkciQhtpSOHZNg+R58CXx2AopdiJmDyRXGDcD0kOZJQpnjcKyiwYpsn
F4h++4yPKoRo3UbQacvlU8ZLChhIl98IpWSGWN2IhmxyIgnLduxCcKNNVWLTQznOADxRUx7rVOvm
UhPb730FSGwAHYQy07I7iYSMZWI/a2tUChFnpm2YL5cw88NU0Kwq1w1EtNeJQqtHetlWcVp+vmmT
ElzIJHKjNSJeVwrxsFf8sPZlPli7ZFHVz8wlammbxneZfO8Apzn1HLAJutf5djrSZYSXElRtqmId
pWXHFlFNnM4UcvO9wTSk8AwwaIOvnHCWoIxJKNF8eTBMiGTm6N6QCktyY1WiDYr1D4P/vJr6gLFz
U76ITysnV6DGHyJ7/vBFwsUXZWX3ID0nhVb0DfCg32Ws++MAIQGrPUVfhenfJHbpYNAHACHujfJF
lSicr3tB1+Q17jbz3Mc8YnQv5qv30P1qLU19APfUAcDmpnqqFMyBr5YgMf4qcsS4jMfD5MQpS9IR
LgBl4WUz34nJc2OP6vzvVwotpiGxKHNIs9yrV5bE/lUqCe6oLvgODltA5oRhHXfbA2pjAFVXlVCY
vtw4msZRJ6Wlv4noyynW3i6v0doB8RlwNOtMnG0DyfpQVr0ek6d34+lRPsomo5awzeH8bkIViHIo
CYFsEAYmfogUgjudV11xoefsd34AmLLmWx40g1IjR+ZBmG2fbR9x+hC0S0hdY2jVM7VrV2am6hy+
gkcg6rf0o4hIFjmnTBrTRvxVGhIwEqhu+vMmue/H4F1MtaQJalB9gmVdRE4YizxLLB65YTF2YUZq
oS5eGxsDAIEUiGXWZalK+ZCLvt0851li4VO3Le/e/28I0AQx8znu9vuMt3QCw38wfsncj58nlaMY
/Ltzu2v4c4UXoLbTU9/St90GviNA+JSPK/VDNewVfzkkoEkUp2eNcs67CBm2Crs2hWDBNz0x0j6M
7aeUgH3RcigIZB0LFE7tvwouXJiMhzSoMpZObtwJppgzZVAI7C0dlNRl9xhCdRvp76rIKNZnQJpD
twTaFaBLjuhfBe5A0aqtysC0PoXuqhx7/w0cpbJkDGlEN/GjdGwoKO9ClI37fUK4dWNfNz3eq4Lx
2wyrykIWlzbwm353INfTlOM2xXT8YhwD5tEQEbJabkRp4+vhGuJUFsij7vul1oj0gLOsFkuLnIvj
soBZ+UsUlBLSahW+npeOmcjwOSziG7OOkCITt5oUtmM+LaBqNts/9+fHXEvdqHXaqTTCkYp7jali
axlS+ColfjvJUL1TO6nwVSOWvohwSgkTNl48LJI4xjc9q0kcxIwKe8NKPrM0TArWb7hGYGl5/yXe
kg/38/jDEAroI5aCaJAqJmqgGrXnFQcVmcIsO9jr3H6EzKN+IIQmA1z1UBFH9Ta0ttRqcsvzn6TR
pWFdyniO+MOyXXSvKPBiv4No8mGQ2Uv6ooqRUTZBKbOum7z+t0HFjIEnDRB5CVj68f8vmabtiDuK
AcHExHg69sFx1qtPjD3NylGTeNQtaGQXRNXa3nWbA1Fix1YfvhW7mrDIvLXUwFghkr0ZtUDdmLks
9NKffvGnKdRRKJgfp1h9ZzJTGY4jFmSeB26KZJI+6Naf7poGH3yJnBINCHSTajwQE0PB5Ovn7iVd
zhgorAd2tAmGgop3sSwCkABbkrKlTkw/ypja26ZAFil8jNTbQS4kkOnPTeKW7BBM+9uOMxwA3S3Y
MdSVF3Q290yVUF8h0wxFyf8bAqNzoICDqxJcuXkQ82TCykc+P2HE1xcCN7ndwOOXQafegKidn2j7
yES/wiWbWwwp8w+DC1D1p1s/xNowSoIcfCMSBPGXVhC67yKohnX9hXkZ7XzqfvULhSaWa2genR0Y
onuy3siOdfUZqjPhKPSJ+W4Xf2Cc1imP9fas39QZnatuhOKkZn6YljeqcvE0Op6yESOIfKBDpngn
uhYEJoE2NFLYlT8jHLMjFTyFRGaHV06LAP3SYRxgtXWE2pJUJ4Zk4iIkMo9vJgbzoX4jYX1DuIuQ
ifmNPzv9Y3hhxd+gAP4t/5ya8jEAU0fZb7pZCnz9j+hwQfy0grF4uBwM3m1TN0JIgmUveTd3Nq3b
Nd8Xy5I7OqKUSVI+ivqUhEbCXUjcrAjUyKIGMVJS6aYaCMgKhDDbXLIC4j6DYF/d19YVp9CaxY3U
p/gnrwKhDZBkcVNts9THhUflZI1O6B4/eFvcc5UNutiJLtOSk+emGslhwL1VGd2Wlw3IKKE0sC19
NmKesd8RHCAaLRzMykn4XyIrF64rSuIzvBmmj+U2QV+992Jxj7iffaov3ZilCTGvls8RhC8ePoMA
jIRiv5hCO44Cw41GgtGKiktd9j76T417Oh7OMHNQz9cWuXj4nYk6/XXrH1WLUENWiV1WvnQSHhvi
QWqsWFodoeac21yqLciZWrlRHh624JQkXWbalTWOGBj4pjvJhUJOOX/dx9xf0OiS8Dn8QdBorTHr
0321vjoCixDEg0iqNyDnNY2/5hwxq4mYAZX2cHMYwijWlewErZNZbB54er8lPYCUd+TAfympBvez
0eWeMQeHAg59Y906Pfa+qeHstZ3+xBogkI+Ylj4IDIgvr5MmZEtzzu5NGlUULleiclUxDun/V3bO
Ml2kYgv4a8wkOh1U29Qo97jhh9Klk7yN/mncnijA6UrrQZaSynrAMCiRnJ6Xq0kH8d4ilmvnrSCA
4J4oJDCzQQGyWM3uSi9O81ua1Ww8oGn7QGglbz1OBwp4IIVvKM8klYsxBt3LJhdOISLcECK+Fops
PA+CsmtqyaB6vCmXEjvpqpv5enIVjt8652PZkj1FpTdnWYON+s9p5bIFwinbJxOT1nIfT4sAOMsU
MUWxjr/Dq76yY1/TP8Ov3NDHYhAgAECuLx1Pbf10Pie/yoOWnbSSz6C0GMY/fM2WyeQoJmD1Kspb
TG/z1+ty3cuw8O5CVzY+uqO4yAW+x7eaPsnGuPXm/IP2Oi4uZnnRDVLsZOEu3tsDznMcagwUPcvW
PJUBISR26ptbwQnYAWGHTtVRBwMVhjjASzkzmpthbVUcHT+FCnYZPjKstP8VUC6Mja3KailfpQzO
NueEUoqzA605YnOVaCQLfwVIKm+502uYAWNIcpLj0wMbW8+3blRDecKkX/geUpMr60sz2Pthw6Rh
A3OnQMlyeshWq/2AnGxCQW+8GGQx7pld+4mTMjSGi0PkS9EVsymtoWjJ8OF1M44xhbH8L47tGlA/
14zzSlbNAew6t4k0J1HBHK4xPw9lzld7sxV0EDJ4n8/XFbsMSjjTbKFGu15qhyofim8dk489tLTl
hzL+XUhVt5Ljj60OSmRG8aewd4eOhQhC48mraEik2XPHXts6h6NxrEDE4AqrWel/2ING9N2FhT9R
OHv0nxKgFgLSwX5QTOJiQFWLijZI0w7N8n35VZZVinLllqblqHJx0DKr23uGnb2DS7jowufEOokw
+gXcPKEA3WNKRv1kTFdFvdV2H4U5KB1hyEOww8holr3RnhcqxDOa9ESjwDvEASb7HacWiebvNrgr
yYC6wDM+Tb2O5G/N++vU5dr+kVVZPdfdShZN8/eXmv0QSWp5+soA2zWMWDcvn8M3H/K4enJWfZG2
9iOGNuh83nTifajLKJQOw/pGLVpKxNZM2EIBxOlMZy1IGeY4faKgaem6X7Zl/tfA34vSGabX7hE+
dzK7E6KxJwuZcPCkgFB6lbvaZdQ0v+YbTR1r5HwHiRAlBAh0G33VCVMjhy7AmdyXqY2c5Gx1lAQm
yFBVCn9sc9TMmJ13vJM0zfZVLtJWTtcVluDRpAC6As/si4siChPA9JJ49BTPShlliEnGAe5S/JIx
vF5vnRdY83oh1GGJaVNjhogdRyLvfl468V/d5z4mxZWt9F/c31MeD+13sKuiPgsT7cVEnirAXXl0
WtjiwATpS2CNneCgHb+cLG6doW7sLcD1xk28hhJIiYO1h+N5n4/ckOkx08c47zj49I4RFgnMGt9q
+pMIckh9bh6Mx4t1DlYhlwI5NCivKsezZA0btk3F4O7D7QS/d+4jH2nqtmO7kXB68Kj9KaEodFaT
ARY9p/QtNFUhCloImGI4a2Bdx8IKCdr/dVDsejWXYGi9o92p8pk7y/rf3DAqw2VLOASEIo3hTvQF
WnnW0YRawOrA44h+6DXOzOPLiea0DppzdVGptGIoCcIpbqXnZ7+wOwKVvqGYdHOEnGZ3/PldnyDy
WaDcCPg/t+TccP8Q6KuxEAgDRcOOXVv8iTlkGEfQAqI0Z/9/UcAvhzlqqP/4FI0GlsGKv5Bywwfa
Ki6AT9AsJfWKtOaB8Fq+3mbyYoc5+rbScaPIkEQRc+lmhsvRY7H0qfGUMI9CD68tSkRSu6B98e2a
qsshrmjZ0LCxOhncYF/TxJDLKLw5H6iz772hLWGuQuxDrDFYfjPThuJprHwChhYQT3HDechsFlEj
meUM/liAwDaFbohq48BU3auA1pWYIZmwf3tT+3VLmyzrjIpOYburtAoBIuopOxbv3u7f+Z8JjNfd
8rDygk/iCY0ayktVsryjsOES1G5v/ikAIkqGO4TZdUEwBTWXBE+N1xYKQbWic7i1uj8rQndES5Zr
/kL9WUuWrmiyVB/FHw+huvFtgRaY9alBZMLxtwo+F5354utpeh6/IP7B63/x5Zx9xa+avBOtwn6V
bgXaDPcn7KXKVFJYtnjh3GgKRdAzuYv7y/x2YjijpJ9m11hzqrOdun5B9CtoOKMeZQlJaucmJU/E
nQ2A/h4hjy7OrEg/3iuQL8Xdzth9eLsWQBizj93dbF7+WU7BdLMc7L0NVxYSoyfYiFA+p0hWEnx8
Kd8pZ0TbQQlizoJwkEYqoFrM+WzOuE3x4sdzcAQMOk73cZaofDpviO5LWlOsPxaL2UQuXrZ83FqP
hVJpumSFupYgIMD4ispSAR7RGaHO0xuSiao29trsI1y/GdKqrMmUnHKlk9fwJucYfKEdmdIFixi5
tdptdLS+MpUia7b0yHSrKZmMtssWxNzKcfS0BBF1Do4aVOQqWL5qmaOD+/o7l4jppFlQcWwSIiof
Sq81UUshcgb91mk0haNQ+PK8f+St8yoIxutUdaXTGqhKJrHda9qfn+WCIRYI43URAIjShIkGwe8N
y5AbAI6hCXYJXVLi0jViva1INk1RD+DYatxr5jQNKk1T+HybLVQbFAMNEs6l+N43NyiH8Hzma31y
IqIbc/0k4Bd0vpSQc9AaTGV37fhe4KuIwcj69vnuXnjduk1roS+EAxJcovOl9S/tmBhr9bdhiK0t
RODP0cGVbR+03gLPmHv0HpCSvedrQ4G2NUshsvNqKo7g3Wbul6w/c8UEe8WMakPyNixLVqgEWoV7
m5Lmm3HEcjGVRFExLd/3O9ML75uajQBbIh1Jl0Id0EsMTgOCx1WfjvRZ7NcZUjKuzG2xhJOOWKjc
mLcOmNIjB9Qr+X3Z6Bg18GOX8WcSZNl3RYrwTTJ8jZpc1sEmoLp+YRCpQzCgy6N9WDWiThfWQ6EA
n9oIYUdJDs9Xn9UZOPICk/ynnfkoKKhQwzQ3jGPaCwez8SOJi+CNJrFKbj33nw20GmT6b/LdFwss
BGuC3NYH/Ryj+eiS4FiFOHc5tDjVXmBr5zV8cqZWvoY+0dsS52+0MStwrCi5sPl5i8MjoHDwBE+Q
Cg2Zh03DdfcBPfIAvHN5nxf/gEONITw7liWYRXJ5j0fo1NEiSpKD98VVB9pLTi8eQAd/GQUI/WmI
3GZ6NhjGJqtgygsSg8luLsgCAPJhAsDR7NqKKbfyEqGtDkKXvB7WEM5YbJAySAkCqbxB2JgjSQeg
Dr6PRdk3wbRNLQeWs9K+OHdnEZGu/61G9p+O4NBVWs9p7fkXgjiZwYh65IyJX7YJIAu4ieLSiLBx
HCjGVNTJfrEEDcapOw+rXPrTIqnTA3BYKKh4SEkSLoa8hASsW3Obwd8tgW5HlZzUrJ00T6vPZuhZ
eAuqf/ZxsoYIiLD8yLne0+5Z6hP8BguTN5PR8cxQsdsv/P9cuOSUb20YCZU6SCuik88vcegjIl7B
QMxhcsPJnd+bk4mprnP/X9oKVesase36wuAzytmQ/YSGWeSvPuozWLp9UCAir0uDo+omQYfT3Ct2
+jFIxNJuoGyaENtC1045o6Kfj+qVazkhmh1WS2TdDHWQC1M7oQK24CPPQOlsTtWzWUDzt7Knac8X
x6KNbW3alvjhZuBhGvmoF0x9TqaxECu2SXIOgppREbqjQGZ6d6YXJIo4ZpfkWNLCb9kTUiSIJOlO
A6h50Ay2vk2CekEr4XUcSFROGNeBwBj7wf5EbZoY8WAI4f6BULnltxAlVwhw9HXXICT2jJEgg8CS
5tC/83FpXnqvX49xst0RKnxT3qOIFx2ANFl9HdPzgcFv1M5K9awjH7GOE7r8usls0TWEgGNKmKYg
p3vmCoFnCEDc2AwIDXA7eOhUheP1HAH9XqR1MKQNMOyOalHDBd0GGsNet/PVgO6hfduLZP60NnVz
mU+kvhyQHrHfoMfw+OB7EApBDcxv+T7lZrPr7Y9TqHxaUXtjmhPnuX+alNQiz1YpgzM6E/Ri1Xcc
JyJucpU2X0eVhz3dnNMt6kaKekKIdEqDsGxuB5dApyT9XQyunf8jNUDgowyw0U6Z+lsABKxrUPk0
ajQL6+fJAhlyPgzrAe5qQmjylLyXhO/smNmKhlYXZHcYhhhCFWGMPD44ttOiXujT83JnUK4TeAIU
aXaeanpjkkR3P15Z1MW9I9ufoGo8Yqbv32oBzQoxAeE/DQ2NRoidB5qZITGijznZMO/0OZw71QGL
PQeg7jfbfkIjxaKy6EdxeIXXo7zNxwKCZnzOkpTY4p3BPknrg3NLFkmIUAulNdqNZ4p2sEzTaCt+
ZHdg6wZo9jiQkYeHEHmoG26AR5Z5cIjJR0EYkLWGvbFivrNWGhT7W1NCT+CyAraogpd2hPNTrHe9
/XCW/RVZDd4zdqaY3H5OThMz/jJAtHwMipgxf52n0npAHgmax6MMExYIt7qnG+smjiRbWdgsulSz
EZgnuXZ9CX6qtK9TPO7Ub77vQ5CIpC0fPVPZlaOG6ajIsNv6QiQV1nAoULkDG75bYB7D5DzJCjdO
mQapsoUPUdLzofYzoJ16X1ujr01dp9Sd04mAGgqemnEWpPi0GOq5X8OWmSJ3CJeM0WLu0cHzYTvc
nWCThRgw4AqUS1jbFq5ee+c6we8UA9rcVXlxB+/1gVcSzm0AeuyqGhF2IkZlEIGvxxWnH31+4SqG
D+XhTOKH327HiytxQOmymtB4ZEPkY+aBld9snckv7Y4nKKcm2WEQ7AMzBU3Ae8r/aU8UWYQ6efaE
pPm9eJejI6hCWxQ/SGThVi95MVp6QIjzcAQLjVYDwgkloxV1yIvTf5fxnDdk4/00PRaTEf68g5Ob
yqeni6JQjewVUFS4H80Ts804s2bmxJTwq8sC1UDPpUWsNXXiDdHBa1k4bUPUopZqrKk2dN63X8Qy
WGnGQ9Is+USKWRLSwI6csjjbNrPMKRZ/uCnhesjEyuxjblaS/eTpdpXORoKOvYTOpylgT1VUa3Q/
nPNnqyM75wKQWHDxjb2pV5V8aA7pyrgVdjsEOYy0d9xAnBrRTftr5GEkyxIUsPRAGslCTNdSJk+H
AW1C+YWa+vq8qGPtzI6YD82Lt3emq4AARkn9rStDm81nlZcLp0JJr7+jflnAscbFI2NISX8aH/QR
iZnvn2dFa9c6ItkB6Da2TpvQmjI2POPTywMnlQh7m7WCWAiWe9L9uWHr7IE9Uv67TNM9N/vR9dI4
3GywIqdWo1dTkvaaUvlK/4OBMimaihAmGY0pn+o642u3d44A+3MGqGbs8qmhUGuaI0XkwanWSR+L
+afqGQoimml+KT8YBVkeu2h8BepHgCKKxmOBOZNU6vSccUx5eEwLtt3kVEChv1Y/AB2bYnrgAud0
33re+APjIUBIq+PBdq79ANA52xgjW6VtrvUOT3vshKnd6Hz7bj35JGPj2FNWc4aP0lD+9CEDRpFc
d1B5Trf7EViobWYyXbBjx7nnDhoywbKvt4LAUHq4FV1PC+zxUe0/FEUXOxBeLHQYPNgxWYY5Qnob
MIm4zU2vPk9A6ws5vOo3eIrpXiH3/VeZNyuU/O7ObOI0I0DM1hkMBmdTDpgAmTl+QDCxUqDEYAah
mwRMDltYBGgeQj67twqNibmdqA2UOrnlIdnULu6tWsnhIwNwK/vOYpkGFs6VbIX6eaqfp8aBv4nJ
yJjFnGVvIMH3mFLApbVAyEUaSVZADTySpuR/aNuRJLSsyReaFr5IQ2i2HG9Rxh96X1VzwHoSFvGi
IIV86A8q7/v/Y/dDrjW4M1GU1qRLdyMBOsdZf27q/oq2t4gLSR10WuVwLibhW9jSYZSVWPC/t+x/
beUGiSHYvqMwF/vcdril9+HRUaXD8KBtNyk0zJix15IAo6NcHFCFC2tOR3WeqguMVrjilh2CMzHE
WtVr6OJQEtG6/BTHlzrnmC8K4kk+1dGTTjiMYdaSYA2muun7KXCXYeQdgFfPgRWTlv2vhB8leLMN
7P0EZkjmuro5O337YbvLFoHYGx0ohQJ0Vlqxvhg9zvA6885kRKYnKapSr4Hr8QM7MF+n8UaPTq0L
rZ5DSnLT9pEiKAsrF4H19hqJI6DHIr6e1CS8ZhQYJ8x4GQEZbtyCld0+EvNACblOpExVNDUrKcq7
OJ++g4HyFWzRSQNLsBxFoHQhJvP5lfnwyzNNrSo37Qlcwj1kIFSdnXroPN2Cmwc+orfg1SlRgYeB
JGpihycDCln+4scjLDZmIyz0/HBcIWIID5HeLpcYOd3rgd39e1COtD4wPLco0UrAiJoT+W9Sn8gN
cVfqFD1FKSzzY8TrzCac06pWTL4SeYbgchdWgAmG8HciyT1nGmkTk9xpjPMZ1C/8vk9hLfnE51a+
h2Z/Mi+pH0QUhWiidMN0ahWHTg9bUG6OxZmNQG5OUMe2JIyeyVKyuSJZNTrjDt/MMRG0ca1M0Gio
+QlaP9pw8PBtKKnRsvr2e24IsChVANrUUs8TGbhPJCFJpzt3GDChtkvYRUhxMMmkBngEUJQ6bVae
4uqdrglZy1E4YyMyTy/+p7DL3LjWwvDGvhqGUDAT6ftw+E8GINeIG/Mrm4I26+2vP8F0ZX0PkV0G
f/PdCnHV9Th9AVHS1Ju9Bhl4wYQnVQb+Cky01lFVTIprg1cdmn43sSDboHKTXRfaun6Bx2gVxYow
8bNcKER033cg3P/TDRLnH+adPDF9Rvb2SgsokHQLefuzSG9dZiJ7KOCNqHyK0m7KF1xRqDUE5HOx
zhMejJt8bJWoYS1rEmYk7LDOcfwZaagxt5io2GF/B4Io/ab8kkwXnLZ0fJ31W9tgn51k8qs3xS05
VJxDJckkJNR8f7rpS04vM1yuANeeeSf77iEnhlAps2x10hVydHZPBr+G4fRaNG/gix5D1P+uZiVI
l06qhm4fwqUGDN30W+yvV6sGqFWEOmKNOl15mjKtMfTmFTwnkcWUMrl3lrpxzaky8T7dnWLFuVKL
p2zti54D8Fyw4TCt4wsk2Y8feM7w9aMl3Ryb9sUcm1jHdbSGTazgQ/7lsgPo1BWf88iBSX9PIG4P
MpfEc/c2uIpT9NnhnsY0/l4vJDq4qO4yhpbB93VDVbubfP8KapfX7sGBfQ0yLxFTY5rkK0UerQXB
JBDpjkntVVu6qMSMU69ugnl45YFn9KeQxNNnMboH6JQNVRqgp4kVosP3rdGd/ZLPF8K0g8j/CqgY
aTHnO/UYAnbz+KRZ63V2+oagUtbPbKv58Qsm576BmzJcljT5hvHJBmLWMtAE+IBA9NifGvP+RP7K
CXVYIaxSLuNGKUv3KnLuWXT8pAxThdMcavKkTYcc9Jw6pktvrfbRF/umF9+zKE8JvvPYRQqZlbOM
yJsKMFtqaeTPkIZvM5cVkfPSvMQ7hWx0I2GN/dQGkxgt9cvx0Fag8jAsuwAXkf8vsrwv7dd611MF
uSIja1gEGpKciGKy8JvbVYusXncMuuU8SjapDCdmrFeDnYufJ13+wyWqghIHC8U2qHYIzES9hKjD
ljjhM/a/xRqtVRX11jlBBjmzcKOF86xnp/4RB9u8UPzaosuMcOJHJCAqIRv8fWRaMpk7cqIVBLj6
qJgWEXhITHEIWjP+8Pn0GwLQNOZBq3OngAvSLhpoV8pgHh9Azdssa5tJJ23Vca670BBRHwk9sXCZ
byitYpYhEfTcqHFvsb2+kH89PAkTYwaNxbCh558bMVpwezTMDxvP4iak9bhWWN74d7zPIRUARZzF
iD+t5vOObo9EAkHPCYW5AXub6X9awLengHSqrKU8LTa1dRzCvuIzNDBqAlOg6TU9SbWLUNB2Qz2L
sg260PYE+EAJacuiYwLTZmEPuKrWxIlepy0BUZZTLtTOiU1ZnKovJeEnl1ToGO+qDJb4LkEvnYya
Jy+m3lWYNvMPwJKxlqKG+F7mp3+BoSEWsI79wE+M7Eho6BbrDQlFaRuau2tlFJ7w9uJiQKDaGH+r
NCZLHUlOiCC6xbqSrNdeUbaLp3SK2M5skkTR8agEUJrJZL85xNpvbIN8tzau0VCOStldYwY0w7Zx
MgY00gLTCxvCZ1uIT8+1t6pMduG5DHYodz7fnfyWXuiUwcK3tJRc2Ub1hQ6UbgwPlmJO86CX7Vmr
I73PmddYS+gqkorx6aTkC815BKoECxy0oZIOaRdETu14g7IrLTEueCpKrbzl3/nORYlX7HjdVjWK
W9EI5FR/SSLbQDrk0EHuBP5isCD/pNCDk/bptANzMUdqsaFVSglY8Rc/Kv2cVM0OvJxdg4f2F52Z
bHGSfYgIVD8nvidClY7uCNoL5FTThIfzRRASxgGCMd+tb/3Kqjx23gBJtJKPZ5qH8bAxbtkZ+PyT
oPAoYiYYpOJr6cUu58UtUYf5Y8W18sIVprMIfiW3WsvaFmVZK8CO70VjUL+IWFpTznc2TkhJ4AZp
15KZnHWtBnR1dqZOnSr9yB4T6JKVShUlnREF0KTBvHdaAQViRmlo5SMYBxOmTjh3Pcf0/QJ93zay
EyyLgQFaw9CMObx985SNP+JKNAZVOP4UMU+N2CHn7zoZAs3ZyZY8WomIbnYAI5tECmdxHxEopv89
Cn0YTWa45qV8dId0KhVGDMoHwFlguYNxbNPB4g1Tj8fYekynOGdwNlDC+cLiAlgZSqmwN8hN4Els
/4yY1j40XqwTiLXKRWAlxCF/my5uZm2s01ymSUXEIZBuHxUDC6xqzRjGCyvnsnJ85NVarqWiF95D
TXkDtxWjCyiKXJOQLDK/mkPsWnZJ6eMFkfNLSopdKJA9TJtvkbCekcZtGDqyMAiNua8D/9zEALf2
UJ6eTzuA0HK6jfKqK/zxCuFDkMxXgedgtrOTdiINpbXbDeIExd/9/v5OV0yAYRmLwYYVY13CfY6t
OuQC/ivjUoK6qfoB8k2OLf8nom77mpgZBjFb4Hjrzyis5gflueGDAUETuI644rqdhP51qy7TPvKH
llhLUwsLuiDXjwzQcCwnW9X2qSclxeOVleYOxNshrUHcQ08EiyO1jH0EjryZEJ5hG0EMIyf0fcXZ
qK4HsgOJSSYNUwSxxhqx91ltU518RxD51buTZgH1ORVUbsYr7DV64Br7RgXFDWDcdl2qcsT+wUaF
KCrqMMaGol0OgrT402i6yQtkT96EqPniKDmNpzhRLjK0HlRxL2ah7r/qoHQj/587BOa5TBfg18Mj
jbZ5FNnyZAhV7aK7qYHkOHZvH2HBzB0SHhRM8Z6QtZb8dXXsxFND74uCenwa4LYpktVpwcDjsU32
H03P7TdQVHlnkqfHsriLaJMIw73YRVjXYNcdSWUAq5tLLlIWIMvAD3eX5Z5WJ7rcwuS//QaFUQi+
Rn6WeDOrYgNNrrTdQBCKqzzU6TjKZa9FNy9PVzcCF21Zdl+XceIBPrycjACb9t8OOAYPr+5CcjJ2
zeWGylVbp0xP+53BYE6XOt5j9o+phKdaEX4llAQ3JkxIJxwuHOBGlTqQkNGrykqlanBSUT3ukR67
6cueawldYOHde4cYPyu2+YFokj1rMLj4k6We8CkjqzuYG+TqMR2q71l0KsRcqc4XhsSTRjvfX7ax
3U0vuLbMc5c+yIgrF79PoUi+WxrG0WbOKvle9yBZR7UKKk8ewpSDQHqVfrDv5tQoFM0Us6ja70Js
VAXp9x9yPIs/nZxb8DXJaGW/pLMB71eFmovtilpLxFuoh3vvZftLgW1zT+ZhVnwr6EsSlxQsVASU
EFUy0Lf4uSn6qgf+SIJoIUVlAyjR8y1leD4w6B4SnGvEobAWKthmpIzUIQXe0rG+8T2PbglTD8mU
9TmvUt2LP9HhIt6V85mVgc2Dmd3uhjUc7slXC92yUSimA//f+FA/XlE/plq6mxbHzBWoQdv0zIQ6
QK5+si0lWWVxJ6k7UEFAmx+tXzZCybwJIHe634mDSfHw3g9icVpmaJSlwxHo+jXJbF0wAlDZ58eM
Pmu5HOPNTpa7VgLEW06m+Mte1TLzwJ/H24xjBiIFWOnhzRxl2AMoJNMNdex2+DqLk2QVoBV4pPdl
KPPlf3XOqZBZkvir7+2/nviezYbsidSwD7T7QoV4IOvmBKRoE4RdTtHc+CnedL38vkxWj5MzN98F
uC0x5Zg4AIKjMAQ4iUxT8giNYz1ZjXhvFv5q72oYFZcQRVddrKdgnd0mhw0GCGOwfuYMyHF3ZFZc
wQ6Yvm0catavh9puKLFtj1iVqkZhYheY6cSEAv7Fw6X/APoVHQNqExPUttwDaRdUFIROUbgaZoyY
w//DhhaeiVwc0dgXhV7TdKEjDgeWEbwUVnFbLQAY/HadWKjUgPpSlN9OEUA42w9chi84y5vevH9S
7l632LH93D8hZQ6ad3KTa0nTL/4DtsnRa97QaNYHm+g9nQ8g10NTyg0MA4Q89hM8HgdSZLeI4jPB
GENEZuM58w53egaDClG1xmCOzizqiJXilHh56lrLy5WZlEdHwM60Hn/42BkFGtjmltYPs9LKi2BT
pBafwtfMH2aG0v8jE3c8bAV2cHCLDXvDmMiO49cWq7YcPaqZFyxx+q/QAUrdGFLJe0WbUZ9RTEWs
9FOLVdqrkfErwdI1/3c3tfJPNvhV3Ff/Ls7a5gcdC1Am54erywtplonKGcJwF5cDieYD1Dd/5zeJ
WlniqaPdotK8wc5b2XMUuIYqfz0aKoBJUg2teqfVOFgp24eaEPEXXz5qlJgWJOrKqMYTPv9AkXLh
n+gBe6uRLNJGhaSfTAZo+Bl+XQ3k9K4CFj/kzm4c3c7P7AwDQKRAU69RLUXSpsIDga/ZpuSLQ5Uq
G8nUL7i/w6e0qsWMtdUaZbjxMzqkgLFzz30oitJjrNm8hfKp+EnjcWYZ2GFLLtbbSQKMn7fg4DYi
keBB+q9ImL/7eImLnDBiaLwetLI85VPeVNk3/buArM8a0/92ts4tG5yIQ+h3i/1cwDfVJsYLi3ij
j/T7sH+zDmd/tMKAlp5QyU4y9bDLDiPdyV6Hb5crKIYsXJl6lAOnq4xYZwC3/hJV1XzCWe78mDPj
lc+KLACQ8hTIGKfcRjM4XzYwz6ML9BK9rk5NkR2AQgJvuhAWghZHMeVnBI3FLT8chSqOb6rR/7LJ
MbUOtOb/YIGqOdTuGI4yr8VlAPXY//rRv3PbjrxcFHOBjo28YNLvls9dlUcVnQolwq4JtaV8xcC3
tJLCy0VK+9UFF2uKJbQDTRhS7SD93u4Cb5GY4Ruu7HBfQMzcI5j/42+EoIKXzaui8fnPqLJ1eJjf
WMi3QKu5bEyaX77zxSaHyf9pbaYrWiDqvF47xcY2m8Xz6caj4XoUTWl/+alVv2LJO96aLhRgK1Cz
TIlgT01HlwbGsL9wLs5TxU3aMiG2yJUWEFHM3apQ2lF1JqoVLKQgiQB1SFVBzoKmrSb2N/Nw2Dxl
5giKi9DPlk5vOdogCnH6NIhsDZiR4Wro/U7Z+5Y3UuaP+yG2t+L8fOweBCFZrACTWrm5y5qrzsHt
34G0lts2fojS5+3gOLKGFSywHC1awkP1LQWiKlVh+tPHTvyB8nF0rlU/7W3ue3zVd4jCMHvjMU7m
5aSnOTIbyPWaR3U3TfzNUqg61V/iKyMQ8QulceT93mhPdPVFYKf80e0qRXsMtvkNneBtAAcQflt4
1q3yHbO8v4wiF2EDFQSqDUPzL8ZftoKVj+TIaEtgCGqHYps8NwkYOvmoT6mliaxknvhFxSMLbFjf
2teDXygMMoPYAMLS1fBnJS+XJmySCLAE4izRy7JhtdpqLUvXNI53OGmfZMK2HL+n7gWp6WODqiJ3
Q2yCm5W2lmSIc8kHL7CzgUc1o1/9ZT0k0IHhARjJ8a4ePencGGa6ROs/lPae/9Fhp/g7JmjeR/ds
JIqHY+Gf9jz12NJMTrqXRbC+Xp+e9B/dVQrR3KznnquJSIrhonTuAt8NdQxfagG+RHJ03ZJQClJ3
c/rXdqRLAIU130lNZf3l4cxfpDqOsmz1lWXNhTeyXjUMmIL8VKrzyZo/2Dp6WWYK8VZnwF9E/dXy
xkkCU16X0l5fmFTdvmwQwpviRQ2orMnPj5VyUx1UenMl6ewTAaQkYr67Lt86otofW9eUVVPGE1Vd
S43FYRjB7+RIy+EuRDqgkW2JPYtRyust2CY2lBNSuQHyMtR6/Lm3qblaOE5laJRct1+QPST+6/0p
SpRG81znhF3Ks8Zwr4YlqHhQu7MAcL8SXdZJ4owPB5M7Po27F4ohNrFS7+j+Lfcf4I11AMZc1HAP
n0eK5GT1Rr7UCDz9Ylh9RUI+Rk3TFvFi7O/6+8pftVAUf0sPvLobmbzjgzkzgccBwhKl09NM+MbR
05z7Lf934MVwLrT/xcY+/sjHOymcP0b5TcvxQqv52iNcryUFJ32GrX4wzKFkcrAe38671jqEw0jB
0VgdfDD/PaN+3zfa+hzfLrH+1z2zaXuXzEVB0HcvVji64DX+k393ez/wp+G2H1A0+C5VoFNGG0Et
tFxctAixO6n1t2WH8aHxCtkS+4yFfed9fL7IKsDInbbLRGMadaM2mfj1QjDKu5U7Gp/Y7zSdttab
KofKa4T1WroT6gegkkRHP2hJzl7lbDyKPtzRJcegvx/v+/d4RdvA0xk+ztMmzJC1x3Yl+viVbsql
MULuLVS/S6lCzQECdo/nesW1WCqtYsYoV/vCBfiCNOb421rQM6QK2+/5IX2qR1QTZyDypJN3BKVI
5NZ5P3H+cmw405qVAx/c9seuHoGuuS60RLux4xidUdNJ/H3zaWMDbJKGB9jaFNmfxYeFz+Si4zrM
N/xG9hA9lJfylyujVPSij6sd5QIZ7ABNGtZcnVmEiHpJprawAXbT4hLZBd7FglrW8ZfSnVa6z9Ql
H3qdMqpcREtY++6TkAbSdH3jA2bHsAdYnMt6w1J2NIuubcAlkoqdZH4lea6llP36WmD+2re+YtnR
nYKYkasog6tB9/K6hdR1HtTXebZ2Fpx9AJO1hjTz3WXTMKij1OGn+KDsWAYBhiaI7K9s0DszgVWW
lOqKVV8enRJNkGW9kJzd6TlD2VB0smdWbvLkFr3zCEOWrNgdMATP4JqUo5X43gQnbHORpiiEe4aW
+4fxu277ZT4w6roDI3btL12X8mq1u8MJzYTrdvcsFYrze7TNVz6inkuiIJ2bzojCKn1ZXRYMXIQA
g4HRmA3RJMddyonUiRoLRPIBdM2sd8Eakjf+tuTZeenEpyIU1WmzLQmQ8LlFCdJORpNWHQsfdQXw
vGnbUN67mNf7fTysOKXdbG7wd7Tyc/unQdOZKSsGKyUg6umNG07kl5nXYvaTTtZNh5wbelDnXT0e
+698w3DfquDEU9ztmEfcBKTu7nr/UlASmhIIlKO8smhJQFLGS0zzJdRQqmZ3kxx9IL7sMr7HlZ6F
9LWIYiLb2LmRWtMA2L6gtK5rhI2/+Q6kWgSRQr8lOJ8ZfBT5CGAcUOHCFjoiB/2QWHVDKvIPptsw
Pg4uUJfBX0hf7omiJKAeKdCzT6IHOSXzLp4+P7dhw2WgW7GM0RegN+BHSZOBLUYiE+5kTqqB9N7X
kVrrwxLWqDwlphE2tKaWtYbDPpNTZbD0v3YRC8lYwkeeX5IU50vPUibojFTdYnSr+Vag4gjN04W0
W3Rb/4Oao6ehQgiHaaeSckHGyLnQmRZPaYrnGkMLWg+G3kqDCF+hLWv8tecEBAGxnuuHfK8SeYE+
uUuUSVxq6EHIp/jbDSQobLg/SN4RMg8VJW2ohCU+gVD9lbxjwqBqZQ5O/HGQcciHS8D7s0b1e2Bv
3qXIMVxgMPnY+0LUy9zwcVQu2VBd9QTIVZz6Z5ur1UA3c0GPLGehIzDCyJOLxfDIaC1vgGVTOtWW
zgwxI/i8gj4w1zOYGoY7PrVC1IUI9KXytzJKygC7xRIQKt7F/LSaUmvw5riRMlW8VFJPyRfkPqPB
iqrIL2+WNnyAlwE66lqBXdsVfAn0hkP73wXqEaPo+yjKa7qsM+AaFlYx6kGoO5duZba0e9vLnEon
L0bZCq92P1cilGf2/kJf2c065JavhZiuzxbKYLU4G6MP8Wm3rRduvwJNTJzmEaK8dh4BG70ndVnJ
Euppiq3i3sa12BirIHcySlkX8LB8IY+Mz3fehRG57ckVAhmOAw/FwFutV7h+JMfA4vxoWqExkawn
S7VIiUSZdMnbNAN3NXSL6rGAbPMtukWSLaYbjO6wj7MqUF+o1b31vBCMrlMqrCiq9oPp2nFdCXwy
c7i7vsvwksAFAX/HhFbJVTskPw2jNYe4dAzW1vl6fG5EJs/YfUJWmih8d3F1BqHdOdWLpem82t+t
8Wp/JuL8JR78GsL5hvGS/+m6l01V3Y5SiwZsaBJ28NBU72RUYSiQqbPsgBsaby6uIWYlI6P2Q+0G
pWHXcmzh7eVvSijqtiCF5xUQtxX74WzovmUvnypdket2IxW83W5/TqWxVwsX74Xr46TRaheANA/q
uu5CNpIpcmDI7mfUyL8VBp0wdsywthpFA/rLGIDcRyxDN7S49LYDIgNhxe7FzoYjpfDRwQPHK0Fz
54U4+iuy15SOj4szYhlverrrJmvLcNEekM5zehKz9pzixJihn3ba5wlnmVp+eNJnxKe32R0cAJGs
v5B01f6IGWvIMkvSIuzFTQv5YiuLr25Gka33EaytgvZDDloAnCu0yel2gOE/dgMh2sTMyD0R40Q0
HXCTz5Jxk09NaYtppbkE9a7SjGIzu1blP4l1O5+YqLWcvycfz1dgHWqFBjJ1chxKjjVZsXlUm0Q8
vcmnk0Ugye9r6Oqkij9yQ5jNbzvQLAclLcLOIMBTJq6srre82u8ZZlmFr0H/EjeL8LYqbBUm7THa
zq0zteSzbp8bnV7NFD0oXoqdtGpClADNPGH9A9PDidoStonP876/x6dnxHUbc9xLupiPBs962mwt
0WsJlmeBnEbv9Ftp6qhKQ3AHjx9KfBTJPX2FP0Ph8neQLQMSBgwpg0CCVV1Y7YHfJk72cHURVly8
2iNc+To3QkDzlxABqjyyV0odilxQJRqV9B1u7+ek5dKINRPGkDKi9TxGZoOKdpgpxCFv03sq2pXp
+0S/BesaZT6coW/fX0hROSjfurws1dMtoHDOiG4M/mv+LUsuy95pUc9/iOASyBJQK4Oxlc7yfL5g
rkQWWrxsmweQGn6Xj4Z2zz+j+FiG0tV5vSAAsEgUcH+oxPMjNZ6lYVc7xDbWaOyZV1fPcaOIznj0
SYu2EkFIlkWEaBC+4GtUK5gdWXkqdvJ+QWfI6qryXxg/zv3xs6CVQsAigClLb199PyGyCLeVyoIZ
/ZS9D+Uc6dxRtwWrnhNagcP1j+9tUOK/sKS2SIPiLn7bdd0z5Rl0WwZNvXIS4mj8syn07tPvDm0+
Mp72EDtKy0MsXpzu6gsdMC2Am4CAGGSuA9RBOTIvWXqzxis2t9qeF3bDHPd5QPyNEjdRGOtm4fqY
VCbZHKcolC08bJxdgCbLUW1Tct0h2hlWoLJZZxmGwieoL/6OMYJaGfWtLUNkx5665OJUk0t+9dl6
RcKX6pR0WJH3mBoDxEPDFLv5xpJMsY6/kz4C4KlR52Q2qeel2a/b2/dBIU2auuYGmu7G/3QFYXjJ
T68wfWc/smHXPIpwVH+Z1BUr6JlcLr9zpPzPQv2mKm0HT4KGFPTsev5qXWwTRuEqiDpumAitDDiB
3Ger5C2wt8enOLlHqFRNia/QEx/03hFmYF30uf8xKvSoq12XttIShjWIaO0RLDW7Z7+R6BqeD74y
REedIsYlCi/PGfs/Ra6HUIrbdPvlufNlTWNQ6V/ovTX4ZerCxLQIgL9Vui+wIP4klAS9t1hG9Bks
bu0NHmnyqoHkbvOyrrwAmn30sBq0A3Mw52zHnmPBzGKlwyoXHZiU+h2sj1B7Zu3horhlZcCm4K0z
+yj8kN1wJrNT7ypg1gngnLcnOZyPD7u1MS5iO6VyPLGrm8M+W4YiCgeRIE6uk2LLeSO3I60CMACM
ri52tukMxTLh7pbmzflqPpT7eWm9pS2LDo2zY2apPpZrP9QrE58N0mHBQ8i0iQQIVHITJKta4jHf
JVPZT7SS1rTWmfFiq4H+jw1NB+Htm6ziGp3i9/qMzqRxEdMRMXFYiJZFFiOWaJhT4ecmmCY4l4F2
ck1Hu/lxcLGHR6glZ6vC88oi/FwKP7p4/rXw85KjuOClFUN0vDFyo/hCcAn+KJ+NmqPrCXILKlK6
PXOpLWSTFeTXGR0HxGlc3B6IBjbIyKn/Gu7s8RVQM1ohRYGPLX1dmuo8vBbx96UiTHMOItFNOGof
LjictFE4LBAkvZ9INipE4LZxvDEqbH04gfyCNCi1yuG/bhLnB5X0ZXkspQEX41M/sDjdyIw84N3U
TWxCF1JOBuKEBagySJr4lbY8QwHZXovMCoXxjCazGnsBzfR6avhklp4bSXyhg0oOvx6waQFm/T3E
ogKHXr+kPvjXz8w7uJMryKLTixtb94L2qQpEihb8d3E5HdhNWnQwKeaKEuMUQB8JYUzCyRgrN5MT
sHq0kn4w7FoEh5qTykNtZfDiLjGdtOEotZKyk7KnlVKBvWrR6Wl4vFMVf1DVbq/yMlFfp3iymaiu
nU01L4SnsVrkt2jcw8nc4na0FJsu2pl9/vFcq5ZVqSubxqopFD6z/D3oaoDapar216erhpgkonYB
Oc/kCk6d8jb4bdbUHML85oUOJzDL0jeuwo8Cj0DxlboK1udZNOuIcZChnictDFFMWylJ1SXSGWcI
W1X4X6b4wFb5ejXocP1J0KoW35szGcYxOrLxqdGQzbvdDHptcgfZuZ8K64jSnRkM4Ho2pt0NEuUZ
G5UfNTTGL5kkDUhshjDSWFmDAslopTbYeCLQZmTHiJpRD8hbk4tPjajVgvehwV34/RQ3p8sxj73S
D8l4qp7xVm3hUbQFlHcMaN6/uh6l+pPeoNgP+K7Q94ugdqaIqzS59WI4R9tOwocYEi0Cayj9fr0i
yw/RF+r1TV0DDMJ5yPIVngPjyvbYujvJbyC2GxQtoGEdUEy87fX0EH38uzVvMQM4DE06YhcodVrc
kABps+c+Xz1L5Cf/ejEfJeMbUdkwJo1jDM/Eyt0pe5quwcbx+0eQUONF+OpgIRuaroYksuQmWsZu
YR3C8wClNZhyj9vrUW9j0cX4dq3zc9o7LTQLJPdRDmlMwoYHj8PPKVtBKCgCc0oPMjdzfpAZgRcZ
XaJSNg62u15wdUobK2JA4wQMSQcBGWbfIdHva72FEXIQFvcRaHrcu5A0cXUYmcolpLytPEFvsdfa
gcPyV/HPVnHEdv8L/Qt+ZIBvwfwIP7f0wLd4+fkDeu3RhiHE/1MQ+vhzEeE0CWg2Es/sRPCbvcxe
U9J48NkPKhWQxdIK7v+SlSS3y+4AlKMNM1GR3z14RsbbcaBCEnKit4qeu3PDUCFlYriRws7zqmxN
Ix4jyD4JQshGbnhL8Dxf3zTQIvEtWZJXhrSaZX3U6hFjG+pQoIvH8wgBfLbzZKDN7aya1G426GLo
1n7/bkyAK/rYe+jKLPJG9rzkpOj8olT4dHPqg1zkXi5iZtykSQYPma3XoAiJzZNIvLdNt9vedaj1
he/ji7ynGaZMlQZq0xSolrYCshMw48nSSQ7g4nI48oHlj9ehhij73dma/AnPPIRWnS1PPvDYsnrX
vtikPTN8g7+ztZD2bxLB6ML9KLv2SDUfdYkkH9eDxyg0eHd44RmJoKhpz3bq8yod2jxQyapW2pgA
Z1U/d4+m3KobaGPamqYxRMTiokZ5uY1zZ63iRJ9Oc4dzaJfqWYE5BKduecgpoL5NL0eaQmkEQ8//
3mRUeC42IFcY0ZllJU+/FhhtfVGiuT6rgcy8VU9PTeOY/lA2AEhtFgTA2pRcfSHYtZQTDW8nZWQd
Y0tyW0lRA3jYid2xiNzxsCwPKwhWkVrEn0DA7KiZc9vNZRqp9Pu8Sm9qpUFX6wHEvi725dykrGgS
sULLNCNU0PCkXpP5U19AOeIn1qXpstupSaSJrgSAnf+bqyWOvrHVPhve/TKMCpmbHeGvDvSCE5sh
vzMWywOfNQQAAcO9GLbkZw9Kz1rLZZbffK6zZnjq/RJQB2orWD1i0AXgRnwGK9whkwxplLw3mCB0
+tBd+ZqNOXlw+iv7t6YA/doZ/l1UbbhPBqY2id01OEWRA2Z2RethcNo2/tyAPWmEEVo0NOfwXxv6
D0ftXC/014uzzXjP6scwMyJMBSTH0jXzw+qq3fLvYf4Z2fo6mI2rNiIFank1aiAFIzujJ2bLJ9GO
xUZOE+HU2WspGQHt/h2YKSKTbkZyb95Nsts7ZfrA/tjZGhy3zhAlA01fDIal+m041GOjxeDTotqG
NMQZDPI4Gr9EAAJ5BQZqoCrXZRfwAD1TP/GdhdW9np1hTkhjphaxSuuMZ41aDXxEyYZ2a40QXIqz
lDrQFKzrbp9upYOjnzpZqWYZFD7ID8TLeOWNDmIVQasKvYz085ICgOWAanwy2xcOc6ORysbKp1hk
Hukcj2zVU29BIRWYdjVPa+OBqraQi9HwbH6gHFr000M22qDZS82oTdGA1P+Yxn0BBp0GnVw3oScL
0JBhAggOGeunomM7m9dQj4hpZZ6oSZwvslp1uX566LsznITASfRuQxSDe5B9869zVN34l0fHThfZ
33pgW3ZG5+6JngU+QIg0OKOwA5yJ3NOVTdDmv+Mds1Px4OJtyHAIWDIc2sshvDQ9qs263ruZWkCf
gTh78OcUyADxzFKt6QPXsASMA+jrq5MUon/B184x786IBgvP+K/1Rmpddvb3tvuqpXjI35RXc8wl
3cLqxkP46rhVUEfJUB3036OM7knGtId0eP97PQGZssqMDv17oMmdOmOFhGrDS/vqS0Re7aJ28HeI
+VBZXQtIoeGNNBU3O6JiXPEgsXLAWjPLP5t5h5G5Gz7UfjrmB8RcPEwzwReYENk20V6WH79uMDuI
+j7fWIyS829V+HKNK+HUfLUGmsbcC9lRaZWVH3Vm2PNLZ0logOBVv2z8ZkXvqsjM++lnXsPSYf2R
SttZrRoBXq43lqCuEQQmU8jdiCSnPKiKSZB6xx72fMka8YbIPMws22gAfjus2dxl8nj6VMX5xq8v
5+0YV6raH/GqE+ehkvPmXX/WYN5fkO1arn/pBC7nqX6mPWlh/BA8u1N06FZkIovzourdupUlha+R
/03A3PcbfbKRKUBzWRfece89iLWWQaUdRNH5opeNCf4xeJnZU0JOMJ4WIYjrd7gacYZdoqhtN2aY
txfRmzIO1SMRRwUUcaxM1fhxdWmolNK21DR6bM1ihcaeWymljHqZl5vkb/bj6T4VM2J0Kg+5S6dE
WFUurKlCksMQio9JGieFW5okAxp9DAYTpf9bHkZJ9jPnGHGvz2iglDVzfZ3TjWopvFfqjbM3jgh0
Hqy/Etpmbjo4Hn2xPcFLq9ipcP2D9C6QsuD5JX7+30n1SebBDYsvC2JcvB15ywfBQ6j4ZiJyYDgm
GzTqc0XGN3dEt4cfPLIpVKuCQI40/Es12J+oBhl+LwUSDvgt8pI01ex4aq+ilHQNqrAndxygJ4rr
glqIu8y8n5IMQmW8HXzaC+5W8dv+FVg1lgfjGGaHo1Fd8KIOpt6f2nmiyd0qLYpHDn55K3ll6olu
rQSr8t+pjcKPca7Or3R1DQTWJ6CtztJJyz/Fm9q8mq3wAZGyHyK36gXahG+kvbZaTVKmd0jbiIPs
6rL6q4DwL8kWiXYh9sKFHtnCOHSWZifQwdS4HPKz7L9SI2s15NDO/AXPH3t2G2ExI643uOeqisea
z5MxUxss1YSF8Ws8XXm/BNVMWV+l0pVkrp+c8k/s6g22wEDXe+F6AVitw040Wu68j9np1eKOfxpg
3klLNmjTgVXC/u4zNvSakGh1RpT7hkNdcxQ5D4D6cqEi8gC452qL5qIIG6ZBGpsoJS8hBrS+w1u0
ENlN2UcbeC7ET8zY5Z3mtIVpXqhOCuQhaF71WX98DVOB41pDIH2YK2TAUCh/AzSfGyuMQDdQslGa
F80t2G4XHG0KvRCjaAA/EwSjxC90PwyT8aVtsLAND4l22w6NpyZlK7LKTFDWoQAv6FU9EQz/n2DH
mLY1TSqRcG8ZvKIHF518DpBpEInEbx7zUUqibZQRSiyrj1B5ZZjsFh3ubA4SfCfbIVw/4H3VwB9P
m4tbECGFg0HjvhutYPC7p0KVaotIBTBT3Vt1WgIdfjwniIDkWvVTBWSoRBNkCSkMg63IAKL7SJxl
VI057Gj/ninYmm0dIPX0tpvIu3wXOXkXmXw1uuwObV+CuwDr4J1tC4Gq1czwovWFDW6hoprviSyX
x9/+A3R1iXN5Qnls265IVgopxo4/0Pn0jHU12LXuT/vmhaQz3OUalDx/oSHPKnj3ghYYgL9hAn34
rJU9dtJJABcZ7e1oMYl27ijDsok68PfL9f8rOQKkzD6SEqcrPVZN+gfRilmNp30GJauu6ftOqYTU
SC5EPYfOvTQ7M2N57vCbyrWVqegKMrUIQ4bHMHmftJ0bwQUtHyVlfQ9FM4MD9C6Otw0lscANeRuZ
VbYA4cdAv2K+eB2H8UeHBuA2GYbyvklf95VFx4lJhPormX+AqFIbE/qxyp2CK4EovqyBclkxEgxW
TRyvYrPtznRASIoOWWgx85sN0U/1R7Oh/1tsUis5KdrokpaLc/dKaKkDB4A/rZ4xvuftKwJuemfD
aUj7BGi53iaQV60a6gkcntSZCJ3uHHo+5lyW3EiWOvOhR7gWB8K4P+QjwYptyLpHOwKBZNq0vcp5
ohZn7N3CP5HV5orxSsUeCMtKld9RtzcThQzqYVPjqtmERkuTAv80d4tUea8wsfRUA8qngswisxOh
zl/00Ah8rpDZ4bprPTOglJTOrM7+uR8a2OQMVQO8fLJKJCyTtQYxL++5dI4GtZ9SmvXjts/0M5EH
zxITqARtQ4vwsj5AAdvqrrvmgVI1ObYsyVBe2Hs1DqaW+aEkGDurFA0E4Y7FVGcMIsPni5SFJv/P
+IMSHuASE6ejq4pO6gh7zN7cnthikJl9chKaddIabAPxdlAZUqCYkGgfejr7eUkEdbAnf2nZLsjZ
Hgp7T1Cp4xYxA6j2dKHAqqwrvAQPTzAhso4CRHyp1DmMJxFoEuLFQsi67vwJytOYpoSfTiJhdooB
CF0SSxTzUXgAzyzxz1twghLAe53I6fr3EII7McxUW5y3WRfI0mARTyHmxpu7fnG9CX9mNjoZHIj6
7QtEwMmHtyQx0XH/hCEokl0WosTkiJp2KxV4cIqd4nM76I/05U39b6tFXvC6VQbiLsIc5EtoRTFf
J24/RrPOBgoTZ0sTYAgWv9IFi4MGBPGcr2T0wPQdeENQnQUPpQuHANdsgLgdm+Wx6n5NT1UwnOX8
rIqTBia2Wb4sVA6Pf2d0iFwuIQV3yNnOVg3pKdtSZylKkZhOpVsoPUuKvGHY4pid8rYiBLE4L3GL
IQKy1kp7d1n24adMB19iY9g2RaNgf4qhOH3SvFJ306t3HpsrUSHCxo6jT1G00yXFbaoxnsQco/SA
KPU9JPBw4nrQnp8Wl0HoT68uVWD05yjhspo4qPU4C6peQHipXKzPelHGrdH+so8KpApUAmx2mhQg
NwhnCI6xxmydxuEypKHTd/4lv0/ANaYgG3E/KKtTFaFsXBC+iKHfqSnTHypQUavd/ion15Pjwvvj
gsRwcBpLGPCxyvH1TUZtHaUjE3PxT8on7IMk29fCsP3QgNRGvoaUnbREvjklOUxeIUaQgLhdP9pc
m3IAYCkuBL1aEQy82/Sd3myCCatrUfMqF3n76L5pJgmrj62cRlMetASD1udWA7ogY+Jh2gsKsjsY
GowHnO9B7lKcMF5u0suv27oESsRQ2weKYMMygt8GK/Onor59OJuqV6HVyTDmiDyj9mdVgTbNMwXP
fx6yQVHQcoCPrAntAnxjqzFi1OESjbl9hmQOYkhZxOW4DQ6FbtLDvUjUmk9MdI637BR+lOXPBsBA
CpSYTynhvV2r/lwnAjlQ7V8lXIITY/sjtvP/swkbBE+xqQAZgX1od8bJoh08P/np0FR0nCc/c+KH
/lz5OjEVtwHx0nBaSvTw/kf+qpzhM6+5EtA3GSkLeaTElHotknHFDymh7yxhTXVJDA6ruuq0FcUc
I5xlhdoaGoMCwmAXmG4L9AOt8o77KzF1FfUEbC++eyunSvc5Sr9hOj+t/S+VBQ2HLG0tFrDZj3KD
tH+tAOIfEiVTJIQUfZxdbVj9nldHcSkQShDrZwCjx9LhaPXSpIKFkwciBysYjTeIBVF4cwCf3/Lg
SMjTq3JBxCFXKKTKI94hMq7UbXkZE7tx8ptvKJE7x0+SjgV5M/6WXxftDDAJ1LPoG1JcXVDKRLb2
hDW3e55+E4o8JGUtwkZ9W7Hl/RWYtu4OnB/SGAHxRyDhAW8L4c2HyU/TK/zESpXuZbH42MoqYACe
SlyZZnZ9yhjdTamzKPwG6/auimK4cjFr90juJ5dQp/tPdhCQoK9E26JPelkzYDw106hqxw8g6QIj
Mhat79/KI8VAgdrxrzKC72mabtNJNH37bWZ9T4AqjP3V2PUTCI6ODbj59h5LnAAsQT6r3YkHIp84
QDgRc58lkw90l08EjR999/5XteHgsqysRWbnKMLIXwDnVOHl9wuGBpkK67SzgrDEFGt9221QYj0R
dS9pZ3Fes8+y3pTaZLxDneIaOlpCTbvLxQ30TsxAWqgLdfwImhb0y4Ex1tG9UDH4lmxTtJsTOthM
bmT1bxlayzFPkKtIJD45oHh8xAKHbZByenpQTw98U0+pSEfqYGq6xJTy8XdoecGRCD8L+S71ecLR
u2Ax1/o79hhh3CtgWGfE7lBwnvNvCrW9CpnCI2+BCvFCoV9XzXLW77gu2WHPt/IdEtZJ2dWgvd+B
ggIRoBhlDtLE4VXrQ1548PpFk3hexLM0A0NOzBr3BXsFDTbLUEYuccRcg+s4BgMNmC6aFGXovDHQ
lJ3mDB9043D3wxZrOInJoaCoO5PYYfa3iP1XiQlYEQljg7rBwwuYz9rVMMXL46g3r4/3VioGkxhE
krqlsrSJx18uqZJP1CQ8tlQokecRNc5nJdDf2KVMc6szvQWzr379Xws0DhCSvvNHNyUGgvn8xgkl
K3TMtG/IiftIGnU+mZFxU5MM9LLZ0c2E50zRgn7AbXt2hVAhNS72OFCVStx3n8G4A0gjWaEPcsrg
agCDX/FWfiDgkVSaU3VZRpB5EqHAJmxGRN1oQwMg4ykEl5NdJwhSapJfs66ZQDMFmNiAf2Tf+vX+
23s4imob3wk+Pn16PVpe+vm8K+wKAMg7P3rUEHeSu8hWc5CE+49ml+SbcFf4NfQ17tZX+4MjDW/o
Is1kj2YHLbBscC3bijEIhgw52xDTMEmiqOouZ/DEqSmyJ8tH/TubsuyMnv+sl3AL2YP6XcIyWLUs
SUWShBEGiInZMZDQNXDz0dz5JWPzxS1jvg22/ih6S1wqzjhRB3tm0N9PGQn/6D1BnzXAdh2rsXh1
TRYByPNjUP+ELhyhWavQTEKoXp95z+9vgsK48bgkarXgduGxxfC0TAfurw9jtaTFczu1hUJBmEFa
buPHZ+9H7qzkGqVGG31rzEyaTYLvOK3ck+F8akJi7OjpkzGKCKp9qoFddiIbKAvVS5dGd1UW/V/F
FIJXSFamWS71gmWVfPkI37HfPSEUuVzbVifIJs+l9UBRWatqIZlTGHzJizOYePJDkZflR5wgzVkS
H0ckBzSnEhGlQ2V+NeOH5MuPV8fP021TU8yI/sJCLuvf5zYusLbE1bMW2MQRcB5EYV8TePMV0t9f
lcC4wDKjZz5oXgbK4PE9zMWcr001ym9PViH3xmeUVLIdCwGrMsPEgnNPnOgC0vnzuEg+OQwHwPHL
gJk4ULUflUGPMnY0liEb6yc9C8kQUrqOxAl4ey5I6Cc8BCfCztbKLXR2Y4kNTyXBT2EdQD8sPTFn
6ToAVhOmFQT7Ev3qSqM1OriMwGxRLcjNa5VXrdsCsB1zlDJk6hkUvGhgnS8U54frC0TWVnL6jNgj
zY+G5oDjOOx7k7FG1n49UPhNniBbVYN8Gm4/rR2qAiJ76OjB+WNR9SpqVHig5FyIPrFs0pZ+sBmo
3UTljht5ZZRbM2ZqcQB0UlFUjrqFlRSbNh+J4Rb+AmXrgDwNlqbdnE9DevX97UY8qarRDLB0Rg7F
k4yptXpXB23vH1SA2lGWgET39Zc2lbh8sTyNqmEKbXnAIdx4RQ3PydLIBc8A7XwilWZQuHk/gaAp
krae5D89spDF53MtCmfjkLspf3BLRTVkLULlQlUMpuBzBTp6qA78Z22RhsJMP9ZS4YLmkjAk8I9f
Vk+mVxoCd+RyGKjXUxunjfiUKaJA5Qu0bAzY/8Krb2k1JMbYBWiSzJbVgmCRe/+FlEBjsc1LRX02
O0jAZLjlHXNg5aPKWGVICdIXN4tvj/JO7g18TBgSPf6hxSDJI5PW7ZHsT+vX3sR3eZlIMA/2LigJ
9YqGMgJbAxqrdlVRgTKXfo326TCs8Fh1hRmPp1KSgcx5MR9IuNwUexEcVn/c0KJOL8kFfKqkl5bH
RSeFFCgPXtWQBjz/OLknEzD+8DkwsKgiHDMusmJEZ8vJXG9RWs/BpPLkrNjLp9upHozm/xJ1mBtU
6ArEOtkbr/vQC8QJ+JDV+JBFUDk8muOdunGSvq/xOkS+QEscbP+Te+LOtFM99aK7tog058XRflNn
wfSqJb8B++fTBW3PzVnFpieSQ9JY6ELgVx8ZTx3RnCH+zw3xisx8fgBNUa1+C8p1mkmk+WdvWdpC
9vEq8Z138zonkRiStFGHxIJrSegzf/iegoiQzxTFadsFnXjVdJeK0ZkV3aJMTqL4YGZNH8Dtryjb
SZbVV4DOV372jxqWi/WtaHMbAcipa4bHFKJTo+1iA0Q447Fc893F/KJ4soM2LHBGboyOs9Ugkh2H
wUjx663x2sJlgIeaQBsUHEUcrTs/ErkpB/tntoOR04df85TPqlGNaYXZSZHB2br6lfv20HSw5hdZ
BVI4g73PucD33ZC0uK21Ir1/2TilR4pN3YGC9KOqoIKpQANGysVhh4fVqqwH/IPdIy6JI26F6LMc
+OQfrbHqu7NnTrcjESofOCBNm8vwtj51suxJ3wkuBGs8omsJT5ST75rka7/Ib31J8s/mbZ1iOMSU
z6XIRJ9PM4KbnDrL+mhQGGkR1C13OCRfzqcKU/7gpgdWps3qf+wCgrPZWP0Ty8Swx1w0+77sfDqh
Sjvbha9H+gvb8qpkBUEQhLrBtHUsxYo1do2LEjjlqeKCDRFqoxaOJk/qvBq96M7MD+lnWK641lIA
HxXgivo6YGK7fr0JRE6TMozcLCdgpicEMIp+Wb2MHm53GgUWqN5B+ioofGcbfmdkfKPWM+bdipqL
nWHGjoNp4NmkP0FdDoa0S7HawAKPWpUeThNKIYVOhX0wXDxnqljhHgPaCrGOGrs9mtoZZQmVq02D
9I23ToW4vnJoXxL4ByhcsUC8SIlddxoGE+h+u5DZ1mGkmuIVdgiExS5RtdcNeAz/6nQFH0HhNjYf
SqVbvlXachf/CUnlvpNtxtMM2JgWSiogJr8+svCdICSAOQP9R4P7pfFX0LnW0eFiksZjykTXjnfZ
Ls4gAiRrVORGfRPabCu6K/yq+Uo/0Hcsj3sn4Llc7YBiOTKcxed9IgTG9S8tm0wBSuLWhAHU0y4a
dDTIXx64NHKvCsjN8gXBHzQ6t2S2mscK5ME/owNeRMoVjLr/oUhvg8El5CndQ9fsXfd8/ZZxBEJt
XP5Lnk1BVBMqxaN8X4H7I1P5i48UT87bSjiuJ41+zFFukEDgNX404ItW/6z8L8FWqvTuxQDxN4q6
EN2u3RyH6TTm1472ve1altJez6eQC7JnXi1rYpv0QCJZag5b0txzyuXhq5zZfVSR7ctntlGj+QqB
Wwat1HXTh+zbaWOqMnu1gPVPKrguCBLbvVydO+8smvMAJkKItlZJFHbku+tMl+j+8uWU78LYL1UH
ETrwWG8QxtklmluLdcS6sJCaFh2x6DqPBF/1Nnj2BN3gSX8f5CfmzLXVsv0S6s/+PIGMopPf/Zzq
Poz5KkREok0UvQTwpbKryY3wvo2bNOWbAXlJkBfnFv4qAO65eXnDCGLjnC5HyUS25uYx+NZiJnl2
bRQhkAG+6H/v08+cRthYcwodRMTCZEk8ZulfCQc0RzIRu4Kq+cDThX44cfhvacMxANMVxXI7bkbM
hTWrKYGWRovB09d4mPfrrPNSM4XWrKTi2iZaRY8Qs3VB9i9+gciv1PreI/qwdDt108OFqAbOY27X
4VuzYIckEaCS7+zpcvXEQ95RwRWywlhoFyyHmwqIFQVn6DkP2fS7FeTUSSI3l7YORZTfmuTcFBaO
jG/NFQH6JhQ1elc/fHUx5W0Avc4y84Eb5S8y2n2REtL6Pag6YI09kESSYUui8Zh9aj62nBs6VTOw
jqXzbl7CF7lUpr2g7Hqu9n6TJj4zAZ/GrUhJGNezxV7oUPvp4Vy7hIgEhU7HfaD/HOlirDwkcfwO
f+XpWNijyoXoZZcWUVvJIV9GZBJAQA1Ix8LvOcrG9WFIKKQJBGu9+jxW2mCNCpwZt+nFM1CHvXu2
neX1olPm7Zm3wDEZfyWjjjGHUv+3yAC3PUncQ4Vfrs48jDnOTZ8nlO6zQEysjyGf3KNpV8Bwf6Cq
cbZr9LCQpyXY+mhfHDPdcoBY6DB8pru++nU+OiHuZx2dWI5sZkQhbuFfHBeJzSCf36+L+vAGLzf6
9vaWAgvc9RLmserymrPubak9ddWrFXPrXUGZOpzst4z6yMstbyYpCEgeAuUh06A+LGxlOOxameSY
7WayhEy+f/FH1RKNcrhJBFCgzPVj1wasY9vxgr85ogzaB30yGn2NwuyXU3HMOUtiqo/HN0oh5gp5
Xwox9/0tB481WnQkSzbHpYQuh8KWxKhQ7n7u+tcNf9FruB2LT3VMfdscbFke0eyv5ls1nB3ETest
5zV4z8/c8owjoodvT82HUCkk+j35Dl9URcE3s1AWCa6v7GmUT9jlfp90fiyYUg9qyPsn81/emls9
29iZ14j3dH8aowTRsJcg03Lejq1I8qotSOHKsetk7901SQwfIE67Uqjg4kycCA/ctMu9R5qCHZD4
Bvn4L1FWHj0HbHKvZac/wYey8B2u4VFM8yLpWbhg65kXIqmkg8uojOZGtf5GEIfBmnZ/vCQ94ce4
JXUsdpYfQd9rbUyZPDQC9F4wPscOrk3lJ0NozX/a8MiExloFwGW/Z9yt9u2VFUDZCLDV39/wm/iW
TfQ3ZT43hASQu1+t+IxTLjno4qRK/8KqMY8j86PKuXePnGcr3Ng9/EqKuT6IRuQVVJtUKP17cVdo
JaSpnc88SdcDJV6MRf/U66a4zTD0TLaGDA4nMq/NgLWqBT+OwBoE7aBNspVEY0r8Lg97m6OQQpfw
2kVkAUkGQ7T/w/e2EsFSzpVrDdOBEJCFCzCYpXGcXvRKQ9WYvaWdPFZf+Uwu5vSpPSARRdrCxjfe
33RixA5jLsrigLiHcwyNlcwMdqB0iLsAxyfnkGjNvdHvtWzWwRiTCIRLVIp8/Id1oF1Wht83gNbW
oMT48P0dXg6/ORqHnIjunr99MiRpWU8augFb10Jgm6d0Tz/sLQzEcgUY5DaepeSuk3tnqeJbi5l/
F943AxGZL58I7biJ3M0eGoeSmF/K8dMVvA7y8D79+m0+C0lTk4DtOGRFDgFPnX4q8Qi82eET0/fD
up2vM+JJogk1Xvj4akFk0wzCZ0756zzbpQMFqexyFeeOpm8VQO3hc3+7Mk9gY8MJvU/VUPK+vr/h
R5CqOZjyU4CPc60IFSkODX8gwVS8A2JNPLkJlqQicvamI7r99GSsTJzdCV9srrHcweEa3MjeKAsE
9BUj47ZB5UkYJ0vHbQKAMINpsvy4E6dboLVKPQbavEyTnsXzTNzJMtoVdu6t9BFxuJrUseqaG65l
lsQ063QRJB+DRk7tnABMQrv/P89SyUwloCCGebQziVHEkjo2CygKI/+xxGMU4KSQ43bS9qQ33ZiV
3eYJdYJZQPG61lI1mAbByP8J0cP9wXtSdGX8b4JHzyYOYmutX4+OYMpVVmNquvy4rqLQn2ImJF9y
ireD3rmww2qs5fv3lza/yUMAMCFy0EinijQzUoGAdVy0RbLKdsoOR92Hl946ZKXxq4k7xo71U2pn
0FVfD7ZTBPcV0j3Utp+YVAsEpuS25eibr6NjsaEiZ3FszYqrfrUvDsR/CP3uaWzqmRIu6q6jG1Hu
TBBSloHK3eizTxT05PMa9fY4fGWMJgDv6l3CH9nlnTsZSVurxAmOuXXYuFl/WrR/WxpIaX32873m
kf2TddFSkqkjzHua4Uz7hxlyyXjAL1Dh6ctrNkA7xPHhnKFQsIvt97sTue0+UCmPUhAtbaDX3Lx7
7YIZC65Vdc9H9ejlMALup9qp5TuOJDQkkodqFC//fN10s+8LDHlBurFIpZD1VKaRUDeebZNcsGZ5
Bqz0w8nhC/BMUi4Qo61JB6lq7GeskjUgj/uervG4NzBMNHvcD2l5/ilS0BJC9Z+Dr5Plyys27RUQ
xsjEQ86fA12lQMjIF4Besj/3AdjyC/AQxZeVMazTBJuV6kciOb1JRnKd8nTlOme6PFJsU4PMaABe
Ab3np/d3ep7hQXsXhVSbVtUlG700kpoqVrNtoHnZd2RbAp61lu7ljozfJ3KR0+5WH0JCVFSWxMOE
fnkkJUDGsO7OpHSSC4IEI4W1SBRZ4GtMJLbiL6mZZn9JK13wsGuovEka6nqAG3o5SYaO2NJ5Ri1q
qMGyPjBAplS8ZfDSJXGRiWaiWXQaFpVdjxVlRQ15mcDSUZDhiylwZ+CmfffN51Rou7J4/daccsC0
bcV0GZa/9u6/YTy5+R5S17c8AHBeC1kwNl08N7unjpN6roykEGJVbIOCH60vPn00WsVCQuJC2nie
C0Cj2KM9DbcTvlFjKCitYWWv03p0fQXQolhPxCAU8Ldwd0Pw4qo83vj/YzRSPKE5cQzJ4SU+FuQZ
6QO7KUd+0AM0qXW4FaefEL8O8+Atk/6wHsJN2gB1N6qugYM1GKQnu/dD4BKjOIhVSE4iD8ME3cdH
bWXJ9XmI/I/gW+1GhD7L6JtcFv4CokFN6UsJcswA2PMrFHn1rcQFe5XwkjHWw00o+5qM6unsEY/n
GmnvfvkZwTz/hg48JPuSyUHlunicVoLCkGUWYMj8286TgJS+lYcTIOncveaKz/fYtiOnMlce9MSB
bianJIPfKkwkhy5bRuLHVDLh4Nti9QUX1RN2qIHZ1vcq4NnWL8r5CLh8d+3LBJSU5H5CqKM0H0h7
XpnL0ZVDYMRgGpFQc5M28nVsIPEOigLcFfX9nfp7eCshpj5Bxmex/F4Rr9HvJBgjwq9wGLMa2OIH
h1lJ/bZZ2X00SvixS33qS+RSEiGz9z5RAOV8pzU0UhvWmDVY4mcIwTIZgT7/RsakMrfcspvTT1Um
l3yxz6UzISXp7OKbGlxxX+yJQn9r61P5NAtfFFNwWrVrVoRdMKy9YQh9WNTLmi+lXfLZNTgP0xN4
1dc/0GzpiNz27E48jYSYIktOkXHcQ5SbZwDGNflkoe8tpBgiav3mDNgfU1FrII8Ggoi7ZqUvI3LY
Simpivf7hMs2AU3SJwvQ8AHKXUTPBZHzpN2qOEQ2SyBBd4riPNlGfyotsrls49XZMl1jc9a3VN4U
20mL/X8MTlMkPaiREmi3bIaup+WzFOmV8McaJttnypLX7XSPn019tCchrx6borRgydeEaRSYvXT7
Ac2lD7AZykihGRlvpShWx+QILnzwXzUK5z8ta25g1ttKPqg24EB53kf59gDcPvEWV8Bhj3m5f90K
GuATlQwzHYCs4ZabnJz982m+Z8cGpWrnQri2y+N5otrr2/S2z7jvRd4W+9GSEFdVHUqSJZk35LAA
oiIFOn4ZPfDO8z8wqJlm9RBKU+I5VKJU2dwjdi1UScR65qsnhafsLTa7lwdgX19M+Zh8WEi+v5os
fFEaRHvFQJTCMyFf/SDXty9QnFqELphMad+Giw7GNRbdll7OjfEdsfSvsXk+S9TtaW5NokM9FZYq
uzezbjdZvwsyvVrkxWyHuYS0s7qBJpwgv/VN3gfq1Kg4/U/b3eG6PPI7jPk6c/W+JIpaRytcnLhL
Yn/JHVass8BykMiNsrLLAv/lbeX8JWU9kdxEHFncFYlma7iLVs9fYHqpzGK1gFTGtDA18UkVU1xU
vNMTXOHE9Xmm2W/21LqZOJk5u/XlAmMuoGTJN3zMM67CcolH6EVOB84cN7/8kpMtG74abQ2Y/joN
WHuCXmeLEXHcRV8r/dwo7uT4VAZWEXqjTWtB7fi73aJKAWNnfk0VH2Za3F1+lpG3u0kmtDiGAlUO
LcvqE8VuSjzS9jKSNGJu/CEmBOAhOVAfWXjBA2otTXHcZftyI0e4fXok8EN6KMvaqGOhAIbXQebG
4leQREmoe42QNeWgOkn8auHRM/Jf+AXQ6x1wa3CovLvhaOulhIK/xiLIPeu0cMV2bTmoWlmATpoB
bvxXvnGoEcvTeDSL2zyvbyE767s/xV65z7/+0sADRDjkyvjTf7nAVtOWXmfoe9+VGqte02D8+R/e
dWH/o9mV2g0G7xDH+qupjM6KsG0qopXpZfI1Iy706G8R35yXzKmlIYC4PatQ9ZkrywdYQQzN2d9v
MBOCyL4m2Vt4RqPtFHP37I+ODBQdY3HYSAOKtznlwaqGgTFWnpStMDUW7H29uAnE8pHLDfGrRH7l
tZRVv3Dkuic+kn99Xf8z1myWzi+dbn8NItOYA0GrhT0nRbx6/F8S5xnMLY+VQTc7+3iXWYLPepln
Y9amUgWRaerfuMBn5/PGRrfJ2k2BcUtIQqhu9yTHh57HoYkiHd6bO6MBgmYXLXSbsK6KBjPBkrE+
NnFNQ9wgUgOAdaZ67hPVZ6IY2gYPHsU/yDFABO5QfM8C4SgdQgor15lGhuXJKWXb4lsI7BfQ5l5r
iZuPiO66Ghx9zC1Hd0VFIgszbfY1mYkCdngXcYlNn3gffFEhBhWrrz3vMVDFi1WoHA6uKX1Mm7el
TbZchv7LkpadEyAVJ/kZuka9q1Foe55CZ1DnJqIhqjMsgYBbugjZTjmFpFyeGKbC2Ha+vAJSkauL
b4CZQXrG6OMr/Fj2TH2URNg4ld+1yqbK8YVe8kE9w0GT4LPCtmFbNMwTGNxLx3gogGxGksHd59mE
k/oP2WCqHOQ+HzHugdkICkIAfYfjbH81W/jm9KIt5VyhjAeJ90j2z6RrAU+eehek0CD6CPlxLPx/
1SkQVbBHIFAS90mCTrfEo62YLqqVSMq+vMxTha6UL0qvgWjyDe6B/bZ8sUBKDl3lAg5JLnPFVSDJ
e8OcHVveEqGkCUlD8MYeQZgsdjZ2iiTZCqo83eIMtrzPdY9p1mI1A0jrGzF/Dsw3LRk3Hauvy9Xs
KhLQrns36dJhfqyrims1Hw1cHaobfEm8K5V8gf257Yci8cFpDYbnO5gURFbdreLUvE1jBOHMtTQO
qkAHcALtMwa5RQi1Rp3WqCDlSV7HxoPXQ0X+EafV7khh/EcPJZH2tBE1XbXL00XIvCO9M0jHoPGR
EjqlA3OT5pq6CkFIiMnrIDnKN693gqDy/cJ14zTiU63N0mtaCNRYm+0uNFp2EhPHZtI/ayn/gmdB
/M+aiNcjSq43bMKDlHSN0O2Gx01JEIQoLONh6A39xg29mVc/Yt+6Jk1NGBQ84vN9mNUs++sG0dAG
yY3oTzRT7OKlhO1Nj9y6d9zP6XIRB71LttkGzRA3kqM62cUJy378M0sDi86jOjx7C8TfbZXctS3/
RmR9X8MTeb2q760WKqcpXKtD/Y3y6Jt5XN05eCb6U0NlW7OpjKtHWnVIHaefltNkzgp8Mamigpip
7mUPfjvzrvU9dmAMjyksTBJA5PSNGe5sRn0yAhES20PwsUFOahK5zRI8OoykXsVHGDlfM6G0vfuk
qFX8MXqIL2xiDfjKFIVM4LTQ0+b+4OfUhC5lFF9IRK/TqypOqj6VJZafykq9O/nZkvOXO5t8emJE
t7Td3y0j5+WWD9Fic+idnObC/LW1R2VOT0WCrSwSLjRYubcDJXQMT4DQWan9rVzGo1yRVrLsnTl3
np9rQyb7ugZpz/09n6KREpvnicMZNuZ5TLgIeUDU6hBH4Ns4ixYaCVLxPIPtFi+xpYJro4+wEu5t
8fHhowaROGSuXQ9qJlkxgfmzRgQb0jX1FIG/OkItNHhhNX5dzAdjK46WU+YZEBbbk/clzCvg+FEF
F9+FOAp0SatuKKLrSq+7w3xsL206snlOG0vLzk7aBTzc11TURUJYeRK+SOQI9hKDrzdMmSaD+j0f
2McgyJ22hqq1LQG3HbjxTeCoJAojDPIwe4XolktgkscSXTLJ0o5ayB6fLeDoPMqxzgwpRGEjUcVJ
TRo8jYCHaxAGKfAwvixiYA/BVYGWlCLNEt8kIxqLUtEDDieWv9mMve+NgW+spSDlkIa90A3Fsr8Y
ij7ql3l7p55CB/iI4MNk3nj1uysFEhsw6PAPYS8FmHtDGrQ8ysLq3ZkVsKvn8wgJDhy0YNhewK+F
BRFAystDxlebFLK8XqJ1nYNgg+3RXy/TrW/Dhdx3tOHpuDy2obnzFsvKZlA6p1uRlmznlklqmLHJ
EZ91RohSTQGaa7/gVniSrg8z3rMVy8h91i1HHsiZnQOXFHWaBcc+1jsCcihcnzkrQnDQY/hrM+uK
JD10ADpTxwdNmRa6Bh1H9WCVYqMhdczdgem4fMu39JjSHTFBn1sD35+5rB0gU2NVta+pmp79fwGR
iMWamt9w+WxkxzAPijyp1o3m8UwA0WrxdL6SrIadPrYA187M7JouBnsiNuTU+HpHMP4ByJrOYAOd
uO/Ael9reSVLvOqrXLZTnT9jIF7Zb23uKfA2T0LMOfJPjvziA+TG10WHEMnq01KK7zzwG5hmmPUq
1vDraULEbVrCX2t3s+ESWmyj0WB3SfdTTjSH8zV65QS2KkNVyq7CtOd25oUnLPWLR0TYcAjzqA2S
fkHeyd98E0YA0YsnQskZnrNE4Tzf6cPgId+jMqTdKBmDdK09GC1hgkTMNvOYeVXoOl3DRvxkQqgF
OKnA4XgAATVJ9NrYkg5NpdH41HRFNTs2xk4mXpbPX/WkT2LFNc589MJoGM00bpWKWM2AsL56IU9o
6675Jsk4dun6zWJ9uBmRtLbAJHbc83mguGJChESpO3JFRrWVjlwYtHuYxt8X3vSxF9j3Lwska8s1
0n6hYxG2mVO1076Y0SdvwOzi8RIUqlbVLNbMsGsyDMQDji0qjeooaMYQRp0PtVTo+iqXpThQ5UeX
pIC+oDNMK72wQEq/wvtuTGx2LUscO4xrxfYD7oLtZShJDN/yaK1/3NhVs29X9jN82THsWePbhBkQ
qjRkUbspzCHl68nsPT3VXZAIReVaQJ/OZHDnYTBMVo/Kxe5/oeoddY8snQQvWAdce+E3AZ1WiEw0
BTrqglQPwKk6OVpL/eBPB6WdF+ykAywwXFhf/0lx6M0VXH6LDWhpW8QnEh/M/O7RcPJG+jcIJ1Lj
nqynS0LN4ty4nHC9BOIJ73mLgRdnpY1Syy6GWc+YPYW45sVIWAWAy3HYf+YLXW1eHUnx+JqRkKUI
qi/rNeUIsXdK/WrCw9/xhRlgzmPNc9QD3i0r0Q3Waj4q5M+X9fOgCcFMVVk1m2Y2KSrVz8pi+xnO
rqfFTZgfci7xzL6MNKc0D0Km5O1wbe3WIoDfJCaCkLrqxnFWFFqYaXZ2AmbMWADo9CDZGV1GIe6h
A+qvZn9Zlz6fibOZJZDiMGhvPNK5vlqbB8z0Jgd/0Y9N6znmDHvr9QavUPTCw8BmX+52wO7z1VOa
/R0av/iqK94KqD4Q5TC/pT5u4LsK0cBSNQiXjYWtjBGhj7RqJxXejiipWllKVdASVdML6LpzV8Pd
pEtOMdoerDSDoW2ey8BNjB8p9FGxdvx8Q17JyEc2oMyZGNQ1cZbp2lzwi2C65knsGxw3BjSSjz4I
K9okqeOmaQvs2xjQMzesX89bA/lv8OBiYCxBRLPcd6oBHrnFjXHaBziKc3Zkh9UbhTEPpbI7HUOS
50ISVhIwW657320o8S0f47Z+6QdE2jmaWbUk8koip9Sa+pm4SDKHFEvawFxCwulVwEToYEe28soG
dLQ+EfLwEzKFBMQW++x8e5oId22wrjilRtlCPWPSHcKMipWFM9UpwQiK0X2vZxFko7XQj6FiK6eG
lqkuZwhs8OZZ8/zKZ2mAF37p/NAI6xhKrWPJ9TVYxe65SMofOZjBO9G/88smECMw5Bfk/pOryix7
hdMLO0A3yDLJutY90VScqDJ5M/OLXGM7GbiBrZaeLx5PZB6sY3EyrP5h87LbgEvlN7OVKPqRk7X0
0Q1ieOYjgEMkbR7M7Jagkr8sP8telOpWD4lFCA8SSdBtVFncb57G5coKRa0hEunmxCzsWr7qrv+x
f0l80Y8eX0OqIj/8pNp+L65VeF4975eR9mQjaLworR17sLUEsVdJhyEnVMhMUBWuc0k1ZQXNP+kt
HYe/+TI4q3C8IKUBZe4Twj4y+HcAlEvmKiV+WE0zapRTqWm05hku5kD/RbOuKdollZStkCcn/0Sc
avd41ww0rZ3ASe+bzESYEgflesshFPx1cX0Keaj/5UMh+l6k4e2W3y1vdjsotpp87Xe0AGtMU5Z+
FYDGJivuj7BkEr39u5h1/nfaUOTYzt6E52Py4S9FOwcrmXAMT+OY8hTwJaWPUw8zhgVGvaGTv3yD
Dz95hoo5aKdhXzwg6+hgj56IQHvoGtOrMA7S7nbeuQ4cVUyFfPGT0fbP5FJi0g9oh7fnkI199GT7
7RtO3ijkZErxsmHUZfFq2TlkYuzbTJvU34VzKShhv1ZrbZ1enT96rDSNYZFmmFJpfKqiiT0WvPAB
vLtiOpHhOsugsI4E2VDkOSoNZtnMgxHnPrgXnQr4zL5TyQgkc7j2rXk3udgJSwrqoCVnPZKkjzxr
H1xgdgRxpOVlGGD+ElVzReZ7rXDs6+Yfjhwvhq9P2hAn59hgc8KTOewPSKcNT0TzWXBKmV/vTbSo
OmZkoCzkRU1PNqcGLaoJhmud5uskrI9hblQH73tM7LUbH3NbYZdAVk2y2fGzXKSMccL4FTJKfTl6
faotF+hZrvczdBJOQIQ4XSdLLsG+ItNsZOzZ/EQ0NZ5FG4Cvy2j5XYNUd6yRwM0t55TDZmCnXzuz
1OBdLMHKTwRNYUK8IWjovUiQ2NZebN57qxLXzZaulLnUlX5q2qMD7D3G9Bjx5cASUs4UTE5848qI
liWFnJNrBR1nk9oTx2Tt++MgBcgmeRAVKGrovGT4nLZIYk1n2xaAcp5MY8BvG7YPzx3q2n1AU5wz
DVJ1Jqn+c7n/N+wbYkshY3gPO522iklzBg64BMpLxA/Id2GX6h82GwrzpnyqYYoq00/yntZVlYRN
SfugMwYCZbVJBvSFXg8Z/ZGBGSAOMjPWUsI9F2bB+7cL836Yy7etLJT5IqMjnAEa0q84RhDF5nYg
h+G583AQoL0/MTOZN2P7oIfktQACNuUtIWsGtRA2+QJ7WGSG7ZD2oiu5W+iRk1evCvj9ul9/75n7
uwQPMeGFA/OjGCV6QoK+f9EZhiEvO9qJNSlSH86a39jR9nmPpej68SspH8sGcdrFBI4E4k4PeSFL
uUoUHkrqtU1bJsRDoMFSHYGL2W/HtQ1IMq3sJPWs8/qZnS+OqOvuCeHuzLFk9leo/viNQjtTTgqe
iP4OnNNCAk9UstJDrw+iZupy7bi9+gHbxkArG3qbEu8KqxhThYtVxcYDruNbeHgBbJ1y84SZaNkK
rGBLbKkkhg5tR6DgoE5iqUqbeSwy8FT1Tzrqkw3b1ORcY/dv9qUu66KfoyA0DsoBv5tYKOyYBEBS
L2gO1JKrwO1HeUo9KXolsre9qN+tD6QTzPpTe+xAQmsFl9aoRfEaiT0pqaDwxsaZg1+BHYwpqvP0
zZ5gVMRq2KpKEV6Rokys9kU2q2ktnjbytkMS9sG1txq52Kwh4+1EqLjTcto0rRhneWk2MdiUsQie
VubcuMzOaEa42sVjBrMAPrg9jSLnIfr6S5c0p9z0EOAAoPcOVJxJTraWeged/3NgpkUztwJD7UgG
lTZJgdQW8grVPH1D3HK9XuUMMeVQJNa6vgiPgVjhR6+zBlEKii23xq9oTE9aeZ8FH5kEmyp8A/Xy
zG35HELYmz3o8qtO9XvLhlt//ON5LbEfD4myr7lvF2N1Vmu7sHbgt95ahxEi5zvQyBWDocq9eh70
paSp5W2VOW8+ei2Wte8YSXB+wg9BhFkFTxVB3nd9sHiU+LUlDy8UCoBuZXXWavMMwDbxSWeNGKaH
4YDvZ3Ic9CPuA38uf+8Ot+vslnSUe+Dyj1chDcyQTdFCZ47k3sfSH910X9neOmmH7LyN/rZFE384
MdlI5695ietVJAwId5IOofF7qfuiwDHfSAbGqyCeo2eUPAhhA9/BNO8pa82RHcCMLOPyX12kQvQ7
0DoVLX/x/9Bj3f3wBstAh+8KyoRIOPLfrwwVumlLpugtDZwi2fWDwR0RAdSTINUYshBed4qQ+K1q
kNiohHfolcJxvzS2DLbG1Yyf9Kh3aL9mZwa6iHr0aww1f3jhrM9GydGyPRqrKpPf4ucWJaA6LMcO
oESCwfu43RWR+erl/IWun6QdiGtwbsQAPpiRH9cXIvd7QM08EpmXd65fMwmd+7tBqFws18ZW8ZQ8
UAQdHw4OQ0I0vbB2DpTY9Y36mTDvLbUBEHkBzVLgODrfkVRiopmgTVaGaGjYH6nv/qrv5Qnflh0r
TbOkgHGrwMeTnb8BrtjTpeNJMetkyk1UhbxVjBslT7zBQgQ2FBtC0+rEPLsX/65G9cSy5TmSLAx9
GebxiVwERzLpbifrrM10paAjYhjP4eY1EubFlbPds6JfbGvcNGffpmblNrchzwPbfCG1pv+JHFlZ
WpruWDE72Qm3h9mtEDIvIHnVs6lJu9J/GqijAtHKoRl7jFtiiTp3Ce5g6kKlJVL2tF77O6bKUOG5
Li2LUeb1Kl02GGDQTDyTEx5+l90HVy5/PtguoFfHNq28h8nPkz1OYpcy7/SxU9EoKZvb8fsk89N1
3BmbgoKiErjd94JWee2HXdiAPDpCrfX25xJLgAws3AIWiDAQTa3SPoain4KX2VRALv+tN30X6Zo5
sFWbuEZPXUDhz29tRdN1jLO9J0r1XFXJsM4GTEyCCyRf0onmr4j/6ftwQD0lw1DfZ1JRW+Gfyk1Z
SGJxve2dS5oXI0S6nyLNI6qXR6MyTdeo4691hVuRrlfAbQOpF4g3HMWHojtGhTcGrtxzmHlzxtIg
gY6jlyixlTvrPV8p18UWuA92qHx5/Hv+IWE9Xi4p3fmYyGfC2xnPnQT+yOtG4kEBscAOlZbM3TIT
HAMT5fo7im1ao9dCqykeot9L2NzGSsSH7qisNtN6JS1Pcyo6h5YW4QgkjMFFh3eFfBKkkRJs/Idi
NayEi2ZbSiLZnli//NBqTEio+cHPHtcxoocM+3PkwPDt9npfJ6xYQzpUj6ecVt5FI51UUCc+2aGK
wDjCkC5WYXadU2nn5YEMYWk0j710ECrPlS6jFs+VAtbibWGdiKQ+3HdTmW8/RjMx4RR+rjvr28fQ
GZokllrbbzZoGh3tqA9vQO+mtP+JqNrB6ECj++aUmbC5mr9baXDxXcfRfz83WQEwStSNY0KGeDnK
AvUO3PtI2NrgtF9I600hYzewRAm+CupSmz/f48DxaFDHvPBOcfoJFyvBs1ul1EvF1yXh77KrICWa
mtn7EFS6LSk9rAJftyFvYTqEzauLeaT44LwT3VeQrJn2MKzKABnNm4maRcusZo7wsIm5CFlbsg0e
lklk39FRkvTM/ABY6sXegMkfj11LNpMgthfGU8J+HGC/8pPCJsWXGttcpa7SZ2MK37M22ckyEw7A
3bWJrPGmyQgPQJaoz8VYrcCrPnrhu23O9Azl9mrk52zFT0Z0RY8AIGmy5iliBG2n2yvcrC44fi8h
fBvdtEon/FkbFdwTsmCRLOxjbhte5SRsn9A6P8mqoIf75f84Omu4EtIvUrt1USXHdSFSEcsFYmck
M+h/ZvE6WGxjqHHFsuqSPdPRags864MRzhnWVjuz1VyFp4d67tkXppIPFaqzH/VRM/ikQja+ohbF
5AFd3q3/8IpwTg9EFsDtTj6S80KHXX8VKgyJtoIBhcS6gV+cojJMZVhbxYzFC2G3wyhajcJKlqd7
Xig2mkBQ5ZYypzXaYohteH4az2fsrdQYyo2e6dB7tvbrtVIUBe1cYbL0jaY5ra7TGgTk2yQv6N1M
4SP+yi8FaV1sqHwVV0S7Is/EcL0aIFYtZd6JV5k3QuDOOkODt0xnVJYz3lXIK7BpkLEsIdf6IFuE
D/mpvO95fu0Fysx+p3G4gkxJOdU5Vi1+5Hj7QOzK8VNyyMc6objZoP2D33IkXayzgMZvsgJvY4Mz
AOSkdPf8Icbue/mHNw/NPdwQeHQ6QMjyS7PaxbFMwYLO/RtpncoE4pK+M+nMUAjbU3IqpAvbY4vA
QKJEaeslhgdlkWPeZBXnHkgi0JeJz1NwhIQU7FKWTuDyXeMNAPZ7pUScjaFHZrBYVomf9Gafvxo7
qtKfvYDsyHnK961GNxQ8HGt/wOaNulCj4LSIUA3Ia2qMXld3Sx7W2Kw8Avtkll3cdKm6zsLjTjAq
E82vQdJmVSjtQVluF7y+vHCi+mbM5XWPvfaXWx4vquze4pyazI20S95qJZcDNIiI4JnWPTQRo7ub
Sqhj8DhAKJffyKAg0fkco5Yo5eN4RPfIDru1TL70DDHgW4y6X5/cUAbKteuJQb2mSQEBG2KOxarD
2zgveLt36jdi4GcIwYp3my7BN7LoNA13HKasxj4cPVFCuud9FXciOdEhC9Ur1u5BO/Wblp4WMSfv
FlwBBxs9H2nWmK/4UiLol4G8ONH5kuvHV0FflgkfzB4fFpTDy2neydxL8CtXYPtt0MVbotL+E1bD
O8O5ijV86kepvJDkYy9G1xDvvSIkJFNXDzgk9Fz4Wejr1bhR6riMpH6Zq04WKk7OXxmet8+Jgqz/
hRxz+0a/QBlAzqI6kPMD80w9jNfZtQJVv/isCMY3OW/debshZzLXmdndw+c4TmM1THLyFE6RK+MX
1gb5nLNxRMF9xMZUYN7FcEEXJgqpQShhDZQL9bxr/EQ8GmCjokr9a1fvgvtXLYZTBXw67+dLxykr
ZcsNLtku5q1YbE9fPan7PYPmLCBMee6becpfTxeUAhZirOtqqOJ7pHr9RFPmodGK1W06ICEJ6J2B
WySf8fS8+nldhbxdAYm/nZJRcbJGc3xER+9tLgMUio2xWJ+FYUM/9w+cHN5xnBmgvjJsfN1Pnw4n
u36BxRRHl7n+1+nZEo9s1wlUNPhBcvFIkIwAmcUyX6HJEKw9RWdi1CZzLEY6qRMdSVCXzJMr86E5
7BWeYU5hHINnYaNZpg5G7klF3DE3sxtdUCHYaGvLWdHiTG5vIa6Ctjm5b+Y7xN2S6GSuye0keiHR
Z3PErlyCxKCBMDjO/2PkUST7c/GK4hlx2iK3Fum6n840mvmTxlLl55mZnXdELms4pMqEtOjTkuog
m27lj29+p6CvKY80zIAacwdfgrG8DMlFQaFY8pHL3C8UMYRPDnSDwc6Zoj4g8o+VW7OHyzlvOPHn
8g48DYrqafnnp1RPMdp1ErN1EYFkYRUPRZpIUJg3F+tbmPzukCtm0v9B4U4cp9zZHXnL8yqovo4R
5SWe9slw6TxrHpiWaRAK2dA6r8J+s5QIECLHSLsuCho41mK7hXQrDSAN3FqcCMNx7bdQOLuzqTFn
MjtI5sJRp1OV3VYK44Cp6hRJ9M6jhVa/8U0NkZ0tr2URldosZIq1Aw3IE/1VAe/zf8nRpNV5v64o
Af5V1LaCQ263YMy5K1kzIhAmU3XYNLELdrdx9H011kMB7pIiDoK4jgy48QEF6msg7aWroI1PjS6Y
vGdThrrsA27no09oQf4IrbOVcBuJsl5fPsuF2V6WMFPqphAewV/BPg5XMaQYoI/tFt9DUB/PtVL/
qYhpSN4Hd4UtPwCcLAemEbql+wJyKbcvPCTxFuSUEUM7XRi2cQoSMB7aEfrs/hYDuYHV9Is/jgnO
2CdZ0gGRU9Mgso9Eddal+YInSkP23BaGVkjP5xhVNRc6R2u43gl7EQt8yp4u5mjP0zvHZo5csd+M
Pv5Jm955LGO3Fsjc9jWfETEiA8npEyqHqa9cbNv5+ZuIN1VyR7HQOmSNVlHs57rBf0F+iyA5ZnAn
VWLRY+UsXeuEfCN0T0uwW/c+v9cowz7S2PP9k0BSXTlhcFbfKpYfY1Fbl0DE6Bo2MHfuAa1WNlpW
Sww0N0mpOWDtPT0aELtLdia3EX6EjDcrY4a0b/8m+xdz6bBlXV7BaZifBD8tH+QvfI2tDo7ogsFm
BA3fPa8wnkLcR2nhut3GIQ0//LTErU1NuNHwGPMF73yDwzeF2h8kCO5/+NGL9Tq/JdkTJ3wN+pBv
yeFakk5aFjpwu40Gz51DM8TeX0yUM/w84QroIKKK80dK5KmfFJPJtE+zOg+rf3HWiWpZy4l9PyPJ
yU8GkVo7G3kXw85qXnLCQvSFVtPjQRpu6UueQRKcBjwUnaYHQ+T0NsA4wS7PCXJQR7MviEhEh5sj
t41RbkPeg7VU0nSRDo7jKLsVWzOd9b06/TUtScZe0mpbl3QGzq6HpiW/30wpPrBuOLkiYixY4Wn6
Tmt2D7kAVSfDzswIj30K2Xg5TkcoYF+aVzYtPwjCWl4MK29LxmwxqIm/Ud3BZuoRURLWkud+fCxJ
J11V5AQn67rooCHW4OwmDPCX5Hk7Ujh05wECX6Vlo1RYbiYtYQbshetA+INTOruTeIHQNVFyxQ6J
7ryoQ6O1ArUhmyFEGdd7XiFaIih301vudKjTi0ny3N0HbOFlCGFosWhHljdUrbL4ZFVL7aIIhOQd
3DKzTmecI7D22gM79PaF70Xd82ZjNw4nFuAL7iDc0FchqjAgiSuYGpw/PU3WNfzZeIbUQqb7aGhZ
GCEj0wp6dC572Nun54q9FcbnpMzn8TdjJ2fhyRCGmVn6brw4W6+dUCXLttr4h+Jim/Onl/ZcEr14
bldksV3zQ/tWfNfKbhhV09eK9jPtbQrLYgVCbfViwFhIWvPUK3UMj83sbyVmtSInw0FNzTRp3m5E
x7+g0D6UsBBuTnx3enTNOsL9QdWqhm6e4GoV2mhgGpUodbuBSWYP+APX4ub0i+3ZQ0NFCmp576NH
krBMS2JreRfkoQJNZxdmjWHMi0ZwBjdsr8MPMhRqboBp5kOhEY6l3eLBLeaA1I+SkL+lMwAFoA/1
cpMhtGfyBnkoTer1z/gIdt93e+GfZUiB2lvmoX88eGk9Z4ldjmACYHaoZjMLvvMEiWjOPmPfL08Y
Z+v4LAC5/eX4YcSzdEoQQC3Fh3gms/s4caf1dAIm/ojyLuSYy+2eSTozDrC4FaDVd9oj+XFPaJbD
Jh9D0EFldid0XCP1t6IE2AJGiNmuiAP6f94qsZtU0ArPzXCYB+mkR/RcHxI040A6IRYo5Wz0QcMl
B08nW5rfgD8xdrLhAqFieshSAk/ZF0kkv8t0kT5vZ56gDWcTBeFcKy6hJGUWIRc3k5m21FjHKlI3
ERXHMmWXMDzMwGfcIH3b6qcfcTIWDEfw/qrQQeJaYeeBZsNSwVQTYoiF1JIm9Kkq2msyGg/mB3hJ
D2E1rj6xoNSRe+A7tHy+Pa0F9yVF0VIG7qCAwdZr0rTeW13j7GM6RJJQSmCzCP3GB0EqWoaau+/K
or2+DkwtisKdS+ASI4bZCqLnD8lApKiZPXMvgy2ro7qr1aOZXN+kafSir+eKcTzfRjHXsDGSyCtd
KhRTR6jJFBrVPewDig1CLaMkiA5xT/3orSKjjFyDZ2GCOzt0VOIBEr1iik//6/jnA8JewgsXzqb0
20CeqVdLLUrGArLN/jZBVl+iyqjJ2sC3siOSu1XjWQgE5mDH6MiJPHgYXNJaLlAINamdDUHPtCBX
juP09tcKrpCREAj+XxrUTCFh12iMYfZ6N704lgyDA1HqmFa56AWkzfYGnO3He0jX7EOX74+S7UDu
JQzm+ztbQ9k7Tf30lWCXazsMn2jKISQLzcb5J8z+pjMb2yMpvgaqyv/XZSmtLy2KBDXjkiA62RQA
wKjIwxSf3/ACEEXga9PuFptUB322c00vtQkCxsszG8ofEGiFGm2cUCq8h+i6qXA+3HaTRp8bfV8z
JRz4WH/XXttdKsjwOGu00kSajWDg5z35gx0nL87nUnc2ADEcvkAv04FCx+ctMFhiz9IuuPLVfrZG
u5awcWMo/JiRXXwhabtUIY9EHmHyvYVWNaag3O9ryUEXYGT2t3GqeYIkQhXR93gIQSii8SHe8OpM
ETam+SU096AsxjMMZjzVK0b/uQQaIlk5GcKZjB7e1m/gLFJQ5ETHPjUiDX04lzHtZE7bSGCoZRvX
/plCV2Aps2glq/wDjV36Jo7SyKFW4wPW/e1E/i7zdnwIWarY48LQ2MLMvzCY5P1X/YaM52oAWef4
5CSzdC8X6DSZuKttQAxaCJXz3XNpB4rlExKEoLAgTyGXVDRUDOJeddqtcJUt9KU6W/UVQyMlrruv
nSevh70dfUWYV+c+4hJM14vgQmZpWNMRudoLS3HOq7Py8BbPMjc7jcMjCP81KIGZW+Vv6JETwL8H
Ak2kvjzKpco+BM7XWAK9vKTWEswjrixN+/YUGDZkulA4JWPvCUUeBiTd+imEABQnZi/41yymPZkj
kPNkXgcc2C/UdO6xmXqPeAptXaPxPool6ylh05TMZdrURapVZtKo/DGv+SQI1zm+fkmTURKe4tRj
iERHvDPG/nACIrO098WSrkZRtBLH5uAVMHsCYoEJexDe3M63MFC9aa8AHqePvypjCZJjHJ380tFQ
F09v8sqc3ulQgc5uY8PmOc/jiVx3sMlZav6osXVtQ/GDFXGVTjjjr7o47PmwwpSxcLdTbe75ybSV
wR6Y5pQR3HolEIrxdGgoC9pbAvdV8qrdjHmAavJlQt3T0kmFBgYcxLe/4ugYtRxXgJeSN5UvHxr2
U79H64mT7UEkZoe/ND8vPF0li7Oh7VG8Vn9y6i4+L3BHTunZBz8OX5K6eHSs6izPa3z4S+MBKYNp
/YRxGePPuXoozcOfwd1ut7gXj7dLvlRW082tNeZUM+pVD4z2UBNdaS8GmF+0pxAW5NQQ2h3AD9l9
CkAUc8WxXilNrjCNMkiCDrYY3WkwqBMrzp+dnSN2PGOtkQzPUjnWro566riotPmEgOMpnUdNjBvo
qkQhIhO8muiP8u5uumaHMyvDszpj93pkVCcMIpILouSklZp/k9MPYnDVXEAEgQkyMBYdNT+aRYSj
fltuze07dIgllhXqGTMuHv5m6m9vujOJXc8OcpOn1qVULIBTFmD7NCuyLm+jTHT0NyCjNRIU46yu
S6vDZSkiUMGt8VscADp2/mzFvQKJQKj4+IvDs7SMyYiy1H+7Iu0s6VvZYMGyS8OWyWMPIWlq5dFg
IwHe4zzkiJ7KEPGCbMfCJwnIS0qVWUCm/JpZk/uj11F1tHLQFOSBwH/7gCuYsVduGfk3xvamhZ31
5WQ4iYXHvjutVgdoggOYQhlkk2IHyAY1T8dfkYjPKKqwiGK69PV51bDYQt1eqq8b1zZJegXumAB8
B7MFpiCvGlNT/3tiYKQpCz7s8Luk53MuEmpD97Qj5Tepk51BjR9yacsCOAQJPfMgRsa3nQvf64qX
Ow3TwoxnqAzqFrgux+I753sBa4WAkiymJU5a366clUwb4syEhkZiBkfWA8lzNj2CxsSq77GeJN5l
xeepYcAm1YQ99GvuEuqEQyzd3AR2dxJ7Q5zJ6IHJ0Vp/f9ZUt6hdBLbYknk4ROyaGvPGvhqWlbPv
buPzF536B1b1RIbw7OSY9BPIDdxjygF6tD56jwV0TadDCHJQXqL/RwcNE1riGV8sTilYLxtVBgYO
byNIqhDo289m0TXRrQkfJYLR1AI3Tpqvv19b5D4R1nZp0JjEP6Z2QqSIuwQzmV0Mi4mj2KAbRA3r
xflFAew3fkbVDNmF2Gt2rO2eIihZoyqe0sKFrcNei8HrerxIJIGbtDlr/ZFdlBz7I8vZ/T/fz1Ej
C4jf9BqIa9QKW/tdhue9GYcwCpVyBq3i5K7lCqrydW7jOb+8gHBpj5wiq6fY/o9/mJiIrxucbB1J
ugFSfgqzo9W+1rsHhDmvNWI8LaTKLACBViuZYXBvF1LvkbPmwaNdwKTxz5wmEPbRAGOt59sKZuPS
D6h0bXqfVF0GAV69I4g7zvKOeVlgKe7rIkSdrvFz6BWpQe4reDGTlcd746XG+x5xre3XqXn5Ro2z
oECX+K8E/91XI1/zXmcMHeVT/IKZzmlTF7gvRduQLGFbmv5w3sl5I1N1XyOP7NEdiPt6ubqKy7xO
hcic/VRJh8JbsjMsZKQVangz81pST+H+ER0QZ+pkNIOeC8ZEDVy7J0gAlUOFqe0GroAfuv9akpJD
ENP+HdiU98WjM4QAIo48ybqfxs5v5dPrJGJmm1ZwtFeH+Xfq2uFKR2T0twAPkcO12rq04ehHWpnQ
8HCYkggm47J8sOTjjB6xotNTAhN7qOvriHRGzlnkhCpnBnFBgr+Spg5ahUrOR6uBfKK6B+fJDsU7
XqAYfpgPYORrS71mJKADGXPOLPLc3+o6JrxAthNFWyKUzu93/JqHTk4zJDIUDwzt/dTFkyaR4ZSe
ZYtBV1kOE8jz7hSYAZGT5oUfO0WzuiO7A2+jfsW2wdzAxpDa0FVicfL23NacvI2Ttg18iXfQ9/ds
pQ6w1s0fgMAGjSbV7Nmkd6x4+WOQAfSOGqS7YSZMHuLpDSFjsACzdNsWRkC5PijXIIQPe8zjzNIR
8RwvVUce4VApiRcl3LmfhKmdVSBNIpxAGpSsEaRRKJR6gMLgdeSSXWNXG/maZS6/+rGeoD4MQPPn
ersq2s2GuYnGIahqzKqeIbyXRuixa0DdW9sqfEmvNyFYAI124PW5fX0Qu5Xq0Nv5ONCWngAPIMwr
l31Ai0O3LnKA80/aSeq700XoZ3u8qtthIa8n6GaRxOOqcTF9CE5sIU9wA328bf+8Ytgtu4SzOwwz
k7HqPJosR205pJpy5JzBjVdugl82y2BC+aWE9LKFTUb2wd9fN4NQLOZMPK8JyyCC/rTFHXX9Cc8s
soy1xSY6ppYrCBqG44CjLAw1+ymscNiMpaMoRGRBm9foMeR70mFMgHsZnt48HuryuK4i07HBuZyx
+4TKJTmf8YEH3EuVcXI3RYCTHPmggTgXgXOLSuBYrcOn0sJsjDr/tHQjAfBFoJx+9nVaZUDdStQJ
lET0nXpBy177UoKI8B3hydTtsPeCrRj8wvlkFHw5XHQ42s33KI/8yABr3+jqywK1re1PUY0hISvY
31oeDxAo0Gq9J+moSwrtZ/O/X9n44HBl2HTrxWAeGCvT6t3kxj5+LGPK9YIgrPCtC7saHlqCtWAQ
5tAMDWNuSbRsPQG8e5i+ezbmteNVrq7aW1IhzRrCYxhat+ooG/0XhTw7WvepMkXeA5dlkzoNBeYC
DzWonBmnT0BAQmGLQJnrQqTHYo33cQuYhshMY4tI9HoQU3gn83Hr6ssuSDPW5Yp1MY6VZBQ/HnEv
RvrBhCtqWjbUXr188F8GQftEls9XQaLBjlCrswx9Nc5iQHOeNcz1z055szYIu1/OMByV7kWDp17E
7or0Pv+Eeu1yZEt2ZuaYZvL98kbcucTcycq/7tEqg6o1wUT4HLCcmi482bpqf55Y04thzazRcEaR
5cnmaxk7pejaFxpzBxUKGx8SBZNWd74s1SNKMvpWYWAUqaQnF58XsSAh3bMEuCQY3Hgrzx1l18Uq
MfCkpUQeq/oRhTtSqJOhAKeK8sjBXs0Cfqoe+p9OdmxQSW/x1Mn6fDTUTzxZJa8VQM2w00G6hksm
rfnfXJpD0vPMYX/SK39yOmm5G2Qgha5s2ce35Z/Tl7WGRfyZz53ForXKlWM2nEFdcrVt3Q0CveKO
b7lvblw3aTvvChAsLWnpUsBfYU6PPZnJe+z6FgzyCQInxHEP10laCCcKu6xU16cPGCVQGv9+4ah5
DVqkjD60UhEocE5cC44X+bsfY5E6lvIUR7mzG7I+ueEBvHB+Cf+m++yJ28wKkIqyNWQub59rUNt+
pzx4vovqtKWuW4QhjpaszQmY1bhcJW3n2zpXYKNsc65H216A+utKQLRhpbfz/NBw6Xc6tIvf9h+f
aNEbRB+6DRA7Fe3Ie+otaC0mZOVulW5YJN96S9nm7sqtUPnWJAYygs8srfl3QGxBVL+ynfBe3vAc
uWiryD7IWVHfYANhGbiGytAvjxzxdETQ50M3o+BfBXm2EPc5IDkiI+u0cKHcxqcfWl/In8zG4/Wf
+fzwVJy8TvKK6k5YFL73vRRxVt6CuJBjSoaW/M3Zd6SwOm6m3jyceQ+HA3fM4rlrxQ1ldYb9zLPK
puB32rhUSRIrOEsF4mq+t/7as7WdhdNDpFkDpe08mjPy1ThWhXPgWesg3sKNeQEn3BVD1Mc9TEsk
UGUEhG9ueHG4KZN7l3J4wTCjAhfHJqJx6wv4JT7U7njGDC7WMBsoxf8LWVnGJuS1HQ/61OxNzFhg
gTm8KcJUGG4o43PKE6mYhC+AFSw5lVNouwCdXfcS/OZL5UJvV3Lrw0c5AJB0Z1/lAs9BOwiBbnv2
1o4tMdX6UlqKwHMlTbm5lTJLznGw3T8eBiQRlobylUm/DYqGD4jQg47TmMtsw4A/plIp9/9M6BS1
/Ji5WOzy9K0LIdcAI8byKET/dHFpggKbMzBnHrFGbYktuNmLxx0cruPTCcBx2AxJgFqfPkJXWs/O
jYlF+gnfbskqjEr0l4xT6Btd5EWHENZc2I7DQThJJf0g4wQVoAP+VTsk90ulWBtnxh14gMRKM8VB
HZloeX2p0p31vgg7AsZv06CoLazQ9S7tqojV4ZGs9ZKSfKzXIBO2iYfMsB6gvgEJfNra4Su0Nhe2
MtHzo72TGpPUCH9nP2c7bEOHjAUYb5h/JRYi0tPhRudsY0sPAIce08tXY38hB8TqaFYGM/LSL2tZ
t9b5S/Zav0LkJQq/te2zA8bBeE4mzmFXccZBZuL+cpcULjaX+0myz62tucDx81juHISCfM6IBEP7
jUt2l69QOiEho2/uxtXj8nacx6078srXyVOyQeK+FBoCooR0+g0JUXD+8qjWnP/iM3hedlS+Amfr
lWqBJD1QoXt243iWzc8WJ4ZLHcevn2ss6zuDVeJanFzJD77i5JogJRWP2emPybCQqh89UlfIBRRF
GuydUqV0Iq/82qsWTIChZ407Mdg2GZmDEX5S0278OvorB2MSZfbuZ5I4EnpWq9Bn36fpsjaeUPq3
Dc0ckrnGN9eZk6Je9uiK4KTRDdqxg7fFvNI9y3dkX2CGE9neqAQhGwOkF+uRqg9K4bBT/YzLJJOg
8D89gDXNKxauVFDvoPMNw+pW+W1atqZDmIKXLziz0N1lDbrS4631EFO2AUMHxOPSILEyGSfEn26Z
EAeNs5LLY6Q3dQcku1HfLUDHqK1IuT150ir3mD83zcBXxU1XbuHz0olfPdft+7sLMCfrIjRGQq+y
uTLzXP6p3VTcCe5vqYZIU2LbAQoViygFOwouMgh8WyUa7nW2rrWCHG5wT1Kvm+HQBF+aaFObV3ng
hI7u+5wD2oSHHm+MoITSdPMnpFriuSJlp8kE6+6KuGjk5gkl/+kLUT+7iEZz11OLXxhUQwhQLtLL
UrM2xFSCSubjtXFBGvLit14YCf7lF0mZFzkLYckFB1zO2GSKjr0J5MTqD7rGQfsP1n4X7cCcA0nb
HU/oKGZZEGMNUNG0HvWItUf8iAm3V1b7Dd+4IztQG9iP1Yuek/6DMeJnLqynVsjU7Db8DGQmTsJR
D8ugfeemTL+iiHyr4lpJPnVhXcIuGykhkmPQLY1FsvZtWeuVDijQTpzUxPuZbcYOgRfcD/RdqzzP
UxkH4X84pCEaQjKJTyq3W9v4IZKLTeCqI+CO2i1BWr7c+iRUQKAw3XtvpkTEmHwH//sHQSTkpfYw
cOR2tprlYj83N1Tg1+mVMtkZ5wdXiW1FCA4t0e7gJrsMwaJiNmKTsXgzSX8566C5Ff9WBRy9rj26
joFMMQOKq4iAkBB0px2hEskxwhL2YqyizGwGcSV+PeGMvWQtM4GZu6tC/iOpX8jEatuhkxmbRal5
qyRddb8C31tUU2tOHXKU3T/No+RCXiC1LT7z2mmNe8ymPEts0U0nqvGIMSckrgAjYZfuaJ8qRtqL
TYkROJc+mu7oRVFhfeG7g2BV+b6xiartd9wuX5UBJhSwiGwW19NJ6FMStlEq6ehPXE3ue/LVD/RL
wFGcLYU74OS3dGdz1DoPqWqU62LmjcB11XC3nBlLajaI6dTngMBvqZpjNJK6qk2y+X4K5nO9tWk4
m6QPsDQ7qLp5EjSqVm0MKOranrExOanzHttvYPinencdMvv2LlH88GMPp6V4VsIm3bv0n3zpN8cb
KInjmIt5FP++6vfarYXd0hIvQ5qjdPI4PquO/UtVTY4c0bfYlr872WzQ2vps9aVVn1/uaC3iM/F7
xDMDXBITL4a6AKDpNrk4BBHG3ZjhT3n5c81ebk2lNfWCUf+r6bvcnExfRNsvi0oh9UCd99NAcl9W
/stA93PCsyynnG5j/N60ZR7bXdMv+0MZeT+D/lnvlyjC5QPc37xQ8FAj1CkpXMPbSvPkMjPEeToT
Zwg0JBU347HWh2eC/qlKkYD13G6g+dTCBX0x5n85zKMHb9nwAoOheFqrEyJ6LIgBYCLyDYCPcVXz
WLeCeg3rQfsnQwCHfk/rPc7QCJG3AratyGlu71HHCRz/h7pR7cvzZJp3VPfqVLU+oAh4l5TOInWx
ifI2QZpIae43CsICpLV7HajOKV99IV0a8L4kdA7+vHdhqJoqOuk7POl1vYuAgardF5Swvg6V9+bk
XQygkqYwP3qJV9fA+e4CDEOjUwLtD83MOzBNTaeajsP1DC3brxWGfWB0qLDp7r0BZviimOJx6HBQ
HKO+FrchuB4kIRIVB2cXNji3YhYDGm+5Fls1fHhkEGUPqgrTMFhmrbvrC8fR6Ts11IHgKbfxJkT0
RWAslcCMhtoFrycZvQkpQNV1gYwd/Htzd0XTQpyswBngFScDJyfcEI7qDRqf+IjTZmaOLiTpKND6
kmNQZcw1SYcI5D6MTZ5kk1/5qK7HLt089CYHcN7+9PMC6Ic0UH4O1zZxpupqIxRoSHMTYMkyrUa8
6rCN90/RsvxvFlRlWZWlExWJy/gT5+/qtJx0xQyC9O+GCx7FWlV2bJQr7E7zw+lgI+hNX5FLN1ri
TPINLfq6e1Xq55E825rj56E6KouhLIcdpxF6hM+80EP3dcFh/KbQXBSJiXvZJLLXw6bLsUoBYHTt
WeWFHQyQt96sZ/jvZnhuCdeTqVZpfh4CgaoAGZ1K35kwMo12Y9U3AexTnBWpYT6MHZukoaC/tqrh
xrY+GkjpJA3MsDlIk0AoCYBL7qwTWxrVMgJ92SLCRdqCZCdYaPKJn9RCk0DPsBh+A/PPtRYJjqhz
naY2rT5WUAGeuu1hLSyy/gR81BF84JZaWveyrWDWCa0rMwbFiPAHvpABTodjjzVMnJFu63vl0rJX
rISZfZ6oYWHTVAkKq1fz+QRUBsLE6SAxF9CHJHKvpXWz9NaFyjnJT6r1Vwmmhnlwg5nZzdSo+W3I
nMJhO/bfgJW6PS6VkViRK45kHWwfwFX7N11nwVeSEvLtESfvXSvaJYUUO6cbeHkUKgGB96r4pQTl
1xWeFDebunUeOZxSHhddfHkCrMOdBICS/Xt9tiXUP1YaG9tm4rb7k62OmzRZwHsVRM5BxpC07NOn
f/+WnSVt/f7nSebGi1xihqOsT4E36+3MXr3OSPqE9KjZimWwcaGsOnHA1nj8MwNAj2D009aIP6nb
Y4I4uu9Zfcas8TysijadGlmUbevpMnG/Y7OaWKefhABUa0/wRrYm3yJRTFH1KgY/MFnYBMZ+ZMc1
mUpofXlsPcKq/isT6eM2S5eu73caxqKKOB5cU2mmlPvoh9MqzLieysQodqQsaR4uvQsualEsJH22
Zom2s2X+MXu3YlWkkMYSSii7uBa/WIHFAc9H1zYti+avI24rMJgAaSNraQSLYEMX51Oqo24uQBsi
xkIreO7ck8FLtQuGJ6NN8EcEtIDJaQbs7WWGJ2/jTXg3nv4gJ7QOBI0IjW9SVRlEBdOiEmpN2ma/
A+Ju4tqEa4jeraymNNMkqjvtWGR55l9BcbflRmkBk4ezlmQ52Rj7BL6P7j61FmHR2qYJZQN89Cuv
hWkgJ9E+cYt1Avc1rN0pXBVMerWAgEBbpMBqFqKkoWbcxj5r/3oGzodV1X/PIJxc9BWE8j3tuX5j
WbioIn3D4VW97l6oRs2c0uOddo40yh1yRis12sNBt/A9bRgCUmlFJ7rFR/gBy6FOu8sTwu+piXUC
E9VLrdnzw3vGDww0eOGGYMRjPCzFQp1Ed6x1kEkvNMFn1m0iH5H5G/7g3MuxoTADF2Ul2oG2JSXc
oRB5uxJXxCinJDgZRqN/gu3hIiwx9vSC8Go6fwZyQbuePX5mW58Bb3JVPBHLPqsYrwzDu2LLN7L/
LabYsvv9bFF+w7YyTIq6iJ5XR8xWKE2RZIevzCUL4ECeb2NR6vc39rLH9D4yNpMvlDIoZqrkkAWq
e9lQFUWDrXH2DEQe1SwlQCHHlMhRliIKX1r8w3YW1Q4WRMP9/BVskPYGPEqO3j3/KsQe9PyCpkXN
JwFKDzdS1WALz5zED7Zun1OSRlgijjZCWRqsCfbCy36AxiWvc7lxXzkKGbjMfPy/j+o7obGD3LDv
31LRDtjtlJ2ShweaAwetWb8EzRjQpbNpZpV/cXXhidFrs0lk6AEuKxU3MRIhJYxqyi75LDHdY6T2
xtyneKK14PW4jGq05chFc+d45X9tSOurqmnMce8+mOaB/H0CZsE1qCx3Benekevuoo+WjCuAWA5E
axBqt2It2G5pv3sDcTN5Ijm22Ug3LXuWqJ/6ldLGLo2XSQmnV0yd8hz2knMF0jlh3WIINQr1wbA8
j10Br9HLB/cuEqcl7HH09NgJPnwkBmQNb8b4ZUs08pJe1eHwkfnqgd21I9Tailr02EgEB+NkDdyW
rzl4+87wy1M1uvgaWlWbq3J+QIHvnDVjmKsT0OWvg353VZ+FPhfhpY+MT1UOGpEjGE3wLRQg/bYi
DuVea/qdDUVOkdB2W31z1JSOUBzHqV8MrVpl/kk37uEju2fbChSDNHcM2L2OET+HyIDtXFEkakEQ
Ucr/PiiT6Y3bbhqUihSqBJr4QBKrVXjv3Ga9AGESVTV+jQsM1X9CGAXVS1z6CuwRgW4UnvejiEGc
JsNxQ8Hvt/17FX6Qox9PHYAkapEucFLwprMOxlEC6x1qAGZa/Stbm1yJ/PpORc8vTq+52XkoeBid
yLNYv5QNZ/y9jjTX3m0deuhEZ7wSazf4enzarv3+MivzBSo0byQIdwwAtYg5KycHOIbW7AS4uYe+
oGcWBYVqfFA0+R5bGDFkElI4oN4AYpaAzrqjllOke0Dn93nYaoZ2wyZ7Miz3Rl8fHNyz6xHxub2P
ylQmOWFziBNlA82QINc1WlfY1w7KgRfasO5ZiLKV/cr5Kj1SZwqG+6A5f5PXrjkeOkOJrdrRa/z2
LbezChPJzT8GLRudYcTmpXJUhRHjoRP9pKu0GMg1vTuH796J9taIK5ET1XxtUwhL+I/abdnVc4pM
5wWwuunOsJHnReW23BocwaWA0b4cTVKqpcK/KwDA4zQ3sLs/9sR+vCV4u1iyaiHEXkIU7/tX9QxD
ujzVpNkHc9JvcjxIJjgJP5nuaJ+cTuJqPA52UFCoMiweHSCoYUQMX/3fRYHfw0ESlmc6s29OHnp8
JrWBaZWOQP84WQLCYKbWOOgU9zntHP4U5sIJiRvto91AjugFD59hB6gWNbh3+STW6iVpnQl6s4Eq
/JDFcd50sNhJy7J23f5OnoNLeSW5UdIEsATpMtAROcaFbL1B4kY6Sp/JJnUnVF5L4wQAFyioWQ84
ft2eJpVZva5EbgY5Sh5p3lSvlpOx4rTj+y7zzmnw++9OVU64yGQkaOM2ncK14xWhxsjRNO7IQ6h7
sSdzeUDysxFAnmmwFBebdU49zhRV+nuci6g16EEU1k/4O7oFKCiiNoCkMzT55YbtPKdZIoSPxJ1r
o4kfPBCjK+QsVHtMuiNWus+aRpKA/091ioKMFz50mVMuTkz1Ilk7PGFjEzRnF6HPMviBKv/VFroO
slTDTdlLNIqOUBKHfTABs/Aaggc1tYbX7RXpVgr96/W2l8QKVMJKPdJJd8qVuLzpfytrEJ1jQeu2
uznThhT8Jxy/3gd7aHSxRcSjNK0ocC4ucvD42oiu/LfxESXlcRqfsOuydDP2VcnpgRPTx/0qnX/O
sNrL63KK8mXeyatgOrnyENwOoLICOzXdABLlN3TH3PSizreRMIRfDztxaeC4U3qDovGpy8DMNxLN
ZODDE8mUsXOk9l/16kNd6R5DhBi33Zxo7mVZsf+5PBoUqy1WSRsepbD1q8EohybAJXNyB+hKe9VS
N3nASklsnlYAxZ6tvyhD1GPdLUWaBlHxW5WCmQGz0/weBOPs6eGmFsobop+Hj82OEWnoKnYM3OKu
+JYJdhjIu/VDXAfqGHNpE3OWYedZhCK7vlO7gJ3nPa66SsBNfgeWE03j8zxr7wUNkksWf0K+mHam
PPE7CmDSUNCsekcuODP3ITaU2NkUFkaamKGw2nTkpBd67AEFv16ScqyL8WHXux8GXqKhjh/iQ5/y
KkMmgbYjdvOWu7FRAijSV5rKdg9+La+oomUkQ/Sezzk3kfn9wCSYJ14g6UHV22xhOs3rHv370VQZ
dbW0GDRuwvUGbPEguyKxyxtLqnijakLLJNBLYwHuhgtn3Cy0qt0OHSpZmhMgo7vgCNU159NzKKNN
Z9PhdOMEnVC6GLjCl4FZnYAogSmWWKdA9W1wGG7hqgN56VoMVhj3+IsNfL2ASTrCQ+WYVlFNtjOx
1Fa5PIDnjsIr9lKc13zy6kxM8gubVjJawK27jl7dBU6+PScEtnyZNiuxMFaTeht2rxIvR12I5XHn
vIVvv2+6/CsA1AR39Ret/DGlAhCcsytjErSnsmq53ysd/SFy3rHbHcZSvDJZg2qQ49v9BQ1mtdcR
lcshDLceyU8cCgIUZ02itMuEHTilpfBZ6ED2cUj/arI0NJY74YajI48KnTRHhiEww58ob0umo40s
3WwMBaCaIUaigU39+If6pSaAyvHOB1aNzH5n5O4kbUuvVWPry7uc8HnBcI2gEQoSTMHyrrCMmDSR
m388ergo3aXxTjWWjzN4U4WI1M0J77RY6AXum4cKBegASZNY7W3EKMOo0H92PR+ov+B+QSLd0wrF
eJT1KimygpYIzHVYO+ERQ2CLRG98f+JR7sJuMeM8ae1a8tT0oXvBEbh3JfUiH84hJakuoo7bh9yv
rKAJQRUznDi1zJtH2YjLvkyabpeVtulh9ddJ+QR/ihZr5u12Zk0QLaM5mnjztusP4ABEHJIoXgTK
5wSliLAOTSsE7GOH6+G/yHxRGagdoMoXcbdijTo4Rcd5nkLFhpC1tFJuG4zJe5Y6WaiMj0F5dt6X
NKTY0k6hWnHtIVKqkFbCHYkDGfAFGGFff3MjxxdaVUI+QyqvERHQzk+GdtyXepQCCfpMm+nlEodK
GGGwx60XICLZVBxTTX0T+PWKFhsMAfMM9hMddvqzWCOcahgmPqt+RvK1Uq+4XhaipoEEQE7xSjth
d85ocLy5eWuFckxVMji42cTqAEW3gda+rXe/zoJDl/70xfmH5jl9QC6y9obxdxC4ORQuTdlSTatK
tK1y9IFz+79fNIdt00o2ynM++QGXP/AOnyNo9B/uFiWOi2YS6ap92Fblc4Y7c+esjhBwB6flsGuH
/JmTbMK1ELFUQ0JGPLGhJZzHRHlFH52LasoTIUqenoKbXuTDtKupvS4+U+nv0jLA8HwUG4eYJaDh
QvPdeQddlcNFQDWLDyAV9k7G92lH8fmh2v98HyCTsgKgNw+D2wF4rDxOZgouVo6yKUHOVYB+eOp8
MyFZkAGqp/J+VoLdUDfUmVBIlGBvZDWVzc15pZFsFevE8yFErNiXqsXwKLEAK7ndlYpqeDo3cPLv
eRW9SnrD9NegGjCkN9m2jxnIOwwVSd916tTXr/8qjJTHIjwinDoQildrBgkH2pd/27XD4rKN8OOQ
fyuIZCrNM6d45h1AiHWYSZuDT5FFYMPQ2OiMkVJG2XtRgo7qpsTacGVzSo/TcGbYR/sUM0VfIVnF
Sp1bbLTgj7Z6lffEttnXbKAWAKKS1i5zK5I4aT0an3SajEHHdMJZYxF5tOSjJ3KI5G+H/zgftQJv
tNnUIpZ+2T5T6C0YOr5Y9O+daiK1x9mzpNPEibbzpj3aiz8sFzUisKuoqnBg+7E28G0E4jItrKHx
oMFqVOPzREjNp2vO6m7x4XFhVb4yfmQrFnIQu7AV/L7yCRVL6ajEUX7HpmsuPZ4lijkChaA7r2ac
0l/YaYL9NIygr+Ug6ZSRLENVTNNTKHa/VBZjcEYzGttafqjyBstbIWDPPw9tVn7A4RZWXsT+c114
6G91pg5TEYW+CjlkPXmmeRPFWuSSY37WdhbnKfkWmQpcpdcdvdjtm3ljtEUIP28jK+mWXpeeIudW
wA5EV9F1nra3EnnDTh6PDNWeE6SCbQRtiKsCKP1B7qtHn75Nb1xKrp0Arp6ZzufJ1sfwv3VfgW37
v0mvn54nDE9LyuZULO/33cAc5LM4TkRnwvhYVJAKXiSDKYkXuvFEKprmVcaXas7om34VJKRss51R
in1kq7kl3Z81fWy0+CIQDWpJhENV1W1b1yIxx3NNGu2EBh2UMtLmYCkWJjj/JrNuAai/psFxFCUb
8x+XSXIxqRyWUO9nRY6DsFfMtv4EggVzH5sr7giAJBHMPeLgN8R6q4K4z4VOpwpuCOYqZHcOi+CH
IfU2s2NmJ+yFN2nOXPSrCyFl4NEJ4dXB4dXcX6GDPazpv4Rm4WVu1Lnxh16Cxo16sg6D5LnmERzt
iMz01jWhgDHrJaGLy08G1io8uhpmvTtVIVmBVXKbQafBTCuP6zl4Y1O8VU+DaFQscm3RduXb/PSv
iiFfnVBqL4hn6DVCcqwtjS5HutszBQiMWVPTawvKaTIpoJHb0FLDnKhw8hYnLve5uVZm4kaARbuO
0SH/HKKmsjNIHbJdYaHy8zuw7mm+PY2HtLFbujdzrx8kNwAhI8TeVzFIGZxBt4llyx0hcm1Kuoee
IFm7K3b8DkaBxA81VScGoeaKKKokJkSlXZC7exWzudnl+wl+1LDLUTey8QoArp1au03QZA6pN30K
8D/I1B1Jy2CHoUlpE2FbK37XGvZ9KhpbfL4odFUbH9BGzEvcNMWJLDixSqzLBbjHqisJhQKBF6v7
gxoUYy4zKDntBCdZGp9dRoNYYbLrniLZ8h9orqeeOy/3YDm+YzWNAdpCOW8z6/5OeJvQuelWNWmN
NvJ37NQ2cw7p3RF7znBpY0aJeU98ndGldbrdD/NM2vIaCpSqobfnQpJvqKgow/O5mfA5pMyXsKVg
QJTcEomltAxim8JoXIU2reVmyRPiQZxEmuSWGcRyu9u3za9Spu+nbIlfKue2ZeEr0GXIaH5vyChu
NmHhlPmtm7z2rnXc1m7rVCCT6tJMWia6IqQmNvSe3rn+RWhhHYZ14VefMgCSByfxr5w7ftRPUdSs
M7IWWriRlsYYIYgt6YO59jg6fZqMTCP8+/UYQ2ze5VTCWIS7I3QLJWEDsUGAmoe397lrm6QOOO3w
fWOLn3cLbRML9Lzl6/dLxubqBo8NyOH2a9bs9lNgTn6fhV/Mynb+AbjbzPOt5h9pNw2W9lAPS8PN
0jBpgqW2H0uAYJyjKyxJ0s2VgIYgH9c4GGEX0j6z7JrlcdlmK+eYOK1sPQv+G9wSRaRiMIZMZLeh
XBjnoGLP73L5aLnXhtN9fDnbFd5ZtiMAetxpOsjUgvIzVzvm7b3uaOdqPx0acrw7qmw6G7aURTlX
Nm1WTJN2LvVSvMtnmVh0GwN4Y5/M1m/jfV/R/VE/NW5I7kCnQ2XPmG1GKYzQpLpY22W2j4/cEULl
hkdfcvDda0EKq4WAn2yHrN4ApuubpkpXaZGy1OAK9TO60gDhHeO0bLlCsl8zS/vG0Tx3idTzcoVG
SNhn/SYLr0fXtH/klsCojMv0uwWxrXXOK4vU4MKqc4GrqL1/o5+6AEKaIa6tqArNF7zxLimKZBmf
U/8ghpW1xwYAggE+3ZCgQNLRv7fRprY8+8hlMWLklovJVD5XJTiWZ92a4nbgUf4vzFZ9ceDtTQnu
TXK/AAbFafGh5ZBRqzMSSRfj8gQrpPNdgJZquOX1UeBepuoxRrB6XumMZ9E794SUlG2FWvHTmq/4
iTXTvuQPyX3Sq3j/InGGYx14NSs8Y765wtZuGwzbzky7kayMoznPYW2f+F1Ata9im17xrCBp9495
A+mM1aDP/ja1LgaUF9u/UB39UHiyjwtVDp63j/WBdNiMLmOhjpLeBP82/3twYuP4ZY7NBHZWmUIj
Gb8cwqxg4d09vyLobatirtlzMPkLoAb9vfM0U5YUyKFgRqlRd5s0WJXEH9y0++17/DQZHd7RwkUM
L+n8fkXm1Atm5+A/D+2tszz9PUhwn0B3BuWrSccmd6k/0JNWUnyieJKiqLoTe+txgJg09I1S76Hr
JSBbx2hXsJDGXmqOHd8O5qBk+1nnA2GGE4pconNjU5NmU+y8VFoTSgiUQPYm61MgK9DZWiwEf/jD
yVSDGdQb/JG/sZQscViq0yj7LRPK1/lLLtiGSeklfa5DjrGuL7mUDNNqColu7Rz9Kc1gIg2Ntl8t
CMWy301Nt/yexAN4pC1pn5sNjTP5d0D6XR811uIDtBWfZ+fB4heVZHmOjtrU+UGJAZIEPdVgz7Y6
tFeXcclD70jptPvTKvMAttkpG/YBvuGZ4jTUA9TJlw5sG8vVtlOlf3XFmMm74sNfLwR2jlL8s9lO
SOmKw5ohu1dB85ZZ7JiwU5oYRMI49s/H38Ng79ABrKBGXjJqPMfclbqnN5wsiStipqQ6no+TKnWN
afWWx53Ru2jEWKB/SoGwg267MEtOMnAI3mxn9b0F2CYLLUblIcSDVPxEysBPevxvSpCTw9NXeR+b
iWp1pfuEWjyV28eYG+7NaY/Y6Znv8RHL721nDVoTmOiXlDjJBdheBQweS38KlK4grw/55G4FnKoc
uP2y/TOKpsCsmb+Sla6jxzBXaek/6PuYvAn3KAS4WqN4HuHhM57iM5Iq7qDZ9vfc+uCCQJAHtDkb
+dGDiIAL5X0hBQXjz2pbRoKF1HuxhlKrESxaP/m8mIIt2l52naVlu3bVQw/77JSeEvrM0n8RDuYb
8vTi5wTYxNvhnPH9yOwSHS8W5Hp4y2lotxOMwZDmmJeVs/VF3bZMgNnVdEzlhXH7tIKebuDXmInB
ewg4MuQBPBHH/FPwJqJOz//Ot1xSucImR+WSExarUT7630pntM2iBDXXENiv/dha7WSXLiYmazfv
EHrDPBESMQKUxPKt0BfAdSauRoAp9ZzidtxUaJYLEqolK6vfSWK6T+9BbDxR78aZHVq9BfiiCHvX
xGX7ysiVXZH1dFB/XFtBtRWkWu0lMNPR2VUFHX2BU1e+MXo4BZwP0qbFmSULgBJXis0a9WrtcSNc
1zZcU/Gs7T/EIWI40WddV/61rw7tMgsQEpaMmkwImXR8opByeL92vKS2KCpcQMf0SK44TYONjWDC
6EdRT2FkRuZls2JMj9SndfncmfZ2c2N6d7modUwvlHUq6sdrzirROO4nYxz31o+i99Y3vdAFvv0k
WyclCu17K5molDS1jJfM3PUWFPKrfBf4QhAODuPYH4Pxg01gLAzK0cRC2RszA9PfxhYUOm2lzBab
ocNV2aBUoWLmKd3RwqeSUiEOMx44gSWV8/4Ro7QsEuEtroeKWLQP2ZFyxvCy/kUDkeMf5XPPtEZi
xnIbvxohHHYcibt8/bv9ahBqUor6dycZTnZ3+zG5B9isDGZ5oFWYYIKPTli1rlywM8xJLk2EchKJ
gM1tTYMuF/8p0llMbs1F7+10sqeNPb3RlvSDEFRVPdr5o0qjXHzj7PXEawoL3Ihk+IaujgWC7vKn
B1VDV9FKCGNbYqccqoYf2cnQFMJVPcEWBZ2K7nF3UXXTNPbR0xn4Uu8PAsrv+bX4e6JaBJBvHcaA
cgVXyUfM0+GOYPv3pX3UlkYkXWA2xeqmhxvb5mG7ZlVrns2tFUlmKos621ROFKx7ic3NzAVhABSa
i5EiNPw4KmP+sd4Xus0GdJKukYwtMwqfcSHYxz3VNkCcoL0K7fMFdkSpTX3ehdjsZUlkKItlvHYn
B27C7827NVGYi1MNtqGYrMf1OyoSh1RfSzk0TT+qJx1QX/URiNurdNzxZLwaX2SFy5iM4lZlp4MN
fn0aZPEXAEEOfBokGPXjtLLLz9K6G7xQAcG7rnU/3Fwr9rXjuvGwVaIf7SILU5V0lGPQV5jVziob
KEH3qFR5xm2reNdiu5GU8sJqnmnoQeW7utk4Ujmgch6DGzh51jMd7zsq0gK0swN63OaNic2LwmMY
rVC/C2R5K/TO+D/0UfBbHM36gRDCPGuZjTUdv2TzRlumJ9l2JURGS7xzVdZ9FBeWpsGsOI5heNH2
z4ryWV2ReMNVKsKnXMwoa6FH5gYRDGojLPqDT0lbwbIUtCTjax6E39W3t3g8NFJ3PPA+oHJ8aqYB
wCyRtQGKTUreOwXnPf8SfnLxbiVInBLRoBgesM8sKlAO7P4wqEw5qZr3JAHJ5P5BVmxvynUMG6VW
oeDOLZQA7n1faRiTNrqmWxmRvc7tQf4qUXx9rDozYVBV3eAyd7EInrozSQ8rH+68ogU8ZhsnY2vo
S6uCT2BPOrBtnMbDk9QvQm1CJCLbLP/NqYCYqIsMfECFvaXfoql0YokoRimEe9C5MJGaXP5NtkNu
+BE1IzP+QzyQ8wAYQSXXJD+licB8RP9X3SmJiF21pOnGnWzdNtRop9SgEvoTqYUw4Fhm9vcL02WT
V+56ldSRa5fvyNzdYCDKDno8Xe5fi1sj7bCwBxlXG+7e7sNV99yxChamy4qbO17adCiUWwovLQBR
aEaDJsuM7GW9b6DZUOiwoJS237ST5OvbjEU9yNhap5KfAV10yx0Z/Z53Oj06XV2+tkYPjqalAakC
PwrCKvrKosr1W56IWz3MQ3+scdyhAoBuo6lUkts3s0MpjRJ3GLdVta70RSXTV1rdH7hPEEqP+rHD
sN/fl8RbKSFLZbI+/W2/N49O2PNOjUyz+U947BRH3tEld6a/XFIYoQTp+0XjQnMLUd+/jAkDEuMk
fRpXdnlqmguH37J/K0fGqRM52jY94y9NyustiJ6enkmQy09LDf3Dia1SK04yfOqwvCLLQjqK5mVk
rAnPJnZND1TvuCZDy6zHrfI43MURTelY+r3O0IJ71avDeK9P9i4hc9MaVQa6QOBadYi6wY6m7lzr
paQLuwv+EFR8JlSb/yIG8f3GXBcLrsnoDzF3cCPmhYcKtPr3H+gUYAbiOAwEaxZweWwG8PeZ0Wqv
6Fb1t6ea+X7oWKFKQuRBSU++OCPppbP5kyBN8ucKQ9MEq5nvA+jf12GV1xxFeCV0h3vGN0V48e0r
wfzEioh0p1AfOxNvxc3aWR8RYX5jkHFN+fYWWffeRTyoVKaAi2zGjpMpLzqrlh7B20LMhtEXL5Hw
6ZugxXCWxQrX3JQquX1plGpKMlnAtNTd38SMTUfrddaYKAT+lkCYJlI6zTleTtROKT6qpa47+MS3
WYv7bU6Jis90Xqbp1AZUKUPasRQTxCI0PeqwtZC0xT7YKeUPwJrstQsQcx9TCXIRrcpNlHBrN+ci
c8hElfdD9tqpktcF1zIuha6HtY+PiUJq1lk3npEoBgU0vCJ9v+CAm/PYzJeIqpr+B0MVi2utQkfG
vzH2Uz5Bc37O0Q0Xsmwk3+ZwIvWt+xwnVRZZzI3iR/UQiAr3gbNmUE+mzXXN9eDbfPvtHHaa9WD+
QR1f46ueeOk4W7SzlFg/GRncmCf68GsCTDKgI8Wii/FCyLHsHaORMGGMNh8cpsqER7gOhvc2dDYc
nbo5ATrbUwADBofwiN2NmEY6v6aiZb8ACdmKS1q0xJhN8Rn8qZC7tNq6QkotvZMiKvmc7E6iFLfK
nacOcFv7309ecMzyGJOPetyqlGzYSGiW2qLZ39hgebT2bTZTJgCAf/dbwepcCFgFSy6jjpQ19oZ/
QDrFMc9C0tZ2WrEC4be3SCjavrOajdPcnCzhfjmwLbPj3UuTKGXbzmG4lNROYZYMegJsbTmyw1e3
5QykOQXkEzqf4x6cKRH3BKUjTr+sV5ZUmBMNh0RuHXSIJH7E09rFlXW1BSmOqLlg+jK608J/w9fM
fleWmUUxsWTPDuvyYgPaJ2nTh+8DKtgBze4lUFRY/eX0r6wRVqUd7NQ0PxOtcAinO9FAtT0rC/T8
POiWZ7Muy8fB3hdQSQOM4RefqzKssV78ThmaikeLU5Gsyi0CvDbbR2ZhRDnNSIcQnbgJ/2YydCCD
Mn9lex+iBL9gE8sRHmVXBxzdTUcYGDwMAbVLjFQ8fYt9TsC98+fBbnuID40a3Sp8XZZDQ9tqx1mA
lnGeEAZP3qwUHCx1rvrAiiEuF/6Mlu0vmLsc7izKO/aBWYVdKGPRZWcaYfxCGIiQvnvfQ3njNl1v
8lDfAp0Ci03ygYocW4pht5dtaOgd7I8Vip4qA6Ejf7/EGFAH1G34nJhW57pW63cj8q543uzz0xW+
wYrJRo28QorPAd3x3aXM7RnS3C6TR5p6qAOleMjzepp16AQbEWjwthzD/Y3Sy4h8CUDbjFzFpqPi
I6ejR25F0X9lvJVWr3TN2Rt3ND9CD42F3R72AoMu6V/geE6QmSec3ofLIbGiRjel/F52HiatBYgo
5Xpq8/qD4BrLwLvYdq8svhxhJdQym7tpigd9HSPcbty9JgCaxZC/tpv9QtCkF9Jnc+cB2QohUiy3
ao6vdh4E7VcwTVv99IGYcyNDyiClaFseitw9gKZ0apADNZpXg/kefr/OJ+P5yR0Kh03yQsRAhgP0
WStVt2iNI8i+6vdYuD60Z/AmPdKUol/6aUJRK8G4iC+1PZR9hTwrQ1C3NthN+VVlighJkKlVroE9
P5RZwV8Qxp6oeQVZfVg5tikM8WD8/9/xYnv/AgIf0fhGBKnUjtNZmtsswmuqSSMTBL9JSsU9WU5W
pKxmJcXdtZwU5DfVzBhw0Zkn7W5/X4z3WP9qPoNlRsVLNNqc6VK7PDrndCw+zTAmjTpm4xEqkglY
c6gjj/6Ai2bIPj5jHJbdGshqnBTf0o0bp+dWZVZgs71eprupyeD5FKJWtq8l3TRm0GES6yXgjryV
PIxRRssT7ivgnOMQmp1vkFcpcicxppgjWjPXouETCPDW1oWZeMx+EeUAUsxDlxQJsXBwbtDau+9z
bJl5fCRAtswEL4nNdP5lRkpoDXzdDbdqfQ8NNOWbI0i9NAJDRTvIOokEAOe4KDVfKdEEbjTN1Qhn
5M9xoTRqszSXRoEuq2aUi8gVm+cXNOgygtZGw3sVhbJ20FuDfINkFCA7Uq8THRCP/0AOFjhzpXOv
Kqppsszktm9ZLi+Bkkc2GmZAGREVyq5NrfjM6v3UmsJw2DceQjKX4KhmyrWArCFUuYFFeRoofBKx
d//qvSfajruX8QH/JPjLCfgzFPSFIpBRu2pPa1W0EdFn6yQHDLino/1irP3axyyCxV7a9R+YtkJd
+uhpcTTtfVVWpidTSAM7/S+0/2bzTJgAqcW78k7w8XG6XmOoyZ5UuRJ6nb0yznT8gy8LH8OGB16F
zC4Hk3jwvOpLcNuETP1xmK0TKLVvnKEy4IWSufJ2A47n4LdUS05rAMyXFaWr1+EYjZMUa0EW5R8i
yg02C0BxsYqAP1q0sRDSNssFuh5/fdn/iqZleMWXQsj80h34TGHPYJzOq5ug8Y+yAfg/+Hcz1A5R
h6H/QdXAaRdWuCde0L6FDh/U115ENGvvMSRopiKIzrmOKp6I2rQ82O3KxOXPOsxvMs47qQsEqGOj
AEbTuehVKz1RbXXD90UMWktm15Ltb3wIT+UF5Mt9//nqNi+sxbfR5ADqIKmzDXxqGUpAKTGr+7Bw
nZGD0khfOQSYL+30w8yxQgEolwJg76eK5QqvYvpbg0jsVB0HS8mtvOdiyAE/Jusnq0Gqh36yckDJ
4o+QqINnV/jWLWx7MyKL7Kesj/VgQPFYh0byi6z/IAvTm8V3tWIL/QOvZCGcWDBPugkWtLk1oYNz
gkmMX3r0XW5RLWMBduLA9OLGEFaNoKgQACU9IQmvlGQgbX8TBX+BmOR8l/TEtQQarNgE/T4fXOXu
IYcDhJrR987b3bGlccqVivSj+XEqN5++niTr2gHm4kIO1o4/jbDc0H6/9+sTH1FzZAdWtDPb+tjM
fR7NHa5jN1HotTaxDYSCir7jYdriqANt1Td8Q5xD7gDChXexDtinHV1yYX0B7kkyzx0YU6AgL/Ug
zD2xW3dnAP0FrK2M+zTvSStpqfDDlRFqSLq0PhiL8FBJSqFbe76KdPZW8nbNPZnrZi6JFV8QUej9
MbbmDnJmN69NqTMCEyhYl0qqDdI5eGQi3xCe0Dl/VJXQP2hKxC6xXPTmwoChiBEvwxfQBdiye7OG
wLMa1stM8vxZsJPOi0QB9v8ClhmE6M3fl+PNwHhKp56LuWmBFDiiC+STllm5bk8b4TJ+KdU12yig
ZXCgiQ/eKAZ/Ylw7z0Wl2lATEHQgr4k4wd7uZYBwyNVEuUB6f3WEP+7p3/9FEL4jANtTkifLbUu7
uezwl5E0t+hA8dX2krPesh+8VjenY2QYs9O0MihlzIR6j9/ngQsdWfqKrRnLWO40K6mAxIDhw7VR
OKP9tCPlsjttTKKD1jX9fe9t80rlm5HL2QTn/8jj3u+tFra6iVky9yCEDGzbGECAKHHKlnfeU5bb
OnCZaHNHlQ8JpIvriXoaD8WKpZVepHyB6EJxZnENYrvo0AV7b+OG4Pa4YLQLHCIRib1kGhDPXh8d
AukTaKJxh/1YyM32/T4Et25s28FpZZ2XHjaOvV7r3hplr/5DdK9j0uhUwaqmsfJY4D9x0PaCXfel
0yYyzzM9lbv9kzQSnbH01K5Yqg9Sb9PDztYBL0UQ3EoUIJpgX8jzExMw5vGjBWE6CM9P2mYGGTHl
cWyYQb8TZyRIC9w2ALm+4l8kfKy9MuYoung9GtWyp5piDlhBdDghs9jIJegJUNmAgRoW+CdR43hs
ByiGQdn8cUfp83YrZC4Bzq3SxCMTM1PxIw/oiR+TAElxSc7yiKeqqsU2bMCfmkr47JfkiVNSfBEt
cOBtpUV4iWDh5exaWLrIZXA2o27jC4ZukhVzibjJPBtkkx4AHJ8/gx9YUXYq7US77P2x7cxaChRS
+8J6IeAEcxrt2JsJ7PLXxlLgpd1zo2OMDrHy1evk1o/jeMAy17KKB1JhG4wfKVomlDBJ2Shpzpgd
tjrZRtHfpr9TqJYVwM/v2pclrKqjvCf7RFwQewjow+2cIQg1/23cJTqjjZTgzYUb5QyIYmA0O7Ai
T+hha46rXpBq7h4Y5cH+SIS5qqWmZODK7impVLxQp+WqlEEbsZY+j+mORyt1thOQSbUnGmiVNleS
VzGVnEnVSnnKdN8b6s4LjD+zw7A+XJxYQQe0IBKMoQy3TYZsBnDEUGZYxjR3qnSyxGkug1AjwEem
1YOPSfmgiZFO1WeSu6aN7RKQiviqUFYTjlci3sA7DZUXRhFC/0SdQDcdP8dH7pdS1RjUxQDJFhaV
r1j+0PWYoJxQ0RGM+5giwe4mdK9de6E9Ev6nrGWGbxMNSXJrBAXjsF6XgYTo0nfdhHhsD/U/P8IE
VjHHIR1OTo/xTwmEdHx5HMoNyeFB2q9qHRX8RMjxVc05LJJa3h38n5VNuoMrh1wzcyoVTOgEERc0
yJoutwbhGjAeTJZn/06nrqJBACbep3ZoOAC7Zf1EIrfSon6cMOGNbX722+MXPC5cVcinXvONrTzd
10/Lhz9qPiyMSE+Hz+lHJYRTQZVQi4XLbmym9sHPpksS3f2BYi0v9jJ3CNJxRgYf/ud/j6UUWSTH
N8tE9mdmdb6X/qYOJCnkKtw16H49apaaLij+F3zt7pzQ/eMURrBUkgvIp8IYb5iAJTEIN1MZPSLZ
tNBFNG1yavOso7dSYKRiJtdzneiD/ZEM0nBZ2lkktHLo05F5pPW6M3n0lq+3VR1rjipc+GUhWIZV
0+lvetAb/FNeCbuxBzQH57QmsdFVFXtIOwCNUlWc5mj9AbocmWYNDcYWUqTsHl8yqggqKdg5g5hm
613S0nFWoRKJA+gxPpox43zpYIIkLPNe5aLsoXzkYjaRfW4gKl4Pce3urQyeSvD4HepQp67NxnHN
qwkPFWli2Np99bgDjcY2M9LAfR8LH3J1bQ48xI0iEqbetO/I6rh8LUWfkJRIi0oWsJCtHyQSzLfr
+dS0zzcLSjPh4KgKDUsO3hB1VjnQ2yjNy+IIVM6dWtU/hlOHWde+yKxgRDNxSvKu+ixXXjKJYL6D
dy5OnJLXepsUu7pqlHxDJ+6IYPHiw/tJkb+rJZDtJ5aBujsC9hhJ5GHWGNh2Pi2hNs4aZqJCk2Jz
c45KFOIXTMqRpSWCz63jOKroh+QgV9kHtop6sUY7/S+8qFoFmGDjvh6m6X41SLO66GrlKo/IyiF5
JTPLspxzVqfQKFF9mgR2j1zN4z4kRrTNAotCUP1g750ds3r3JL0fOYbw28zXA0gYUloAZFpp0j3N
bHDTOE2srO7T1NpcL5Sv32WTZl65pSIJ9/oGKqVM2MznbxX+faj6PkUnVVsCZEXYEZLEvDhtuGnO
dsP1JYtLPJHFZ9kHrp+LJ13B1lfDQs9HxyDsZ0v4u1WIYad/18nNTy0q/QXuO86GeeciL3UbF2AQ
17kG/6HUCxyYj6XadpDYTnw6HLS6jF0bg6JA0aPuYt58i7ZrAyDLIK13sHsbthL7rr2giBOWddxg
LANUniK3jSFn9VsOIhLZ2sfl3rHKuM16pFMQd2uKesVi3+PU+xWPk1kzvr6SQ4eU61HyCrAlNJxS
X3bEvUBXizzJ3u16e94LSIKTfQ1T1uJeFj6OSyWMHIG1447yVQj4G2HqoHiyKUF4mK0zc7sQpJg6
CVZJPfl7Uxvsy14mtbxqHoxHWkXYQPvt2tQuCTOmeNYAhjlv9knKtgR1V2HSbLQWm31SHx0Xtftd
nHJuF67XUrtQ4j3WUqbOXr0y40/tOWKeOZjQRC/gH8IAcLdd5c2ec2ezIDGaEdIk/s+MHWWk0ciR
2EZVElj79As/QZIAIh0Iag/fk8VOhu3QlO8/cvPxswPUwOcFHJOVFV1aPYuBtDUOMxaSQbsNRlbd
m8eB6bAwp0zq2mgXPrJZsjtOGrU+ODzOcVe6ZbqQV34t0j3jBpIIIQw1ckg0GMNDc8lgGjKqL+02
5BTGuM+Y0Df25UgcptTpmGKrLplkyhaQyktnQu+jbFvC12Aeytj55TijYpUu+6lPLGOOwLcv6j9z
+QPAbN0oIMHcSn9i0mJ0capBZAz+xU3nsBHUA8rpiivEy+YayTAkdjn29nZoelzbkSHgJfqOIusY
Wg+t2YmMF4h0m2JWIeBKQlFu6a3KkiSAnYAPqIwAJ5b/FwSW8zhi1FDWAnarDjPoghpI3hzBlcAq
io9tUx9j8DfKyLT6PTWtAhAAWT2lRxSMPdVc8h2MILv3e7mksrSUWtQQXgeokxcEiExXAzWttNNX
2TI140XtLh5Tw9wEcOEvalQOabjukYKJ+wQfDUEUv7aM8j1YUxLbjJ89dMuJZY/1yHITPj8N23wj
SrobwTSlrfkMOqOGwWq/I/5e4n3tfgpSvB27fmxehDFpGPUtELTvjJaGnDGYP9EM+4OT2SVJnzVH
hi737niScMfUygJW00lTLEkmqsk7a1ak9CIE8CP3L+R+VoGQlkBQssqKBObbQIr7e8kSvoSsnZ2a
5XpaouqeZ/BLQTqZM4VW6aBjF4z19lNut1ScXEHn2bujq2nx6BuiXsYTDwH5TKse2zWebJhl5cxf
Fxz7dAnEgijnQ7iVj/P+IdYncQ7h7hj0C4K0mZA6WxDMwxiKXTIoKYftBZmLSY+/JRbQAq62UYbw
OnXEbmpKkqNCzB/LVvvE4OxCALLsaUD9Pzb6Cq4fnTFrB/Xj9m1r2q+N7B1rSqNgkIP53Ft9NdCi
hDgNu4UbLPmakPOU7uaRRiJTaJlcv/zrA5oM8OAZhPypO3fVaI+0DcgtQ8ugDbitgFDmijRHl1nv
9PiRnCnE0gac7lRPzLexc5cfVD0CwwL43XbGFKc0ZepNJMb32TMFHrFopNHwZeh7/+/WyFrc+DZ3
27JdUSo/B8l04SYF7SeA1NPJ+vjzt1uCWFvFowivQr+8CJyy5+MUdJbaDGr+SDjCVL08bd3h3vs0
vfhs5b6k8dKkRToiKVKAe5HdMWONyFcPspdo/VWCWnqU/DRwGrlVIm7QSK/JYXxL3eJSSv9T0in4
RrHBUw2w17fzHk5UcaF2w79d2Csi+fDQrZhZFGpwB3lm/KqPo7wNpn0weH0tniSn4oPn+HFGd/WT
m6Ywnc+BarxkdwypUR7Qs3QlmvMdnSCluNVZ18x/kPDfilH748tvVXcPArp63rElu4bzPWRgoTMc
W1IMupw5+DBoQhlJJP4LfkYe7/j7DIkb0zVmnQXL//cDg9v1bi1egtYqr8WdagKm+5cR8c8XGwpD
iluOWWnyC4UTbFnvNe+2L4e/Qo7z5b5tpujkhuXVUa77tWyXbSTZtX6XUQQgcjM/2aPjmNW5ptg2
AM5c6bcSROlSA0fBbE24O2p20Y+YFSVwz9CXX4rp76p6Gzu0dsfFc5U4e9dAIvMxspidKFxDbI3n
20keO0AguRhMb1rPSzwzVgzrKifG0IxsTIGf9NQha2lZBQEvD4gHfKPL2ycZiOZjq/GlVTQt4Xg9
6QLOassJFD8l8kcRMFVgKEQODwAdNMnTL6sBoPyUCSMCU2+7anKO8GP+LmjgyiLd98LqGJEEMSLq
N0938xz/BZv4ZHqw4SCFceI+C0XUFHmAnr99dMEfpGyIdp90/g4bTQzjh7DHV2EEC7dim6PsyDPA
p23GIz2ZoLFDLO6BmxnfBSktR2mgQTc/QVlUu3VhHPAeqUwVeLd8WF4DTqE40uCXr9TZ3JlZJm/e
0L1lT/EqMrQ3KW0KapDHAjYyyPPCi3AuXQHS2wWhfJTl7REAi+px2bKY2KUGkC4hz5GpJjWWbutW
68cztBEt0sDA6NBR3qNMZUry/jn7YDIzzm7w07x7x6qE0wjcEGUXpZY921oNQZumzju+bQMNZLCd
UYo0rv494DAQJWple5HLosldTHzCkfrnTokEhHzkg8PCtwMgpFouVufvQzg3yiwaNzaT4ToJWIa3
rcojllhB6V3UaOTx48TEGcTeETaKrJ+mUF/dCQHGzgofgQ/VH+2dpL0rqOUbREAdFtamHmCkta6p
F+lBWfZJGL48XcIq67uGUotX+WlpGW0LDvOlMDtwoJcW6eve+JvX+/ZpX+Ba7bG0XFNeR379WyOw
Apjwbqrs8kaTRz/W4weDp3q4jza1BT3EkZXFBzSlnLVvMI79gEsVZXM8/Zy5Soz94lvA4q1rYa0D
oRJacgfc0QtU/HaTLwMdmeUY58ThpJptnQ1qNs75aRmH+M+1eC3Os12NjYsGwhQ3WJHEyNqlihU0
Z+Un9HOL3n/CDuu++Uo143U9uqEduGoua0PqKOknw74coGY4RYbHv5DegdIo7lRgezX4HgBEy5Y1
C8n62MJFYkmMqODO/o2tjoVVInWuvah2LY5jQ974UqmIE57MCIDqinxA71Y4iWCU9++dK1yD/7dm
e1+SU5ZwMYMknsywyMPAp06fnyFYP6xmRwUpU9c0SvR5KwFpZ0K8MycNfrEMdE5QFTR/sHnuwt/n
b937fKuTwwt+DesyxSZgHtsY4mQO9r3C7TibEdSd0MlN5iDgR3khnjCfdj6M+kc0PRCxUr0oilxD
lI99hvgqa5hg0JP6bHx/rXMBMhn5iGp9ySie9xwOLCe3JIuKIJTbfTPhXZMHDKdQIgJzisIIQGjW
8mwiSygr6QIJi83FcCHzL8ymhL/udtCxOaqdGEg5s56dz37Uinh8S/9JyU0ZedH+LToOgB4S7Lyq
OhKPuAa7SUEsmpc1DiNWULz43vc5cUGlu9FaWZNXntxuEOWoqa/5sSTFFy9AHwwJYeBDzsEYcPkx
LMQEI4t+sfTqyTYpweptBFQql1RDEs6c8JQkCje8wnSdp2x2pHCT5Wl6gG+NnK9vFVZhwl6F6It8
Q77O5MohuV/0O08q0mjIlUyJpMecrIyo6qAyE8p05jJInLvc8LCnmbCq9paUrhWrU2ukRPcVYJvO
tf0iigfSMNKDL4WzK5I5zQcRjOr6MsSVoywOTIg4SYSP+DF9SzUHMGw2Xt5xNOqU8czeK4xP/ryg
5CG4WWJ/Bw9JKctC/M/++OK8FHEowIsiQjS7uk8ANUn5YC+vEfRNP2Lce3aGq6w0S/nwDA3fzjTD
l4PZFCwlqEj/L+9RDIaXtF+rzy5kCl92D/u1iVI6jLUXOi+zHvKuXNH09cUlRd+MgV4AhFVnQFDK
HgGS8Nz6/rhgLFSLnDjNAkAC/9CSYOgtn9++Ck8gazP7c8MlWtOm3CcMxGuU2u2Huf+mNHN0SrcR
SEBRsKtuEdGyad5ehBHUQ+Uxw0SrMAR853YLEk1BMMRQ/7/r4eUdW76ZomrctHf8XESiYIOtMoOQ
+o+JIp15p0E/OrsKEjECb7F0ZPlWwDO/hgx0WFNgp7ai8vqtBsgM33DxVMCIFjcaPXSOJZZLbF+X
Zzkc6Urpvmln12+7pJj362I92DblV9Jzt9SOHh6FscjIpb1iORzo09sMLnZL2GIWUJhNzGL8fGx9
+Rs4g8rbJ0PRUH4PkMxag9j7Ee7dXGAy0qhhURfLQBhayDbLQFt8A2UEIwFVVPCK29CiyX/pyJgP
qFnbTtY5npkyYtgMadpTJFRvBZjMe/65mopEyJMcjL/9iSxqMg0JP68doS7jK1rxAYDRuWL63n1T
F1PIYb+AqJ6XbJpHprnkpg6bDe9m0LTXa5csckMGxEiQz2slm7UDR1RkckQLQTQZDeG3sPvA/hiA
xhUShXUt0HuCWC6e7Wr3HhMvMy5n193ndFWpCxOSICav/AQ+G+7pMhXTyv4F0nXChSDZnO3/T/zK
WBTiqBy3Mlrou4MIealtlcrtNLOrwYfALl/lqOUCW0ULUix1kbSoVGcbOqdaFv5CIALTSnToziyj
3H/zh3sU2kgLAQRpjt+wsEBaoYno5ZsnvvNzgoKMIBh14aSQdZ2A1/WeJxFw4Ky+1oWLCAWN3d5X
4/ZDrgbcKecZHyxCbYFDAEl/4NteEMMECVo2a+IxMMszoLKCICmvUhBFUDSNk6Ag8dORqpNjzr7K
ffY2ehj5sOrzEGPZv2tzWTy9U4rbYute3DYuRCoUl/iJ2BvjNEh4ZHKY+swQzmhuzkFE3XpAZ+U9
hQT4Nxuke0zY6PbjPFhe1qBB67cA8HpwvImNHEs+BobPFx3/vLj2K6UG1yoetsZ/AUIwBWYPkc+y
dJcmPi9mqzCDxcOd578pKmohq5ndOrIqFa1xgzvZO3+fKezzUEeRFWGhmEHjRD0cCFbQHNd8CTgE
v/zJQ2sBtR/cE8hhACwDp91U76U2Xp4IJ+Kq9ikm7FIVfmpc1IJzV7w7d6iiWsYOsEFbdY4ZSOZA
oywk6RpBtybi0eu+cnv+aA3hLl+RX0fa45LAcbt/yTrwf65jI34om0/Y0Cpq2jrIIyeigKRwE5rk
BghkiAh3HwQAKiLL7aJFSjJtleEs5SsoDanwXnxBSUtCGXNFHYRqyAxyRqW8DyTFzQ59CqT9dVPj
7/H20l6QAPUZozXGDD+lDGRYsRLAm//zebzY3fh5knqlDkkx8cifo9T2yUvQxXBmx+E6W/cMOY7S
VZemjVWyZLUqQ5FFz3grdKoDwP5gdc1pjUwdbWiInLgULoAlVNNvPEreQ0QQRX5jRK2VFeynyBkq
sYhNiiYzURfSN23mX1VzicTkJ4xBqRJqngr70wT+Q7xXHy3+ko4T2EV2W4f7eCHzOftg6TrAFMl7
UgCyIqpESNwmisP8rSse0W/8XoqBU7yb+s/7Oo73bmm8zHG7XJwD16PZKr1HfEr4pX75u0dhW6O1
EXvWPdXYjAEyZcw2NR5wr00/kvVH8zMvI9BrFJBM+3zWino9EbYKlqcBFUxKvDMeQ7rel2LMd8Yg
ASUJaIdO6uw7s4ULP51YVav2aGAmSpamLU++j2MPF3ZibyL2S+ZPPp3vWIh0qvrKPze2x90WREm8
IASoJnrq2FfEN+1E2bTPZPozsMZstOzmM8LhMb/kO8rkeUfj5K0KUymliNga0mVd2uxy5uRzbOpx
f3IpbYRtcwG8kwVNcoHTBX5lhHp7i6klJBAL0LVoLKtgoBUfIw6sDqYGyE0isuSTiiN8xDqECYnG
RFAEDhNVc6L1Dom+DNxnD5l3VhujMwXR2Ifdnsl58UErsSanBv/l/gQwNQo9PlEENL2NpxaXq/pR
h0ZxtSVTbJv/NrBnv74WB6xZi0N6jj8s/RbZ1kqEJ9iylB4nQdGi/oq4RgCGp0HrhOv4R6Z1y5QD
inh6FCi0aVuDS18/3X9Ix3PkIVaRGDoIZ8pOAWj3dptwJVHkfRj/biRQFDb82oRDjg7aS/uNdKQ1
iLHCzjwexggkMRZlxzt/nPQY5CabvrDevPWVF+D85gt3eE7GrhhYvZuyPY2TLT/PhpzK6H4LYdeS
XLyn6DNYWsQ8bCCY1NqXhpPAwm1rHQNMKiDLT2rTE4gS0TQAFDFP5rz70pcZXVa37vNc6G94Tlqs
DEsZ+qMO09cE7nbhziKXUuW889XSgk5X385H65dmGaB+bP7ngXT7Bdg+QaNzF+z/MXpBzVZcnCPy
kkuuRWFlfW+/Sub8UKLVSsnkDTFNaiu+81XbC4tgoo36WbCRwLlVQ97xJTDdGi8Y6kgdQd0GORDR
YiUxCfSm47Bx/6qn9tb46Bh4oDxYkEhfAfFShGIYvzfeveWKOTZhWX/6oYKKkBRZnSr0utRZyCU4
FNHItRoB1+7ib8voQQAk4vnem0nI/sNU1XXsGaZCnk4hJQvCq/lM6IKWskfAGuNcllVpRR5YhTyj
zEey+RbgL44BPGjdGENxS1Xb8Qemo5fGIVo+YOpGoLu1Gseub87CwSjrlEB8haYS0UfNG5xDVRzf
x7NI/w/89L1CxlGcAvGNAv1L+HZZxsmWLumpVfr74ljLMi8uiH/uEjNAnRQ2YhQ7iq1vRd6XgKSY
jMumPlO4C3bdEdLZ97Ffpu56U8UsBLTFB1jGav27Tq4b+RrIhkNNYD7LMuiqPiEUtI4xzftgC4Ta
51vlT+ezj9sbRQUmNXi89NdKKG3Q9gPnFfkBWf8J+ozgmTVuDJU71R/dPm5dxOulWfKTDD7LqRWl
7yezB8KHy5uA+V1F4F6sIWx0jB7nJblX7lIbDbIt3Q8IgmbEPIa5gTWeDEf922+k8aXBXc7cNR+q
B4nFtX8yhKZkM4zF0cQobCQGW+4aAGyYK5369Jx/sIIh8ZsbTgQ7YteZZaSScQdRARaq5vxVfgN5
zBDsdYJ/xkbw/9D6sZZaHjzqYMepkIjTdZoR4kSJzMUoI3TzQAKCEi0dVAqdJ8mYLwUhIph2B6Y1
GC6lrMGHdTNCQEuF8btwPrU5ithgYCIKE+wHieINPuVSOk32o1D3gXez/vsJXAfyQrLLYwWiRV3C
IYuH5ZwXqq4olh0Nl3QpQV+93EAv3jMBHzbc5CCDvsRac5HCg7wby+FzUiORK8jIm/IfTo544Yv/
mCzwE5LScBUDe1W4/fkc1rk4iR+AYjyp+PN5riGex9VDTzaFkAmupTzhy21ux0QfuA4K7LbAzTde
m0KO7nlrMXVSjRBpJPYB+CQAqcS+P5NbsR5H8RLDke90oHEhM/MAFln0pj837zcGsMCBHc0C9oDl
f3f1luByEiHi+bemT0Jy3qlCCbwNAok7hJlI7duW3l/Ui453ELzEGOvNkcrguC3on4VVHcCYdaL/
iNBXbiWvWMDkqLXlCBROHv6Xb18l9QS3JhNtDQISUFJgZQRkY6D0hZhsaG0yWuF5+VDWdqTFfDZ2
08Euzi5xaLqlLr9Ly/fSqGMBn6aFdpomMeJIPoIAqgoZXZANdVY/DAhxnZMlGU3wxYQfJm0A4/jQ
ASxM7qi3Kgv8z5JEoYiv0G8FSzqkaEGoqcJhXVW1hvlyJ6OZDYhNH2BX9z0ZSgi4r3xVdC9rQjF5
9ZXUwKSWelqDp8yk9m8OUaYVAl8Ptah91H3lRVbeWqPBOlHuRnTUxmmP2Ns8KGFTtGXtmgC6FsD2
EfiQZVKBwaebFZJ2dNph/W3cOpH1WfnJV45l+suPb8FUaP6msQh8zFHuIikmZh30Xl+gAa+5l66I
BC05quYyC2l7nMup96VwbLxQGtetPFSLko9d4gRsoDeq2VBeymgfmt6AGUFnU1z72SURfd/CUgSG
rGTT6oI18tpcvWIe0AjE/F9jHJAw1ZE3d/QWk/98iqgjvQbtrhm4b51W3ftLC/abI5n1bBdXr6/Q
sHKsaDkD9n+dAjN7Kqf7nkn4inoVFNtMYpid0g+QRcB0GhNv1Jg7Zd4yI65ig+iIDkA9XzyP+SMh
2MBk6rKCPtUEedPCOpcSCSoJ7ykQkCF6IpKaJ5a5XcZgaZcfYqpMy91whgCDKnIOr1aKWOZvV7NH
MCUjX4As4UagWZDcLAjJVWa/t7G2bjsiC09VISsPMhjnF8R3N+lv4KIbW83YO1YDUYeuNEXh8g8y
8Z+DsmibLJu/R0gRZWdQoAvBu04hBLLR++vIa6IQhfSt0YbouGE4KdaVRTGa/bzvoKjlN3Wg3bhC
K3kL5ZaiRsSzooBWVdYFFonXKEmNvPcEmt8OKqjG6PFuvD0OfwYfh18tRXfj2e/TLqsS5eHTfHik
8XSUGV7N+0sA/vcH/c50MFm16k+AYoYFvvnRq0vS/fTOlMP6u0RettPMNE4aQZ83UfAeZR17dJ9s
TqAqaHxonkJi66a9fWlhbMcy7rvZNZGkeNvd8LMKXxGLfqUyO6Dqpy7ksuHJVq81ONtqvFQbq7wm
QYfSgK2RcS4VwKhWG+friGCtcKBqK8R6s4dXBPeQdPBCpD22B2twqi9pJHWebUE6AklHpFkVO4Sr
IHYMzSw72GF7Tk3QJ6vzjjZ3GXF65bG68MuyzJIzIQwT3Se1cgTiFOe6papQtnoJmI1NqvQBuSZl
a0mABZJkGC/3alcRF19wEFqOnXAaI4BvZL4F1VOPNEJfV62z7hrP+3VYR/0xPauurrd6pXYIwuev
5aS4ts75qHyM7D1rGd8aEOxcsANjxNv8oZ0cOm7HWa7WNr5+jN6oSQh+2JkXe1JWm8YkKpD/bBPY
bvCDEjzii3OIt9g4HmCCmwiFtmazHa3W+cWSmRLNYxzJeA+xJr+SKxyAVOiPD/g8GmT2naxexxnY
8VvmxA6s/k/42wmm/4rxHztxGVS+ZnwHhoJru4mYzQTWKUkOGkypmxGfxfga/ZGtpe1fgJm74mg3
XZd1UfgdQAWC1sVPbUH7oI8XkuvAbL0wnjoeRGZL2AUwMxfKUPcnc0QOJ/qZs2/h+oq33L1vLF+3
nFwP4cHs238KsmdG7YdnbdBiur54etflggmZ1vL1CF8znc/cd6hE/iuB/vy6B6djnN0ru8sPoBGf
Hv71pV3ObTWiY+Hks3B83P7qdODULjjoDWBI9b+s1gzgNpa8YMDjAmrD0v/wfsfnSditN0TVTwBe
j8Y9dQdqk71MSD5Y7dysIMFHGbT2zhqL56jOn16UDQKJcFQvFvH3Fo8STHegc/lwei/qO08qV0tU
sTt8DwCsSOjwr682gPkmVSHhF4BzZmwMpiYLLWVtndxHNmeWKcsCwC6N8+HoKTp8P7CrKgBCGeJ+
opIFt0wSveESQ0hqHEW/dogiKgzyoLHk9Xph3mYA7IkgUe2+wBQd6lVH2h3fOC+apNbx8wt23UvU
WQMVKALzJexrg4FDv9OjSYXwmbOiowTV+KybjIkRey5loTbnl68umKwxcjOf715/KG8zaXUPtQiO
xAbo1RPXe08+hzF0XG9u43WSq+uy8/mtj2xFrOrWlT7IVJ5t/1PhAGfd2FHR+cDzN/nNIeGlDc4U
vfYOM5E7cjahn0u8qoUCmEL5A2IRGnWrMj7wVnxsJISbYfGsE6p1Nw661GZyVqG/XkuDCmFKZtIy
nCT/F79oYEGlem820vJODBAaaPkOMgiueu3sOGUuap7RSo0mrndemzTOAfcqiAMvmv4l4a2yvqM9
nrRzGTPM3wsdhyVeudLCi3wR62cFbxweZnhb6l9+xlA9iXVEXjMzSYGJbopxCrqdMd03FbwtUMkG
ZCuW4cNeK6fyLJumsySq3zmLfhgVHwvwVdCqVsPlOyitUr0BwGB9vSk3t13k5NrWNKYJnMSMi192
+J168FTcvEbALkME/haz/dOUwL4czg7SKhqUBo8HdFuos0Oqz4yZ0h1GHXgC4NdH9XpxSgvTx/3K
ov80fZcx/Rsscsas1ZWgirt9gPdKPaUFl3OrwUk3DNf16eb4kdW7da6Gjl4G09KmefNv/hJ3YoA5
I97L5jEGE8YsDo1xaijs/H8T2J1PoJ9Up2NnytqkZO1MgOZikftEMsUkdQqo49jRvSHT2qUivl3W
3oeyOYytejqIOFqISGYhtPzltYrRWmyZJ04Lpk4q0FvFA+amF9m3om6y5l/kiGszp3FewnVe6Udu
5ZpIMZDzEtCqIXc/KDtxY03+9Mf1Kx5WvJXO4r5zp5Df5xSTaQ87Raw2+xwvLsV5wKWAvbzQd3oc
TROya49BzLJRGXg86jC+djrjDYtYCbpLj55KFD2ruMqP5eCxkQCHVBNwn4ITlcTq+5HH/0wk3aij
X9T9mFSRIU7wd7QiY/YAVH77yWkAwjJA5SfsTs8134z30o9Bk7OEBnlAAPvYc9aP2nBossToK/2T
XUetNGrGdyxDrkOzrnpaMv3fCKnf6QxXgkUfdzdjbru6SPcROta+QhmUZuxqVi9Cus6JNHo97Wj6
ycWL98W5UL4Dsmp+3K1YdBvalkwy8AcKqhe6cxAoi0x0OZakBAuvwR3dRIwv6jCG/ieWOa3Xk1Jy
tCfUVBm48r/G6+VOoTmWhmyobLOT5JYHn9dRE/nlZuj72JsvYYHcknxA2xQXT+8+4BVh/vZU0EhJ
ka92zGUttNoU0EmRpav3QUEeiPJN83CrgIaXc6E9vqOtY960M+BV2Tm0gKRs3Ljqbsx3JgasaCvL
A0a6EgCf5izxnqi5VzvOXQm5upZAKlz+K+bzHfoKuIkSdI5V9eDM7H56WevWZobsGUY2Jq4exGEF
sGSRFoAeJmNXN36NKavqxGqTClNoTt/jGHpOkxzJQPuRekM+5MB+UyMaK0NnHG9Ff7TWdY92OjlL
wHqWS60YKLGt7zxbqskLgH4zjE1x+gA89O25Y3SYc5wRBJ8WRxapC3DpgCxDUMBn70kLGmp/6WjL
arhUp+da4OySaTieA1tDKLJnM45MNq/wXhG2P0DfDIBoqaV0Tz6Nv0pXGmhkyc1RxqzVtZu7GeIK
jaXdEPb3VWB+gARTCfa0bKw1cupSyAwvfBDop2gdPSvLCh9JFGdBkQO6hpNYyukOQ3I6JJBMquqQ
V8XeQ6GaXYgyXlg1qHikqi+Vjj7zkHbJXE4frcq8Jf22TumJFzUpC/oKUC+LXHkimyab5osAWG+G
TzTyEUAbrAARXuDFc42+QlcgeFYp9QVwV5wx0puiJTqgd9os1NjmzUxgKXE/jXBVzEbiE2sZY1s0
+jE1qdB7WEcGDNz8SK0+cml6AMlCGFDelcXkxEUnS+BAnp9XPrQ+PenUYZl9A+cEBoTH6FhoBaiN
0zsH1Wa5YicdsH3hF1ovUIpXZHQwEEwqylrFWqfkfLx9C2MiMgr+UklHfRHG4YuCvkDNQZiR1FfE
DqOOPJBRnTT+hGJFcrs8u22sfYXFszWLoDmNRa3TBfqOIdwnbXXfhEeofPyXO2oHhJlI5svMg5M0
N24QvY8nL1EtSMR2mfIL+UEp0IlRd2fwA3z8cvynyal1HtEI2KryIYno5XIzQ/dTTTWsX2Tsrqaa
ysE4gpOy8SPzbuZ9g65+w5bCDKpO9chKWn3XOp1QsMItjefmD4/AM9VbowqMaKE+6mugPNkxeZtB
sj2s4z8KCdZEXxSP4fqSl/uqcgxzJ72vctag6CSru6sds4nZGIp9UA6b/BGXHu9jVLKPM30wZIf4
ljvsMp+d0KhEKM9meB/rA05Bb5jmBKaX2kzshd6J5oq/445qsElvoaMUt/2E23WLtjgFbtzVPPGC
WAIHiiwBg43fTu1sJDJjyb20562eDw82ciyaTfxIXzUMnwlzzkCNWxKqjimt/u2Qo2nMGUrxGvXE
5eH70wLwtCvTgs/DozED7hsn4qcKJ/s9QpHqgyTJWmKO7jZg9+XveMFslJUVS35KvNHAP0tW69FW
MPDASpc4rqtMd3qxgr7pbHXDuJel4D53LI65VnvgaHKv5t/ohrJ12VafO3JL6P7lczCa9ep+AGc3
FpxXWC5zwLtJbBb+5Q3z8ZUy+hstoBw9+oJjshsD/1DdZnfRroLbt7YcwNBvuoBT9xKCS2Ex2r6t
6iOQHjhI8uaenGBEGABodkkQUn4UiVSgl4BAz64tgtBRXlWoSJ30fTOzssa65WjPTU0P3FKIKe2+
J6klEKp7gLp0NYsMshpdk4zgnp5DFK5kUvSfTJsIu6xq1yHMJuy64fjwIbiaFr2MrDH8jRIyJUPK
UVRVwKySV6Q7vrJfvB2Q3OSDTVvo2bRWCAOvW8Fh/cQmpMOKrfCkOAURzCyXvcKtXMypbmzFWTew
26gozu6WJ9rLJEq8AtJr3TVKLYIYPHUHinL1VAjfof/D+wtCS3XXynbSO98PP8oF68JnzOU1r5eg
vPO0lNHA3BGP0mC9p1h1tWt/zGxehzTM0Te4a9vuizCeQflBBKXtoppq5qRT5w2M/p+U68oyMjEM
aeO3gSDJAHDbhCUvX2HcM74e1ROcN47L8YkhaYpVPFGthnZN8D3zcKRqGLfsqgIbFjLaM/oMF+S/
egbIOoXazeRkrGkuQSZ+vdv9q7IXqF28EtxqH2pZDv6ktP8n1WQIwBfjlk413XbxuZRbVRaa3G9Z
q3dG3WaEWZCONcOCoGItzHFetsQg4bf9mEguiCTttVUHRuHef3OMdYiuv0mkaOED5aqkZG7rZxQ/
NR0EJt0HGZdrfk/TfgBRlPgyURqHbEw85M2hDjLY1KATxNq4TO4bs3wgPPEjSqOKPDrf3MGI0dx9
1fmflNKwQIkXjXsQURR8/QuK9YX4U34OAHHd4KZYHdvPRNk1OCEooQEOAPnGBvUactHI+8w7RnEq
8rNKwA2Tqi7drDqKliDwW8lO8KrojyAztXaeysiLlNGmSEnZnpzKbuXk8JBDtA+cf3SCwSiSXQDz
orGDITYO/doO7DXw8OMucFGiVrvAHc6awU5/9rPD2YJah+Ou5ulzegSb7qB5Cw5cc5V4XIZHUYYw
GpFzvZIoOv5Cg/oaKnkbZM8ufz9PEjJda/KvUnFpKAoR+2fCFSnQm2MH7izs9ZIuqYTuriEg9trP
vB33jgNqfwo1yFAwa1Wc15Lf9TJwbGOsBrY53ynKlxUc1IijKl1BHyszUAAD10h3IcMpmuRotE1E
L7Gxq3mVhN2E8WLtY8nHtI8lSzHZGerRqSp2wNz7TcaKHs/nEyzWgM4HPl9BCVJvEd7YqGgvS+Tu
E5C8HFvU8UgWS0pyKBu25gJPWp0qLRBBoMWOjgD8Asv9noQ2YaFct+oHPryEmckH/+cKSWyXei18
RptQ3ApsBJe/L9JlTGx6fDlxITBz4MCE/yIDFD1AwRBh5UucD/Li+ElGNyLuk7/92xr9ayfR2nyJ
p52Bx8koQyHOWYj/lCw2TPytVaNWT/Fpt8gjeVvGdU7/oYJKffQI65/Xhfqe/qIG6/kv3LAznUMk
YD6GmYqk6vWmIa0D9fKqm8GQtskQFP4hVVkwikiF0Vx5ZIwYvDP11+NOBp717Dfme9IPBu8GLE9d
QsUPSGjR240iFo0fR22McNpxDo3GX98blSjzUrBEcwNtfmiCWrOIHTmwCLZ1yoLURcvf3DEfkZjm
GdSAoR15JvAkrSG2zqcTrULOCMSSMHsgyXKzBsLcVhAXeEtU2PpIr1RioKu623Ey3++sbdKUe1Rq
0PPq4HcKTcex+WqZtpoGW247nTQt4mjRogCLiKbeKo9BDmwTMsQjE4R7pIYKvpXvzPOcq8YShOtI
hKuIpA8OlKkCjjin6o1tAkhSsDl7hqrjoV9fznAFhhjGnx/S0k/HLvcryV3m6n4Nyi0U9MHXPng8
MuxutafzYRFbaMiD1AtzDdzU8pgr6ZQBjfrCZ6SE4Yf8xKGRQAHyVw0kNMZqnYdWugfw34g7C1H5
8Od3KOonmENupIGtwXZBaQ8sadTQmycsQ+3wlCrImGzFd+WW2LEkToS7gg99EzV28Ir28iPUKhO3
7fXhbWP80w4R9aTekP15kK6RrDbgW4nu3Zy1Y+YkxmOj7HncMwSxN0g8zFd492BSuUzpX11wlozk
O+wbO7F6NSFF9tQ8RsDmkRrozmmNMyu/Cx4Url505Av7rnLxQ3ZW5iGkai4XcyCvMycYHRQYI59P
Gtvd54LZmTX6LXpDu9M1Irpbz2KjiN4NmyTBpFGB8XNnbUJmlNGhujeZGCqXi64dOa6zh825djar
SegHVLOx6wpSTH9Yzq9bkL4fs3/PJ9x/8INT/Utj7hBY/o4DMWPuwhdnFoneZbgu7amGBeur11eV
d2DgUMEzIroo2DpKKccoBB8klIwgAX/pPflZRY7JoqtVzfaiMTdzPJqKWtpptrqFBfy3maw5PSuV
jjBrHX+s2tc08zK6lzALMdzeSmnqHs8ZuZul2pW3CiU6W9Dpb5CrEUy4pT//01S1Vm/O6TDepy7x
Jx/ihZ8471frT5yRQ0TPwUW9dqLReEn4zAHFa7Y9d41PXJxzwxEZpPDz7ZlR/lrfHvXK940cG2Bb
0IKLF+3JoKxipfQv8hdroKnyr231zsij5Bim60IU+ZzgM4Z4NJZDkrkw8PjewVksUkq5wSq+3Mq6
3xAugAIYP8yB2dgroX5JAighUGcvGnTCc5zlmpMpCmf4no3LPJ3gAhUsZJ+roY5VBFnbf7xseRM0
Ez6ZWGtsx5UiyBXv4JpT+fZkhfP/Z61dC10L9Vm9+syQWKu7eV4OWPRW22Jg3vGgqiIFfNz67/Oj
/DP6nDAVRgcNk2nXnqZMXxQNaGuFWd1g48XCtqbtvKZkv5d75WV26gdauuFu6KKiqkYxH4BfBYfT
Q2+soeQ7A1lS6w42A931EEXL8Fw9xXLVIAQ8hpl+0EWSjrz5HhYvWk4vsFiSIq58AbRy78zCRgW2
QTMh/bP76tYrVLh2Vsrd/K83pzc0NTMDFuC11FM3D6CPMyAGUEk8TJLqw9gEDclZIOBk/IZ1GOSF
Cai56eEzcjsQACmJw8W/t9OM5fvmUh+JEMtDrspbjTxWP2FfPH45auJzSqSgY+4FN6W3LcD4C9yz
sfIWBS75iMNa1/0iwRN8DsStEBlUUHfUfYqmRokhpM4AEFhDVmiVmKavsB6rJY9TmAL14r0oezSM
8i+IC68gcuJ1KwjUWWjoL0uZozvpqd8yG3VErVG+kpEvgcFy1+AOQyZvYvOQ/ErScY4CitZWKZ0H
H/mN7+JM1FqoFKEgOgYXc6nAQ6H/nmfPH0yR7/Qthf0+d1fwBA86L1PKGDuAPiOhSSGebtHJyhIU
VzWoH7Ycacj0HUJckI+o0ZfoXlzzmI2XrKI3UOfl8rPYgpIg3ETjX295jL8SnqTKk72DVsKqSESl
p0biwuIC+cvW7WqqxY+7AC0XJE/9ePGfERWNEU1UZmKirG9M9WAeyU8jTjgFtxY9cczQce7y/JSk
gruL9cwDq1dNETymVzag3ImXoh9PxlrLSUeoFJEKmXNMirIGuRvvf0htOm6X8//Oft+eTnso/iEj
CHHxMMcVaH32GmhHxq25QcVDKj3n4gsUV4h6WEWhsldLNtvxUVNE76vMp3N3DEeG28riWdh0MUdV
lVfgU7HKU3h556DfKkg2wWiaaziPmsxVJ7HYuYQCtzf7rLuqBM3siXjR6vxWa1pmhzldfhbuyVHG
UF6Fkwx+HHinqmd8Wx7gk+8Aewt8JflEkl05Ecv7uOdYxMoaH8qY6fjOBIBtMi+a1GqfeABjJloK
8koZNSofVo5TwpaqwSKNFigoo6dwIg6UwyB/vcvuw9sX3bcMutT6wr4oYndwjTubZvJgdm8+Kx3c
Mb2R+U5uQoLP5zRo9i+0yorMjuJW4dsuzdz1i+pgHN09tBgm8vJU+Vnns+bSNuTwS/NNBibBb7KE
IPTae5jsn0fSCLXEpD/moFwG/ayzYSADKwbQJEndASwGklCk5zpr5bQxTsxRrcK0FLAVjeW0TKh2
Zn2yxy1IRwfy57WGtzYyVUSfmCvt2XSWHj4Kmm1v+6N3RCsqNpzHNsRByS49Uwiml71t2Ae1Xk0x
8ngqEPxT5IsaxOwJA1CthJoXPxStaigKdBPYvN4tOtoArxowLnJe66W7LNEG4PWgqtD4gZV4r7LC
lXRuAsCqsOvc7hceJnkeNYp1C6c9b/aEN1KuRwIC8eiMBe+77lJP6m7h0Cww+v3MULmhAemyTZK/
GDqZ2QDiE20xC0ttbW0fXWimI6/kx2A3T/az/Tgrqidt2tMw++corlCQXLwJWDK31NpTvLT7oV9+
PVsLaHZrUcYki2ex5iOJP7wtYORm7sUKMMDAuQ7654v2VSLpPFhIwG4z6xWHP2RiC5LosIWO3QzV
7Hkb7q8Z9ArfitKt5/HVyNS/4eOBeGzMBqNS+dVTJmJ8Us0YKuYSpktp24QRpbMyX9xzp3uJXczY
cJyCCoH9ex08E2VvG6wipXgV7ST3vP+Ji41ixVOJTjB1XhsaPW/t66UB3Z/ef4qOREqFROtcJI3O
8TUViAgkIsXwvBmfIL4raiD3lafuZiHB1KPnc64nLn0KJyKuztx0VO/WR3M5K7xV7/LL1y9qyukI
bSEYivQJXmCJwOLU8heXjL+3wrJ6d1WCXd0BHgbGHZB+TZDLJJGHJ4r6/cKRxNU2x//hqYFvsv1h
0Cv1Jl6zRhgFNHlUII5OdLBXpPsD/alox0ehv+BxB2Dl7cHJOo8Tf3HCcM8BA/YVe3RLKzgk282h
W2cF4gUdEohWHwRAA2lZonDNwlY3du7AB0j23aiEGQKesomeUqA7H3V9TEZK0IkbaVv3KNYg7GO4
zVAFTc9ttVUfBLqQRGsBmnTCYW8BWHKzj1eIlz2iCvH9O4CmIXKc9un09gXmHeT88njLLra3qFjE
nzJM5b0tnygnkdvmI7Y921D9QmpQ2fj5oUaop+lgoGFhH6zUdUSMxT5e9ornsaeYG3pihSuVIkiQ
QWq/uqiZgFYCWIlyp4v3L+e1ynGcEOVTLuLVTyCfkT6tMWAaHXskm0ZHElC/SjOzwoKmIXwTN61W
90xfLe2va4Uk60AUT2nAeV/LqjXBeTk6yBWgtFwa8AhtKsfL3SPsOU+EuoTHVqLU82CgpaSEFgOy
tsellT7liiNe9iQodBGHbCZKFggmUu5rweKon0qu2QD2EUH8Y3OnL7IGItf4jPGwh5KGH/XBiquG
pcx3X/BZr2jzcyOKe8qFKmwbEP24bObVAspfMMMCsJ8LzceOe7SAHwNCWvMoIjFTqNbynuiHB6J5
s6UodjrLC3i0gu9H1AcsNjITDQctXyWygraf0rK6zZRmDvDiGjs3QKasUItFQGdkZ4U0dw292FvN
Xv0b/56QCH+9FooJgiU5LI6C3wpcT5nHDCNmoGoRoSxodes69TlmkQQTlBSUZozGAt/L6W6jlHzh
+AYgBc0d0BsER0GvU332VKJjqn5aFeld87rTFQaxBJP+hcFXhMCvlgtCKIu20LZE720D6Kwsq5F7
ueADBhXCOvOwlnQ3I9ruY9XSH5vt/3PlmU8BdY+wtVXWj/nkLnlIdfOr4nh0wT4hiJXJ+dAiORMX
buq3Vo4Mz1RAb4919A5KPecP/9m47Fcyf8/bbQaTJVcDRYzP6dv2FQnxxo+4OqXmYu10DO54hnxp
YBcg9HLRL6oAkvfGgLaXHYQSe6EeyqxlAESFGfm0FKF8RGA21wGbtxNygnEj3yrJ8Ocj6OaxadBV
u43v66zXebjP+I6el3fUp/e9cKFlJoQ6gZ7vHeMgMCyHCQU9lRH7/KOWwnlJy66mqoTOPVRkVy/+
fL8fvuzppclNGWq3PQwT2SeAGkkpOBWdOak7yy4dluV78scHD/F04ZdhMaEe9Z7KLI1NcnqZ58f6
lyVeePZQPPROa7Zy+4LgVpaSEoeMa2cu/adMRhuTLFPlmzL9slPpYKrtANWVo7Q6dpiRFR7cujeG
n32PMXBjaOierjArj19StHf3WdC0odG3VTkLLizULOhjz2R+Y6EqptCQZv+ZWiy2aR1uHQ7vOls/
YdIgzVP8A9gWLYD4yQL1GNJ3KdEvavClSb/Q3QL/PixYiYFs6WelU801jxF4wWYMp3jzXD2OTYOg
7b7LH+LW9ZoyyrlkfMuggWfsVbQVaiq28bZ6QA/lkIhpjk9g8pM2dbWaMgY5DviTRXuIyuZQQVHH
0WNujfZPsBNts79L5f/+tHWL4dy5cM1PddYp9Vs0sN0TVB5b9q9vG7FEWCYsdGOdEEEph8oydMjU
Jjo+skxcFB55zdzhH5LfHphmdIS7IFjyH80u6KJV00Bo2wJwgBfmOeqoFzyRM7n+A4XmLPoWRWKt
GKgK6blQemIo91o16CNNZ1Wg3bNszXsC7fBR4R5sjo16AhzqTASDcy+zm3+XnQT1dJ0j9I/rGzFr
t3H+L96m1DyXBCH9bbjLc6ExkC+hLVfgY2Otb6HRJept0mk5VtQYBzvYnHedhhz/sMIkmanySzOK
m9tlKB2yE+PsxqycFVOnVpF6AZH96nGktw6n68rNROz6kiiiWQGfiS2kbru3/Khb+NWY8C0H+7AY
o05BntBhgFjvfnKjw6YCiq9SjJUQp6J6comlL1xWTG8CDKjon9jLWpPhrdOvftFYntklqYiDnhRm
VFtr2VW81qhS79ZzPsfOgLWfDYhJ9xbFhlEgbkoiAvwG08eRVUmCpCCDcz1Upy/PZXGzxViYRZ0A
FDQvAbV3MZevGh8GQasLVXfYP3fCwahC3X9X+u4R45xCeYQWBkVdKh863NptanF2aHGSEW5f8IXT
95eVssE7dF4nCeFHaUd08IBoxtDfWvSbebZlYdwyBUNQhcS2UWbaPIppvtD0ZL91litqrllh258m
PIKAG6FiGk0vAFKssaUe4sdP5V1nFdWQUkIcX6p63Gs+34fjZGuAeRsinCqxNMBnHVXON98qhb6v
ERuD/mQClWIO8Y2BQmz9M0hUHupSXET7qUV303YR7ztuGXBL0nYFWESMKhfLxQ5CC7t7s799BLLq
1XmPu3nBCZi7ZfNQEnoDnH4FaBP44yQFObanjeRaobo8Zb7/Hypclyo2EClRSyDCxkEJnhGk5hF+
OMebiZIz3VDJFoeRgM2cmgmqg0OVZOJGGbwiX5lxByBJDk8nnLSHHRq2VPzuRNxcAC86kOMSf8L8
u/IAmKFK5dj8ATglX/AVHIqSOEHeF8KJhXYPeRXDw8ZGdqm4yWvG9IfCjjjSptR6nF8u7DkP3hPw
Df4GUZLbEIn3AtRbJAFULel+MgZ2DTaUrWYDjJC0e4LJSy6fdj7CTFRjFkkvLxnMmcBDRVI0XCL8
s/KYaQqz5aYhQ7uSHWudyrLQPcwm0OvXHvsh1kB+chZc9DtF6uaDVBzShYx2bv+XCR/yHPlbtwHA
pEHsl8cGeUHg6bMMh6EuxCS1IXUS5mCtRW6yPqd56tYJ4Ha2P07iVqtAi1tIG2k1b2ohWLPjZM9v
UsRs1dTQvmXjmKonxnBtZTkJgBDXqNe4MlCVhOJY/SphbbYVRZ0jzyx5UVuj0jqwRA5vyNJ3n11b
Zk7TxmfD1ijfBX2L11lDyUguyw5rgt6rS4DXK0TSuWscA4PxxWaneIn9c9O6qHuT1vAGjm4bLV4v
1u54mbvSoUElNxZh+BviiOplxKfSbXvgW1lPghRS3Tbpaqh333EXEdvJjgS06uexy08RJcbdKM+n
2iPSY6mfRFxv4EJv930hrhvB5TEHQrxgGEqLu14PsJu0Mh20+BoseVAF+Sf3od3Up4OF1NuChked
TNdlu7MqmcdjnJ5xwYprfRm2MLb85U/t20+4QTaEGKCuf6ERGwv9mXKbcc93RNr7X7TWMLiD0okV
cJkhF3dRQ4ZG3w2BhadqeubZCJLjr4Ya4V/0kbqHez8sTaxCUucFEsBIHMN2DxQ9fH+PJ7BmE73i
zNhjbfM1H1mwOmbjBLs6YqUmr1eK7GKBIY0c5I78Ri0oS34a6e4RJ3fRV5ALG/020QtXLrI/CMsC
zlpBrPYo3K3Wpf/X9BB7rI7gKF6wLhO+3F6zkZEAg86qIxoVAAE7n5V9T6yUd/WzmbN5lqz5IMSJ
RabIp8grHTs2/um6zCQb44uaw25dggsI8diPK61mDNfrK2erAN6sk4NfAA7lXL+o7ojoBDl4p6YU
PYqcZs7Y4BBRYzalR4jXz/mibPZMYvbtN7yabXB7nfrG/xgM3yyVsGF1DctgFIDyqezeB1EVqb+T
KlCIBj2ZzMGmrxkXdEuBKSG7PFPkcyFfFQ7Zq7KltyZN4p5xu1iSvwYlAj/WFAZrXvjU0PsQgAz7
DAqAnoGYtJeTRxiUsu1HrP6ajtvIHLt3DMfCvD2YsDOqRf7bNrZGG6tHgB0XNa+jkRAyqDwQOWIo
d5rRpNO/9Inr6fAm2IO52sdnBjT2hkSvo6I5r0WHzvc4Tx57+YaN3c11Y4PhTxRIn8R3HTjZp8Vp
PT6kzuV7i3n8Q4pORYphNxY/UdbOL1HIvUE9lXU8uGVTJ2IEpfLeBm8uvozWodxCg34WxgBs43GW
hVyzhFVxd7VmXZdNXQV9ED19oBBEibRXMrGFPeQkvOPaLVfI9hCa6r5a+m9WogtFv//g6Yox+xJ9
abfaQ0Ld1USBXXkCIcWA2qLoA0BAGQBLxae4f3ImwuMe1nC85Gf8cxDNLtRMpFOMasLe2fGDchxT
HF1PgirxS0RvUNEoy3rk+b/2PnZwA6JqaoVQrSY9yospHG4DYDQ63+hKZiIMb2KUj/Ib38Y61YpO
x1hzODJkJtoNvTgjLPCEJP6xqRibul0BkYlDBvhRzjn7LDDXgngnrJh8jWqzuGfZ1Pwa7VKnOhCL
RwgcWicpSZMGz6GVGVCK62Rx17GIbLwBtyzYmTECk/R1SOoBlYMzQcuVzxOeSrdoNOMwyR2sdrYo
7rvqxGGL9EcG8J0lH+4Lu05UhqehK52XT8vcAF1AQjRO6lRI2Ny1Y18grW1ZBwIL0OlrPYH8AYyY
ERhk1/W8s1WRcpkG52meSuyDTfPM1bH/NWWXgB6Jafgg4ZGIxTNCYIKGCleet2+u/FzbZxkBM/kL
CIeEkfAIH0dDBrRwMVyYtCeL0vQ41K51CpL3jai9CgLDO9Sx+6tlxC4tTCsOCBCluoH9lQIi5r0s
r3ZTUFNMIAOdOuxtbf7dKrYfF0CIgJm3mC6BhlEnOoLxYqIwou/57/LSLtNq3ubbRlG1mVLOWxvo
Ze/peLOEMIsYdUyIB0yJPgSy7gGKRVa+lgxKxoAZ/os5FSdH3vQgluBWCuPiFLzI8CECmpmiLzaN
9+8ym4rc7QTv+GzIUImALHd+bGTF/qVb8B3HTjA8ZP3hUG9FmW6citTxu37ia68RE823VkG77pLX
ljcgTF81ifUpuuwsjR9XbMwfjZ4m3m48QTpVnOnTPO+OXJsU4+ZGbO8WFF77eNX8n6xGhDWqx96C
eU9101cQ2Wyv6fqO+2vzo0AD/uMZ7WWunrKDIGLEt4eRggeSTnJGGyAP+EHT9MQkvTxgWgF6uo+e
VY5XuRIX9G9oA/YMCbOwZ+QCwqL9xnsCiqczKTVEzvVKtjpmuAdzC/vKyg3Eh22KnOULIATsWPw0
ErjfTCwvyU6qICzNpGgnCe/cc8bO1xbr3bL56l0fwUzo6kGiGtgF9oKCFGkmaTbGkmsk7U7FjF1o
PnPZz37JgZInzsAWoGV42VTJpE1/+eheEIhh0hi8KY69bepS7OvGainuMRGsieooqOFn99V3DRA2
4OvnJBzOwiUMxxPRZV5w3dLjNIkTnlAq96nyHeebsQCIKgYhPrls8AzeyHw9m5zUTk+GaSUFiDfA
LsQCm4Cztrwgi7WR9PcVcLEsXShmppqW8uEGn3230LffUy3g3xhhhj8ZLSCaQ2jgbLEsBh2eXc0E
t+kGZOh2d0ouRLmcmLKs4T054MtVPopeN9e4z6QdBd1G4fn7lr85/fSx5FMMMsKtqd0VC1THuUhO
CrcCzdPXcB6rG3TAsoGpJjlqgs2aHamPI9UErxORMXZvHy+YUKUy3UpKMM9QNK2gNDPufy3kIV93
idO5mhf7VxJCXoKqUU39RhwMllmKbbLNbtDsmOj0zU4sDX75mc6WqX9N0tyRK4J7bkpIe+mq1e/1
mMiEvWTKwzTpBPGZcXnKiZsSHZC23ilBAxkUnWwBzUdUpcMlMfvJkqeZcTfzszE+zoKxoOowo+AY
YRMgfH/jexGZAX/TGyqj/znercdlKTdw5WJ4ZKwK6MOX+UBld8pUyOyu0CtJvD6o4b0+D1thwLX+
S1GKzaEElbCHy0JSxLdqIJo0/QpE6QEvzEP2Vi/VMJRSnQQfVRFV2qalEvH65WHpYnt4tLk82Pbj
QU5nZVep8DD8dMMfSgkwRSZS6Za9EqnC8pbszKf2MUhfQw0dOlo7mUPI0WfI0W8dKSKHW8Fad0vv
tMxDcnx0fbSOYtwvVbBxvSdgqEtLUSlr70cjRO6r/VLZPVODAVzljQh4cxMdmFO46TDTGzUUsdM2
FZn6Oeoiv0Lw0wh7HIyeYHOrq20Y/OoDfHZ11X2p9M4wYGKn6b7850z7mM0gjdvj5zigcXPR871c
A6TmXgMEg17U/j9k5MwxVF+ezb+V4VVvZchWkXZeXue2dNFPuIXdIJfmXrRzdKDCpFvt7eXfrKyb
5v76Jn4OhM9sR8ib2BGz3ulmw91zeAr1d+l0V87uyrsvseOVspUPPUFRs+d5qxgXAOGvr6vrRhhv
ps06Ett+ZNyG65bnzuSuqVDmR9ObwIHGwv4P9pl056dnuYAtX/hTnHnZZiLtgPUyqtiQB1PTJT4F
zmwoNWLXhqRP8u6Ztdh1asWDStyjBlX6IXtlHhbr1F3BULJ6MwlqAKxEb2cHTmGY5ryhCYvU10dc
Y9HSu2Ju9P3BTUuk2mz4O3FcVAf0/pBk4NYUO7gNHwgMiPhkgwoQXeUGa7gLBg5zHqOLG74tT8eb
ZfiqpLPq7VNKlKq/QHFf/e64jEwm7QB39urDKFVdprZ1ZYA1c9O4Uj57dpWJpsoTAyYGK3zmasCF
c5tgwI+QalLWk0JLhFQqp0HxRAqFQ/Kk795RkJX+LB/AfxUqNyB+7bmaA9u0v4ACepTyXVMMblBW
Tt5J7mmnfyYHru8/xOukwo6SdPPiw3vIh6PCAkhviIHEaNwjRhhLFySkJKLDOVkMuDFVX4I4Y6eu
68N9z4ujMpE2QTI56umDC5M48/WsxxZ+tP+xl4WVAUM0dN7NMmkHWpO2jF0GF9/qidWBmy7fTZQW
K67XOCTkWWdW1ATmwtYVdNEN4pN/gHIHFm/LzjGBc6LM2aiYRDfhz3S2wUQ9XUMkWVIr2ajc2vn3
8NXZE4p+KP0jUBihVwJ8IrtL5FfgAaskZqa9IC7NV12Z52IOkLKOOXjUrMCTjri6otrJsdCeV9pM
ZDhnM6cPR8MMcBBSPivPJ4AMeCfzlJLNPR46hOt3arEdOJ/xNb2mUqAXdtegdKPCWptw7gUiiGmr
slBJC9e2DAoI7ix2jzn865ibqVEapWglK1XJsA0eXoP6/R/AflE36ls0HDbNa23PiU/vb+hPL94M
hDX/wU9q5uWlZK8TPjvwvLF7Xb1Tog5NjnUILaa5ZxRCZjCqnYvQZzmUMde9jhzDYE/UBmI9jkOK
xW1n5RRPmKstP6pP5Z9LOn2/vS69whupgUVSCpzneGpmCZfOOoVWMLA/26bvQV/AI7RvzWzyp8fa
+OtYM4dCz6J/+ZeNFw7lX7z9CMvIqVTOdrwsjZkw+ODaKwuJ7K3C0tG1FZ5hEvslzVBt6OhrsYG1
lMFGrWmcl7pEkdkITS+Y7vdwGdJp7i4E5oozRZwCiieD5G9SBkqMrCtWf1lfmL0Xn3jWT9DSlC8I
H0rUXsNcr0QJyAt6nvRlpqLOLxH+1AuBXD6vtWUWX6m9Oo1h4HJ3ZEkHvcnRpjO+AeG/1vO5HB8z
4Vq/X6txxEiiloIP6PZPCpH03qxKansRkj7fyTMouvajofg7fKGeB627EB1LRfh1Txzg6k5BwCJd
jEiceKnh+IwChuykYxZI6YH9DgGnyX0q0uGz/Op7ntUp11jrx4GsW+ehID+pjy5bPZsn8Yfp2rLg
TK/N+U1D1qjwKQPBbER4Za31tOzD8/av253NhZmdWwmDBkawinekwkqMoM6EV4ep/Pstm1n9dFZp
2IRDH1MWw2vYkJekeNFWe8glRjsxQ4gJqL9CBuv4P22N1BLJsqI9267M68TslltuYSqOH+wzojej
1nXfCy3Isw5u5PNBK8ilLVwjPVdXcFWIjaex9MQgucHpQjc4yyJOu9YvYs3ZZ6aGMCpEe26HWvHU
m6g0mY/6bAzKcnF+dn+PV/bShY/UZflkyRnoSGIwdOlQtRTAwo7QF29zOI05Udan1gsEkZux6gaa
WbQ/LfCtxkv+LRJj5Ut+GP9ZNqMnuTHdCpEUk0FbloMiOaz/7y1PxCCNlAKa00UzQnr3N5i1Kid5
tpssYgaeNFtYJzS1uQYa4B07FKykx1AIFTy7pxGza4IdQ1Y9sYUXTEtLP3ESvi4u2DSnLdUOXzPr
DXcihSGi1nXE93izj/+xCLnJK4gDUxETJKJapIyz0+2K1Og6Q14cU+mhVibwulCK/3Q0lTq71Cfm
5hCoObsTnEkdYUyYnWkzYk/BWGvoFrTq+eaNYkMaU/WwB45RRw2NCZk6I8/rON4HptTR37uY/VbI
+7vXm441z1CEn43CJ1PnrDgwR89MTdWV1hKVbPy5OZeoSH4K5ITN0FkVr9poQorwEic/Pqlj3MvL
kjPUJSYHZVWKDp9XN/Sw+k87X6bUoarFlWsonf/b8tcTfqPA7tT5E8MhoMN525WrqMfQ922lsiSW
E+CwK8C2zRuDuHfgzSPo0aTDMyNt8r0LMpZmp9N1aHeT3nfV0dkPGcsXS108SkcQHP8Oi+ZZUD/l
51O0jgweS4AwdjoSg7CHYuH8cYnky4o6rYi/aLEd53AuCubrEkpTZVR2WVWrfySUabq8PA5icIIJ
YP7qSpiJX6H5LVJvDBxiEbx5TaRQdNnMFl5ETcOZ09noTJpKMHQRd117Nv6IHUSvSW5A6mP4PECj
3alZjbM+MgVNO9QVNqZdN0HR0xHiVpUTJ7MRrqRL15EY+r7ouMOaRY8AiSy5DwPa1AvyS9hxe1BS
ylRP22PiAEh3RMuHiW0B9u1fYX3fyQ0+fXa2kLkfw/O8HwJu2YM2ZDMt+WJSl+VRsKp5W3hi3Z2Q
YsFrlW/Xar8UJSLZrs6XInD/Np1okFM6amFQ4hOtsD+a/cuECAVgN5c7HLTB0Jj3OVuYAwqjxM9l
8giunXsZl0Z2VyJDgSWit2uyvfx66MZAOhEKQPoaOwxtygrzCMPB1ppWJy3bwyBbPwbw+q4w2YBR
dXbDL+vYU96XmIGdKKnS9SDpXg8mWV/4jLliugbmUNSmjfY4RFD30DPRMyhMCtMi12a4TP3Jm4H1
zui7gzqvxuJJfSiLGnSBL+fh6sdkT03cxC3wZ22TvgksRKIblSfwty1kPQGx2ezoz1ao/XN8wGr3
/5xHzlZbWU1DTeA78c5IKiHshF8d0pg8XiSsHl4w/5t55S03XcWIW+bwhpMV98mf9V4NgFop+ryC
OQhrtqukDLCJZHX/vM86wNCUZBMmEbZ73Boh/Q7p+qAJrjvHajOSfUp1tDpyWKGJu3z1fJT7m0+v
dXF+BmxMcoAFXc3NUm5USikomQoT8RK7bHTpzHOAfKs+g+lAoCImcSlKet7GlKgHKZkk5KvzpHqy
CW4IrX7ye6jQZD88CuP9qK/bG6abqXh4oIYdjNPMYhsyyMb8OugzXcw1Dy+5h1Lr8779rXlIaDVU
6pMa63r3rikKP2ciMSGVp5qB3UzDcEh3VMMjzoQiiyYu5H7UBIHG9az4I4GwX8EYHhfk5SWZTj5J
JBWkIETAhrwsPEyqKoY7F3BMgKUK/oI5Q1ZZFhUrZaTp2UwdVV05bRuVmsGKb850keegxPJNmlQ8
mXTGEhLm+jYvmR5WuTo89GaROGQ0yFjHhxZh8Ss3EN0JO+Gy0plKJFuvv0tOtYB9h9oLnkPVyHaQ
TIb7XVLfNmb0EHgXjOlSt5nVBD4hP8/9vUeId5HSPrcCm6yYDyMDr7hl7IqAb9XU5tz1hZG/gHCb
uGTVME5TZAPFqQ+uCWaSc81r95wA2p7fL34tkiVR6FthkjNg5noH3TqnOR5hVOcYAMVJKEFN5fNk
i/r+7wsJrsV2Bos+Z1KB2C/6sdfu5Lzl/4vUBUYTecwyyOZSfqAgrrFNvv2hdxRAAMdmhANTA4Lf
zTYrEt1i5nZtGLgIK7YNhNOHvvFJvm32iQs9wB0UZFQUogvN+VRDyldIHLGCr/4veaJ/sgJB1tnw
pAySGiGiHab18oRtQoOLrVgPNaxoqDuWzbk4svNGExlUrs8y/1Dvik9KGhrxk9QhHcGGbyHrOgAW
yOF4BQKc/RJuwLyaojcXxNKs62qye+S+7bjk6ov6gzMxuFS8B0gueHk+AMxvWw5kxwjHq6zQbeAx
881HR6XVIaG8KfVGDKeof10jZDMD4d4FCPjtHVbmf1i5NzSkRcuDEiHesXQC5yZyqcPowfscu5Bh
YlhuSa/5VME/K3aegMvvr7LyC9Izoi/o2+bdcS/SBLLRHEPtBc8fP6QKDSte57OIfeFzX012tD1x
F7xvhYMb2oKnqicghtipOYqNyqFkc6YIexcLQKLOSzwmLB1ddeKIqHjVe1FF9iDHk46EwrXI0mBk
83yS2t1i4nsmy6dg1xdcvPk9qfA2RjyOkz+z4Tms4OKndzCifQtg/M6BmHwr3ysBTeAuL2Ya50/g
EVA+uYL5jbFprH3RVmI9NvXTJ1VGD67101MbU/2n/dqWK4uEPizW4CK9IzioAID5xs7Wd6Gz7ENo
bXOqc6cYyUBwVSjWhlBAEPg8LoYGYj2B5gZk84+qJ00TkA3KNhVEk2bvGTQ0om0Hz7005/pN5cM0
wBLEhLL/bNaoYRZnZYMRo4gLMm4/xOKPJqetqmC9XMY7WI9cmCMCh3WQLVgxX7/ENUXnP17W39ym
u19hk0Yeet98wDMiH5DGTX11aRDgwcfGdUwWm80VUPRBh5HVJ+y/lpyEQtKDGWpHpchtSUkafaJM
R1JZP5aJ8DYgZtU2EtwRl1LkU4Sbe1j/nFm6IY/K/F83IcZwkyJBFmnPk8n9bcy0QQKH8b1N3/3k
7cc1ZnT1d9IQoki2G4ofkKHygHBx+oDRRuCm9C4bkIsXPs8PCRNlKY1HC2DtcNmCwkEwbNIoqX8d
iZxwGf0JDi/9PoQxU15zzX57ppGMtKvnijkRAB31slz1KfLZBhPUQHtGrnj8cdx4IZniMxfw6+63
P9lBbhFpsU1ONZJlxkjqXTot2Mw9h7ewL4+y04Hyu58KGzWXh0VQURfdjq1zsEu3GZsoLehsr0w3
TMHamRAdYwt7zBnV+tCp+mI1uQfY/tlCDZfzm3pWEAI6cAWU1/VbW0ZILzNrJrDU15uIs1Y4tzVK
PsWx9KQcBUZxnGTzPbUckf7H0y2phLC/rGechrQdvz5GG1Npgf4ctRMJyp57Meu/mtQg/vmTSmu1
8gMT9HUy9k+vLleMEXZf8ffsH8aYHvqfpmx0YNK9FH7rSrCuR69NnkmYqGfh/4omj/NOF5IyVrpd
urLIP7LVEp4TwCDo8GFNI/Kpf8z60zltrSuI9qc8CXGsVb0xR8dUw9yU7zoCe6QmqzJ6C3yTFr+F
mpZcDrxDVF0LrUUpc6I0ol7N4KJvrQbWBCeuQsz2lQGOAzFHbDuO2Am8/aeMUJfGAPnQC1i9+Mze
QiKo1CTW4IvMvOhfI++bmBbIBGcihDSAOzgZQPPkVnwtYOXX83PTGjh7sQFmhXAbmDiSbhnBlkq4
R2gPrcfhc5AEuxBcroyt9B7QcuZFRXTFAtgoQCZHYYCS2Gm5Nv7ynkQpQP5GGfhb+dk6G5VLDB6z
ZatLNcxQYgsdxrzmGqDAdW4Guw2ZFNoq3qghTUu3a7f5KdaG7XbyEQtbLIA/gYfP1WjGzg3+H4E5
jNv/YBriet9QFYP9+wZEvmZejAH41MO1/KbVpO3jObnatt2VDj+w7x5Vu+jOaWsqhNMmDnKDLW4i
bXyfgfBC2jVa5c/JZBce6OqWg9WEtbwSKeskjKIczzu/AKTRbPp2T47C0twRZ8p5n1XN7Xu5MTtL
PrO09YhmH71SEsdt6P5J8KBZMLeIcp7WUnvHvIlHhMTGXAgHYTEztzjvCQMKMzvFTToZTm+zPnzQ
rpmr1S1MC8XamtkpoFikj3BesCIH8yd6NygExPxVz6OSPlmOC9jw7+/HYHxn4WeqBLEZ1rXJj/D8
pPDb55RII+Ceug4ye1tXWH507FXoMLu32hOr0vbc4upz1r+o70WqiUXtaYVRzzNVWhz6Urv0k4ZF
CggEsthbkznQXWJTmyw0SlbnZGJ1lKn/hlM8bS15DCQUVxmKIPW+366msXzmzwPqxpyzmX3XNEpO
20ayRLDBtyfKevgSaF4r5RrKkk5mbghNiSUYIqS7+KHKxabng4lMQDqHGPzFA4BEReRfmbYHnRzm
L9A3GHb/VMR66QWsncHQGzyyedwBb5FkLNtl4jW8P1AE1T551b4wxFh3TGHGpmYoXGjnQo5wYaoA
HKQUrTgMUWk/VAWIRzD/cn5sXP0YgwYcL6AculBLpQ8FKdVDd+qPOF1uYbNlrq5JyarkMTUZnzoX
FyW9kpgb92y0zcL/DqLSfg0nxV9tc/M54ar69z+DZ0tFifq2X8iiFVmXlLb4eawm62exDf611oT4
/On+Qb7kzUhXhiAXEeAkT7lYBMddVJI1fiCZbTSLM2SZsn2+BxcGLsb2n2IsYfl3giK6T+65kfty
zb/wwbGofNli205n32cVy0BngFbyVzXuLDjWtlcxJALHkb6Wq1f8fviSOfV6/3b8S0BgWhFEk9c1
yKxQatWhQRAyD1evY+sRGRbjzYle5bs1K5otW52KKQyFMbE04H2wDBjFzXOyzMgMDUakK0Y81mE4
moq6sHoFi5RXEptTHcdMABofmvZEH20eUP6j0rgz04l2rGB9JrFHo8H92ZEawscpXOp3JKfDHcMl
Cq9/cMysKckR8Qm2Uhdy7W860NKk1gyCE3wGizbaYEj4idl1bJ+3Il24QhSB8PP/isDKqTi/ez13
E89LCGRYSem7kcDbJuAXfnvip8D2bGHYpFpSxFwdPk+jg5eerdc1rgGZiCdmvpf66qjwOVduXy7L
T3xdUN/LJ1iyuWO1sdiUc7KaKiz/gPNeVRRfmZcfugQYVq17oBBdpYHZLuOCOI2h/sz4sVHliI3U
N1nvl+ZUmRc1TkAxWdp8SSa7wNu68vkZvIFixzp/hyv4wjpWbxstpofubiLiv80k3ShgWYHMxFRb
lA8RuOY1yL2a7d76HSbFmFa6swXSx0LjEXr4B90pJ3ccg/ojVXgIBehWkTXmj7F0HENixi1Pgcy0
IZtCi7MGC6fdcBKy90wZSL/VQkmJxB3Ucr4mBJGhRCHbWs+u/430x5Ot7EYCDWtv6qwzmU0VTjlp
ce7FIwVX77GCGL9GlCLABA1gxRTw4+/ahBLKJN3dYFNh61oRVl/Kd2rl/1x70QrLa4CeOozHMqD3
HIvdWJnevol3AKqNubodITZVg4b33DsHUqDbAvd2whAUmlx9ZQQAkTmDB6lgGfBQdkINqKYwoRNQ
4KyLR348Ep0XpBnzjJ4rEg8wADNBLpYo3kP8xVs4Q63PcdMXHD8R8nBgyS0bXnyA80R72m9ivwE8
oRqy0glTn+PcDip6I54PclN4S9EM5FBpuyeYj8ae27JbwjsXP8fbbJ74E3RW0jO6fjR3CBUoi8h7
taZsGoRwPCCvvBOLD5Lwe2cWqSgMdM6ImN6sAxK3oVwrJmZc/DqLVPK+7n9l3e/Pnu85+E6i8yZD
uQyqJWhAfzCVxo1WLDRbQ9Su6HGRqfHS/bOil8W2Lkn/9rUfuGgakD+qmBKS/C9PaBlvH3mcOccG
zx3zF18UHwM9be6Ug6T0709IhrK/0cfWD5VtVqOWypftTFDR+JaJlt4ze5nndwyElGpGLFzbBlks
Sbzmzc90USfLXdZcUALTrehA5tQWGuJWcdZymkaV5Zgzg78jh0MO/j/pQ10ZTvHMfniQ34sJ6wD2
ybywl3lpyLevQjurKoOJiz8bTULga/AcWVT+263fFNbbWOR+E3+Z0jcLMW9bdmw7e5dQiqiNuUmM
kCdOJj5AYACp1uMDMepSQcM4QDSNp/kHkOg7HiyvaaFe/bCBpdXD/sHYun1Y8GzXiAIZMyLtiEHe
p51IjVBe1+w4DmYDhmRTtFQpPs1p28hIhLi/d2Ej41QQrAIZsz6sTRMbiNaGIGBebVsi4OUGHZKp
rGwUT8sK+/dwWY0/tG5ozPzlC5HvaUByVDkXovRpPr64T+/2ES6NUte5A63D5wGlO2Pa8Ef7muR/
/1H0SCT2jhNpZyWsBBUAQjmsp+/hO4awD2CkIJ/6SIA40E1DTft7kH0ZqTGF8eUdMimnrnNHZWqo
S/om+hpYSZoBWYht5/8Nkw3HJ274DfGzAVElk9JxJZtvhX7TmHZLoWTN8DCpbQiwKfZ3Lrba/pJ3
F0IdekT1h/m9M5Uh0M0FQHOAq8Pqg7ljQPbqLxxs7gVazqy4lg8kGNf7U/nwwdifS0UsTnY6cYe8
iHU9omI0oGlS7WvAcJZX5e1Mmxb4yf2gnONZXUxkvTmIMlPEdlCD+UmhBIViIFpZj/iS3jFQpIQg
6O+sV6qolHcp6+Sa+WvILDQA0xpNk/8v6bhhCFLBCvZ4cCKSi9aU05iCgwZWWDZTBbu2CIvvLrXW
/XYCEdWVoA1EcJMp0vqStAKTGkEDwNKbsvQvXBDBi7/aSTRis5vzjSCuTetU+hwtSF8xtga3LZ8h
WyPUBsAolUp1uhPhZKTQuFYC3M71jO3P2zWAphOFf3M/cWmpRRvb+6ah/rylWqXnhtufrGHijqeL
dbDQkgtANIX2Q9SDPFNnyOEwml6Zh6YXunT5pJiestdC0FHm8jn+ALQbCkamolE+hycpxhdWjg6J
+kz8KxJdba6c1aE3oPnkSQnUX3sG0INiDt69RHzVUSremxmMUtSFBznD8y1ADZgM1eCu6Zeecsl2
N/zV/jWNsjbXw9OMWYt8MIWHWbAIwiwWgy2Hm5SSw6T8apI3INMaCZ0GMIfoqdc/4VRP05F5bN7P
+OuljW+jfdFYKJl69V2fGegSy/5pwJTHdajsIqlXAxHgnQUIlRvq0LDOtYKLQqLDyc6ZN5VKiZ1z
YycNUHIhRGXbY/yx7BHpNXhFrqxLnlkmiGmQJRzRgCllghOeJ0JD313IBEPbR/XmARfddESbN3zw
Ao91lhH2yBiDXdlXpoUw2bKPw2X328GMhxjGpbgVJtAiZ0mywRdFZ47C+fR56ss1e71mwSjnTSfC
bRUxSaKMTeaeZQXC6l4VRZlkklblk5JyWYqyvSjYkpX+u5daB7DCD8NF+s3wnbXp1ALCAPdilu3P
DO6cS0Y+Q1E/ymDn/Z0Sj5mc2VeMX56PvO9xmzM6/QomVAsnUHaBLT9Is9jX3UHrrlaz6modSH5A
HATNxcOS1a98/riTddlXYljMmpflQbEdvHual3te+Y1ihlN/XTXOZ5XRYZPW51aa4nHkNoWIKYvD
M4peDcTSxJ8YvfkmhBlyGMYuAC1v+tLgXN8/WkAxuBdJEggQe+RUC7Ge5LZxHNBOeX8jl0fSzg0F
xYYzfeCilQk8tVFWFvK4z3EnolN+ESsSW+k6nMB2Q4zJN1h7XJMqTstLYBkwGeTIeou5GjZLDwZi
Ry9CNZnr+hnehmXqw07IfsbS7hOCug+p6Znbev6xWn/9ZI6uc+SgnNbbw+lXXSAi9JBloEtz1TRf
dSpyKPdike6eYahQXEccNwQe+eQeIIGC8EiCA5YReDbgRvOnHUk+hPKDrJ7ub7T2IK1e82m54Ohd
Ub66tdvb+x/kazvHZtpRyvuLm4YpTIbUu5UJmtNGaY7K107dd6p25FcNHHHRTAUDlzt2gUojsJHP
BptgRKZL9VJKXfuK62MI5HG2QTCNLlEqNVKMh3HmCGe+UIW8H++0A63nUxC+1K/2qAlfy1/SoBpJ
ZUuXlyTo4K57dtt+vpNjVPWhxAeEw8Q80Qhb94wFre9FqFuhQ8WvN5Ftd0ojp5fqTZeRkyve7dc5
VKj+yZQ+7nxNXgg8uIK0+BlbxfrgaKsvUFt/JnjXA/dFi8oTeTw6QI95PG3++qXVNYKPw5zS6f9S
EjjAknCczFwVMhgC0XUA/71ZbmkZf52h3FIYr8n5TGk/1vO4XTgdrlw038qo064Mu8VL5YVoKR+i
GVoxk/vWAsqvGJrnH8RHM6PypEKkvuvcFvQJsMlHQvUnj1MFhNwky/AItW6Fq0GkKe8TOc+cP1Pd
2qKciXo3ai7Es88586nI/quT0PpU8xHWwsbXtGPVRglr1NHHDxcFbleUEL7dQ5aaXqOeJJJFaL+h
tpCcp/BK8tkCDKaQV42HTd1Z/kJHbyHdP4BEKaYS7S0fXuzgTWKIiOIYjLP0ojAcZQrCSzIEjPSy
2c7PMiaTyF2LPJOzcSIvFkARa2GOuLbZ2eYZFiYhQFtttMhePSvBuz5fSl/FIAYdOVvyZb8bvYMj
5fpl+u87wol1N+ded2xCteDcZu5TPyYhZ1BIy7lZBPVtwWRxBT5AB99zoIxCEut9Z5OqzKR/bcBn
AfyuGd/7cthsrX9+/ZD3I+9wQsczp42nNcBZ5RtJOhwgO9y8atVZlSKUGmRcO6MnAEY/lQxbBwk+
tQ6lCrWDuHHrHyE+G14fFNgAdguu7L9gaSmbYnqEmwuEaGz9fw3IiFqDXJ2oYsTCspO2EiBdDuoJ
luslyVRGPyS3dskU/+gVn6G0xCiDU/OzAZxvhDGWQ4LA2JFZI19q5NroI2r5Vhv2/dz2pXrCVVv8
QkR287W2VZ5ZUmoyqrtjeJ8K8cFJbbrbjjCDJDNkXgNwxpK24u5SQoBZ7JKjvzor/CbKzSRbR54S
HkZDJje9OZBi04xb+Ps/HrR39RZEJI4CIHUEBwBs3J+JJDjyUUBjxAXuyG4pXtrgBqbbEgMoLI2m
lr2fdI28vvml1Hfou8KxocLIj7+dfokRoroUY0kGvl/xjuS3TUMTkdIHT5cjH8wlyM6PqwF9r5ZP
veRNdX2xWM9F7MWdy3U5qBR0ITHmGjWSWGRZc9bv4GwIrnFguhuPZWP5fnK1KoSHUT2A74aOK5im
5Uc0TZzmUxBiEB4BBcCIOQ0On5uoZPvy2iB6KowMgwaIW9Jk7BjoBc6EPbHw5Gr2pcX4P/Htefm7
Y2bosuYwsK8CzKTKAXZAf9rpl+LKcFm3m5+l3IO+qOFiUpSrP3M8J9a0D6KwYXixT6DMhaxit+zv
/LjV6IXCsEwECQyj3Ww5qbM3qm5wwNYpTkLzwu/zkrBpAt5sRS0e3eK+IG4cty1U2G5IXJg3pbFz
dkaUkCZMWqAyZlQddVFF7wAX1Eptn1261KrX5QyAj3kYB9dHUJJ4jcwXMHAt/LlwT7GDAKQI1Vkt
1jJiFNqT/qfCWuo+qmX8qqstO2JURm6rwqeoMn4atS7hJKX7eHRC1eX6liHbevIpkCyJAftO5Gvh
BqtVS3rcSvtk3xjZPrSW3r46YE85Iz7P0c8Bufn+kP4wzvhsujReiV2FqnLqbe6VSlntBJ5pJMFM
0f3hkDBGKvnSdU7TTgwPUx38svLskoeexgkNM79cpnmvB/yNX9qBSwg2NxB5MNU4SoAWP8JkWmVj
/YU/GBr7i8+U46Hl46ae78vzgzj2OE/ohOYNcDSiJ3UtjzVCK2GnySC4kr5F38mBJUqYDWKtCqai
DOd/AeHEzdrOvoMXnQ06czoJ6hXDql1oy7xFg7fo8dPwAGw5wL2l7K7RPmtH5QX6a6TvypGs1Zx0
ela0QrnF0Lw1CuPXFvbBykkjIu7NB8n9T5Ni/XvFx6w0nqdZDper4cj+ImRW4i/A0U/INCP2Kgfd
uh8tqGFda3a8SNqaZQKRgcepw/64dVicRBBc2caz5IENU12p7VBkbV9qHKZ4aA1EkihT27rcqCau
ws5Tz6MHntuAm5Y/PePY/ze8z604BBP43qhV5EYL1e8M0UKURb5F9SPBC2gR2QnKYtqbep1LUysX
+J9VZANrKo4K+FnE1mN4oDdHnFVCXdJy/t69MIxXNElcp812kJsSJD8GXMbqp9CK0ucMCw2iR3HI
ssapO2e8LaBSd8vlEiMbmqIQkJFXvZd2VQ/eVszAyEhKPCvTrV4jr43dlaLE3xl2P87jg15TrniC
EMszSVEKp0QHQVXXwsNFUW2htMLrsCrCryPM7DLokb8C0rszrWptN5qD3cFVBAJfa8Eg/h3GWVBa
mumIUTG0ep7EYOLqDKuhkDLBoi+ODgLgRRMTXfFJTCeOp2etd8ng1rUkKo5AmCc+ZPy3UeWlfMa6
WwHjR+osRMiXSDLutbF1RPGw/GNjjB7H505pZay/OUod0YHNfG5+KnDpdvutqhRN7IHGm/M7oiRp
cfwjM4hvLji/CcFxSuaIS1Bpj5Z+rriW+QLNiyee4FgG131WTBwtzX191Mwh3uQlGnUmyWtcql+x
OGvGMSyXF9toNqrjTQ4yJ6QnqgHKpHGe5IEWeYmlpRsgMJ0SXNELbq0PK6038nMlbr3cbg1qYeE9
qutuGH221X4rkF1c4GVbGB007gZVqzHgUNGSgvJCOevFJKmo/dEUh2CMEJpta7+Y8GoroAvNuoW8
3lmuxxVaSsrhav0agxw4HMf+dgBQsfw5F6KwCLN3wKOWepkQeGhHbUS9lkHwb8cdjMR7fs9B9BkC
JVmD4aa3vYUAoVwQg1gBXIAUr6NNE8sXLh6dzErBal32xGKgupRmVz2hE+VSmxtHZ4iG+tCpKsRp
yHsvCrFjH6nNWQMjuqyElniOJDr47prNYGD0SR1S/SJncm2jutM8ldAyXzjJg49pC6+4+9yeAvuG
QyB04VFehKVWLMsO6JqpHx/9G7hiLkfVhZjsEfCEAF75n2tmGmEzLRYvAW2WlVtJLPsg0hMZ7JrB
fkx73VLFXlT3XpKmhao3cvmhRxiwvQvf+o6bqcdPD03nj+df/2LspGd1WH5AaZ3FLNkITfw2b4XB
df3zoYVCxXGufHCNoShukA4c8BEaQiI8fm9qnDFaze6ucOm2ynfgYLnmS8vwTJaXRGqkegScX/In
+X2hUeigXscVvtmeYfzGwHh1DgP9mObWI6NnmNDZNGDeoMj1fPRvf/qFh+AeXdVFUks2DCNWj+ks
auhzv+oF5yGCdJv5uoBlhYyvbR+u9pBlpwbrBFney9ZF+fs1zQctx6ouViCeeGfWw+1NF1dx5Etw
wdsTIWLe7yPiDnU+wZfn/2Umy0HTN5t/gAwdO2w6WWNLO6pBjwjjSKQayKPdBPEJdzvsMlFcxfIS
JrURcEfjqFlxOFXQrwXqpckaEWHgqqa5htcgd4HDdIhTn1uaGax16JoJapplNIrgsEgjr4dIx8yf
KI+vQpyqKCz81OCeRWIt9fiH3FJ3XeXq79EEkeW4JTliYPwn3uNBSbAFxOYV3DCM7lTpdloHGFa6
DqgWNAjAPp4Or28e0yAsSVZabdvdQH+Jr2OcImjHkoZ4kJumYHUjeGAuBvffRHaeJNGe3Wrhms0B
JAj2q9qUPirfC+GP3YXohei8s64J1LL7YD+Uv1A3D+JOUNtcP5KgDniaGZuhger53T69GSzTJwel
6KBYh9TUVXM1F1GxobLJIuXo4s8Disx3irma59balrV/fKHsLk7wnQbQdgiqvyzWIqicg0we2PYk
PHMZv5G76YoDY0abLsqK8IhogprTPi8DBlnHYm09mKd70LSjKX/9qiyN0qg5T/jFTH4xmzimfejx
+sQWdt2viQ6QOIL0WoyYUxGCXCNLxbolTWQNxEUNSTEJ+PH/2gFdKqqETlOIXlw5HMme0ikZrfwr
7/5Xl6f0KSF0FkjIqcQlKRvvjFRpaPm6xBoBk8p8n3rRlhXlbSRNIZCoQ/hdTF8VTPadaUFs3iI/
fbjI5mUMqX3TZPQlKGHeYmw0tipbmIXO4nlRXg+GqwzxbnrwGtganqsyqfz8n0V9M3lqnC2AIgSV
1Sh1gaDw1q/mbk/BXMneg6mgPIERKESgEa6iRArE9pSPtKfzMWzKBxyTOejZAitEgqPF7X7VWmyH
9PFJFeP4ySl+PY4DfcjULrR2QHMMl/baSXzQEywPvD6xZXc6c9mlQPVWUHVf1+Rrl5skQ9HZx+K0
lw4GME60ftfBJZyTosgcJy1mqJDtSEvQhrFlog/WzvDcnY6UEc+eXZudhvD8bOtT6CFh28cQkZ0q
GU3JX8iN3qCoYu+z/ztFhZ25yHURNhZ3LxeEVi+FA4xfiF6Iv8UO7WuqMW1mInMjmEgH68QkSDMC
6hNYizOmxedB8B2oqq0pDJoQ5lW64L3wFILHawH8Jw/DWgAgu0zNCsvi7VzXtrmYR20hjXvQeDtc
A5bt4/dM7WbmIAJLxv3wkeynoCseKWgSNHeq+nQdDwwCa/djhlJHmxD5tG2MVGJADXqPaiBURt37
bIHe2uzTyGuSqxYGCyZ+0FPmJ3PXW+3JA7sxdNf4aUVLqX3mxvJxing6UFzFmIvzKVq9l6uz51Oz
Afs4yPtIh2Y01bgiN+rXfEEpzlci/+vwLdNFn8NEkN0iKG0pAD7b4bclD0JAi+DEyP+0vNUTagvh
O5qjmpTWmuygz7fNgPYGysZtHI3rKJ3nZ1pS6b32PdYu/U5+X9ExI/6nU+dTrVeUnmsqYoFj3rEg
OsxTjlW7uMHqZFyT4iOePuDNPGRT4+vAcGJ20/+RgCXtx0sLfReTzs1JlVb9T7vftme9wX7gmIPE
PoHjawnmseTep1W8k4sBeeOA1RDCxE3xsnGXmOP0Ove/N+Zh+M1jaAJnE2QT1KFKV0VYfphxFw35
bmDZh1ZpFtEfNMbypaC4P3Z3gTQYOahdkoryxPCe0YcvYqYOpY9v+l5VhKIO24PMF32zi1seBM+K
CLG/LNpzO0FaEa0GDBLkypvkhWYU8/xiL2HMgu3nCXhK62MkSoFmp2Rm0hpzxq1LQzb4PkFPmF9t
ZolRb8RketmRKKD/bNtGSOk3EFqG3XBhEtGwCu0K0Z6JWVmNtjhmUnfMGLKOR/rmw2KCv6NE48x4
hSP8O9K62/xkdLsvnB7RzTaWN2vdKlYMMrnd6qFGZ/+GHEaWvqSi4G3Ly9kkcUTaa3LOxKeYDQUJ
Nrvq7XOpv59PC6YKqtQ4+wmnalLr2/97YDDPd1iA8B+pPxF3ErZZKRXo9DFgGBUETMKqVisQGrNf
cllgvrvee3I1I5gz6POJEjVmQIycmNZ08ndDWqR9ygDrjgxtin46J70hEVVMnI3LxXd7KhA5KVyu
OEODHj7s3fgjAHRtj1w9N0IXQBJTLFBrVYt+UGE0XLhjVkbILGdz3r/W80lELeOmfRFbyj5P/50y
porIS59K9BGDwlJostKq0CoRPfJ4DVXUnLw/Z95CfjF0km6/9IfFi7sbl47VqcrB7m78vTXv+fPQ
kevboZJFIg2qp1BAGx7ZTRTfcywL1Y6BHPSAk/Bpop7CTbhX29B87Jq+Ng684ETdJdsO9VsUQ4Dj
r3usBVi3bvkWrcxnkmFHCc5Gpz5AVGrR+UQf3sDZGoOZPNE0Nogi4+OcSPGMRKASZvEVPI8U0lRL
7h+YDT/eEJRa9QjDIY4JlEC4gsvtvKda4vhmqy34rF++BMpWF+Gnb82QG3B6Z7U7JFMPdmfjsMiW
dbflp8IEv8kgOLK2Ej97oa8GILLeYRs4m2jl+sd521AgWrRRsSe0JUBIx3IZTv3yjezDZoFt/q1G
5NEhXwkIgoEmtXoEhDN5PR1vY0oUN7gZ3yTXoxpbTOsx0TRmb5GRWRduYSevjfDl7/CWGrfzQ2DS
doVrnxCIR4GNSeRSNh4PATMeTvIY+oN97SkuIBHzCMRsib0zdlhKzNBGMu1EFOuAU15RgB4A7N3K
65eZi2g37GLEykw0VFxW+dk5dL5KUtcjLkIR5f3Nxv1LElUBnO5Ynz736sePyghRCXIHt7lWsx7V
E3oJnGb+jApWQoUmhwsmgAupf5RWXuE9VCw1d8q6gprqZL8pp6Vyud5ow2/LOMd3iyTrESzB70ah
OM6yZckRyYR9n+BTfbflXXWWbGsydwlcgrpVHD9O8+ZAqZvKUw83bHyxyBB7FfeyAZQ6ynHyczgS
at4wIEenDe2S9QMJy4ze3mn3EA42+gxbEG4CfBabRlZk4Ek97SvZ0ySY3Dz2RueuhFxzEqfiQ04j
g8ln51Zw/aoM3SNiHqmrkNtR09T//M71Jbnkpw94Rdxf6TalpmARm3i80ZO7WTgFA7M+flq9AcQA
aPjK49alaRN2Orqce5//0m92AUeI2APdo0VU9Y5/bPol7PwfTAhk+OtQ4ynqkOxZZGUest+oqdMl
kHGxNpv07oqTHq/2z2RZ+5ah7XDtPnLSa2YU6ZQMgrC+SmestqFT5HaawE37u6X6/UALxRnZkXyK
IUrlyHgIgBcdCTBaLZNwr0q79ptE0eXDq7xzIXB1MEUGZHdl0FwwFmCqSL9wscdbKC6rFd220LK3
s0vF9vgsZv4j8vzXlmDi/ip+C7eZEpweaRw5Nf8KUEZVEqVy/AxEjFw5xPBuQot/zOUtz9+JJc4F
cu/5SaSUYkJo59Yegvm+HMKxYoDqNMli8BO8OITo6qqYoZan4tW9qCu9TSvWGooU0pr7h8D2tOZj
1ajGmBi/Esi3FYlnj6lNF9u2H+0/BY3lKMlcB3UBz8T9Y7jScO8YkjlVS+VAHR1hcqK6dbvxeC8V
FFmALcCq+F+VZmpLaP2lZImLkgDOIoekQOVAOj2jVZ22cvgO+j6JYgkonTpbpJ3OEAUii1OHfSL5
P80SuEgh3c0nd0yu9ZDK0WZTMevTJwV/cU9CYUcbaDZjZNvmBV9c83Te9ExkCXGloYcMLh1J1Jw3
F3lEexYiAW5NMvY9whNikMWOtOB7JTYjUS4gHkXsftLkaWbSQ9DW/qhxO/r1uZFnAw0mk+iv/gJC
Isn5K5jZ6KuUcBP+xLFM1BTey1uCrP1fI99bF/MqcpW5bs3SbwbehXqdXDmdKkpiJxen+KOzRmYS
jJqAnfVvdAw9gIy+znJAEQ3pLK7llOii9eVhZZgzlu0Zx4VyhOei0cfgMlclV6RktkLXyVTEMHni
GxjjcTXhVsslzEYSbRH9+7LW+yYGjea5G6ZMgbK1aDo8zUP9Z+XEAbU/KiJBHqzCjQlTOmqT8zlh
lDuqV3/ic/D23UJKBVYslDlaAZyelndmT0r6jPHAyUnZAQPnkyXaTHeAIBT60Pr3Pa1cx2C6tSn7
1tTpu8eD7/anXN5n2k4Y95BqJ7RX/6D4NYH6oDbD5qbbtb8Yefl6WmIMmN+XCoJlsaHZGt4b8Plf
IAB1sWTWqamHI3q5YAzrs97CvGzGByEzsj2RgZpUACAHKMvaqK+Ya9NUUAvRwWExQehqTU2KNLJY
zL0ywxmcepdxP2/1RHiIwye+rJZyU75/YS5x8N8tPii19NPOSmAkO6qnutcvTYiVNq3sDy62AD9H
XRzK9u0P3F9GwaHInvCyD4t920T4wcgb6K5BaSessp3XpP9PDWVBPFY6odrFiMMzylyYtpJVRJkL
FDmz0MSDAvNFsAdAv0EWfzv2BLJN0YIVu66lmcv+dLjTjvSlWtZ1DwLZ4VsASlluz0kTkwnISsqd
h+RZnOxmoKpTnM9PeVUK0Q6QeikvOSvYom+rwulKVNtP3dGo4pkW6zh0m9h+YZC9B15wiJqt68DD
X+scQ8qbISZglCpexOcSesIA2N4F/yXxBlEI3D5SLEU/Kw86z43gnLKPG9aY8FaXhLN5D0p/2jXo
hMHppxShY35rAM1UFQsGVIKIhrbqsJF7Ka9wVXn6ChG49hT41x+4l033Etn1QDqRZDCj+pLQWm9V
hfwEeamDaJwUTmt4T5JjUusMNPYgGUPfmZUgQInVeDSInfSeyQObOpWZt/32MlD7XlHlzt2UvXOv
eReMpqHGQLsEDik122hAkV09pGt0SuoG8ME9SI+Jvky4chLxHFYghYW5HS5jR1+X3NgALVkZs0W7
iOt5tHaSrV5rbOuy/5BOP++r64qM5me+srCzz3bNBm8quWrGoG90AlhKGLIIezlzYvQ1oLHW+pD5
mshraulq47caLMR371eXnHOfAtU8wIxekyqmC/v0n4Wvak8ZYv//Vojk38o1kdaJK+BR5lNb8GxG
ZAI9SMhubFqB+3ixd2vuDs6I4rDPA+DVSudwngjjLk2dvMHGX0c65BynVC9AtWzIIPpqzH99beef
ZHpZJ4tYtMWusRKeiV5GO0bUQp5i6JlbkCLZn1CQe9ieqVzAkKkR3UthyaR2l/h9VDa4sGoxcAbe
86ITlW6bXm88XiFfFfIFIsnWJVXvG4I1bNtUuh457ipDwXcv7SMtElwj9Qhrobi4Joek/VjOWr29
6tdlPlBT2MDi113BgPQsFZ3TOVsC/oTKdenWT14oekY8syN413w43Lkkxhn3VewHYV1CwqccPxtw
w88PSh0rgz3GQeuHfs976dFKY1a2cvP0QxP4qrcS/sj6o4tF9BJw44TjQQAlaBVx1mBB2NOaZEY1
K//bhS4ViJjR861M20BxxHji75HpaIEKfdgsH6Z+ybDl00MuXQER8NriqOvHl3e5u8P4H5egeX2S
8BX4hNp3hwWweKuyzEWELtOOgV+xcTSfUtR5drWhoCx8eXLZmEQtLv/xc2IKMvjthoAqs6+sI1f2
uCkr5cteWECLC7u1S2/p+nIdr0kJIYHqnh+nZ44hcIy1tCc94U/pVTzYrgfJ2gn5rPAYSWIMuRvG
GsLuaYGVPjKAKgcUHsJfhlw0eABGnqK3R9x8mb02ZM/uiJZzQTd0wU0wG8xkd/RaRnjtt/5S6DdU
eGkGkdrd32GHWV6yawYSf6x7KOKib7En0bmnHAZ/i+0ZWJeP7sXhRu6nNWJBt6yk+mEok24qGtR/
brbxIt549NH+zjiFHOvggzaIS+WGYLK1CIyXnLfyUp00tiAQM6gHhLjqfNv4pckqE3+uwmY7tweA
DBomsMM6oMnoV8EIAUypveo84mnLQnqs4SvJ9Hj+IdW+ZPkqajoXulkJuuTxzbrYXL3Gk681HWJv
o0sA/mWF8iO/RAbCmpRH4QgcYFZ757TCTKnXTipAQ/jKmsDUsY08fYoGkBI6OOBM7OqSIuHL0NDY
0MeW3vH3TCno9baaIgjC9AeDcN0eVVHjGGjzHzLlV6h74z01C1HhIFyVWKYPdzXAMvY4L3SDjiOW
dm32OCbW/lUG/qBICKUo86DYmQTiaz8Rj0SslGR+4NrJdjjsbtthpAQWIq9FmUeHw9TZ6kOLgBdF
syE2j4kTvIo930GftgqhuPVn0apsh5EnujMWR8JCzLV3tA+0g7zBUc1U/Vh22QG1cX/mam0Xxoqa
IVKkDVFdXsQuNrqZif/Ch4PzNVCydqGC8UWCaM7g3JI5dFM5nyMTOs3ias2faJ56/ynBIED8pnhY
ejqIMcv7vGkhOEOYLkJG/bkQ9hPnO6C9buio1JFpis6y+gtJR9SpbeajC0soW8vINUN7S5aCD9Fm
1GFb815I0StMZ0Uu3VqOIE6e6NpW0sPJg2KGcgiEdap0lCkEH3PRFLV4zL3ZgKcjEuqqVk7BqDAW
S82L7+o9n499uWGmX08+3zwjP9VwOvgvuOn7Blo8hxEEIVGHefPgIODX8VLRwexMoIjCUNBR/A53
aiUlgsr0Qpfqj9YHflAXbQpga43Q6vK/TPra44DJMz3U0ktbGBr+17xzgG2/i5jyWQKQ/59i1T1Q
bkiAoneLXLcCqFeVP+HnD/Jh3lMMtMyQ1cVWlXY6nKSgtAdkp9u9hc2xGIZxDNa35J0n1iLGVXrW
uzfdhizZ2JaC9ZX1NPbNyJlQDWUBm0KgsGbBGhrzcBisEu8uEX+6rVjX8RbApm5tp8+WHJQgVfVG
fc3GJTQpLGGpd/TQystL8EDlNT3VdpOxwKnO8pWSSiUI+ZG1ef/ylySQklTT+ZdksAaiCqgk0CA6
sDjo5OWz75Tyzi2wXUNJosNEYjM1OpQKh+jWP9jykxS/OdG1TEQYl3b9DpG6BkrvmTVoNGd9Cr7U
l7Nlxzb7vDLPDhIl4Soh4JSJbFxnXBPzeF2nnHxhz4242s+VaHwYV6xu4eJV+PPsrO2VfvDdjMKk
Z6PUN9z2/5XWCTI/57kP1NVZZACRvpCou7szfsmho6MakTj6SmeqKCTceG3D2slk8VSL22NsrC3p
R6GI5/pH+bp6d+0cGnGO/nCkm1TYTDbqRo1hhjATWECMfCOH8i3cZZ6SyzkOrp+QRf/qwa4k0hX+
q9ijpsn6ZgKlXtYgic0SM1fZRA376595u9Ytyq2USmqLONGzHd6ueZiqacx5I6+wnoxltwSV2n5E
TmAiGw2ojRzR8tiHrWbLG4+5ppuE1FeDl1x2+Ex8DrOjSXcDFhd88cRIo+L45DSAuD33reTdmzU3
X6lUynFs6HkY50zWsEXDDJA+tqsgEVktBYovvjMgqprgLwPTZ8qVqzBwrqnhnmLYq5t52l3QHJs1
1o5K70nY0o1hHixid1EgRB5l3sflhOxhKTNN1UJnxNkjZau/jsAl+0rfs03fs26N0RDiuxhYy2ef
UpIVrILgwjyZBz4YO0V6AB0GNJY2Qc8gW1qjcyCszIq83Jp6fDJJguUfequugvPLqZyYxmc+QsTO
k0cxiSQORAr5rULL5bHVU6do+65QdLSNUuTww/YPGyoQodU98HzDvHcWkhAeAXaDA6Gt0eLCikre
QaRyYi41tI6bVyvcGaJfPNut3332qki5boKJljm/ABs6nFey2IkWSa+JAjH7GuXZThClSojro2O/
nAJ+GHsGpn+NwfCZZgm0YfNWLXpCxshp/Svi09kK+U2wFQTOATLcUL8mgK2ecqjj4O02ctZJgpel
Qyq52sZsCefNPRI/XefpkCoG0cSBWZGMEeQBHUx+2OOrjXOhVjHrACM2lOquh864VbbAPoxD3/IK
2x6XsH9+wDJ0AMzFmlGVbORJPNaj/RiJvb1scS5v3DynBnz3Dl+KegPE5owxqx7G6ZZHcQ3fx1wJ
pM+42Pa1RBkOdgL81t7dns8nQ6mXkXT3RC2IZOupuscyL9HixjsneVY6TAOaNjFvai/jU9PZtfZz
WHNYhRGpEk+5V9Lqjv5u7DQzR0cw8xcswPZfgKu16uQBnXeOiPO6XThOWYFGpvU1DKehaMZ0hYac
u7qptfJp932awMnHBBjkqpMRDaKSQl3LJ+TKSkK0xKKUXKeQI3GRQ6pJLkm2KgdmoENKOg9tGiBA
mkR9Qr/rLyDnDlnh4qH5p2XMSBRPBeih4WvUWx7dWYiV7EEnsAplUPPqQTR6+73sKSdgi4D3gk1P
tw56LjqMMGmQiA3EYqNyJkyb9cvN3oc/fhpGlAIMH8lB4DaleGAYbLoL4+A1rdT43qDpFkcpIjGc
Arpz/T5CBAPgSY1TLlTSxQ6OJIZ5XnUIBN8BPbfddFgIfOp3JpRswTzT4rDuQ+Or8RhLEmTJuYct
BI6N6t613ACUzP2oltdiWPTJRwq/EnSkF/ix2+N6sG4dL3TBQ76xfwmUqUv7njH98X7tHt6qfL4O
d6Xx6I73GichgrcQ5bjuye5uM6zVFK3PR71POWoMjNfZUYiFIVw/jBbm5buoI44dMNeXU5rO617N
Ebp1NhbGlNQPh0A8H50VhacQbgS1KprNFSC9RgkaAHN7dyDnx1zT72s2y94g0www/36nxQYBN2nR
+8Mbdxj1TLYd6l5L5Mfg8z3ps7J0hLZ1d9SNr1uAlG0F/yjbzRTNGhPjCNocusmjRKIQOOgzoLir
OIyjJmKz6r1ticmGA1gG70ibdb6pG2KGUOuhFAmKQ9q+zmg/UcxVk6L9QcvriqIwnAy7N3Zw/598
cS1CZUKnQegSLYvSavaGACVm8L/hQAkIJDz6P/WFr1AJ0xAlir3fz8+FMLIH+wdyrDpBu25HikxJ
Ksxk/RAJHdJEsrtvLJl7aoQBXGv3362RMc4SG3tdjgOBYt3WF+U3Tn4A2XxaLPXdwQ/xg/DsPOpU
wAKCz1edfxZ/JPZZWjwO4xDkP6NUVHGy1j52cc2+BT87rhCJeJJl1kIVXD0j5HyWmMkI5rHP+Ch7
P0LbJRR310qhKpRg2wY8VdgMHYYUzWgA/1OC2wDX+XviI556IvOenJMvIOO9etaAXOCSAIIftt7g
tukCp1SRkQ7Egj/7lh2pMu+OsZUPG+OPmn+RiGvuwoTP3Zu4oj9iVipNHqHD8uycktNkKJbfCJsH
vJeQPLpw21pv2D91RDVxqryMOLT7beKJnYSUBZq9TzykQAHcnjwrnsh/aK8czeG/50+WKbc25Uft
8DysmWZ0Mw8tTVRK0jQs0zs4dW9PgXQAK52RSDR/hmnQj2opEvQ1mvWUlZjeqztjhh9wYmxoKebb
Fp4/++Q0wruu2H5iHPWH+T2kxB4JbmEu8ZasrkYwUmO5uLlfhig/K51E4sxkDgfFFLpNuwGrsKW+
tJoaq/auhkUwssYuIqIDafUzaErDrCRzMe1raJ45oQBifRIzfrOPoO13cCvzFWYA/1778NWYSzm2
geQw5qfC3lRLUVTz1KNe+NRl5/1y8K68DjESXVS9yO7gCHtJYbEb5bfRDKZ20uDd1mbyaSCNexRg
CpkqACg0aUXpXpW5O0tqFG2EeZ5Qq+CGNlaxK88uvNzmHSI3bejWWSyeMG66LhBuzYrh9lq56iok
PDr0v2TZDglRkf6vbW9O1hzai7wdncc5Wk6SRXOYpMuZE8O8IxstZ47UpGk3mYXsgQItb4/6GFy5
ZoqB1hFvnnHCtRz+m4yTmgTNCrXs3+vsM6LPv4zjyWw8J2YPZzIvf2HRUjwahtubQsmwZZvUITwU
r87X73AWrks84praVDVm3lEnb9Ht3c+zTtT7cCp7H7HOGjHmu+qcQY5vFHLGfa39dN1FXKdbjLwW
/YTtG7sR7n+QlQ/uZJdPKjXhiHnCZSGPi29htv63Kc+iqM3d+1o0iqmSIDa6Gsvd/xZQwp5HOYJG
eVqf9Mgd2L030SRZlCeYosrGK0z+CI9uFaCryOT74NHcDq2wwB38Ft8DJyDGyKLlIeIF/N39LGaR
b34Pb2z21BpaxY+XZ+vSG47ioMz5yU8s7/6ypndvP4iuWoGFl2t9frlxKRjd1t3um/nMtAEbxoo5
UJLde1CQCd1p75/mjLd+Su71uT/cU4YygVAtST9Wntz3dZLb/niWmz0Wn4pi7EwacQWiRxHdC8HC
DYVU1uI+Lo04EVhtfrRCinBQ6sEKoXHKIzfLbEajYuY3gRXHTgrW39f9d3xxDyRIfIiDIQ/1kH/L
RG5k/lc6XGNPDNa77IyU9kdnrSi53YdqJqckTOqHmWc3fmUMenlV3CLvrjctKLESAO4xarwMRg7a
FnuOg0IotZCEroLgkGT3KSD8el+7bWm8KzW4stuKaCWKqjS5A9ct89kuPhwDJ65MDwfU1BnRhqu5
BfZX0U+x4Wf084rCeBL9AQvY+i9C8Tw6seFK9ETm/HmTLZJTw4XeqCpY5nZjm9nCvoCJ87bm4C71
9LzxdOTBMdpO/egN8HFXbNnyn9L3DdyjhraKpx0fmeaB2gNHseg0hy1IaDnGKcBkRuuFsUQS9MA/
GFXhRDzmqgDtTk6HSrFQXiaiFHAdgPv18h80e0ovgF+BcQTWgv13KsShfWe2jgAKJwlvlzTIzZV0
9sKbbiu28yip3m7Mvj0RQX9sfu/Vyw7gqcJ97ERQC5u56QEFWt7vDbP7YthH4pIeByINfv6IHXf9
TKRrX0w6bVHuMZH/5NK1ZXSH4OQQLAfyNaiVstpofhN8QwznFaFLHx+INfCd5SHDY4jIEgIFvI8R
+9R28Ew3FIj2lF2G07e39fp/Aqq3y1ByF1W+AodOEd20vWfxWbJpkp3yjMCbbXspx9N2SDoijshs
WntY4JS/x1WLsPPXdaZHsNrrcAsZp9JOruGigt17uM2CJPbPvHlYVrBH0ALugG/uwulNLi0/YtE6
sUeyKzpsdW/yXMlKUDfwJYRIvSbcq3YL9O8pAuKGGZsMTyDoPBpxpxwsM0J2eIQxq4q8SsRfL19S
GIw25qGtp/PEl4qgEncNa8imCoO8a7yE5lb15TLKO0aSp+xTtge7PnseLx2SrvbYqvUljmr5QuYW
+u+iWtqz6kKZW8kEPkxRqqUCPQNmPSOwScfoeeMehyTIuWShWV9vhgx6Lhv5BGnB5awjosrmazSJ
0ALX5QhgOiT2PhsSbvAVf6DmyYPA/8vkZ3O0ElILlBNDF9aN8G6LyLgw5YaLyvhTFT656tyajy9n
IyTWppY5QQIQKjQOAb9c2xDpYE0h26ItCR8sSXweO+Kq8OxAveYx/bIzFTE+e6lSzfEvKaBNxKo2
ll+MgRqdUCss3BdJqwGz7NU1XczbtBefm+9gw0sUcfye+tn3EZdE6CoZpCFBsU6JraTcDp5yvq1e
EFC+5eq70zlh8B9kacS7n2t6mQ/uSq7PPndk/B1F9B4ak09OzNNmdb0N91IRTddB5e1cdIPkMob5
sngGi28Rw6YQWD+COiKJQMs9Zz7CQxeJHddGeVVqnqsJYW8eRdw/4Xt/9srbm5bpPYdlbT5rZTXc
2HloNh0xCZ8IlJn6xZHOMEuli2oP87dvdV91OQG80yhWR3oQBUzx6P1fkpL8BAHX9qv/h1dAw0zG
AJ/mEzh0JJwhD9tKVGfZArHjrPrQ2QitEYm43KYi5eHW085kljtIxxkyHwc3N0JgNuo8TO1nlS5T
w0n3IbS015VNS8QTBYDGWPxiwuUEXtYuZ6HRm/qM0fsDFJbtNjhrGjwsIYrpLqQkUeha2ycSbr39
sVH1maHV1nlsO1jBIuSBjEK7THvATygKqAG3cBwtC+IRhwi4hNHHj3dsbsKnGK20MqnfZzUL0uf+
m4RPjeCsYHHxXDjfaqmMvP6o7SaWx3qR2u+2nMpQdW95MXaoMFojmtw5mJo+hPimUYx2woSmGmGw
Ib7SibXHeZ31va+hTLPrzH8WWJ41Z8A3NLy8AWkSVP8xHkoACIvTPsReGPTYIK9fsOl0xOiuwm1N
5ncVRMbmyxVrd1nXdC4FkxoOLvLGPZWMoaGL08UGjGS0vXqeCnRlE5o+EZ48hrozhq0ftEbqAOFz
KDe6e+9pHEFFWQpQcn2grOuuJuZbOmChKN4hXSqDOR7ZHY6qE2YRBy5md55FWU4Lh+zlS7gbg+8g
jAp3r59mh3rn7C6wJC+4lEeEigvbLz5Aa7AYPbNtDJVfkDBL3lDzRPj8MGliiT3/AEeqNE3g0q/f
Z3HZZwkULuHDnrE3pBiKibz79AYEYl8+e6wmm2i0xvBhzYJNQa3J6Xz3FKbD5rmbdGSEUe36ZD2D
IjG1d379jL0tqtdKfQrKNwLB193D/0Rf4TSeWQKW9xTswe2H0lxKfohfgNUS0P5nKxh4N3o/Gx4k
XDl/NSAIdfbmIfgOnppJlsGGWMok3JEJajGu+NxYLZ2kk8zcSNibcl73FvLZ4hgBrUDZL7yhlXwo
P+XUVY+XPWVd8IKocP4ySJUc3pyBVQYEwUpRE2hQ41Ap27R3bGTAc0BQHjjQvdSTEnx6pEmo+YPo
3+4I30R5MJtM56tqroOq784+BqhbeNcXrPiQaL82oh+bZLPuqWNprvEyWy1R2rKwsd3LjcDk242c
RLHwIAJXo2+xd/UCv0baKWk0wLuMnhDSaYLwzNvKgSQv9YUZqtraAXaNCN2Er2JaMYC3zqF95EUB
Bby71sIP4g8lGfd9SNJUPELVsLR5pKf7xakpwHzUlt6QCGvI4/AGDxPadA50iwGgPu8QXvTI6CS3
u831mo/pXmMC981+PsKuQWGaH8H5CMbTE4U4reG5NTilmz2Eu549rh8793J74C3TTMxCxcXFOAFG
QDtSwxXUgdo1u1P+OIMD6hGudBXPnYUZ5BJB3GC1Tcge1OPrWXbjQw9Zfr/DYJgQ+uC0ljNNy49o
DHOmlKzydYcmyVasGYgp1112/qWeLso9fmaLpxsrHzrXU9E72G3a/IpCPJKVcYrB/F3c6UD4eGUa
T9VcYX969pHsAR07GaYh6hbpXkEWw/rmLfxSQrEqPRLSPvw2UyDZ73VHF/jG6Lq8VjRN9J5lTkYK
AEwE+bOOoGeDH9jC6iv834jXNDQaYJBEj/KaUx7bE57ZL/vR/o7widsXfgcnaULz0D0efwFhrBGz
vbLfO815WDjIZ4UMGslp0nJTXHZManZli0B8iJxXidkCMMBK/pZ/fL0Sv37JblPCjAy2mXo1Q96D
vlddhQDVxZh151qBwOn/Oph3SD+VOP9IAmzOQdH4coF4LEbkw7L/6R7qBBVD46Q1Ahs04NHRYdb2
APQ3RgQF1R7CfYyTZy4KdVMg1boRKiJoo/XnzhtSK19hlMzLjmTjcBj9CLAy6BlLRDlTWWj0+hZ2
0TNmSm5ugWY6r5IfSnL/TqykTWPlxSdfZJ2D3Sn58PoPn13jmOnxzf9mMo4ShXq6Ou0xu1NBvn/e
DOFNLOus52Wp2s21UaTSE7kE7b4LPgKqXomCXwUCbdDNwF405TdBcrhMlw2fGB1aEKT3eBXR61n9
a7jOF6CROND6hx0AAmInsw5r0BkzQJOlTBLeffNjA8vWZLU/Dxpstc75ykcJ6cGQWsT/OVZJ1lzX
w5yqaR3dcHPLAqqiqQSE8QIFn9Jr3BnX8/UpWb4A+Hijrio7hN4fE7WNXVWH17fF4X2nJIv2Gdpb
5OdyGbJcfyQTzR98q0iK3iv9fMvAmYsJHzTrvrxRSk+wABW2lOTFv75lvG39z5yIVw0z5x8F3mqr
eWOcRTeVsLPa4H6dB/LsvbEh6a/AsEftDJR1B4o/AkC+ECZ3G22GBLOrlVjdmjrQDQUsbyxW4BSj
b2G82+6nO4XSf8E4K0xT01m++gh0achYKJp5t2thvtcj1mxZY7uV7UlDR0JU7Ex3xOfTBxl7PYBC
0GpM2ppbsXNmNurbg9kkt5wBUbfDzISKnWexq0K0yuMwSlIhVeOu0hQ90TlVOGQADrTRJwTOR2yT
rYXdwYu8OqZ2Cm+Z0yPi2a+zAZwUylgGhIDLwHILmv0LHiwWsLmAK8UNlziaNYJ0KZox9DGV+RpG
C7omdnnxd1yoPBShZSrDkM5ys6JuURvrEzbKZby+BClZHEZSs4QL6n1qpU7SkxspK9aPxK7BV2+e
DShjz1LH1Z27Oz76iLL8Gi2wmYqGXyLeNbcjW1Lb5vTQhsq0mVNJyq44SLCyxWG0EwXw95BAGV2f
hnWI9vNiD5t/tzYLUmBfmDqAdlv7gsF+O3YbeqrAXgk0POxRlzF/pH5jrZptuTU7NPef6iEa0WyS
NY6XBq02IpXDA4d0YBACS3p+fe+W//eWLyRWMHphcHlJUdloaAXq/sMuZi0/t0qROIuCzkz40+CQ
LPXw68E2ZDjBmvAPg+nkYKxQ3BUrt372Qfsg5TAWmZ2hiCuF1/89rg6llUt8Gqh77jORSOZN+JKG
DvG+mc803l22tkToh9C7S6aYrIase36xsfEAdXJXVWy+WGLWAi9ycQEq745NggUlae0QDzIqZhP8
SmxLN+rplvy5BkkMiwlHcPIgyuWXpvBscXGJcVkoH+bKSdX8OSIdY0PqskMoWlquKhmABUt+ymYh
YOqQaQnY4c7fHhU7cSiR8s3t7H9u7U38Jblb/JNNAgmv5m2uVXXtBtgj3sVx6mJ5VQ1B3Rdv7Rto
mtzpXgNZugLiFIB5Xcu8XIj8NufZPsJgETv8ZYT6QjwwbCVbAEdwONiHcVSoQgyayMuCojDyafOI
L4iXr2wQR2+LU9FB9eU+wAfV/tDD9QKXVCwVf8fAIrnk/94ky+wtGm64+2JbMbT+cPg9SuC03626
du9a0K0N60gbTMXLXB9EQYyTLezNZ+IejVxF4aHPc1G7/bS3gvQLnUg/sx6MKnNNRN9ki/QWRIC6
sJdHErvAnRM340bo1VoUjlZ31WLb31kbsAdwocrbgb0sRjWsWZE7afA2egCahKbUMmQ+Q77Rz68K
VF9KwIwY57iG7lXBqJh31LMbfWgyuciLxkZ57jFWfU/eRqiIX8TmA/3yIVv+kLhRWTrIlUpSTfqY
RO7HYVpGp6B6zI5OPNSAJLfm7mcy5yNSKKd/xLE4xFbK3Bg2Knco+Q9cbOAq4C1Yio/Zqi/jm/lO
ANksFHTQ999nO0jhyw5lNO8OwASYZi55W2UsOvvw3XCwECZfA/biG/ZUQiDiaLIPaF2Ei0miPV8u
8/+kaOVSAUHiwMHakk6PplP6RqGOdVpplfCW2T5CTES/PCUAC/tCCAKDVBUFzus7jetExdsXR0x7
IgjS92iZC/kjHPeofeQIqCxCRtA05H2tiCG1fQrkfwPo2K5s2eeUlFm4SbCUqCUa9GzDgCjhreQc
9eZazZXqHSEtBZOgOWGiUG4/XTCwP6XUqlRw2DEzpLKFLqbBx2GxE6s4RJIklVniV5BOjlpaoW66
prMxCePx7QEooNjuHQx/P6lrEeltnEVAfWkmrBJ0GvlaysgFrbVQwQwUmlh5c09pvLAmuDvcndVK
9MCBEUiC5g/kwso6zjn6d3HAdNGnFutm50mHnqgvuObQ0OTYYuWv9ydFxMs7vRe9bGDLzZMv6sUx
TXV6bohPzeuq67tsMQNjAPfBVzAmP2fpndHfqcfy0sqfql8hqUiOxLUpGOISpWm2RLcUzkyEaV4L
7WXwHaGWNulRVyMPkj7f0sxhf7JGsi6tGbpO+Es8QciDFKCokvoCKbANLhdY8EyhkmEw3siIBe2T
FcFgVvGhn8Hp2MroQOpJbLAxujRb5FFER6DFrK+Hbo0VB/zj4SP527779Rk/jpOnlbnuXl2uTWIc
JrQ5/EbeuiRnTBYj5UjvUsFuUCiTOseK5EUhywZII9ZMkGEpqfiOFDGKoSX32qwRicYofTKcQwOy
lV6OgGlcQpN03lEt2AjafQc0aanTx+RGGX1xCvqc7+G4gJSEFFcU/LklT37bDF8RVSbXAd61xJBR
svIkFy2UwlFcjONZwquP5C2+524csqsMgcLq+npcU+AtP2y7yLzlaFKyKed3rMcLozLMtqONEJ+T
Atu9t48Wi4iOjxbOvg2f/0DxbLm0X9z1h25vrWi0eNc3hGwsWqF8tf1unPpk86XHG1p2TG7rH8oZ
6ibFzcBh73ADiY0ZfKQDr1T2yfnRfd6XDC9h9vyUolSvmrQPiyYHa6u1i3VMsvUDSkLoKPSxi+0m
mWllT1AXzO96j1VZZklWy/OyhpjF/RikztWPHDWlEMqkSuf2ShqXoNb5CeV2c80xmiLEEV6ENJ2U
hyTTHuG3mA2KeCsWP1piVGQFy+CWmzK18mdc8Jeln2r+khDET6StWtCD8k2W8qsZgXl5lepruHvS
8/OnOMcJB7BoQTFEAGd4PGkL3rEX826shX2KWBPDlMIaB71t/XyNcuvAstiY4vYs0d3OF0T+crXO
qHUf/3m9pAaDix5NV/SftdKfgZVfgC/0jJqj4qIzbUMJBOA5bKVwez7WlSINLDQJcw97mKmNTUcA
MwFKiBxYHeUSozhFAWp4af0F/fhjWhElnCwQsjUvRvPRVdRi10uRoAZbxQGlWF2tncQU+woUiW/m
ErxOMlqoiwwgu30BMx5LldRiMv6Rn4SYWIICDyi59k0tU3svtiHX8rSdSBCB/7UDb2IAnvt5D/KL
cTIrF63I5lB0J7hr/OoG0BpX1KWOJA/6gydg9Givrn7KxRM7DC/cSdgMYe9iOhVthK+1XmD33gjf
NcD+OqPYf+F+0ukodzYNfkOSw1ETMH1MlAxZepP38em2rMmOIXjbBrMVLQZ7M7L9huyYUbvBSEoG
sm2jZ9o74RJ0zD/ghIQ5LB59YIrsilzQyFIJm9VeRHStgtzcteKQeGV7yahzk8XFR+aSslx6FLDT
xyFESMGu/sGedsi2ukV7zl4iIA3TqAaVlN0PMqHM0wABVzFacbZiJwnvkPsixqsByx7QgHDsKpEI
dTDRsDwrrQjqmVKGl9icsSQ5tTCr1Lo0turMMw7jD8tet20ZaIhGqUKyuAx+LfbNlGfU0qK7Be4f
aVyui3VgTFtvjG9A8k7MG1V5kZOTBRggk0G3XrqF+dQ+CJe1W9g2QHESAono9GvyxfKYCjr5Mvp/
/U5skvf7jjfkq4XJRVoCrGqInkdNYW+5CckEtmTWGJdBMUaZQXB1NXBtAotvDbOg4zkLmOsjVHwc
dFdtiiL623qu4X+6EBWwjh1i/Zo1+o94IgYZ4k410iF5HRo+Tu5c/5ICcqC7oBffgO1yOLYmExnO
hWydnLwvmjb2XezaC/uXTEmRDuGH4UVhffAw+ytAxlNNu2233RsT0OrUhTOZ82pAMcZDVdevdhE0
S6TEeJAXhPciPiIkcpjSVu71DLivCxRXaL/geuQY682wNzu/4X1nTxR6hxn0/23jHVC3bahl+GeH
XWoHXvh/L2ChRGhhjlTj3ku4ZCBW62XkMHIE6p/poTas+7JU/ChBs7QZLj8xLVxBs2Iw+rKGrSKk
zRTXHG04pjzzN2v7CSE8s56FiY8GE4hgTwm+IFXW5M8OHAwBgwwSGPOydP1ha8WE1isAuMDS0Fv3
McYw8aMUhuczUn5ifGAeVmMTXDvUzZ5QkU0kyCVHfzUL3MgEpx6FFLsXZfogc3kkC+dAcwRfteCD
dKBjP8YXg1kvQFEhULzf3UfvZqYqjiVuEqXF19TdTobO4mKfeeS+29nZEyibWahbHM4bfm/O2P28
KbQEjyrk1PwBSE4yKTHslJsWlw3TJ3NG2vUjHb39OQ/kFT6mLfLi5i33d6YgCHZ/3YpVGoXhuQH3
s9752rwCy4x45FykezWlnNkGWpqtVspM5EdD4redsw/dUsu5pTieqv8FHJ9h/cgadsqYQamLMxdW
UVkfRpq88PPChKAPZua63y4Zc5+c+ljLrP+6FNFAG2nwjN22h+/loWDg2kZL5j0Jrio2OGBiOOu3
wCM76v7q0E7HeMlmMq7jpshRm1brCey5u0cncbwKtylcBEmJ2tzDgQDtTYo4Ra24UPtQ479eXLuO
PuR4QS8cSMrtDFYNM6Iks7Fg8J/7VFVfqrh1nZT44CN7SU09zF1/wCOcUMCQftYBm5pk3GATs9Ic
Poc37o50RsvlKY1dPDIfU3M9XuOUDJ8w77xN9R4rLncl9QLeW1y1aRzfg0XEpsvNj/nzWMg966Ep
LQmQ/nHBPFwZl24vcuNS2LKGjJg+ksEnTYA62K7yihhV9apPE/M8l0dylUVltygejKTcNKqy59fn
fwzdoXCGjDGPinUM+7BA5d2QmNoSR2bIAvTFSmPUQQrNvU2cPwJ0kgCkvnCDcHBn8jWA5SIJ7ZSx
W1amvQ/lx0lua7eutqLtcA3HdneHi8IsOTC8CxHNZrNPeeFvrtjNMT+Xlef/mA4qHfGxeQl4w31z
HqFMIYeR7YGzTd3aqDRcnhwdV9ydVhmocwFriTxCfBXrEQasx9J7N68RSSUD9vgtsJo3Uljnsh2o
tIdL7Z77MQxWRM8z5FMTKdfBxoyWD6zZVBmY+1/JiBi7rae3U1NNqBrBk5emkPpoViEuH8nFKKi7
rdJPyOrc/TEjuh4Vtp3J+dJGRus2Wmp7Bx6MX6zX/p7laa9gctuS80lTQjrlZa7OZ6n7lXXLW6H0
t/xF+9ZgjJAIDyiCx0dB9sFAeMvLxgyKvr5BTF/mIwZTxyZjf2FAHKYJ2DKPYyr4oh3dVcAC70UE
Ep55UHyoKtiWFLlUgoWXkO7sVXiliUEWOhvrAlhZbqHn8FJJk8t9iecrCelu6MG0guNObt06X4mN
3fCrqulOWJLSjTTPRh3ue5Ybjfbsi31CvaYr5BjvpcAfW8br/t6GB0SBDCbGajWS3K1vzVRZeEAF
KE4hH8RcIhsiVjbIHyU+bdzsIPua3GNRSdot8JaivzCVVPSFzlyu+QeVVbMWvotq8Mqwml73cDhv
NnBVK+g+rglV6QcW3kr9O5MgMhcHDrA+Ll+RZ0eEH2nsc40xfvrVo5Fy5LQDNMjSj/Nx2KXDA5Bi
8Bo+BOSxdOQRK57/A3/dZegWqi2dXSdr6pao1TMyXCdD4pCvGDXEB5XQ9Wdz6FBdYVQFnxuHsrqP
PUI7ETb9aNymnuUV8sFNP6FsqfLupw1CgZaWN84vtsvDdmGpmJmpq1pEMin6rxV9Xz/wpof9oPYG
ZpeLJTJUf9JbBJY7tlaJCXcnUPE81Jpx19lU0hDC+PStnauMKXUCwOmGK8SKrLJhHv+mxoJUJBxW
Ldw0//8F0fhiRESJMvpJdRdaG5rED5DsFUDK0D7U8G39cQYj+IZaGGOZBBvYxrxu58sn0lPOs6VN
zgNyLK5L5N5ihtxlW5WkW7RfCMj75NLTNR1ckFylwF/MKI5Zp11JseBXR11OAkfnpmdRIS7hVa9B
n2gTFe3Ti4w7i1K1DerVtL4eOJyZ59iwnAwmDjm3fWaACuRXLcgi68XW964spX7bel7miZMOC4J5
faydEhpDzM5OCHf5YmQNR4HMol9o+ma0de/jAGlurXpVuEPsPRi9CqJwskTapQhH2EwH6u8V+tG9
YzRlnn1ZaI8WKWcxu741u2vuHQ5zbqvv15ACb7w0FqdF10p1zF2pyuDDquhZz6ENhaNOgGgO+c4a
USLx7aGz+lS5vZ3PWgs/LpRRjL3Qn/PfhiDhawNN7gogVP4ZfSHpfw1dooESUZBtD1+qU+gwUIK+
OxpQg7x39eKgdYMCt0y1UMB2vfXMAHGwMBmP33Kvlok41ruUwVwfxUw+orZ922X0laed0bta++lY
Fe8cQtFn6WIftkAIfHjlSl8XNwQddRAJOtAohEPvS4Zy6lsgivQ4N1ubXEo7xKZsLzz9QOdLyJAE
5ovKP3fq7Yyy2Q66IQxDDY9IBSzpo9BDMVYeOWfHxU4FPKK+cpFypy5LRe0kNetOgKDtA5wqo8y7
CijbLRMXo++N9jC+48nGjSVHCBZQZxk47Ed/qKlp1sB3zpx0Lc6LecL90tf30m8bdWaZO9/Vy3f3
F0997E9d+LQH+FWz+fvkiPX+J3fRwQXJWBd5BJDUnL/op8td2GQ+wSVQPVejSmcUSMyhHN+fTcCq
RYL0+6WRfPDYZBOh0yY7ZxwBnSBcP0TSqi+gANn7G7GUwqYf2zWaS4xO9MG2X59IkxHaSzgrZFIA
c/rxowwjTlJ7mtLFFnmzPQK7P5bhObatXxD93Wcuphtwof54cXqYCJc3EPPU603AEpLDJpPOqCab
lB8NesEn677NtfQg025a84uxku4KHRKlRlwiTZMIiRd9KpF5PWiDl+0tLqA4+z8BkHLfmqeRLA97
u5cNbRZuWrK6g5bCE4sE+nK73S6hJ+IvfqYAf1J21ysCiKeOBdYxHn3BFRfvt01PHCzNYuNrGyVV
mb06qnBj/F3PAIhw8TxbUwSaXkbKqbzW3nvV3mhu+98Brh6nH1clpCT7VDQ2FwPfHjhA4gys4161
Be4JVofq8zmsNnS/zNS2+QhoP+QrSWynNIEByHscNbMbmHoPngzXltKX8HkJqWlBASAULNWM+e5h
9Jwz0yq5DIYSV1Kx6CGweOBSUbLFT301b3FonpnenG0+th1GTsvLwNBM2FEgTsicgzaz/InEl10u
sSoSj92LguZu8NjY1MUR5nmfuuhU8AZmbsq/1RqKHTrpb/XvCHCPgwuIpJkNW4SX0ZipBHACOM7O
8N5VLGKMxovBjsc+CS4+NXkZnf4E/b6N2FEAxWfminXB2CXd26Lt87Xgn+OHOcKhqxsjDta16l90
YL8UlM1jFEvT8LHJSByTO2f2SZkSh/0HybrqsmJIKy9v2cCcredXyPew2Nms3KVtDIHj6Eq8BSSz
jStSTww0m8GYqfqrIDI9OyR5gck68BMxyIrqiOzFiV+NjqP6fNUKh+79ijwDDK1ZpZ88lNal1/5K
+RcT1bXQVHlnxaLjstF1Y5ShpqEBKN99WXRDcN2Rcqbm1y7Is7BRFSAYkR3O2Cqyg0WD9BSp//q6
WMLw4sDnmzChVSv5fOwXdVckfKEeWfDT/2RlksPl8vAiiCZc950ZrjXDAmhRKbGpBky4+8OteKUj
XvSkN3nc1vDM/7w0iw2RUS55KlPK30vMZtXkzxGRZZ44sSTiaYOIMAIL/WwhPsgRsu+v1PJhn78c
ipo/nRa1lFSgEw1K/V+v9bLC3jUaonk8TXLkf3I8i2HFm7uJtit58C6S4vaHKjpY7MXyMRKnpfNA
R1Vv2pUVgJErIJFW4QEA3j6rHQfajzOSdpHfAlnyUBu/WQ0FZX+w3ksxHCEDSNDG9wFcIsZKyE0o
qO9KfXFcVewBE1n5H88SEODDQXg6nz3ahJM7Ndj7DV2cXHqXBu/5ey9saaMa7X6Oo94W9vzzub+a
2aacYbgeHO72TuAgjpnFF7lPDomrS/VoKifuM9wUAPTeHaxoPkphIqLlBp+vxPJ8z8XzrKgOHQTH
P/WNUNpB2RdjUETgDAIvYVBSWjeqaGdIkLI1IQneO6P4r8/VTXqbIspgwGbilXp4PlvBMXZ7bfKQ
5K5mdEAyhdwanlgPOk8yR1vzHuBxx4rdTPEFfQ1/bKqfXQenEbSTwU60SYHjK29TCCpKoJwpndtZ
MZeJIGYp7yRTX9GI2lWd3RwEHa/WsWvICSUYQfG3VmK5WMtJa5gptN4026ioWRIq+aWuYuXGjBVa
ToW3fz+/KSBOJNKPOH64hD17v+d45hAgNHE92gAEQwJXx1d45SrDIpFk0Wx6XRB7aIz5Z5ki1OrG
f2rkgfviz9OyAXqw0/UxTvAFVXApNuH+Oj7OqHi9yCuPfOMYytWUVVa6kK9GO5m/CS/NJrGXFoXs
6iEyeiNboPwQP0/zPX2QT5eBd9nLe3KfryPv76YEBELMNV4t8PeCTFrdCoDjnaGPwEe4TeLlWs1V
llsHdVv3D5shnlI4AhGXM9800KGGcRhrNhNP1RwGZ7OFhf82qF0qv30QPPOCfVZd/wbLCPd0/06R
xeyjrAXdRXqrXZyx2pwXJVwgxi5EaMJVa5B8YEA3IPd7vFv/u2DZkIJIuFNXLL2jc1DkGssH8HLi
h3C23reLNb6yyukL483csj7o9oa/zZBLqgwLiDWdgj04ZFXPfXsker1cWZkN1PmN4VHPRe/b+9Pj
Hoy92As2Tt0+V70IhrJhZ3pSQFzj1ecpLAWqMJJzGJAfnuQzsC6a0bN+NGQcJqHUALtrW4XZ59Wi
o6xyUzoPZNZ/qyBEOy6wFINrrBVSVwxN0yO+jruhGNMVW6r9/hF4tQNL/xm4Mfxc8eDKS4XFpnch
z2uTiL19qg3A1yT6Tch9905tkyJwnm5Pacp4AJRp4RBpsreBXf6WLMsY3fynE2fbjNj1z5uIJNYL
ES+9CovwPz0RE0NNjyWpcS1l1Z4iBcXkwHmyIQa6WXp6gK09z591eXkZn3QJAxgveH8HtVhAKVwp
pJucB7okfqmuLrtleGYNPEj+3+oRJZphPL52Q3c0zjDCDwZ6J10ST8If/kTtiOu6lZi0+gqV9UJO
MlJHOCs5rypNyQqRgjblMDgp0rxxXWOsUygSC+dRcjAhk/raC5fxUvPHID58LeJZkb357aGszckt
kNgeX7bSu50H+w9hLb35En+lGAePG5x/k++W4u6A1dLDUV5N0m8YWONzP7lEb/BleVJxKXcaZlUw
h8u8KyqTO2yRQIZQiTiKYpSibGMavISHJoQPoGv+ahUffznsLUIdDQgvRRGIgTGrkjnrf6KdnQ7x
G4uvz+bSZloinUOrC5De+AjdPwfycDphrIOVQ9hpCgAym///kT+4YPK7dV/Dojtj9ivcO7aIDbkb
x3LkfbxbnH9p5P+U9uNcCwmRZhY57mQrEVxC+iezN0zi+oOqyZx0pWaAtJDDQefw58Zp8xQqntZe
PQECXSu1bbY7XzYde+I8gRYKbZfFN5ihL50l79eTmJQxD2kHCcLO/aaPe3+ZYDBQklMFcoipxQS4
U1Ce9Q23tY1UveIskFmtJx06eVs12AIGPIlFgvW+sT3ptcGS37UlOpPYoeCZj/tN/r/0qDDF5Sf4
UUBjKoUKjOLlGkQI4qxZ2jsfDk8MmVLHTX72TDw2+gQFPOPinxFCF8Bu4eEOLqi0iQeZcaRskaJK
hZapUbbTra1u3Wj5l383bMZIl9jEosSO0nj4JMY/TJleI3n+1TwOYa1naL8VnxGG+BJMfeRcyIpy
KL5cB61FMuVQWY1afWniyF3Ul0QQG49d6M1uubXL6v08nKPkR7JwLhTbjSSUxki1i0emJQ57sJYj
EN6F4ZEhJFMc2ft98P5QO+Fc+pryODsOR/gqObxYdejYfY0ki2Xm+b7XDapLGQGLA24u/U+i+jz2
iWvMVyo9xnQKDxXJElTHcqax9ojxraltxBQybZnXvzX5N9kQoDxFL2dCZ2YUBWI+HwnFsbqp0cBL
jmcYZAEFwIjc69mnudFzt56TWPaOZoObwXivlfYD3fEnEdzTy1KPDZrSkN7thcZ2eyuiWusIfHgr
z/fH7kqbxIgCaFVDikTe22YirNGuuHJjTbr2pXLdNRRGk4BoDWt2mV1Yn2oSrMQbjHxE+xNeYFQI
F26LzfHpkZvw5kH5YQXgXr8+wDFT551mGS8PgAFfBBrEW8BI1uEqGcH9OEjaJjg2tepCCtzaylQO
n0lDBC8yUbAaHNnIqaqw6pQzUvI92+ommFAqMlobIbfXdNIMdq6xqCwIaBIgitG7jd3YLMWFvmAD
uqChyNLlB5Hb6IWRDNTfLQCmuoK8u5pl74wFB55l/uyQ85DzcHhE9KMbVkv/6Sn0MazQVzX0yZie
wjNckInT+HDPd/NCuozdUx3WSIE1nEyugZlw/FQXewRlfnQ9MBlHiqL6E+Ar3J9QSAnnTlbLfQn+
uLsXrbsbDIpmOybtle1uFN2zr2MQY/sfpRPTqNrqmfK2Nqjfy9Et1LyJJ+rBuRR3FMD7yiwSqHv7
tBlJi6gnxHk2Oj6f68a9S1g0xTxN8eQ+lSjtGsYowfey231oT1oJhcDkRJEp9RlRF2VQIn19OMDk
lxmFu419OdIaD8hyO0N5AEFwPhGQdX3lajplKYeYvu6cXE/QsZMfGt8be1gmhUqJDwTRk0WlF/00
XU/yegKYzuygOpTlATVSVSDzosYyOV9DCI1IOFz89+yn/zgDpcYK9zegVRvaZPeXxKgFs8FKkifv
p6ObEnItDtSZT3ocCYOWWNpuUaBSOJToBchkazoWnmzPu0hFt6GIMwHxdULT+xj42HwOk2/I+S/j
qa+jafWTt2YYJG6L+aCEortXyZ8R47hMxgEVTvtnETOuuIHvmKFh1iXMLO2DEBFa9yBIw2F7eMVv
QYSiL4eXCrq91A66oSDbyPOIkL2yG3E8i/B20pWt6Jd2ZVKKX4ifK05SYn62Urrgut7FZFrkhfvf
eaplY4FiUPj4JuQKMgzvNwBiPCvPvZsdh0If05wnbCOTozDW4K9icgXNgk7waY5AkQVqD3hgXFf6
mq9RaojcI7gRcf6guJImNRkO2b7LZa1xd+tm6OAQGJ79OxivXrx8Q60i+t4a9efAcVt60nDtfun+
RM/aL7enM6UEDZr+d9Jtafut0hOXH7FU4OE2P2NjMsXuVprthGOXQGJzEvzFIcuoe4rHlhErdZC9
pFz//15/Vw9t72Gb8vqEGqboIueVZpl0rA9NqmgLPSozxKCtA/jHyo3buFtVv5vWi+r8+E0H+j2h
myKEcpEbc0TnTuLtUFFOQo81S70OGPERMWtu0M9DX4P55GMQgj2HfotoyB2pz4kgmOhj/ghzYiss
j2caN8D5A1TA3kJvJpIrMdHeyyj6IMyMfNMgjtC8AiAOOQL3aWgqJw94APLIYiGyG/YWig5H2TXn
PqIntpv6CfP74oJMZEWObSZAjBNz7ZsgtDfuFD0uBj1m0XEpHxIZpBJtsbieuvRQA2s6pc3YF65/
xNHzTFgM4ljdW7fWAVfneecors+FBGNWCbL3lVlnD91LpC+KwGXS9QKC1RAQLrs5h7qNmRZvWXIT
r83bIKPugRugW0h3B51xjDZ420JAyre95AXaeVvUrxcE9FEsU4XP6lLuKxn2FersX2TTN16Jybef
UcnYy59Bs/duJ7bxCnsDq8jzEhadk14/kgzRFjl1aCXJ+PCItTSfZRtdvdIFp+QV1G228z90AXpL
1yRUferQslmAVu+8WbuM+T1sBPtry0IIkNTT6YnSZ2QD+jHAFzu0qdbEzthervmmlPiPhvg2jA7x
3CBWRu+dm6F2v4X9Murtw228RCSrfLxQKksYSYsFe9xeyCPkCabqacfGlnMK4YDPl0WOp809p4qP
fW45I0qGWeiqWPVGzO7JdQA7e2+SqAUluG5UxpUgH3WvOv/wgJnqd6rdfqdEdRCji/SfuG4PmpAL
NBl/wZtPRskRWVE+mEaK4NrOEAUfTQLUa5qBGiVLIdoV5XZ8QvDjQnHkKnp2zOSEwz09/JlNOx4E
/NrnLHegBMFh6Y+C+8fiRSRb521/OTLBiGoedy9dvzrbwg5sCf2RxM7LXJdXX9Zerw2YuTQwvOl3
ujGoF56BRPIzzi3CIT5r1p03bka35cp2QyFDavTaeJ1X0dyw9jYboBu0IEctZWa79N/+vulWLAdB
Ma2E04NpjnobJFwgdduH2AZpiIEuLH3EMB+BUucdzoQE6KkjcD2/nzAXGhDJ53DDuJtzKPG9AbrL
GWXpCYc8wwe10zO6M+DWMXaQCrQ8bf0pO+M0/quavP3Z7BlbLvgS1Of4l6Jee15QY3KlleOy3uRW
5AgFtdKU83Zr38ZA+mO6dJn2PSov3tP1HyDpaeAuF1P4kvCKf/sq4BH4UMKsI0oLuPhozIYxIbll
odNFapDw9eWKwlSwlHD/sM9Wzy1Ou0KG7LrH4OeBhFJrCY9WP/RnKCzALCqkw/vqVHayQfrvNNSK
teftaqSJ5JPFS0Cxr/ohjTNCmORc5x93XHLLbhhOqCZTnXImpQejDWrSgpaldyH1jtLt7uZAwO4U
B7SugbV8CSOxMvBxTVRk8Ikuzy8cJStye1zo2T+Rk1gxJoyG8oq+HY8q4DMb8tUjHVbjXX+myxBr
WxnJhSHkRZtuFqoaMoYwn7zKQ69sRYfa+AwqMtf75RG+5E3Iuk+iCUQ+z91W93J6AkUJoZ3+xK/U
7d01WIfrM3N+CHhGNinam2ggnN6NIVKNow9MAhesIk4E7+eG97D9/4MZkP5QMlVwnr8JvISkmFi5
aVXZCjNrXH3WRtR7zPkV6ubR0+A4VwwhJkYkCBJsNF+Cl3ZypcMXwLb2n+8P0IJ9uztrhQnqqpp9
Nkhe1izIwOL+Wqa8IH9Ynn26B1qBGIzHLkPV8HP31cnzPCriXZQrJ16+FOyTou4LYKx8N8jX8eoh
dX3MVMeXFQCjOzd774GkwR8CwWDtmuJpX7m7YoExjX9iBdCBCZoOR3IAkZj9mzgj5zWYQ5iD1xav
x2eC6Z6ZTIII4SOrIySiGf0be3wGALgxc6CY+sqs81N/I4eFVxwewhXSz5RC0SQn2dDhamCc7XNy
cjs9Jw4xyo8X99Clns677m8vmdvN08SP/YIrmu9xMUT5atZU5vCXuxHkvuPMZPRkc8yBiOHp6WNp
bjXrbimLos1557+hi8sTeajHk/TuDAefOCa6Hmik1Lbm3/nyP3KUlenaylJxbQzSMeN7yakz96NJ
Q01dyWBqyKp9DBc01IzoCg3ATF43Bcq4sl11FduWvXCD2ZzGe39yKKQIfZR+B6DWF0oqKBkzw8+n
gj9L4/xAAMWoZDS5fv58+TWGZS/evOa2/xc096mIYwLD2VkBVSs6fXnHqh5fzB2vNT4Xjsnak2U0
C9UqvDVSxV/zggjQl+pR0w3+wWaT1awyyjvGu0+Pxh2C4xTQS2qdMVBCGTXB3AMSds0d/vGYysEG
g75NOHJxuMui5UsBhyVfQ/o1xLXSqQCtOlnJkWVyu4TUsFM66IXLnwfjcguL6RgoiOTBDMnOlDdk
JpPEgUjpEElxthbIorpKEz3eKRdbOH2HdyV28NY31KPTr8ziGsV6a2Qj8Gf36lcGNjQfQ7u2GrYZ
lsCaD24NY/gHDrw8xAutrPFmAEiQBrdCCpji8HeK1xwZmbeWTaHOihZT7uBH/0j2LSk0bQdwTPNm
dPgYC/7b3hA+4bKbjpEgnpZEtasX5q5hAjLRBVOvsygrZHCcYECHh0bOcxLVzrn501mQMARzcz6N
2t/UV8nShDuOuhHyVm+raxY4XkdkOEtpdhgcoMcPLrAG7xLjSgqILcBAx3q16KcF7CT+xpVQMhV6
OgFYunkmwggSrtrxD6+SmI9RUjrYNjg4ed2ebPCyht+BqmUt6jwXwO/2PGnLOQpmb8Zdio9iQa6k
P0lOSdgOsPRnuffWo9Db0ChAd1xRSV2wy91Xt+6vCrINrJxShe9j/zeTy0US7bpjctkrLx2ghXPv
P+CBVXm6JhfE0/3Trxg/9wvrxZnryn9tGbcczfJAoh0P3w8ZkToFOGszNcBmsGxiUtXCoR0H6dVH
8eML+j9ff20ebNlKvvzONyJ4VznQWX1TW97rP+PGCiDjeIctwCQN5l3t7hm1YU5J9z5J0vbAzJZD
gAWr7IVRMXGn0NihYzJhJwAxDdi4nE+x0L/V2PFMVYTIXQvLWnKuS4yI2lebrwioiNTZ3cPBOywo
UeVyM02aWqAaVF3p9/MBfCkberp4drwC0+YACP6oD2UFewHWTv0vvEtbPp6qEoZ3Whbpdc8ifn3O
Zx/hWB7V4YFgYhL5x/2Yy/My4ORS6gvtRs1slHrpQ46VC0E/6OYayf89zAlf/10FTYvQRTzDP4tZ
LltvTjSOPsStbscGXoEklvWgQlTpGopPDtyJW2s9qZ1bUPWFTCDVO/ULKXrgsilDjHVVQF24dUKk
08ZlY3vFIHfqM+gtzHADLpGpCLOOkXaOllQJgxlgwAQFqRM9kUwlp4UV3FDFuPqvoM+OVxHaQeSO
YaqEtKjpcOcEy7olEsYp7WQAundUCcjAocW4VylB0uJDEA4JwUzHOd33eub9F3qjg4fQbZMYs57Q
117kFrUgpZWKjfQpXOeVxLT4WQCKr5zSNouwaF8+FEtPqCoDc9pMYQ7zrqS/Wp5O6KRPUOVTCpCr
fQVU8XghQvR8ERYWiIehPLl1tsqzRJgCI9hHIv53en8ulGd/7dh23O1J5iPHgPWls7DXex9fhIR6
SUwN854iAGEnFcAsM73hWVzh9l16OY1fv4afu83qxQpq4ZikPIcDdHtelKhWjsCszmpm2qCc6nUZ
3exSD+M72Fz1FRwyekkzZw3jTccD+X1X+g2c6Cy7s22j+TvzlQmuxYss29Y+Emex6l6Xg6NrlOnd
zmYLSwnQVAG8gMuKD1M2awvIYQdegelkDCp+2lYxcJQ2HkmSYHVsAJSScAjIFuHlz8v6MxZfbYzJ
OBrPEaBHM/dtbvkixeGjRX8xJ1z6gMtbyfn8LGkVIMnSU3DtZLjinGCqfhnIqNDiZ3DFc5T5DMLP
KMsncf7hixtpaC7Fcd3OzelyBzHm1T+vqSQQlINTsRWdzXsgoi1iJo4ePVq7tK2sDpqoUyZxr8Ki
AHVoc5iPv5Az4cnwM+oSQOua89+MXnawZ9nOfr/cfgn0YAwvnTZnVD+K+fzU6ZLHSoN2T8WBxgGF
xdWgNLLPyq//jEXJKur6CeVLsBtlbc0fR3JLIyOLMMvIkdMQra6At37fwfSajHDs5HjXJI0lUXL4
pSXZHd6SidIOBZEoRSQ9V5NfMO1MbPA5qcWHYiy+vPtPQ9q7LSk4wKBtTXelp9ql8Alc9qCnvtXL
F4i54Hv1ARRyksVq9Es1cdIhH7czVBhKNEzCgpt5VS+TqN3Pcq/e/tXp00m5SsmqlGHzK30RoaQ6
lFWxVqnm2ZkrKTytJb/VbMZ11mL2DbfdbC/A0EnGAv8sxUCG5YFSMRPuh0cKeoEMNx7jWzgUpehD
xc5L+jzqlYN+lgJPck2vJrgYhL54aGtoiUHTPf5eCxlvLosaUK3MhbWgSBWMSdXXXSKQuTMwm4yo
Qk9lKqvs7Clza+sb5EZOTn77+JuVHvysEBzu+NNXU0FBIXcUlG1GM+EH7of0BoSUGPbwBlHpEDBL
SIvMSrT9qM0ZcqCExaTELG3Gci8o+KjVA/e/FdFxkzJj3VPfc1R30/EEqidsHj2YKugmb7YQWIU8
fgPqlTP0lUfdi9nn0Iu0ncx7oBh5RFUgOE1sgijX1FYKLcbwDPzmJOp2oRHRa+lGiPv05g2/zwza
UHjb3Ca71Ug2lpZwGdGiTD8B31BNS69dbAhNik59zIfXNjb20i31KcCmTe4z0tG48Ln3ObVJTweH
HqMRUsVTxVQiiQWSywNfZJtoBg1uUXQ0i7s90gz4M+tV1VnTt5GHbexSJAVOltqTWvilZGBxT4+X
FY7b8igQvY5fss8tABjfcdKQ/qwVKropcSS1Hcy8X8JJr55TDicJHcqaD1NK6D7dsNyIcMN8HO/k
/s6iUQcn12/Ts4CUHr+qgDl9hE7skY0r+35gBfYk8kelLQwxM9wZd9wGUS0caIfl7MrJoiT2XmmO
U2TY/8mnPirzwpgXsck9z4AOhYrrqgDpFa5uIjoBl03FmG5ME3jLa/RuTawQy/N13GfIs3L4RXxC
NaV9BMfE9SO+ZD3iOrn1sXldKHFBHb6oX/S6t8Ue5trJGCbNNljtJkR4E1gkzoq474tWgQ/pHpxr
uARgoPLw8FBnIPbNeyQR08hy7/1J2t1Z9kUb1zNFeoU0O2L9zaQ7Giwa6dzHXRnnJKKEs15jvuUz
ZyULgJRUO+12SEhQD/1+luHyBnhuyQMzFCfsJvkz3/9faZO1VqXDSH33yQo86V6nryZQp+OAqo/E
82Ofb9GxrzbUiUxzh6cSdK7i7KbGJ53ZpsikQaBhFG4ig6SKPF7KgizigDhjjZ44CvnQ5Y0+ziKm
uzP9kTrRRY2klT1G0YdeuNwiUVhdjpQRE49dyKgaJ7s2BW4+H+otO+ORopsSqQfrSNLfmSy8jndh
leKuTZIFRM2z70CULocBmxcgz4WTIwuTqm5svy88WyS/n5J/B8wh66j/m9OGZOwaaaW8DlY/woqv
cxiaDAWVn8GRjqYC7z5h9OvBegIHOCj5XIMGw1SXDhfDSCKGBm+YBrYRvxrOaS+yWASA+ABo75+Z
IQA9rZJZH+cGE664SYvD3s/CBl37DURymR5Leda56sxk5K+yzHYp3aOzMDM2FO5Z7aPZJAkyPg+o
i2rPB2mbt9YKQQgxVE8ekt2YC2WwQA4PoUubZk9p3a2Nt44XYGwX9mb+u5G5CaMGgFy8P/k/e7UF
Z2M4t6RAEkISB3y2lmMlEDliTxuXx0Tswy/L4fiSq8XgCpQD6Dp9kd4xpdXbaMtLN6+QNMwzapRy
eNyLuKkgpbyTgi/8OwdPoqDAWdAg+eMsOgYRo7gfNTf1lxa2py6I7d8OJ2X4tMV8AsRLgDevuMH/
HzsAKgO1bOmWYOmh1rV0jAzVNlykF7XJBuFTJzuMIc3B8+Ec1uOpmyGHIfnA3wLxdzqjlaa3wlIw
nPyJSTGhw2HL1kzoiQuvoafh9EP3Hu6jQArH9GVGQEcp6huO3VmoovX+NM599BfuBA4V2QbK6lLC
SfXS/9p/weTHsgmV+oIj8Y9W97dLOH+377S+pnbVvXELfkfEPwHoQLAptZnBfUCqBu3XhBwDWAnZ
BzISYI9GFCPb6VCY7nkef7XsVOZ+MWqzpcgWuseHTpEoFzHq+HK47RGk+4baYDNBrAEFO9AiHC2t
ITc+6Z2+zWZsGEiPtj4Ruh6kSHV6LneMRopMnY/X4hNca6lh2yHwzTKlbiZHJvTTiYJIL4SEAOdI
w6SXcpJ8PIkkM6gvgW68c7ps0+arQcAmB8TpU4BtZ0gqoiCZNreiMsiKQgCUoOqOWKB3rIwA/xFS
8iQ+ksw3cxXhtPynb2kZivE+5qHE6kkSeeZe0Tke2IFqthnjfeFGGuJBBU1vXjXihUAptm0v0JAv
vPvnv0moqbD4qw7PXuQlJKeyEK0mZaPy7Ww2/a6ixAMmo0E3XolpyT3y9HrKwPzWKs9AUmFxL/Ml
/vwDVh0NRSNyikVTb/hxjOxNvEzx6QNGtM5g4IjXT3cU0IYuP/gAPNvD34S5y8MtQJhrIB7VDDj6
lcjbYqsWZeg2UQbATQLQokG5xx8fFRzdhOT3YTqP25UCGDeiI9kDOZjV7RiDNCQUwU0U27XqX4hQ
Zg2760I116juT9km8etRWN/FvucOb+afMT37wnupFx72Dmn+vperL+QYv5CL/Gf1FR1SrE40buCw
3OzNSMu2eFSEw4w2jit5XwFQrws1jU/Tmmo1xvrwudht40rnWsXkag2wh3PNira1fQ0kIyyw4QlQ
MzlT4i/i9kHfK9YvzBaN/zYAuN89mnDMWBY7rj0HjTa+PmGQXyM196sr3ee0IvzPXSKCobc+uAZ2
zpxCPwmBs08twY+jcBCRRA4+wwtbtsa8CvRQlcVjTM1OX2BSoetdahDVmAjvtHoXF/vzvCJBvii5
H0j+FmAkkdMXD3FkGzkZr05KOjeJI09xRIKcCOfsDF3T7IbOJNvvT1IDmA/6SGfOWyHfd1UOO0q9
j371mnnAouYRFjhm/Em3Bxp/GdYfEO6H9jYFx6FEoiaWXeR6KAKSqN5UnXpdiGMUZ6l95pDdvBez
Kg9nPrBgv7fr41gF4ADSuri8HU1Oms1reQrwG75BVIDwzGLeXUzQuFgfm5nWRlGQl4Wn9OSGlE8W
DVWdyT9HZCoV29jhCWsF/ypXVhVm+Fq1/WfHVgHi0CcaPOniCGuf3EUNafytGhcUJXdKHj4NNLYA
1seR0Xw6bvC77dUzMnOBIQnO+NtL1qLBAXzvxmVmTSmre0gfsm0CJws53vIb3YALGy8vTNeVvuhj
5JEMrpHPRzlgtwsW0/VbXyEFLp9xtGmM8OLvOAqtbQ7sF3kyDDsku2t4nDngKgDG1pKT1xRzh42b
hBuqIaYT3MMfTZM+T4wsg6IZFC3/taomjWhPsw30HbvtWMh02wQUduUUm6Snsor0XrCkqMJDNDH0
cnleNM8XKYiMjQFFHyRGmEjed4HUAOew4bN+uQ+MQIE1HFUoufGxZMNSGNYMGB5o3MrQzgbxvpgJ
smvmWYiR3XiJhARj3O1vRM+XMIr7qrzuHCU4BFG1PNQDeQT6EaDq9U3EzTOqNJd9DlvOdEKvSPJe
JY8lPjdXA3cBaZcbTrhAnpBfDft49k+VIIZWJanZVztxNCMpWl8ntmchTa0nYGskYbrNLtHBHdMA
JnyGaf54xIbU6r6GXnz60J7SuPgKNUO1HJ0wqkgXjl80qb8udsAlXbK4DCW3W+1b5Vh3/6bOYPbC
SuGPbSprrsCEyzhV2hHbWCUjfo1mb3c4hxytNdI38xlpxXAHnmi3gnI6hN6CR+cRsIzE+FKTMYHv
9RbzdD52s3qbe3cIdrBXIEBy47XfkNi7tc3C5IdZrETKRooQ4iFwqNULd2A/1EJf7mF0iqdyCux8
r8WvL04UPS/5xqCHc7n8cRZYsgNh6WSMWoVKIUoiHzzRMe5vpZPnzlNKkbPnpWQ7MSXUrCZWY9Cf
8svc3hgP31zY9RoEWXYcPA/OlkKvNSeOPDBbIL6dgbY4s+yqai/umT9MM24hB79c3YKYdoBHpKGN
bmjEDfMPw9KhE4onWVpsjgVk5wA8spAjvO7GDEkFD+jnbHM78sUqIHJLmQjG+So5BE4+6M96ScQi
Rq+4KomFdNG1pil4WU4e2n/gwo/E0lPDva+Mlrlv4LQJCTHKFzFynxkEizHU3UWlo5hcvM5j8vnl
/LIdXjjo3u11zUy6myqhx01VFOQB7Zm9+amgFWbd0jBLG8Srxq40UmZVxoX2nQdh4skKoiBoaXoK
Js/+nP/6udWXr0MSQ9r6W6xG6+YDgVh0jOSSjOglxZe2/gCGOKno3NwF3WI8jYU2bmt5orr/FhnX
nv7lCGfV3B0MrwjeI0Un2ZLo0JtWu1IHdVes9XfdqvZHiZvidiUusOD9EzppWC9O41Twx3s/s1Du
8LQLU5Nd+NjwXh3e36ItptoVgMf0SKotdK0OqdUfEGBr/qE7kU1arV2ynGjwjm4PRzVu0dBtuk5D
UKRWgjeKJbiOgk4OOFMD9IxvaVK9f5wb2Fjh6IDYRk8gmepL5GGhjiwZ0eCqLCos3B/FKbRucwTa
IKDa+79jDvguCa+3/P24SizatobVc5RCM77KOkIFmUbdFIMcnfMZY6FS+aS04DmC+RNd4DxQBilH
OXjSUcpO0KrOM7tTgzezzvzuQleIQBiIc5hRDca8zRYiU1fMOWrggLlSQcQPfzfyChzb4ChbE38P
l/iJS7DHnG23PO9Ht4l9M2/uOabu+Z+HJAG6Rngr1Dl/E7J9M85NArR7THM8jurzH/ZmGq3Z22fp
0jfb/nI72nLksGZPH6DXecaoLL6soNjLNh5JT49z8NM9QltcS1hi/5Rz5V/wjaUSjrgfonfveH3r
xem4haTCt15CLstFhf9JDg1pxWAN+kyFSJIsXxxpEYGdIjASmXrbGPLJh5skLc6be5z1SPdZVb/K
LbEcsOIiRhyin9cwqJkxIaKPQMgE+U57irwwd7lYG0YPhLc3Aa0jvuStAxqfz2QCLtDM1tirf022
LpSBNpvctJMtLJb+nLJ9AwbjtqCBvCm1/acUa+uBWf2I+X2yoAonF/gfARORrBEBb41nuRM8vYzS
AeY1AExmrBdYbqABF3Rt18gWffdFSWpQELL7j+PqjPiP2ySGYWRGMGGmLUjckeIqH2xj2qiOZ/kK
xFKFO77lIKNyljGwxGmeRwhhIezL+itSYwKKKZ1BvKgbdZSSwWVqjZFJAKGv6qdp0Lry/GdrUfYI
ip2+/yvpnS8I50mF1MwVypSvj2zr6udE2g39g3X3arMfhJIE9QCaNQIclPZnEn6dvFTcOIDagIgz
NC7rHKLnTd4QQdFa8x9wEhPSx54/xKG+ORNiug/fW4PPtHrUNrzckYxF5yrijIyjhXRfbVYTZtja
ylbw/NZ66rfpcr/k71YF373ga2e5JaIt1YN8PmGeAYNmOUmeWeceVTPpGKjOwspJ/G7jS1YlWljw
FCU+r2tsIKW4EorCTt2QBhaR/DiToOcMS5rgVxJMSIGKLy0hAeYLSrnBpau8IuY48jtE0o9Uor15
NieI7CcNZj28YtrB2I7HdtSMdV9ABK496QfHD1iKexJbkPvjcnXR/2Cng/1tzSvolQ3+pQdlbwiy
7CHZhSKXMGbPooZ83uu1cu3BNppLnlQ0rfUztwB+89zO95izFG+xBIujz/lP8DbhriFmL7EGkC3A
hwPEJiyrUASEzl1ZS4mYPULhmcr3xjkRoqL3vJ2U3GDI/RlIpM+I+tgUr6CM3VAdrOkYthrhHRnB
i+oEFU2vmxowSBIFIEpsGjnn6dZb0SLiJDe4F8gH/Uvu4UPTOVWkhFh1ObR7ND4a0M1BvFHAY9wC
jskRA55Pl3KeOPjLOGu0nzRAYW9oAHcL0P54ImLfhsX7wwGAy/uGhb44RPzn9J4ydUsJ6brbFime
NcfNOln4BNxgiSci0IN14W1fplNEIwid/qOGnIq2bCB/vvOkSIBgOsG2YEEpXKHY8zWYhxtjWlmH
JPZ0iz84Tnkjx4h1GMuj2BNAXZzuil/OSIDBckGAakQCZNJEGZcxDSMW5aaiLc1l0F+lCcxeUOf9
sbKWCUSUMYvckwa2tW5l6iLO2OO5TulLy+H89PzuYuUPnKMnTXKeCmY5iKF64FvYutxTbWWBYQlO
uWtIpE3lmGGH3fTMbPteNvHIs2HbuDrWxRfq8ctxfqlPuutBoDLAfZlfecGz6g+IDjvCqxlWm/pE
rH5rwhsOSe2lIIxoG1bP8KcTHJzQNp/q0HHXccmU7IRkyaZz5lFmgKq9ph5eGsv7iPvMXI2Ig1A0
Wea/d3gxAfi3BtuK5/7iF3vknEgTzGnzjNxM5NQc91eGPEVuZxLE3WcHmp/ar8mnc7+Q7r7IgzCG
ksXjiR6tDBz3uKAQpWg0fqSaSbaUyt+l04CMyKa1iyz+8gISaC6Zz+ltmGCEpIQluVtgzMbtFGtm
myUmam2kBab7v35vFS0vLGMYQNxei2RMBNawTPZkM8UxVSVHi4PtgvKShf02Gzla6tYxCCnbAlHK
dwL2g4R6VtrYqydAhBZuEZsSUHzZ6/WwsUT0xdigk7um0OTcjUmvZAkvqq+TS8Kw49kc0CEA/pG3
YPBlgnTaqXiC5qbtugUuuFId+5d/nfJvDBQ/GEPAwD7eciKVHsOirUw0qx58V924pIXv5IBzg3aU
X6f/sxZ0mbYntF7tGifHjwobLXHc58ZMEA5G5nj9km7x8iNodE5Tsf7EkuXhwL5RDqVvKZENKPKY
25TAZXP/SEvDme8MLXf+SMCC+RX0y2YCxUEmcIzZh8vHTqxMCi9XNPFNYTmrSY75bxbDrzu92jZz
Id+thhp/ReBjsIaz4JZbU64AxfEokWOF8kMITPkY/TpO2fNX+yXTbXkTIzvALzSsySpjPhSGGi33
/3lzEQgTEhVDi2HO0AbVaIG0lYbG0UXHd2ToQWOKsZKPrgIeqyUSvlyJxYh1o1Zp6KRkt+W4KKDX
hdGchJJ1W2uYIe9RvZR014avD+8iX13X1gUiXsLV4POUaAp//yBfccRpwm9JaLMWac4LIXzj1pdS
ASyX8qhlml+ycLS+cbwDJLZ8f1PaohgjUPstA7Xk+CCrBHMJ1BVZrEwSH25COVE6PKEXFU6sRj51
LZ2sWdzSbz1hzX1nRwIE9Qny6+Lae8Jfef8ICKz2Nc94rV5ELmGBuczHBYiMLy0Q4RjgobHPEVc3
iQ/OWZxmG0VncNMbAZ/NsyqzuaidmS0tqi5gTfF9btz/1IIlXPT0OGlTfKbhJXsgKZ+J2J06soCH
mQ4mO+V1ks2nCirl3mnOnF2Fnf/yiJ/ujoAa4MLmDVvqBu926dJJtXJ9Uxll3BtqkDwuniNuVok5
DtFAsLhFvv9/9rpPEKtPAXHQTiROsJBkmuUZ6R8SLDlTrV1TimnwqA4Zi+qdM4389lsOlj7Jn+aa
9OgRHktIsdaY9B/KVovlP0C3LxREM2Sb66nqqx1skVhlcuBRVqpEXR42Z+wGN/vWXwwatYxks9vu
lB+IilJJf9U85sgV/SFCM5IOfTvQV/iB2rIHVq9jUwhydWspLqDbnQvTCfonppMwyGRvRklrtapf
VZSzUDtU7qhnp85AE2fA5aVDiWJLIPtz7qrJfvaEmcAJx1zDxHyrAiUgJJB7JTBNGTUWpYkKmwXy
yTGbJMWuIyUr5RsokrH/5l/hz05PcEOb6AXn1mwFi7rRhelro62PYIzBBnX56b+4tLedSuh8mEvw
SpTGayj5utYy/GP+J52jgdrKfiMXN8fgT/4VS9Z5ZFjiYzeCiCWPnbKlBUXjBNF8m1Nqpx6nXWaV
aMMhXm7O+purLh0QYuV6pPagGwkll7n9cwfZzbKZ9rKfZpD9B9YNTsXVIRKAP/b4eJko3ZrxON0H
g6ZNoolV5isg2aEII1pHeuQaI1PNWC1zzi5vqk408R5ONAmVcKD7ExRgoclDaivlzY1CBaRUifkI
29iQGvBLzdPDYZCPtiQguDvd8hvpuNXCircSquEJFVRzlhFbKTvSrjh5jZY9NkqUR+JMG4+/Tj1y
G/+dVy/Ln1j9+kKOUftwnjSxQ5lG143uySczTSo3gzSoim2eeWiUj5itxeMYdqv9LlHPpKgSpEue
s8G/i1V3dyI45lZoX435G7IykP7kXUzEvGq9/BX7KabpCfNhdDEUVLnN5+3o4Q/lLeGTMUhyptKp
Lax1NY2HxSZi4vvO1W6mEHMRCjp+oeeg1LsYz/w5Cvwd6CJWJuJsbgCcxZ9yMsQP7r0AemAquDm8
2P1BOPOjzrzI1u1NzGp1syQk8/NjVNxvpWbWDTXfFa61DG//ASVse3kdR1uv09UpSC0/jZHL4kEV
EMhTONOE8ipdETOFCi//LEnw+/mknXzeCnkldbWjrhY36kAEzXbH8pdAImUPYsd6He8Kds9SuY5Z
vEAs/q7Rf5cSCnH19a256rbw+fotkjZUGt2JUIllDSFQtnLUcmJJvMdAPYKnj/yH8fsw6bwCCAIB
ffLNzMnuvXF5beDLsg2J+VIC/wh0nt6IBzaire/oGhVSBxOdQioLG6lZg9XQ33CT2QXd6/nBPYrg
CTFq4ml1zgCt4jsHNcspRcsLdeIRTojQ4X8nQZCcLPKILLXan06N2n3oNNOO5juGDl0iObTFi4nk
AJ2AW6HYEnqcBbUTB769Ilef+E/0jTkOICtabAnWYe69+d/TAN5BK7aiB3sUg9vcLNd9gt1WvwnI
vldUJCIQTvPI1VXpkGxdQECvE1gQkvjfhN3ht8615cLNlBXN89GM863d2IbU49YSHsTXL590wskV
NEL8YN4vE210/udkw7a8jK9UgqSC59MCwTPH8cfUPzSAA3KWFVny8iIjvMk4dj9PV/vknIyWXn9S
F8wGjeo9n5lqv4tnrx84tb1UFi21W4Wub+GGEXXRy/uy0K+uzEd4OwzCvD6Qn1bi5dqu+us+ywx2
4y+2YSA/4t5Q5x3v4oK94UzDUgDZ3OUTLLw2hAB1KmOFYLvxsE9GmCuskiRSrunAqmrh2tsfzA0F
JVIBC7OcFBtxi27+ndWqcGc1m4h87LFompngzwaAw0OovJGpe/K9C0uixT24J3NLRC7TEou/8BbT
vf5BhR5oePrw+7kss5LZrRsPREp65PM6rVeH6sM07fyhnBQN5dJ2FpbkXU+CVoKDIaU+m0wIWT7U
jxfCGghUFZFfWKzkUvvzb8sEoVKIu7GNCb7jk2K9DRGdSiDf+2Tblz/y5EhOHPFDNkOJ6zBHG01T
zKXdi7zq/lDwX3zYfbhzqmVk5Uqrw5ncMTKSyjQXlWyUGvxRabp2jfQ5O3NcsHluadM10Hhw2eZT
jAle5H6GTiyP2e9Sh346/AXLTxvbFmzz9erdyLdwjCdS6EvJEh3hJyqtvTuTSY9NMlu29d2VUDhP
w/qpf9QcRRwWCVm0V4giVaiqWsUtHZBRN/Q7g7LZIgwjMNznXLOlLhvV+STEhZLuWkOSo9gxAWBW
L+bomvJ7TAvT0zClYjp5mKWwGhtdPyOW6Ke0SOoNkWBjond31IgA/nIqMgUd8sggZbSmgt9lFedS
xRN/+5bn814AYeS2Q+EuP/FH+6EfzZvrNIXZcNSEHmsaI6u0P/w/PAi/+4JVp5TF0Mmbjx362bbx
RGZKEd41GdYsAL5taOPidwZANId9LIlNk3nCBrBbgDgaDzteFtluov6ZDg282NJ1RnRDsqfJd2Wp
gSxL9LPQ6LaGKPlA7/rliq5DniUppdlWZ+PXLyqH5Yz9RtOKZgWKfbGczrT5Wy1OVbMzkSKpI4JP
uLhGiYz6KOwu02Z+i1gViJKCBtPPj0MF5ItwwRD8/6LUAdP3RbqsmN0vLiuUaGBOdHdbtedboWb2
JGyXn1PZQITjyp28AfW7AK6RTzaFIg9vFPEtevrXeZvsmStDeOdr8HlBq9abU6VAH0kR6BL9p+4g
vHK7j82KmQ3aMzwvKdBjaFlJqhCHaHIKxZfaOUWaXBuTOc0t/swcTd98I8uG38GwFScDtsmT6CB1
yoUQ8k9pVNwvMzEyTBS1m98eqHuAMqvL0O608YCJaQR3GHQEI94DQk9IEVj29wrv1I2QhQ/A+y4v
UUnYY7Q8KzlWfu/yCjZYYZ2EevLoA9NqtlruXcp1MJwoXJrC/o0qAoEA8Ot7hpQDe7LYXZIVYbW4
2sbCk1BIz5JkXsbD/btZ3YeYdqfzy0Jk01fMzP5rxsv+XkVIaPRmhNfgs0RGBRLp/CaEUVj/P+iE
mWb9WYzOwEoxxxyakgVOsUgNOQ6xF9A5w4VPtXMxqzGng/yFOJvKragnsQr1fzLePKKTUueYBzQx
hHJOnYpqNkjbyUre+HMlsVG3EtCAnstmuoa4OfSMSu50Zggb795qfjZhRBG/kIOHp8sak16jP6bS
9KzAIiH+pNI4a/I+BCxVh8wota8FKEvLm9Z/kem2STIc3NbqWJtJ12zCOEBKiF4ePE5c8muoOGqY
yjYJe+QVFbn35Nte1evpNCJVIllNXbpLlSuE/klwAOj+ahmsOtEb0z9MH5ou40NE75W5yK/1vfad
agHLg7rl/YP5MYGmFnLjyl+2ZnMe4EKt+vEOlX1BcrqJoCUMx8QjiQ/+SWJ3wk2rOqgX4+o6k2as
G58dIHvcHEtAE8+OVhw5ASngRr57YHBZSUMCbuCITjNVKE6Tzxfkm4OVpzeOaRo7nP1lv85I4T8B
syLFbjhofSBUIOO9ygthm4cT63Trw6ByuGbEJa5HEqsQX5ZtoirSrHwNDloa2kPPXffoiLTphUdY
89jaLtgP3TxBherjc2/U8QIZEVF291XOH2z9stHPvZSANs09ljsL3PD8JTTZOf6HutUqhyHOzdSV
Et8v29SHd/tfzJVxLlGQxsU1tE3sLvNPPxu/gBLbDmWFT845m3+mgkdOVFUyO+vkjafEdytsexwl
dn9EOEv/moAiyk/JyELOf89V8X1ma5AJDh1ph9SV4L3WDaOnL++k4Dbalmk36zZekmpwzN1XaexJ
/boeH7wWV/8q9gSG2b5hysyYnFSjIEeNQnwwxdhp94aKNZW+7DV/MY5slPqcdMBGAtJQf0u4gPi3
1f3TcoY4iXEIEXWcqF9BWmufNDggxVp55TJ6kya7nCFP3VRXiXdS+2bmR6/Qrb0zaFIgbPJAzlBl
6X8zNgnsonaNZPHc2PyXcSgMDKzQdzimZanXuTirdK+t4TrNBN6TSPlpDXYm6FemmEEuygUmcKMp
wOXHhplPU7hMBDvWwiEWBREZFDNnkksdOtrzsTS6LiwubbLw5Lu14GBLA69X/5hzdmff1L+p2P7c
1pbh03lni0gyiv8ryryb/HxE0BF0BvBH9wKuS0KrG3zFpy3Cxpeqfuh3Ehk1PAlhC1u8Zxh2sJsl
0p0Dh4JUGPnxOw55KUE+A5xUc4X4ZVWZPILKqRMAH6Gpe7cUmODy1QvK7VN0M0kSdhFWreeUQ4wF
YUm2PaqtjKCLsWxqAzY3DtHWPHDhjiMs3mMmUoJXg/HzWdfoO0qTusYI/POvteEg6SgXLgEMF7ZM
KkZn9vVfgeybNevZJ74RmOkp+VWeGaPEXwxZmXRLgcfjqRHja5TmJGrW36ds4IDQaDbkCMjHEG/k
wP0sTA4i6Sxet6b5ad9ryGKp+O3XnjrakaKhLLfEmDH5TZ0+SJTZmMibMSyTs3RWbFQJok9aMp3l
HgB73elp0T8H+GtJQJfxt0qt0zNufRti0Mr+Z9EyWcoYkZ0KlmRwarNDjEe2BaES8TfE2UXoyl3G
PZ3Cdf4hMSF1A+jcyv0wkcutgAb+XdofXX5AmM2NZyGDuGkjtlMXQZdAvhJ4YvYEylguXbitOQOf
//0m/QvGiXfzmURExcdyhRZ5gWfUbewT5NVOobj9iMEdUOMeYVCK7jKHnfBKwIB9JL7lugWplQMV
1xIyWlTTPFQCWYG3qjPfFN2lDjV+k9mE++qlMb7rzJ4aEGh2cHQl9P9xqmpuOsKD72EksFQLyZCA
+KnZzYOLJB7y//xvq5gss8Cw33HhFUKFItwRUeDDnJn7jxDqDREzWqJyNPZYt5LxoLF0fdAo0aLS
USobMgQLH660k1RXngrk7tl1OMmZxXGNd5/5mvMwY6J+nJnfrNdRiclNq1X/ZIcYvoRRwh3F4eEa
SJskNQ2nRuEPaCERLJhLyuspWj5MC2zBRzwEwt3LfiMr6fkRQ2slNDwq6AjYLvdWvka0QluEzFbS
MT/7hTymGKw51SdjYS20bokijdWYChsRHChBqWLKz8egYWJAjui9QhZe+hON/GBtTFYrbnnF6G58
XCo5HTqTuCK/OBG3iNXpc55tf8S6lxno6fq983GHqzAso4JUdWazDf3+8e3LE1PmUpm7kWKN52SX
6dr4+fZ2weIYF6RyRvu4mBOG8TGg6fYxax2Rd2BVVtHyZ1wf3RpHKuBGLX+6Un6N52IL6S7fSurr
ojdGJloomeLANbkKEXWS6E93W3i6USlOwjRQaLs4puOu6Ibre8l3Qbaga05OWd9IeJIOl/kWZBWF
mHcXEp3g7fV+q9ERnAhWh56AnBMBZtgUxKhlN9VHoLi7WwizIggtK1mBimCHacn5imFqMzeV1nyn
hL/e+nB5Akjfv1WXe4YzJsQToJa7oIWZoh870sRTBTJJ3Lsr/H5bNTLBHID1O5Ld5fJsQk4OOQKd
1nwu3KN83ZssXuSdNy+ofXjjwOwtbN/Z7d80izfMJq2hLoZsY82vS5s8LQS2TvVRneXUxJgWIO00
QAUNgO5e5TqIOD8WpiAWBG4b0EHP31hmEq12CiVBx74pObs42XSdPIAWQpPwUQdDN5FVkzJuu4fA
jfXCMJAATLyca9RoRtWfJ1ZcOkT6FbQAAYv7fYnyht8KntGJwkwHFxGt+cHKn3PKPxRkZH1KMoIz
praWfucuN/qJ04bnZscJrWdV5vBZ/TbQmhX7u8v2KpQ+ovBWrabRiOBgUjYgGeJphpyqPCcTGndX
W6PQtlVLMeQCdpVsadER8BmxtIEkol6UzxoirRkdnb6CSsdlrTa5mOyQlusrRIYZULisyzxI6DIp
oYPKqyQxsc4NB45EYpq7Cn77Xq/WiIMVnnSyGjnTg011eTBTE2GbNEUGEMcQ3zr4wAe85t7Mcnqt
ZHSLJdO+3l9NeS1sdNlETqciDpOKJp6gyB7ask8J+xd+5ql43EKFjgR0C7lHBKsuWOJI98i8SRzq
2Fh3dad/Kb4XRW8BOAVn7khexejlFh9R5WMwnJ87pW7AjZqLQWyEXxe7GKNafll3ZRQShRjTvQRe
2z81HKZTjdpOZin3pUvQrw7CzEQx5fJ6hvebM0Wvo1BnLRstgEP6+LSleKef2NWmLeDMbs0tpzgF
WkoCHjZMuLZawUhueKgVbUirpH7ZX3RlKrR+kN1D6aoPi/43ghGPTCO0+ADL1iUQFDKnaB8kXQjR
7Qy/tEAQH8nvKmcBiigNfKPaBYFcCJFNALQ2dtKlG0DGYu1O5JmvYrun5tuaSxlziOIDNasOAS0k
ZsIEDaCJkCLECyoeq72+lE1C55hTnnN9URH190qLWVKDmZYQUocgeITf3Wz0PbPOB2ghzVzLqrcw
x6Eks0iU5GUReqdS7cAdY/EMCzrbr/pvID+ZGzFokSWB+g7uyo618nRaGWC3OsShDbT28hPbvl0K
PI70/xfYlswxitmcPXTqjy8KZ0oR+p548JDLyxou+4O84E2DcSEPjOBDYYDAgsMgGCxewPJkGTX7
KUvj+9OqFpp7GQ2vh6QSKp31fvXkwf8kKuhN5hmxT5JBPMbY9Td7taAuNF+eqNELimWbR4YjFHOp
H4qYq1p1208to3n5nM8IzKWZw4CQH4I43wEkh3eDUAE5TDQfm1DFuYQGQMHL7ONmVbV6/1OiJkiJ
iiaEH1VB5XFkycDvz41/1YcZB5gekY9+7bI9gqAJR9538AL4+uH2BxDL/ofQ63QAZ+f9SmeIcDzr
e4uAU8mHi1CE2Qw9c9/3GdfVWutKBA6l07m7Dt4gjQDJbhE0fQPbF03zh0wDRMkUpsYdCI3TAhvL
eyR6ROg4pVDoX9jfoBfL589GUAPyTsxbcIG6R0ogZuG8MtGnRkQ0Ggr/TKtIIFHPok5s26lnJnFr
3d6t6gTfJUmeACNHjejCh9dm+uhAfhIbJfouYazGYaC+VmKYlbJ0bGbnSjjpOf1omfhWs1ducZ6Z
vKX1k3ZSohGm8DKGtRahWFkBRkkX7NhVnVigg4gel6ROS/9Ll55aRv/AneM/jgfSgA66L50Sn8wb
0gAqB3an6o5S8QuBYwg5YozTicWhY2cGp3FVGayYEgX3aK730T1FEmwkjyV8O3sWariRtGAUxAhc
KDi3ZYAU2qbNLefeK1rRv9btLXRiEF0NXEHzo9NaK6uc7S5gh/aGKgzmgIyJMiibJemjbMqpsyOG
o4D6BanehhhcdkRx0hu0wWFCvRsd+21lv9LJQ0Ta44Mmb5CNJo1y+o3UEMWtG/6r6Y89A6bD5u2P
/PJCpBFzOsPzERzAJtse9D0x6vDTZBkf8Ta4QE2SYbyS26w2dDrA1q03XXv+Zz72kyY0zWgcwsTV
d2sZAyhpBOGnlmWLU9VSYsZcGCPL4hdonDkkL6QrnYSWG6ulITtTMKzG4DACTk8R+PULSMK1aZum
5K/SnqKeUTJTR3ZOOoiRqIdBzt5IZqNUwLC3gk471vyA5Nf7TkV3T4xLWgkp3Is5zrZAEK8sM+uR
OGmMUFZFwNBmQty/f+GcH8aMu0FEmwbEIi7IHdaSk62azVmR6QZD7+CIsoEYjdJc7hHQ+vobXQM5
7oYMm0xwI6vTmrHGDSFjGrkqOh3/K2gdK7Gawm6Glkb8s9x4296jFbsXdaRiNBV5T9BtAaHyTOG5
GQ4TiGJbWPisUVwK8ZbpquP/z8N8/SmiXfyOi1ro6Sf0bv3hmgcmSSacTq07pfzqDVV3+oDYoyAI
LGwehXYyyX0oT9Da47+fNgWy4D6n4v4zpRAHk3KB75CGazKgNcnTQdn0+WDVXSe2QcJvyfxYiV/8
PefvaoMdo6DBOEeYK0IvL/ba4MkZdo2Cnsm1fNjFmGpp+KbRrLIAAE7p4W1p1IBF79nt3Mat07cB
QLJSLeBf/wsX8iqLskFTT08RF8w5vk3ZOM170QpIW4+ltAPxaoFJm9se9bd8mzIRfcYCovjW6mGt
f9Znzmrxx6YhfRCLxb74IU8CbNJ9vUBupwsYyWLTY3JgYzxHs5XrjvYco6/hNilg31KTrgHkLm+e
W1B12pG6KAsQiczGvhYjpZO9xHYb5g3e07+imuXPF7Yvmt/PWi9/KHL1NtZxGsPgvlSCw4MiaOpa
eprVzEtt379I8MD4iZcPcEZhHmw2Uash3NPDex28Jogj7VTAFrMGYu6Oy54GpK9upK4nj/U7LiOe
6sqgMXH/vjsc1a1CX7KqhOUXd1h7DbgDKL8tEH1Q/0/ZP+nwXhOzCfxXivTkrkkNRVw80yID8GSE
BKj00ZeHKnZEKMIeP3NzYCa0wT57z1MVb/rQR5AU0GaQmuBrwsxEXmzfrcOJnKHgatFC6M9lnjFO
XcQOzhRBYAxQsnRgqKVgDkbBPjLGftckYTuG+AsBYtUbDFGNTm5/Ds+KsavJ9W8FQnOx5bFN6EO3
0EOl45H0MqkRKJbmOoyVeWG101YEbf1vEbdyenoqEtAX5LTv60fnXP8ae3hbEbXFQaBBOZO+UnJs
oNSnuDLwx/5zhB3C7dayZ4bS/h2SqpO/5xCMu8YLIlVDJmvpsMyal7spMJzrUL51YlfPYM+dLLC1
Oyt0Od3BY+uk+9WhhcC1nFh2I68kzpCZRXzxkShMcqBFC4D/BDJUTRtxoDEQvQplO+BgnaGjuogv
BQ2W5gIbKXPT3DlV1Yriy8N0WDN4Z2jsxr2E2qNFAw4ikmO/5BOmJ0eIuiROjRuGN8Etx24TAbkI
bU9iUlIggUPmwL/18i8BmGC71x/PscbnbiSiBHBdiHhJ6LRA6SPZzz3a4bAnQu8X6O16WlLQX2v1
nqhS97t2wIW90biUt8xM3xrd1esxTghqxkaCMPYX90ve4QcjU2zsDdwgGudvSugYFolF/8xk+MDC
fu1HWP/jEBcpgY0DeuvCPUMS4W+ltmTGrE4/egtMP+rpwp3mCM8eKYFJDbmH+gn8xHpWg1ESbes9
4KlPyVX3boDaB/L54N2YinL5tUd+anLfrxshbd+ajnxC9UuNyvnwi1LbNHr/fQKVPe7Mw01boYj+
w0Wp1jfEAwvtUds05TMYmCKYyNzv+XffI7n4D7resSoA9f9pj6r8LRWBwfPnexHOuVxhgu11DsF8
QTUBFP1WinHnw+IMg4k87Bng2QGdFHNTuiWxu3JrLRiC5/+dvUTJG8Ra9F3FAspHDPrL0m7WZ7aB
KcW7+zrN0i72ytUzuB5jgMyS4HBOm6KOGODzz7oSBKLRJvoftnLFIWEZcbsMvZPFsCCYKQz8Spsc
477MP4O+4DDw5Ck1I4KkZJ7OfQ7vz5wA/BlH2sijpFU5xHAm70pqCStaNa831xwM8OGmNHs0hZY0
BG2Bars0u1Oyqh6ZZMEUdE8EyrEbaVB+hrXax68R2kREkR29ShNuPV4QaNO4k3emTivBk7LvTNnt
2010QZ131Hl4GRDy/02mzwjhsWR4NNUKiUiC13PsKA976yj+bakMslPZm0GuMF4PJp6J5iT+viFo
MuOD6eL1hzFREkO42bUs2xZ73Wr/6UJ2pVT2JPsAyYYqizPXOPHoMcZrCe5bDPfCArXrHI4nilbn
NAdopW4g0d7V47/gIlleKu7SJUAqpAXqHbQw1G6lA14Dqhx9FnBx3Nl7+eXrR2bZieiku2O8ObzY
20uiKam3VIfIPOJg3lgtSrbwXyh8T+gHoz7Nnaj6AX3oYyiNRfjTaEMIZ848ZkhLFaBMXybxDMo+
MhqTDDCjY0gkPwYnEdXWA/qcNZoIRSs4kakF/PjBUSD1BsK4OacDjQZPuPKhPaML9ux+regsRnE2
7pujDSbVxsTeg4W40dJ7NAcweV8Dt+DamAisOhKY2hr/JqEKdKtuhhSwrMMbWGz5D5A/mPba8kzb
BOI+l/slfCueYV2kyob57WiBFIqiN1ugpLbpEgst8Pefi2YoiX691WVDnBUFemGYurt4ISOKJ0lb
86J5+QQIv5zqCLXZFwx8QvCn8cJTDY4qxEvK/HChjZrxrOE/suWRc5jyHRhl6MmVB4D4ropXwuIG
UAEnXAoab/XPvpJHY+uF3a9TwZ1d/jdaaUCZRc6Q+9rkk3fj1dR/FishlIA6fSGVBYL+0dkyRFAn
FJsfWLeTAUKu7saYNdH57ZStn+JUVOCRTtRoDKVFe5DUC9cr2NwpNsqBj7eOsbXxNMyRihUZNBXL
dnp+rT2OuFxc7hgMx2FIfctuR5LDpy8EucB5AfU/6GTmR5oRFmUfC7GyXq0wIcxpRAI8glBylCGr
EreeAb9TMwAqBYOoVVaC31zz2HL2MrBXe029OotWGmzzPFCu7k8l3OydVcP0HVqgLYlYXPJPuFVa
NiqHWYdmskr0IEsod6EeZM2UXGGUYY+d8bBbjg5G8Yx7WAM+GWUXIt4G0DKVG34S0PTokEhyFUUN
6jCI83nbo075KBuIgaj7mN27wQNNN4RVYf8saycGcKfSzAfYTQrpMksQ/KOCq0QwLpy8BqjVOo3L
ewoIS2DXu6CLlpsK5h/maL3hZTIHdIO87Jud4V+4eUOjNklU81aGfJ/YA8ty1OhTZmYgYlU40hxX
CNvDe8GrXbWcHMJ8tXt1g+j9DeBe3TpU2Zbo5/0EY5HPQ8bzmyxsMDA1vW2KosHW6RxKKcPrFOgn
k0SXG5WwBM9SVs3moU+7I9Xp0Le7Vqc1e1kOlakUe9eN4bx+V0v0XVduvgKUkjfH3plm/tkw2oN3
8zfChXObfQPIP8fxTTIVpewb+cxBb8y89XwNu5idNbTlJdk9EriXC4ZnG3Dr7MBBiptnO/up8Qg7
O4PrVoRN4HcYEPJvuSlTowDbOJh3/fjYt2yBM/Vwax6u/kCl2yVxD8hYhiJcCyDimJudZIA/e6dM
N7bT3TgD+mt1bp4KWgpJwgSGk8amMUWNgk/Qw96tZVkkYNRHStOEHvvIUn/BkU8u9W6YTBz9NVk1
UO4XdCEBkIkBmIwcyKx/UcETEiy+Yu7sOvw1AFawRyWGBklXlr0lNpWLHEAZvLVpEbWWpCGQGEZA
l9dTx6ZLGL/xYHuCZ+6bz4FR/jUaDDCYQLpJ+9lxmrwIRLjM/E57wH5HAw+XsJM9blUfnE6Qxp5c
gbzBoW8KTQ0Ax78e4TscQHPLCodqaBMV92oQJOwo0+8PgSJHgCBfNAuzOiu4VjVbeH7eeRVsVWCD
ntxDkpDdLI/l9KiRbdrnUM4C2rsS2EdikhOL4z9Mq0yk1gNWt6RH6mvTZBkh4bH1kHSCLrqiCMgt
6yyzqgqmEcRjdFO6y8YgZYy++Gez6Wy0QsBnqpdwXkuGtRNWZnN1TPHXlQV4K5Pty8p7/oAD3VcO
1HcUHuO9lpQJAsAkCIZ5/RtQFzDbR5pCS3KvdgSeyExdb31v6FpJxCJ0wjjBJstc1zKNxxNGF/z5
xsFDMOOAYAJkw1N0nR5dnlkVV+6t6E3ZU6HsX6wD2w4JfUwWbP6GP/0qs5MTZPfpP9Mr8n/bx930
iZOiT82tjyotbwTfZbu7nzXhoHlaQkyGjnHa0RyQ6/sqxvlkQHCMa4ksu469aAmjDfFalJ1zefv4
2phSV8oHsoGNvaXCbqx10uClDm4sTfT0AeCLDXScRad/V2lmF59a60HjzaqjSGfMDM6XBMgvmeXI
Ctm39zNW64A9YCe3EZTFcJHgTO8/RwUrFJ4rrLAK48EofhsLfX3rscKNMceEyCupsTMa9yDXj0Wb
+HAaCcDLmknUUozY8YpIoPsHy8wsOPbKd3Zn4lwbhcjEYKR4ju9eBx2nbnWAA46BS71hLLCt1HE9
ucr9gf3V698b4Ax2A+PzBD6o6pd78bP6tBmeyu4idwGtzOTpk8mntPm91FHKjelsNXv7LfD3QHg9
Z+PyBgVH+fZ+k2VhSDP6qjck0qXvp7NulRzdFoxWkfg57EBVLlay9mUPP4hdi5jM+eakY2vSmGre
m0+2Mr4+s5LjpD+nDQbbVXa4sqSf17BkkPPFw6hXcAnLxkwwx4tPg9/6zD9ylmuCUfMf9+07ETzH
xSgizNcIQLyQs8TItB1kjFpB1IncRfsX5BcV+1vQUe4M7vAJghw1SfpFg4Gx3JixU0L28GZLjSQd
DNH5F42scan/Uw5R5/D3tXUoRUFdlPAzI/fS0gcimjp84Sax7FMUhNs239Mh/xEIQlLP2RYVlr/u
Xs08Ynhq5B/RJd4OL2VtQ3Tfh9Qd//PLRGnuSNLzjgLOoZ4Jv3xribn4QodaRpGy0UyLoayM3OOv
ZuYFncynR8UXUS91G/OeXbilG0ppOeft9fpkgkswSaFQ0HBDe5vREkW4v/9WGOgjCWY5cy1DD5WV
E8b7DkLgEN4dD4E/OBjIta2I9tR7f50WWaK66h0QjNGz/SBbqTlP/y8xhSFaT9hdJbser7lDPHY1
3Zbsd7KB270o+wcVoIlcroFU9jhxxXiANltbImYQW7mM4LKSP6syQgGpdvRwBFTSX0gbQtKcwSBt
werEhJmGIq3jfQTQ3KHEGvC9x3A2nMNdsvcwebsQwzsh8pTnA8EuPrF64sod36lx/tgVJEARu572
6c4azvUg7wUXbnM3qwUxg8uEueN/b36PeVNwxSCRdgwg50Qs+GGHRQJrUk25D4lNfjkDcvIQ7O/+
TY4iFyKE4KF6bFrwNcXYinAWMhzl3ZU7VCFO/0XWsdxYOyO7ZQ+JAenQkn187FiZpyC/lIOAFV0z
WS2GMkqVoMq7cmIeh8zua7HHSn0+uO9zi7/hlIVfQxlbi+9w6Iho3ynSveK3H4E2e5yjk6hrqIc5
im625hRzrEswwux0SAbVU2bpH/RndeFPDpfRdXWJvEamWMa0GbW8AXXbUmiNTZk9RUaVoxFRcGMe
zrXkEQBiWWDNvo7YsgW5R4nnexrHiu21zGUVaz4vqnvlR+OLkYu+wYW3bBwAcXlSAvWUssahPp3U
32tirNix9t67yYeFhAjbuG8kMo4yX5TTozhO5w7uYgK2RcE7XebDmI/5ctp8rFAv5eLIhlrGIcQk
+azn7JcYsq9Ijc6ROnUiW0/1Hb2HeeXQKX1iDzRfj0mHwumY/Dh416Mo5EJKaX8HhOcLh4RuaTfH
ImfFcH1IcKbMwgtnoIgl8W/VQRsfsspOaTVAnrg808Q7INF7nStndwFPRzk0lGETshBCL4h/NNl/
1/X36CkVjKDG9PncZof+JZ4CoDI6qRJo71AbUa/P2IyhmDeVZylkgFYkJjhpJwDeP9F4lNsr1LG1
mqqBantqgK7uBSVssyNDv5kCD8GZWU7qoKmKGKilEAHqble44tUCCln4xp2RZLGTfdD9Il58HhH8
jmHvMn/AbpCLj3BQsCYS4kFWHZS9pA0uvI2JDm65iAyh/xw22pVWpjGSmqObdq/qgyH3xgESb1oL
XWc/aZOT0CrL05NZ6tJr1bXrAtPHaXvZKbLv791rpotJbp1LOcaU9/2q+Up89JyNpmoFuESGlaQj
j1fDhc4RXszV+kX0qfRA0+0xrJUKbnoUNG93WYYdULwTwsjj61gz6jtTyj02D4Xavq2N8ZCKmK8I
prtFzs5ulxTTJH9sGFUWr4K6umGC8/AzVtBCadILNwCT/4XfUE0GXC+VQ3lvPWtg7gThWwVC6XPn
ZfcE5jF45UeQzKhWc0eAOQw0KYlEyAj9AzgPddRsRxYxzMIUtXBc6pAMqR/x2eEveExdX720Zxq1
1YKtH5nDf+aWK2TLJttFO4sigDKXpR8cSkqWKFeQjs8f3EG5whs3kHFnsGMz9rtisv4edAvWMG/+
lXdVN1SGoltWgVZqvfqvgijNItrfY4uWDn667/FraA/cbomp0KYq1Y+stLUw/1dQVJMnO1n7m278
8lGfwOjBsgZJGc958tRgZEV099cxs5RQWw87OmHRyCprWMZ0Ev6HDqYrB8gpzLjmH17AYF/DWeQX
v+YiRjfn3jJkdxwO1AYtJr4JsL3H5o5gcXhoYhVDUZ4JxxhtQl9F9oETCPdDCkAxDhAMFN2P2KdG
FuFPBY7gcK8QbZRtlc9zjGtObXyHu7joi18Ma3pEKm2q4sBYeqRvOgif0VM8wLTAM71Oc0fh4OLW
3wNKm5K69TzbiGnGILITEYriXFIaVZ41FUfoJuqDMP9L2O0jj47h2Hcw9EkrSiV3rs6zuGEVqz1v
i8mDVZbn6Iu/s2TQ4DGWwPgtDmN0VL9n2kOBoTZKo6fiUflXw/LKy5tNu7UD1ll4nRKAnk0zHmyo
k6zwJcSO2I3SnRB9UXnHA2zb41avHj/An4ScRHTJiIqDhoyOVsuhWWGLHAVgbOidvRwHE+FSvpqJ
/Y9G0JJOqPYg5igD0/r0l1CO3U81BtsaoC93Vkj+W2a6tQLxkWke2vLDoEqEbvCVSBu8W4VSIYUk
dgXVwKHYObJX8LhViY01sbcyPLjsz1A91CKELrKqBxwYGvmqnBBNCQzIfkTBR4Kz7CNoW7ZhQ8JL
dTNwjwIOSBYnXFZ10S3igBtgbLPtE24ySx04NfF9KKIFeeueQ2jmViOVsH2k2Z4hUchr70jtx1+l
SQ0F2ADJnOcLEOsqyvfGUonDuYxSYVeOEAWv545c554G2WqGDPYJEk7JoYVG/wAO/Jy3G6dVqdyh
qR6vjACDMmuRAURUGmTuhvSYd+l1TMx5rl6KncL6awgtlrLFFJ1XVHN0SBa8//98Tb3wxE5DNCL2
nVaAG5Sknxx9te4Wb8FUXS/8BMtq5gJikXBea0hsITsT8b44u2+SODevLquRtM0OisKr6yiQmt+t
ocWMaebvh7tAmusn8IUjCV6HYja8QFvvBSeQVRLMmZ7658GxU+/7msAn3ReGb+H9MmatTeX+/83g
aHMSC522qqVCJbduUcxJK+5wSEExNm35ZBW+urUOva95HEljtnlMzJvQvGRxf+EaWqIz/8kGwA7P
JlgwlLnF+Xado6/v3TMtdAw+LW6j1NnWH2TCHBnT2sXwxbhqo8DRVBii7ITX5JSm8OML2eJv4CmL
ZhJZezd+RYiyfQf9ZhF3yB6Prg73+IbvocD/2lLHn0i3h4riSxJ2qv72UG9zij0wZdWK6oENcFPM
dAJGxg67HPcKbivtYlrFb24CxgOx7SKbE46pzTTQ0tkLk4t1v77cStM8uIXeq6GH4m4ewmVOTKM3
AWOLlS0bJE38EEbq2uVV8k2+AngnMRFmvkiEztk1PROJt67vdh1Je1urtOnNHzf2Mm4L6SWjKjxj
jsjfu1Da3uHYjFYwHLzq9V9bXwtt7xnMZXVBeuvCCnBqdhyPG6wxmyBpV2ziTQvuQF4D9HMez7O5
63PQNESbW2DOWnNuRbwhg3lo9yIAMrayNqyaDAAsdeO/cdwRoMq8ckum+m25ZoWfVbX0mfRQTjrH
MyapuPdv+wuc7RfYiBnyPjH/tyonzQuHoe+XuRM58Lonl5VGOXOWig5QHMdGw+jbwuZ1sfX9DC+s
8I0OTjexAHFgiKoFrnYjKuaj9Qjl1C7qg4nDp35gef8rMPPOj0hYaHQYdcwFEEaKPfOBSdKYikuF
EpnHLSLKYeaoiUUvF+vUG9n2FPr09hZguPOAeADw9J3N/UnjAejiMwAbeLtpRHtVH/a50WJXLkq0
ykeovpydvo/91asbpASaZnaRolyVWxE6dQrxdK5LRTE6HBWwzZ+EzHN1PwiZ7RtX4Yy1CLFA2ghW
vW+I4t8GOf8UZCokFabTlfnsGfq9ZLb9jD9MFoqAwP7gAPeecbCzV4PWLudCdEGnDjBi1PmLrk2k
mZ0K73t95eWy72U4SviXIpdd8Pzkk53XnKsvPn3tW4uC63pIFCjhCwzvACqiCNm7Iu4O+ICD4feE
Y6sjG7usZg8d+21IBWWo1jOM2zsPgC2crWUq4U7MkvIFXlKSlkPz+if0d+qFCku8HJAL8lrAyWAq
P9RM1RyzRvGShD7k03h4+st8t/XA8ZeJdM8NawKp57lmCp18RgolYEupWQGXe6lTEWAWuS+KJfaH
BYfYHah4T0IvmTV8V+cNE82PEOhKp0IPuB26hY4IijvgpuXAldZyEkf05ZzvVUBnAZkRWNCkuB2f
2CpYOziSdImZ2rEn74Rn0N83aRnoo0374wTv8hjY0KHx0Lo7jEizIle4ujICj2BVE301hvUomZrB
TQknITFoIdknfeUqI82TC93Up8ignK3wDZPZVED94hAKuMymhYvpfe/+Y4eg8jE/IjBChuW3bMUz
boHI1fw2aY622upC1zEybCSPvM5y7ZHlPwABtLi3OcuAeiZYzsGEi4t8DkLQUjaADj8OYcYVRrhf
2d7LWw+iOFTB74nlkKKRzEjbcgTnpBEP61LKebLW3WKg1MIwkf1T+j/1YEh8vOEhMboNdbuIVtK8
mX1m4xb2b9ljPPbRLBR63WvctJltUBbut3oIkkRYnpMJMmbL6/uRolcidVLTv5I7mJlvffg0OmRj
3c6KobLbNfxMjVAGAjN0uHlWMtXwhoHFKiSbUM+7MO+e8WjYGxTKrGH40JMgbwEGDbbpkOBh9Zni
QGkt01H6yR74eEDwpFw8D5M/KSmccgfGwS1ZF5a51rYwUeQMNQJAxlb0aq7aIspJiISr3oGs2zg4
rP39Z19Gxe9kojD6IvfydsG3m7ypfG1GOVlm/4vBqlB2IFdw/YcKF/XIRTzXj2AfVYj33e2uC2Ht
1LDCwL0YlXMcFygCzt1yKR/EXM/OaFzJH5nGHjuV4gFfUpFDRbR9n7GAsYYEdLTMCL6P8MeWJ2ri
oU7YTlkcFE8u5xxXMZd2oCLWUwFOzuxcJqXKO6oCd4YZac0Bs/gQDInjtb8hzbiErNXLOhhnvFxC
wlCAZsoVZrzBu4y0D/Si8VPI4LVf7fBD/FrT7Z1U91vRv6v15hP6UnaAKsx467g9JX55rkF2ZpHl
xttDZv9PgVrCs+l31HcLpjXJ71kEqc4LWWxb6oGdu4hJrJVLL0Ad0BrXDbAyoXzQAe4RYz/gCsIW
l5p8O35DBJnUWx0MJ+Rmw2w3QsLttkG+JuJOolZxA73+5zw47WkqbN245p6CUpqQ2q+kQlnXlfq1
uHkZcGQWCJBbHoH9bezXKfvVQvMJ/WJx1rFCxZUaReCrupOPng9/9IX/wU9H5HPFqFWFNuq9WvvU
lDnOYc+W2jzrAJ98IJxIZaeKWRkKKBd20cWnjYmOFv+A8/tmEaVoHPTM5g/fTrjAyobddnYP01wj
W78dRQ7BxdkkD0HUpM/2Ve5qzX1S6wBv1iBE5D09cuHTBvzifZjjOP7c6U8uxERs8Qpe6V43a+El
N47t116XYuNNlpUc5WHRK4Dd0HZJ3YnIHAPgO/SbhG1+JWLkaggmM37blOhURvCaKQ6ubIhjg85N
Q0v/8fNoQyvqNszmaV3lpnTlgJB/h0b4wauSuQxOm1prjXxnpMYGI7m0rUZnio+fB8GMxs2qXxDJ
hWfEvgUzmyWTGERQrCC1erBkUmEuGu/F0+DoVe9QPK42iR30gYKddlQJCnKGd1gVMdOyNN69ECvL
bXk3dfvoSj/mtIY9f4Q08YJAjWpr7PgLOW66qusH5i7+MqK+r9FRunb7TR6HjleJ6NTU0lCAijbY
WKZ9gmnyyNY/24itsBsekwfVyUxTMwV+EPyz8olG0qp3rkKdo774fURKwf00S0jnIFTdVD7iGcRg
kdPEuO5IAQEjjfQjjS7b3fmH6HFPkG/TpQZoB9KeXyMk/2ZaybieTbKJF5wZ9thfj7Z0SHXewFrD
PDMS6680qAnkZOBfueWlo+qnlqiknSuNx2Ni8v7PBzKoIBeQRrP5wcZfb6GA0TUtTUaDPD5RjX3h
bGbD/Gfi1hunT7Ed+rG9I77Uxjeieb3kuTe/X9WjbIMbJc5jCdGNhcz3syoEtqVOEhooYMKaVElg
ZFEjLNqwxfTCgmOhtp7NNEeO5PAfZtMau+AJ3pqZMsUNYCWsypaonjvgQnu5Xd7/d78xeFfv0C9i
pqmmWm6kv11pdOoNLS1VNzbmyr8sQB5BHO9rnkjn5X3MEA/t8GhCVt/k+EAJCnUo87NhPTYRutkw
kWqKSqs1QwyufPfbpnKQnzLXKswMxHYACkV3Ush3syqUr3Kzr5Dgwk8DqPUdOgCG+GXRoWo3U8Hb
O2BFy+VR8T5VyawY9k6RgbZKlzKMPbpHhV4FM/5APTSsnkq/sK7EkZO1RoGtYmiVfz4TBDJM8HWd
mLDlnAYYDW0B8jywNyq62dTc9QoJJkkIiyPA291bDWh7Gnzv06wGiZrm67789/tXgjREBvbzquo+
Kw0AIobr+6msj743VWqVQfWOyIezCkTVjsuwNGxKl11e2lp8ys1TsvKHOBXQnVtDNMTxZ/rXENR0
zv1fm7cgxinUeJAoUqIqKQTi+qRboFmeWix13T+/6jI7MmfpXtqZ88/2Uz4BbpHL4CJOXow36XBf
Eq72BpXLbmx93e+3ewDGT6iighyEbq0ihO7dnnS01Vl2dppENenlDX8kO84Y8Oju1F+45/rFCiDk
AUr/QpPqsPTnPkHPzkPjtmDkC/+TWNV8Yo3FUAkErhk0qVVLAYy6mhtEIZcM4Dxsy57nqaDAKhUd
HHP6JSbJlWx+IDtyRmdcT+ADMxl7SmxswHPzLUNMqTH4k8zomofnmQ+V/tWd34toqIhVQwVztZJS
wX96mxY2dSlFEa7qghKiEz+4piClGmcmGpfBTvqGnQt5FkeNgLVwwgdkQsYShsw80QOij+uHy2iH
jJo32sa5rwFJGMs2YBpIClEQ2ZbsL8+ituBrZ9tnJQFTEtM3imIJE6tehJXOOW2raCA8mBNYAgeR
xdhfbItEL6Zln+7MXpr8p2urGJl+Ou6ljNLFBZcHzw1Ulsii6LOws50hTfqEmq9Hctzu6LV9Qwug
4wgqkIYmHLhh5M9J+RPy10cVF8Hmg7lNRzBSwvctUgyWQ+g9JqMXvQ5EjmdeXlh/GLElMqsRKG3Q
BLxk5s+Bu0Jgo8BFtUcIIA+zdXome1SwfiehuCvQeA/YeYLBtXBEKjFbNyg+mWNYtrMkBuF/uv/q
JjWGy9jVP155ROLMVEakQPAoYsRbNgcNm9BDCYYWQ8ZW4Rghr8HfG72iOTSqvlkROvjQrwFiwrX8
/oddZCElRQjCFAq0m2WvCULlJb3gYBMSNofsbaZaTT1R0OA9w9QYCglq0JOVKxTF6e499xEnyv9Y
iItgKmK36TcqbzZYr28aHaIgi9Af3DdN1ILCACCkDPCqPUxJ8t6334Yy4gwFPYfHrlbyznq+d7vv
LgZFOJ22sXzLxorI6awVTPaBM6r/WNYYqJTHc9m3Gp175XIJ/8qvfl5SzqYtLtYtJOF77E115F/l
liRt1Sk67TQCIUmqCaYohNjLZ5HreJp+oW4UpTGZ/YUk2/gp6GCMugkObb93aChkE7ATpn5GLFrD
LyYwORs7uO0hQKDOyhExKvczxx4QHZt65YGvFol3nRnMrxd0Pk0874gh0CUlZJGO69VpL+hklDyh
Rg+XVSdalZgWS5Q9ZdS/YweR1OcbvrPzelGUnJffe+gb6C+e9CdHOVLMYOCm7Tc95SHxp5t6geTQ
cgkn7OfWmV9vMMv8wEx1T1BWhoKcozUIMu188HlVBZUSO+WGhNvAmRBJ7eP6JA2y41OaRqZ4Mu4+
J4hxYQXCZNHdqcO2mhqNM5O7paI0ouKP/Wxhnxi4nAFtY94isB/l5DfUfKaOkCP0Au4MoL6ta/qg
95W2oiO/EwNBqPzVxROD0SQ11TAbupU/vvlB8As0ORCy3gbPUuaUVNhCk06hSshgEWbYSWpNLJnM
RNgBf2wc6IGSL/ERGNjzuNuXDCckKE4cR2jTPdo8RE07721WFELTwcdKF9OlrZMVbXmwhRUhopr3
NaZziZ1dyYxFybb/ltBeYvgEkQszm8xuA01zTbQRSgT2GV6lB9fqAF3X6HpBXwazyMxylQSqlbM9
ycFneatGCh6HCquGahkVBYGZVqeIYnqaL+ujPskkUqgahQn1zCOPR5NHhfjXloWTcpPS41YFp9s9
hPjzsnk1BZw1jkiWL2vyi44XDWaYAKS1WejX3cVA7gIoTG+wevwC/bsmJoYsosNKbPKhaICNj2eS
Ty5nH797ciVYVgEtCxNMP8myXq6X94fP5w67ILXOL7AL4rW191c7XBrxbVs+5nDae1tGyqgP+/ob
QabyK0KWtySYRQ4AIgmT3untjv9aQ4su1cGFp3henBlwb2Xbyk7ZQyn1JiebRxyqiLKFb4u4lUX0
8gOH5UDakMEa3wx4h3AAcpRiN4GlD/Ss4gtBtBDNb0pklSuIS+ox1HAP/h08LxK+1VDAE8/35ze6
hDWiS7rZAm3LIo9km1xBVHXZ2uHPTKjHZu7IXe7PQkETEsP0mkY6vVXaR+ouXxZzLXe6hpnePsK2
g8rLn1ev8lLcOBoqRnJ4vEYZnwvv+1OqJ321pdgBv99JIV7++kiUcclRkeVfvuqYN6cwt3X6ub6n
uIlRXYBQpln992tyswxfgYedsGPl1pFNUZQMSOqKOe3ZOeFDmbhERUkRzRP57v7CeLaN8JdondCl
fYCs5RQorcd5kY9SBcYcaOA+D5NtjZ3QJ+UHPPnMOOAajW8zSYGdip9tdsu0dHcHz42lc/mr/77r
Utcx9fWD7cUKmxhoDwjBp7+S9QQy1mXJCTY7qDDGYrUytEAp3SCY2a8wMHclMK9c1xswyzXPWsxy
yzUckISADV7AHfCSVAhnGf3t1efKaMUeCK7AUrNFALGATFQ1OACilIiZPuh4DK1nc+RstfZBx9Ek
psTg29qs+0n6NNp53FHXH+52p+JxdKQlgzkVkE+ZHvznYDC4jm6H3pOfwVKh9tS9ukzg5ah3wIDa
wX/+b6sIIDqmxSzPqU8HTEbw9Tx9WonPVcclfGrW43QB3yqsPOXgKPo8KG4eIwLfJsR7g4yOVFyb
vDOk5niFzMZAP/Z8Kdoa0TXs63uCxvs3dEYldkUrRD5i7j40EODR8EydcvCKelkhFzzDlRfhUE7I
jv9pe/iFJePjf36LWyv+dKUgJZFUpow0d8kJJTjNtWs5CwCurE4z/eOR6eQIJhaz3FJnsnq3J64t
av4w60wzLOFeRiIiPklQsi6BsNRuHFoHCDXOW1eA4wo/rDffrbn4lAExD/6pUbKu0jbtGltIG09o
SYM6cG8nfCmXgIZAF2PO2j3RipbAbB7OMR8QnXT0eYpobBhqod1yZDwI3oQNXrJaDgT2b6wXqglZ
7Jvviih+lhDwYTbHsMlGqN6wHobRKsa8vcbDiTOfX1TlY3b7VFo4tR2VpOEr8FeSwsDJeq5Qs2du
5ckaS1UxjgmnWvfHcXXorqqzYHZ93+7btEdttr3QZxv2xHco+AaLwfP3Z6XcHkstunvP/406yQUh
NNaWA6IMNpU9UufORnZJWKUW98jDO16xnQTrwdR7hfXMOydeSSBzpOhrs4rmC7DigdmbWZz9a7rq
wUUkkbypljZhwBkZHmYAg8dl34wWl5zctE9AhBca1RcZbfbAl2tb7fPTA2dkYQGMOmp5k7IQuvFx
tG338NWpwAjPIfuyZ35mSuOksRKWfApAVc3t050zmd+8c9h2a6n8rEEMDptSsI3Mz+vOq/d2RBUE
CcP+YUYfcaFEy77ZU6MMmtO2wWrhU1FFOfVuSZaZ2HLDWtwhal6t9yLH1sSOvUjMfglrpPJPTS7W
injHxkLPLFLz6AzRa6ZsF2j++fy3eV0YqF6I0QmiXnkHWUuo4Mr3ana3AjJ/EKUPlawuFn/JBOQt
XNECYIPlmLSSZWOt9Q6jSwB6D2Y8yCvWq+4Y9bb1u6OOLzErCLni1J234o6ML1Ql/Ca6FQz4N+bX
xYfJOWc5qIzmOV1tyKeIrVsieZEaOIf0qRzSsX+vJLN8jisTAQoCaElXftt56PxMGFTdh7dHVkj8
Cwo0c3qKibnxpWHCoe4CUUlpvUn2dMYlz1IiS2O+GrZ+ugNabTtoYoHO40vo4rEmqhc3Q2dJEqEm
kd61C/5KRWYUi/TA2bkgDSMeBjVdpCrwZ/AZ6AgxeEFSNB35tJNvn4bQ32F1NZVkE0pCG08WmXzH
aNxDycfh///7FIdr125GQwFrpbCLV7qy+8Jdslpy+dW7epQNr6WSYdis8ZjZzpWSNSpE8ewR8FXO
z2l1mhwEgWZKEPGNKLr8HfpGxNY2t0RoUxpn/sFow1yIx44xv/YaU2VRkxmF83fbYEsPzirLIic3
JGSr52Am1PWaTJwYJvOB8j9Q+uZL9MvBgQ9UT3KdPfjcmq+8NOwHvJi/T+Mu6Nc2xkvwLpHYLSu4
WEpI6I89+zZ9V8kUGx3lbaW9+GjEuY1/7ovsvogzAJ56ranHJCv7tAfUDa4XXZb2w1hYcgEIrdtp
43LPR8MsmPdpkPMf2xuzPMDxKHCcLs+tTedN5NEyMmlAN8PyRBbiZWBt2zv4qGW3ZPBxBj3YtAPr
tWceFS5E62YZiJDI+huQcQj8Ar8Rv/My6B/fbMabAVvWg6m2Ap+dada4GHM3V2jnCIpdDU/DLbHQ
7XpP0zUz1TdPjUpgBlzkg3zea+dk01gpNMJftgHyeUt8+MXao+rph2QRZXLd+662YYMQkPOjNthb
3lVs0JhQarwSf+aWVbwco7yol2SnbMPU2/c1XQD2uglvxhjKp6r8XGqjtzpP3Jxhf2F61vQfZUy2
qcdnyMUfst9q+NMcNMwPsNaOMybPnayxfFZPe6KKqy5eD5sqyT5wl4v4rKeE0Iu3ffheA9JFN6yC
4C3kigqmUBU0cumJXoK6SFQoyuu/ej2MwYxrxIc/CvtTsF1aVudLxbvBotE6G9Kr4gNolkobkH00
R1bSDOtV9NAW1fmAAHSrA1DVe0IFDCfWz2HExf2NId1L1I0sugfKPJ13ooFlJiCZzplnzi5ciOl3
HZQCpXJT5/evEngT6MVzliSuYCpCsi/Yp+jUXhdUp81TMt2uHV7zHeN5RUSl2Mxl1Lx6Zw29TTax
NFPfKg+Vi88Y848BXROtDZwdRiHGdisknZJIZzGQoTS1hb4xAm8z7nLIrymCKVHYfAmfftHclXYR
HQxvCjPS/vSBjSPdK+eZKF09FWdiWrFMqfMCKv1avH8/+CGeJfMD69e7Fxqsr5cbM8wZlTRNATQ7
qWNqQEUa8bU2n2/hPPyfb1VXpLDA4DFzkCDfMSfdYPHgyHSsTB0drJzMLYSwenziecE5Nh9ZudDq
tByufWHgRDHp6SufUCULwdZCvtc5ZCS+pzOeH5+e9P+ZEIvC2XRBzckQzxzMvWiiThwXq0JNlYKe
kKDRNgdQMxnrOngjk27jL7cyyQy/cGofTG+s9gWfylTGh2qNww+T4EbbDkpC9euQXO6szIgXU7qa
dihnj20KpSzbhyLeE8G60TtvDSYfU/FvEYX+sBmHEQxe7UQopJePk5we/TTUDykZhG43VI/wLEcH
ImblVruUTdwJDh67IaGSn2FW/T7kHzPD6CyYMRvQd6Wx1XhsOr875sRP1cuuD4AyvwyKSf11lOC4
VS1bYYeYWKFCE+HXte6mAKydxK4KzfFq6oM8Sh2gvqGVTMfP3p1cgxfoRAeJbCOntu7nz4hLuKsw
DMdKeFTFXy0Jci/WQ2OkSFDRr4egXAnq01WzeVKeJtGSpDo76/KWnUtJM6/RlthBlwCAEhYVdVJT
r8tzjvpjVrms/DB1qGSiTe2xJN2GqWFYKLumO+nbGnfiUtTwuCKwoERESy+dNHERD/k3tMUL+0fr
HaMY08K2bURpAIAWHfz57me9Dfie8VnVMr9kF8b76P59lrHXW1r5sihPqe4vRxBS+qGwphp04TOk
fBTYCvKQD3yLqfuFdWlkim2TWZvjZdauHLwrFqmWM000Cn3GpC/Y1wrV9sS20FHFLwQWR9I54/0Z
AT/2DWNY7P0Dx0CdmiJ3SFWTrvugLrQDHCRHh1zxYlt6rQPSJC8ZQzmBUjlAY9oAo8tRlOSHkN2h
RhVwERa300wdrvDNzjdg5Py3baeFFekhetDExiIG6sPu5T9vsaM03NLSQHLUiUrQKpuQ1A0noUdD
L8fxigENgE70sfzZXUt9K08x529dVIzhyR7Tw94ZAA+AMtCAr8vxiDtv2zOVnH+x1F/Ply6XhIFW
t55J4mzrQLgc57uNqBLEvIIfRLf6z6IjG24LMPzD5FHBCbMHtK4JCNKH0lqiq8w/7Kv+CqySkcvy
VSl9OTJmqv/M/GThExAwwJaOcWEEMnLPwK0sC4otKYOFmM2yc17AAorz1X5Y7SmKChAd1aVmfm9S
sUTct2QxmZjBDWHa6DicVhv8khyF1rHWL6VjFHo1NMgANoxvtLxddW1ZIBg00I6pAHv+KKtZSUXA
R8KwufQmCF/0ueVJteUnTU4DgPp+e0uZquVapQbRJb1+SMEDAn4KrfZxLZwiWbgibr0y77jbpg10
/s+K8qKbdlQnip9tFHXRFJUNAt6yAUZDLw3xy2bZ17B0u4zq343GwCp9HA6D/+FYsze9jXSIB4Da
e8oB+XLHvvtWRb7JTInxslGeZIfcMJ8s9JlVLsHAIR0aYRRf9exWweld9NOqvLysN9yChtUy4dsK
2QOmx+zpFF+XOdEREVFqrvA4Fj83Nm/5UU/+f/K39MEHVBxhy6yTYMyCR2Mv1zwyDFaJfR7c+RG2
3slqW5t3zIJrf8jbDBemgoP7IhM+7DWcwzQt5z/bezRRHTMHrCaoGITljIVMO1SvVRAImr74Zuf3
skGIBNtASEoioMVdpo7ZfcbO1IXXM1CArvM4fFkKpRr/Zym5wO7ECd+ilWh5mWuEPDXIiDrymrPv
useFLu+38b5D9GKtsjUehTd27T7wGSqTRWZDFq9nzmiGjBJwVgFHMIdwLQk92y0ptE1zCROduIwW
3tplyt5zpXUj8PuHo4ViZqWdK+ldg7pKDNRlIlJiRD7nolbheWOjWpPk/v5x7ULl6q/Oz6TZJ7vc
YMoUqG4FyEHOBJulFjYNCVZBM2TvkgE+JJcVlxNsm9ikLVMXxAOPI5qdMRix2pctOkaJ9CiAaqZV
epA71MjKcCdDMTURW0cJpuRSKgJ5xlYBEZwyUxJY1CLRROLAEFmgWzbCQYjg4lBYwDdW9oABHbUW
ej/DBkNNr4Sw0rz/Xtjmb4hXgJhlkVyoRuwJdLHG7rxZrO0Guk/CP1ReGGsmr7pETSUleTP5dy61
ZttU3vew4E6IEQYPlucBzIY/QMM1DiNzLesotvNqoYXXjYJ0Kyced5HJ+eWA/nQ35cenDeOC2+g8
qN9Rm3vG8q0754H4/ISE1+m7fwcjQmZsitpjmsSgXL5eSsCW8ScxFZQL8yVIUh/YA27EZUWPkzB0
YTZhbRTohwTWo4ztDLLEsMpUrd4aDmTHftpHKk2GwMtNiloLhfNCqKFoLYcD8ohyf+eOq2/Dvilz
6Cbd/mL3G8+NaTON2a8RJQdCVutRteZ8N/8LXNBFTVDSBGrGvRIa9+akpBn5FfoBi/xrvjzVZS5t
D0nu1ui8th8SB3cv71w/XY4R2p7pqV6w9mCOH22KHRzvpLrFoa06+o5aVjzYVSm6AGPqFTop8jTW
/NAkfn5X1vlb0yUyVElWEjpG/uFPPBg+JJX6yLwkvUqQ27fMsWPocJzf9UVRVj4GI9XLwfaC+Nun
uA0z1hTZHyQDdeV3CylT7X6+wPP0FVjYt2d2APOHFE/yOY+V15y2609iA9rGe/B002TWHLCiALSe
HKDICg2+N39NkIyRgmd55r+BnF0ztXxaf3zPPTPqM7WoWiME7bWwm7Rn160OIV7mJ9mZ4KhjO9FN
B52guz9DanmFwzBHegk4SLSkBuq1AzszyMQqnuT4MPVOlYs5aErzlRz52OEXkqR+xYdW1KCI4TJ0
gFWHbyZ8eLDwIouudQjvLvdE4IzWre+TTlvuN+KwdIsFx2GvJCEfTl/KdpfJscvPo3ruCGju68iZ
4tB8QfIn+ek/m1vzvHDpDKGG0x54jYI5civlmMO6CZ/BFrAx5d1tHnjLdquyZ6x/DvCmrTmPfBQO
nCZ57M9nP6pzoVFild6Q4DUOkdrmYA6i4/rSqrAF1q71Tv0TsGD9ilaFgcI9ZurFXBKwmkEM4fsA
YoaqR80Cyo6ZmZzoIHCFPw0MwPYLyOa6gJ/OnL5i6FP5G/Y95aadwJgwZJNS46HZA8/PMmE9m9iB
z0bbpskuQSuXf6XPTg4QzF4XSSTmOqo+k16Qm8M5TGtIUk/ynftpaK+NgGJsQhlRhiY9bmNFGC2a
FPUoPqmCBt/WpZaqill8VDjzj3eTUSxhbtw7U9dIjiK+quEaa6pJUgBILDwzLWxT+Q8ymgY1Iur3
6CYXTQMp2FrxTs04D7ksSvxkXeFFLnB+mVy+/+i3u1h7v/Qqm1+mSWxQkn5UoBIa9/K5dDS+k/EY
5S45JID88/d0mcKimp3LIMw8esZOcRq4GGfkHwy4oIz7qWK9BjkDYeHn3paqLSWPbKrklnmS2O/o
V2Kzfxiw4yCj/t/fVpVu9LfrVnxJOacR9tkhFh6pITH4jWeA1zNzT2l7gaXtjP/hUnvH7kiPJAXF
Kj2mWgmAX4+xMoNGjwBYndPlsXIPS8Qs1zIN8mJcPZR4Klk6/4FDEEtEEkINQlXrLOD1b2KnaZfK
KLC0ZbqnSph1JgZcZ+j4LmnAjdkW11HLhgRY9xf9yLD+l7FooBaalcuMRQpxFx0dQAjXfGrElO7S
fOZXP73ALj8W0DVPhuT9pcS5WsXYL8oA1M+/xp4PGA78CUrXmdophAObCN+yiwQsHSwlCXsF0d1Y
BkzqAsPrVUiTzZTlHRsclN0M6syGzZDWZI3QHNiLy3rbCjkrLOV1FKxVOez6iNjSZTxW+pako8YG
TJVe0krM6H0EEF3yzJ8t9vEzbdd9AmbJvEz21bw7Nbeus7VM7drMJ4i8daSwLpxt6TLMGAeLiSKy
/w2MB7KAc0WyEXmYvhT+zknhUY6HHJIWOhRr5eAWqB8V7nlO8SyRf8bW2KhDgcmNILfUtcpdKmjR
ak0cExkESF9SV/G8Tocy7jTsLtwowuwG5XlpRBGmoMNNqo01S7e41xSJMIdY7eNRhnd8AOJ/obwK
Rj9kA5uEIjhTkGHZS4K1giFkx4gRsyBunjUG6WdtHu98CLLsDzqxXG+10ZDzTwj/1cAGG9WxYESf
dh89Zcr9a+VIU5fHeCTCszGGUnYN7hazFEMt/hmzPLXJDqK25/Bp2yRm6SQtc8F5B6M9328Jxd8o
XjrGI/i14VcY5vkNkYPkO0q6y7e1skaNBZb+TugWiqGVMT+eddrNAGJj5g1cP77kLvKaBkoLqIhM
n8htR4MrjsepgBLj7xZJatHF+w+RBeul3N2dwYk+bE8QbT29vho9lQ7JJffpKM3oaiutO30tSDkS
51D/hfuRpM+ghzjQwBlbWYnyweygmAfbb6DFfdwzGotDt8z2xN6acOxW5byfSObU8VhZ+AzV7hLJ
OIXKJTHQV7EZiSasBwYl0v7dqmcSD59rrEc0hHcCGgmvmWSBL/SE0Z6nSgz07TVbhVwgj9g0e5RB
sBQ/u/TJFM4odGFnCRU0V4lavU2M94BDK3aDc3IkLYJrW7x6MNbLuY8EQT9LsOqZsfa0g1SdbIuN
PSkIVs87f3vICtO/0cTOuqYn53Qsva27LOBAe4oIjt8GmtQF9e3IduBw4k+O8phpL5In1HHrKPd+
ER9CJBIjp+j//qT+TdPAbm2CX2kRF8jphhnjTzjNgVzDy8+kirrd3MPksGySDZaV3D7i8DISyBQZ
Q5WcOACxwrVaYiL+qtzbYSU5H177/CMBiIWDuc0EZ1tjdxyAG306VsRleHlkrd3s3QPCHyX6a/OM
/28V3ebV4eSW55MnQyyrZQsA8qQXGUTMj3VDM/0zJsRsbJApcZwjsEnyLPlQVxRmVhF2G7m0l5J9
x2fK7SZ22uGFtwzZBAkMVYWtxprvCMHydShFJ3hotlGnbgX7MiO73WXe5IJ7dlXC96ldbK4UR5Pq
wbt5efZWUA3eC0azNUwpGSrTD5J4aDdqV3s46RQV5z+fwh92RIyOLMJ9l0iNjCqYLxpTzJRr64/q
dNwtIt2hcDGcByUnTLT5oOtPeIraaVKY/MbN9kJ68VaNctGHIaHZ0rTGqijMYwQ4+4eKGnYLTI51
C/UQWs7q4Hi+IVT68I1hWJpNeTQgFQyPmYGHSTn6VgfsCxvYhdLQRYtTtmOUE9i9yCULrLbphU8E
EdWPrJY6FiPGz3FiqoBebZ5BhfdRtt4ZfitU+KHf986QUfBktsrotaAB7wW+sGZJmblPDcq4K+Dw
b3mI0kqmipERkgKpP+W1ptSH7cBaEOYxH2aV32nWP92tTxYld0Erym97/4ZVnL7amFsZDLngbpk6
zQCXkIkAP/bJ11xVFt7zVOY3rI+RJQlMoB42+vX8jDU3ziNU21OXp6KaOgB7Z2dAJrsVJ4XZMNz/
wGlYpcoDyMtkV6lacYUiQ25R2lxdFPN/JGwdXbpwgiFOGUb8BahGuIgdCwMz5xYX5B1yPMkg9ZuY
apuE45Avp6IBtRg8UVB9FdakxvhGQI0l6Q5qanyX/BgRAlx50reQPVNbA6BJbH3WhJ7Sx/LFHnnO
Sd+05LmSqJJLl7a2R+5cT6CJsYuSfbrc1udHWzSJZJuepiSpTRRZG3Px2gh+wBlq3gfQ2jrigGk6
wAJaSW2mSt9WwMPnj/UdoVqxEUILC5OwdRKRkxrY8XbnkYbi5lYXjbVcEDeovYvwPuGKjWEWPGnt
lVrlMr2VXjE0KmnH04uD2xL6Mab97scAQAGcgbkiPFGTcHPL9hA/2U5ikH2pB0Fp60bS1AuEG027
laSWAUuAOZt1QrsZeULB+15EcFli2iagOErRUBZoAg/XtP0gAUDQCjISJMY75rbYD0aqE7PGAs+j
Oe8AdGxv88ReKcp0pZ08EykK2XOZ6p7cfhVAEHi8Kbrl2B/l4kEzslPXBXAoWioMuJf2uwJ+RWOV
SiPr7usQ0GSOYOR19aNelS/Izp3Xx+N0nC1gbdJggezCuAd5QBxQo6PtMGl+C2N0pkfMkQS2UeAZ
T9/3eiTulFbdP1Mv2uiKQ7USG7PmdYkmb+OaoFR5Xsso17SBl4GXgXOn4NcNWyj7JrDLnj82FP5y
hQqPLenwxS7llFiLil3eNwxl9jLAv3jfdpKTWc6bl1ClZf4l2RFF8rPxgPQ0Qe8YJXXQm2CCJDF0
gJaE85HevrUG9I5ROXaw073rXqH7Vwy1uJPwQeu8/NiNPc0it0NHeoEhS/0CHA4GRlZQ2e6CGkE7
KcCvRNpiDvxoBBEkXgYoL9RgxXE412HhIedaRpXiygyryKN9a+29NhgLhpygrX895z3CSYS8nIAF
8UtuA1QS3i8Vl7MYA6iNMKRZPg5JnEfdgry/MfQ/Ny5BnsN6SfPb3jedCNPNGUwf/3msInFF+m+K
PVbeDUN3Ba5xVjOfvwsvm14UTZyR37hMpvdw3W8i2lFMQuFnyAQzlT3tFhVpbIXdzCHt2wTXsibn
vSFeF2tGyEufwbZExfOykKtIIeAfDQuBlp6eZi81SIxuGLRRh6aLKW+eM7wiUCORoizXXtVKi6az
f9C/LhiT0ihnqoWGiS91LOS9a8tgBeiUIka/LqbrAOg+45aXWaeTy7SZAscYVnfykGAVqRpokAf7
rTPaBbwFBlfoe+AEJEa4Mb5/5aJLFjLI0qqZcE8Dkv2gdS3jRUpvUvFf5KC+7H678pg78xH3x9Zu
k+6l35ikYFvU2I6mv2ZKribfS38vvgr5gQFSbEreW912M0NiRwuQ3ciq5uIONWbH45YlWZGmOcF7
O7itpu13CSdsiI3PkIXMyaVZA/OciVkhRtOf9GEpgIvLUnfH+5UGosCcuO5xJy7BKrRtM9d7pdoO
KD++gyKBjPMuge9oa7pruwBFXkUAcz4Z3tXR66/8mXguNNSpnqNEpHuk+FSeA/K4pwM1+NN3qw8E
WcwdpO/n6q0PAN8e3ucEK2FoPHV0anGkdTA9gM3jah87Zp5YGKW8f1cVwEebEbqb79YqX+HQtwyb
CDMb+2IAfpMN0vCHSIWnfpz0vQu/i8+vkGjao0fk7mIrNchmwz2aIrZ7uhFDW3yzu3yi8GQ70p0v
AC9xZs8WorrSQIN7Qn1AWnroAREWsHeiHj55qFp3ICP4Unh8AmQo26+1ywPJCKXVbW1BXwYof7Vu
YfYBWFndMIGI6TukRYYIN7m6T4SJw9TnSqtAaKYFbdI7O1KVsN/+Ge8m+MFVnMcss6XASMl4nA0L
uOD8SP2frx828Pgn/luE07QCMEiw6DjimbAL2dZ9TmsCGyMDljHwk133Lr/IpfmPYsnqetMNt0If
OvgIyNe0b5S3EpRy+G5pJZnjWxdu5I8cOXCXboik/LgPaBFXI9pWn58M7q0ZTl5UFXVIy64DM12i
a+ZoTuZjYrkNRdhWZnQyOr7gsgRFUbSvs/fn/gHmeMpK/SrPC+RuZq04Qj5e25NLzw3qS8Z9vagT
dQ45dVEOdZTxXPIz3BrzgMw3dOOvAPHtwVedzxg/pbuYnZGjioD1u1Oi3n7cBxJb6Avs3XZyW0A8
2RHLGggA6lOB7/67Emm2RjT8H2aZA/Ymyi1pOkXVHTSUZzGcv5bsviNokZWJ2mMN8lTYKWoQTfIg
pf9jkwAnEXdZfWRexffPP0mp8olnHhasS0ji7DKrVFbj2OyRYkBjt9iM73KgnDdZ3nr9tYuTKuQU
cuwvIsSkfabwEICGRrmIQfAOBwVIQFqA3DVDddPQwwLWHjFACt3r3Qvr0TaRcd63zLyeO+tFoMuD
uLsmI07Y0pGlLJTaSBXWmJTuvgq4TX7XusS+I5CKI139kVj+mlCuILct/fBkRkjOGPtmXtXQEG7+
EA7MlSjzt9VYEdmsdSXTXr4y+bEZSKdoOVgVyWE0uEGiuMpijYvjVVMS0JY5TsVwIRUp+Q+si5bX
C+t1EwDzT0ogwiu/9qhWuGp9cQmRXIXy78arVN9WsArR4bfiRe1VHaXT5MVZzBKtsq1+g1/4hR83
kszNV5S9iRr0RUQ1T1hZdTqfohiSUJAZpSaexzhjI7WoUt+IhOiPw4FcYUBXIfR08eQMGakZVP8V
M2NVnKuqNBx1rwX42H7Gdvsu5xE+BjNdXSdzMwMkXbfZ1eHlM/9O34T2twDCWNMt7pRTDACQwOHv
vHretoksEFAZEuKRPrDzUOI5hPmN2EpinDuTrbaSDobqHvoBpFLhA/HmRKXWw+RiZbiozaCVOl8S
yDjERHIG7+R5KAfECTisrp/BeApqYuHG0qvDwSty2BTbGcD+q4k+zfBW0d8YWns2jCGn4mwvsrWI
0yUhoMKW3KUUkhOlVQd/NHebv74LQRwDi4LlqQgO9ghgLLZoRoO7AB1jasJppI0jXVjXeS8SOFJf
Y8fUxOV/SlFQ86YNZcWdFRGyCHzU28xAuXCMZuaDHIx+ZLJt/Ay5+Mnq4/67Utq8FvBhsbH7ucdO
Jlfol5MKADhvHoKImnXUrVcJgWH9Eu/B/q0NrqLvjXlCx047hkIg4sJQDiHzWl4lnTL0PQ56Ipfl
uvNzxm0+0DtS/gOzjEOeONH2VZCYfWE7CqUmEWNKurQJehFHJeNQT7Zf+A5ZKWQeMTP6f0tL1LZj
za/h/LLwePMKiN1MIJBhKHyVfdm9LBhZmefNlOioWAjzPMp6lD04+QejJMdfZmjQzNfD7wP2TmU1
kY+lN0ixcdA68GhwdC23OFeUVgyk2kX0kHx2ou6Eq8l9Tz7qciYYa5nHFK2t5/EeKj+SvKmyEs3z
5ddXLCmfXzaEWZHN26knNJRGfxPnxOwPDI6JZmU6Z73DUGHFvgrIJJuDhitDBazmXqQdpgzxB816
My2sXzxfGIt631nNwZPqC/lu3fh2c3tAwexu/hWbh3ettWciWgQeHlV2iEy6otUVgknDDzlLiQHo
1WTrktod1BrI6gbH3R9Ow5iFwkodOtVfRnwX3Ehr2YBdO6ERM3HKCqm9fCFCh6xYqYH8JxZIAl4X
L/DC90IxdR5tVPSAQG+klXsHnhBEf96ZlDwy76Y9cr0Zekju+ywfViy7KNY9EuAFhJoxL4L563Gw
iltKsToCCO7/OjukMZZ0zemu+gg1nRcar9ySCOmG0jmZ2SJUv5EruAY1gw1OEEJ02Q8+y/W7pZKD
4h5vFVAZScd05F2jyTobzndqyCstbsT4fbqEgvqAQS6J4TfwlGOsQ80ZWVxl2gjCyAIFB+fyL8S0
tQkkRKsaRzlPjiWx13aZOsxj0ScHy9I2CLX8cIceBwJmRwe1zSbiwRDDPmVVqbeIUcayxbpyKe15
RRNrrNAZwzBkSstyvTOCk2XonrWF7cavIo4hTtirmAfklaw23Ov2tbIsSVWhCl2b4fJOrGJdANIR
3nUjuLsOWDLrUEr9XjbXgpTE9uUjIeyM723toHwOPalC9Xs4kcKpuaioauIUQ0SOIHwz1Xd4WQ8U
0yrrKenTxJWdZJGhHi9QRJD6AdGgKh6loZkk6eIO5iOtE2aDJgTcx+AK15548g+dcZ4edwoHLMje
XxGQhDLpEu3e1WfQKUhDZLD1kDUFBIweJPQrV6ZJ+H/yk0Ux5Jf/28AwXF3nGGvhRKYSYAZ63iyY
+HI5GSyD34rdh/A1N45mTfLXJtlarcciL2Mpx3RZHI0GdeN9T/7TRU9yaaHTJXnsh3oqpZsaaond
khZLFWQqYK5LbnlIMeLu3hwLLgchtXsjmNDBCZ2haSRFLOIc6L3WaEwmQvJgya0WxuEW3YN43Hsa
Qip+ONT4G6/yMO8/ayjOge2q3YoQcxnjMQBzwf6rWvCTBG3LUgaMgfghb5SEoyI38S+HoOhRVfR3
nhp4w8NMgangD2rNiwjHwyjA9KxK0uC2HGTtq7JoYmi3/C0RIUh2aHCU8FY7QrSemWpmi1jcqld0
6xMz7CcLkFN5xU1FY0LIEHkBWRGJD3GJeO5Vb+U7iPVkyzhQrB3+I6azfOT5dJ2G93Zyn+7vwx3U
9rHa1xzCIxRfKI3RTMpZBV4t1Cb4aGnhLkSURP8+LX8IvnT0Yf+H/TmcnCl1uHQvkl76QFpIFvPd
rKCmBHEatlfeW/dpKFata8aT4nLzmoo29P97Q7Wb65ANeHqi1VOljMiq25F9A1KNqKtLItd6HS+J
xNpN48Lyw2AFpSKPlKduaWlZt3tzIRRFowWsetqUXrJ/PeC6/GyG+T22MiB0a0VGz5R4F6dbVu6j
VvZCSUOlQtN7YBLWsfGdJdgBgJH2veacBDdbhkFp7X+7CvvKmWFV7foJ9x3t1huDmAG8KChOxqPZ
vmPANtArdII456aIresuTRxiNtTg6fQvSFEB87W0rlMN8NMpKrADOaOgQxQHgtgM1qsqDo4TEqHQ
9zp8JvE5bg1TGhrx9Kges9cKyIQ0svzXS8aDC7Ia/2m1locN7J8tRObZ116CLgpD6tb4oA2UUD3W
PTmO7d87bCaxtprNHJm/37ZtnPCCYYGXJCXUNxFwYrXvUXbFdUhd6KJ2eWpAXzJRbhs44KjiCUU8
dmBsPwj7svSapG30u63syXbouLYq3x9cQGWLa3O+DjrqtozbulEXq9w1MFPzpDrS8bNQb8PILaHt
PB/f/eNupXOyvuUtntMAZ57l+BZm+vIooyPIFTaiTxO8ALASWdflQX6qK6ojoqpfd4d/fQfpuoPn
Y1+6syTr/RE9youiI6DaNfFUo4AxfiBNrcz0YAIbnDFPjHOJfoH4VwBkWywwgBX5WyC60sIUGf+0
8Jgd4qXbHcVHYVZ0DcnJXWbkXZ4K135YaaVJIZQzSq4tJBHeibcpOWntVLHbs8hVO8YjVTTgvmIl
sdm7q70H+qJ/6AfzpD/7VBmono6i0tqouL9o5DTLnijwf1yFrg9H8JzpHXJrP9nBRDILAn7wqK9q
KWZ4x3n2yzVENJaMM6gUivGpJZn3PkydOY7idbl4EbWHQbJhH32QxMTC2vGVlArxEU4XkRi+doWK
6+Hd1KXAz8EH8tb16kjlrGxnroTd/sLa0h5OStlwC4WGXBVckT/WLKrackVAa7TbtlT089r7VbUv
JmUV29fyRJNI22UoHIRN+HtxzTxE5GCE5Ep3lyFqOL63VDq0VxcUy50GR+ndjJCAX1aLQufecAiK
mPSQT7JzSG7Ep4iHKMhdq6sPaeVcHTHtBvVPN+82O8RUL5DC1rdgVS06RgFok0ETnftHjDbcDTdO
Z6s6yvJ+nC1ldf2EZBr9yyruaEW4+HlwCocSRgNZBIbDi2a2qYAosW7tDNSo1kQzPNlVeq8aC/O7
XBoefbYiInhOgzhWVs2ktw2BOk7kfpOFTv9X9f3cY7XtLpogTaKPdJ6+7rVLYvYJrKrBzSrIvDN4
gL3Qekn39a7TzuaJuCgweenOlSPf10ehVndeglNtwO1mQ+/J3lnD+YFtGVULgqKkmMQgS0UhGpp8
0NH2D17yj7jnKhFtxLCJwmxn4nUDrTM6zPGarHvW+qOLEH7NN9iYGoK6BKI2cc8kaW7w95HsOZyB
Ew89wzxxcmi+lygjvz/Qk9GSQplqexVrb4WKXkU5QO6QHbQ+3iPUwT9n4M/kd0jFfMM8WwNXmWr3
hlVVfh/djJKhe0QLsh6HmZwe7k/XSNFgPu4416MJg5A8e6KR7bh8vGCpN6Pp8lfb6zfh0hnvQTev
D2z6Jv/scaNj02/W9i+O6V5UV1bD0DS9TU1SQ8crC2mc0dEZ0zvBzBcc9R0DId/MGLdOiFmZ3/I8
WGFMV9xz6obl6hPqjkHDsAxsHiK7d1ldug1oK8z+WMgHvrtjzUNV5y0M6vnc+49ezjX4SszdI+zZ
1gxicWN7cn/4n1r5Qf5Isc468QqXpvdHqvxedYn1WRM6jvQHkrM6sFx5HK+spb5ZKno/j1S3xwcE
RYe3aAyk4e+r4IACBD12dCLt1Yaz+eynjj4u8dqVWbndu4zp+qaELI0MNcpUJXP0vZJBnIVpDW65
sgomueKp6bKJeIQYM0jbOQ4hlSIPMahRflBcotT0dTnOFIkUJu6A9IJsBuQtN6q/DysKDLDQ+kOq
d78q7y68NNjoyTRu8ekm7FCJAy/P1uo6es3O+kUt93nCcKsTwgNG6RhlgsLd3IZOtQpK4hZw+f7C
ps1itDqfB+74/Gge+XY2wfD3RQCIvQ6pnAhS0WrfOWrAqBY4VPgBLU8Ejrx9znMSUezUziNPYnKG
jY9dw1s/6UtQcL38V2539LTD0KlvrzL4Q7e6R9r0+2k9OkBjAMsbYYME5raSKYt6MTr5JFAIInv/
+e9bkbe8phuKp5UhyFnz2gM85Whsmj9/tK/oXXIyNfyMApRPHpXdMIISN+9AkHUIq1SouaxcX/Z+
pPiumBS/AxsDT3KDap1+F8TcMnHFxQd0BqEBEe86EZFuw3vy+laIoTk5qWjdVX4Ec3ChO1sYBT3S
zUjk//BY19CWW22FGzqYjiMGkJ2xhTp/Lf+FU1+y3kpST0YcMJpcTgCGvnfFhvXW5kwaa1oIIDW7
8j4yTsEzydL7bam8yVNv9GTzqC4t8ZN82/r/w2XwSoRg2XGDto4dw6JBQcGE0qrfb/4783KNHoil
E1SJG1EB2elSQWw+UjpEf/8wpaR7CZGK+9EPV8PsEE/uMZETLtmOuRNXjt9CBvU6aQ09vBQliACF
gkfNMmDo80TAaFIoY5NM6oCAOOR6YcYWrLwekT6nkcXaHCtjJakySTk/9F1KvVtHYQUTcuctnLXm
7TAocLfge4zEGUOW3YqIz70GHTJ/nAxu0tMh9DGQzdXV+yVVPk+X29BD1lu8FQ2ffz18z3HD+4ih
Oc/vCqlvnl0pO03xxZ4+eV2cYGu2WQOI5Q9uWqoUUXLLf+cJmHS8rWJ8HL8pQO5qhmjGfpCfpDvG
UCvnOrmgFDmI2tb6yxThx0cXzKBaibNBnAdzyTdA7prN2L27kpjRsmlgBiAprWIeue9tg7QX0D0v
AcHNA6K6JtOmaAHc5qAPPFYtpo93/rxGO/o/R28NqR0qFF9JOJPmfjV/9DWIzravSG/4psdIjxEC
4FY+hcNaBlgOf90/BQ/tHMOtqYiSl20dr1gflavOTd0DJgsSK6tQ5sAw2k6zYOFRz2xSLjvbS+PA
jRZmBUScVMVyhWAsfjIR8rbfaPwyQCWHS9bJC5+P5Gs1a6Gta0/h1MdypqxukBY3E4+JjntLVeoK
F61mZp7fd1gd7u2hqTcR8NHAnakfoetmVKVe1xZSiVpaUyr6p0MXh5MeGjavCISh9+Y+7xyjo+jF
y6QxqPqsFLdT1gX2Xj6w6ms1FCGY590yHYavfHq9gqDw+N3oHHMs4GswXMJVOXckOFEpEQFZzIUo
r7r63RHuiQu531ydol0xQcRwntX1ubyBDoW3rDWYgz2TgbSodLwkBPgggj/Pg8yiLwMxQPEEfqzJ
rm8P1zmURegTH/pCAY5iyNixqU8bvEqCJnhdiyVfzoZoQM5oQc+BLYqj/CpLNFysyuhAynNGKCjK
oyjd89hlhwWicz492cEMRjBYZ+pUH7V7wMwxvq1SYvhj3OcdQb2CjHhiqakU1YeSwsl8ITjq4dUT
LG2NdmQ1j7N1QQuldQ7pCraqMIBa3/U1qD9s2nuJKlA02Am5AVl1pvN3CMhy4NXcBV9yZIxZ6gAH
CSb7UiN3xWN8tipQIykyitpc6F2U46buPnCKm6RYLcAkDr2b3kToipGq7o6H07dCdMTZDMWPVhbO
1IGdGHLcMlEFUVXkdlVoL8JwS62A2uDT0WJ/ozkJLtbqQ0aLFr7tYxDOhj2Q3X/SsxiPIZHrVb77
qjCce+mqmwunUV9g2jfV3HcjF+EuUXStOuHpcWWdQkaZ2OlNKxuvZbWmO9a1gdbVa91oIRzQew7w
cJTbwCHyjhlP+fGIAgj09jMkSIivZ1s2p1MJyM5H4iIeVtbSwP7TDtZD3bDaFKIQPcv1tk4Fkvpb
b8w2g7eE1rmladY7j7tzX0NF0jJfgcVu3hP0RVIrpuAWIzbazWnH3/y9G1J33/dWLWvSQ2UaVhrv
TNwBLleZNqLQ/m3a6mK/SKT8xBx4I89q5tAxbYths7iiEJUWJDBZh9xKvX/AnMqyTXTA4u/z6m3Y
wnWzy7m3DGkR9jOm8DnUDA2zmvl9zcGf8fwvNrHFqno+VOPak2v1b18WoljI796M7/0hQf74wnKp
BB95wzpy3rH4tNQytOhwgtKmRD3x/ebu2SF0XhD5GUMpEdX2Jtrhk1ahnOiwHVmGZhCUoMaTQ2v+
V29u8R3xYpSLF9xjNHc5zxxaZLPlKjYWBkJIKbHREX1UY+stm0eoqArS5ot6sVPMm3pLiR8Fo0CU
LAw6QhfZwPhTPsBR5c/i9jwyMiMIP3Wlhv1r4Prm1zRG0EhAroH01mxq43SS2OmmT0ND/d5tIFO2
E54imURTgoO6H8JmB8vqybQ82iRh6399bNjQoUNaf5GtIGlxAt8dvPHLrrk+OtvvwI0mCxXNqhNb
8GrhsabU6aP0L8mxB/yABRRifmQdS3Ze/9gOf/aK27TWMATDbZIpFGR6548ZvGr1bXDj0B0JDnkO
nJeZiQ9JgQtN5Inhrz+02cQGb3HN7dPSga4cjM91H1Do5teR3zk+v1bq+OOVs8b5nBQRQUR6EqPZ
+IKw/VrBX/sQ+5T8/uASWnfqclTC8GvYoIUU8ah57RurlxddOtC9BY+THBrdYw8YB6AcfGlm+Aqh
+ipOPrqU8lYsBtMksHRFjM6EzgK5QkFKpJFQ81tfM3oBqD/BlVaOTN7CUS3IBrhBpnrAeHIDzXVs
6m098kMFPCBhcYzUjXtlaV+PZpoj04iuQVflri/YXkX5qVq0horT9n1K66SeKSsQwcGhAmlAVMPD
jyZFKPLHoZG2veQW1h6V6TBwSPHWzAnbj3IqsGYBQiIy1dekqxFF91PjeQKQHmuJQM2437H5LOig
9r6KxX+tzFxQ38My8jVM+G24oUoNu3oX14srIEm17tmxlb1Q2YP9DxHOexmAlQhcsPAen5qNAQYp
PiHUrBFqo8V2qwT7tlwuolexd47FyrWyHKACDc32YfXv0dHqOonuh9E8UqaX2pkEh1Wosy7lwiwZ
53ouowdGDSuDhNvCjHzSsCD7Goz7nVgGAr5WnrLzPiYl1YcvJMEYQcQbg80ZKDo9hy6yjvSRG3Yg
nmMJ41es3Be/AVuMeH4ZEz7Rifs2+R10x/atT1HsLIrlMUu98RJGatAfhhCIr6dbggWypqdAUT97
FS0zIMMfwGApfhUK5a7hE3r+5smXObZWvt+8lMbxO7dwP/2Iy3G1A8yjK63dbk3EZ72SgbSoFcXE
2IsPEeXzckJhSXgYEVJ8yyLose8L5ti1SsvbHHMtVFY0L6iFgp6qbteLuJHrrVxQqglqPFRkfLU/
2ntpENg3o17k/z1RCacOUVs9PZgSYQ3LXkpSfbfdTc8pbEfNfyfGpwAkiPuoHNaLyn6q7e4XVD+n
yEHTNd7UfUsjhBCjYRWTkpipnHhMp2ct0F+A/vwduBHowoeL9qzHK0z6Ev4ItrrdWd8IwtQYefTx
JQeBIKXj+7q0giBaOzJUgYuUiVONjfOtCaB3/UEqvjQbLh9xM4vqg66jvbpjLsD+VtVu7QhbDENe
mZ/SzVC5m7RcubLwTsyNyVqCghmkQ8a6eIetm4Ye3Bpdsm9t8Res/Osom7qYugrfGezJ7zVZthYe
TLYJImfUKNmCXIyJRbR1vHJ2EutyEY58J/73fb12GjZkypzcTRgzWleGzjegMM1pzDlMGqZ3g03C
zbF0VOKaL3wF/Zg+OdKQmTh20hJwrMsEZLU0kCmAMnoZWL2M0vC03B8OhpvD2qMKIh5Ol/pCXc1E
RioEuxUbSmpQbGco0EC33Jl80OOHWKLDGXwHVkc0S1hbDsUJGWrFDkazhjUjESkskesNtC81O4qo
Gflbya/i2Lmzu/o/utIrrxQBgbMDvov+QmnFWYieTssn4TMt3PTfL4qNUWxfzJN6vWxRYBjp1wtd
LuGfQcOdssGZ7he/BoftV5tdHxDWT5vuW3HK7YaO2brAvrBP5nPVP1wIkfyJDHXGG0jW9/JV+Hwp
dY+Be6jN+ZsUuh0u9lXBfkPD3yVx+FjwA698qVLpmOLGM0z+4qDqYwFlDv9UYgUkogCuZdkSdZhu
2oppTAl4MII2VuIXmQUL5mEkyZdeJDw3AfV1eYsKVj576tsN68QItzhhItQ+fcVOxgncKYHA6eWc
J1cLQR22DROXk0NSGMzTcjwwaWXY0hE4K8k+MGIGpcN3p6YjFarBidg7cn6s+0OTqhdHAKjstq1u
47f9FTbGflucT7XdlQb76esU8J2/jNVARAgUmB3ucvpOtReaFtHibwdxu31ZPDH7LTwBHzclT3bG
QIbfovqbC59K7CCCG78TORHT+VV6kIb8KXdB3W00r8+6X1x5S3Mt0YNoKkdfnU7sDLdNVlt2WADF
74BUCXQXpMS1+3dF7AF6hzfV4Yc0L0hd5CA2DnmaXiI+VF0DisIAgtLUa95xXHhfQn17DaWqbKva
NZEw24kP/ZVOcKrRd2x5Di6oumeT5uo7bLxJ8Vggo8mozyV+0cXzkvD4m9vb1PPoHLqtrmmiznnX
DnsD1kuO0qMTKo9du7iiB9rO4ERkmYSw02r7mq8VpYVjcv1LgR927wigKnMpE0aHqe4oL6M5qdoO
FTfFlXgRMiX7Hqy1CzlGqpUv+mMCv6vXS98Cqn7E5+ZWx/DDyj2oM4/DJmx5BISkQY1OSTyFmUQW
ltKBVwbzma9H/4STTfhWNSh2K4drZjvjMuo3P3HbGI/7a6vFlCGpkwP3SLVwXZg7xVqHRrtHemQ0
LaQOZSLa4i+9Q6YAFOKARQ2etKQaL6yBGWL8nOvvTnW+gLGC7ylmyH6NPohHpOM+vl3Z6kSB6gqx
7KO6k8SOKPcgANEyTnZ3AwMhYbE3pKrdQ6vwLVPMtXqOLjcwmw9iUSm0VuEiYvrbWMulgOw+gO2H
NpFzGflX4jHBiY0tT6L2A0Vj5Rs9lR9mw4xIgX9zvr4dylN0nsGSdv9tun1pqchA+2VL3QB865yo
lC6J+SoMJiS/ZYK6gq+2SN/imJ7blQlNbZ3bljInR1UgpkK7LjVAuRsVJdgY3xv9vxMKgpw+906S
CE7hrzaBHzmsUdVe2xVdf8AvyzH+UYHot7LACXZ0v6EL80oJTzye7jAvWKnwe/gUaiep9N0ZY6Ib
vjCibSFHcIP7uKOvuzNXLecjDFz7R7XUMrMl1Ox5tKepk9UmSG8zkYeuEHC8QDhz72IyM0pcuyyF
JMCBT3ytjJG/bBrcZ12Ue1eNPRwJMu+zOCL9FDzVk+8GfDbKhzJtm++za6A98o3blswtn7ESKVch
F+lDpPTDXuufIBpe0FcI9wkiLxRqwtkLWA7wUKRy+G9MTSRRrbub9+97E+hH01tEGahVIraFLFpf
4ElzvrRPJ6XBH19cLWwsPLWTVG+imLOkE4V9inivvF2XYUCVb9nFFTCFwzprwLdGBf1nujG/0rRG
FcoMVuWTsWPHhcsFco+85CqK4Lu09mCPhAiT14Y6GvzyY8iW5IKJT7P2zEapokznTBqu80mF5aPP
G+r0VjeC/aD1pr4GEnCqPmI+gTha2Q2vJXmftKFhSVyBSx/5iFuTatvmY/S6ahbKmZckmlEYoRjg
JvWBjqE752h2urLkuJiMA6o/KlBpV7ClpNimTlzkbQ0Cq3D2A4JZcAGl62lKcmbCyPdT9UgIFr9m
EuJ8NLj9o+BKuVNbmbICn4jDb+AN/FbrTNz5ODDgo+wyrajnP6rFrmyfFyBDXBatR1BEqVSL4N0r
2OuIHTSqpmlDuXav96ohSh4paWExW/iMdGE3SZwQ+zHn4IQRBB+ap3hov4kaN7UxvM6lj7l6oVjI
9pfzjSNG/4nD9hbOJFkY/5IvZf9vSRbHGJhb+yJob1bfBgyMDjnPq8Xm0UZjhLsXuIjxFwsfd6iI
QZph9aTHIhjSjJ1KTNTD3jwdGdsrE7xno3J3MasjGw22hmm+XAOWxaN6WjUXDlEZg4ECcddui0eA
/e5ObPAUk74vyZir2qGesjJhJDWR+mst9apnMIo5QZS99ngDcRaUXowp5MQlxm0s/XNAgrn43voE
UCr6aRDXz7pjNaEwLKDr0R6pSHecdhIIcKT4E+88d8ZZKNE/JAmEhBj2ebY+qflzAIawdh2K9nTl
CaRO3U7TZuDpHsteNMKNOwMKwQhsOcPAmjwFgcwncRHOLplLp6vRy7oIXnUOQC6gh9MO5XgEilCJ
JtnNssgWxY451Y9aXh4tqgFhR5WTsyfzK6idrFvX1q+4+lULS8cZ1g3q+NYPzwqO3WDWro4d1tpZ
gL9WFyy1io9d2OQKVVwUgrP3vptXGhd87rf8vuOhmBZt16WRkJZU+bHl8hmnlY5V4M73U+wZnA+w
5PyCAzrAJFxgitQdTYxxoIEgzFHhHsL2x2kgmpzPwsH+fo2eex29U/iCzTMPpsRPHsuXP8RIgVv3
QHBMDNalFmgYPBSaOskBksFyYYExDI/n2DvUpXJ11JVCo8Aw0p+l2BdvNe4tluycyZZgx+VqNeru
OwXBpIbx7RE5WlkVLGGFYY06JExOaJHBfa79LNvo/IIu0d0AEte7qMH8/T2WmqgtZEonPHNAfeBM
liNoCtmkbAwyf1YTB8cwRCNdXEZI2nVoGKe5Icqf6iD7JoTaB5/WFllJwwqZlxha5Z0ROlSYsGc8
UxQvJLeURjJnCaiRIeEVaNTY6EoZA3Frmc8+J2XSwtHt6f+GEuxMRBBi00EVN9AQKgTGAfGqeqbB
Fvu2uSXLxuKPe69XpFomundJOYr1vR5zdOARAqyL0JbXVYzknPoO98DMxPBxSjxVgM5CsbYYsefx
D2A5+SKBi/pNIh3cJAk8Z4mG7MLUOXOBEuPOKDAucd92SCLPG3TU3YHrepQOlDd2zCRyAqhLWBVv
la5bqC53feOI5jf5aTvaKDrHD8mPSsmNW5BN0eLAJYOuCGbsXtiGwa+mo0KEOKY5EIGPN+40tNvo
fhVk1jtuHrolnI9r0QqwPH7OflJimRd286njz7SO1AV7p4dtV/DnNDC9K+oO8WObZhtpSn0yhntr
GuC9Va/nkeIBBxAXs/2f9pspduhszY3/bTzkIkI9VzbvbK5IGVPKRkegHlbE+88XE6oeC1pW07Is
pmAHQGI5TmazG77Jf2zB67pJwVpC874orLImrydWp8LME+p5Ws8fBRDRRO807EuMnRfKyJMIqr9c
eWb7YbZLimFN1UIAj5+AgC73yeJlCVt8vT5iM2Qk/psOSjAp44RYv07xR3lkRe597rqaZBt4ftNH
UEZbldnKzxplPWGfgd8O9tMg9aiuNevhBE0xw5gU0+4S1x9qkBTfB0Cz7VUETqh41YS6cldWAKqL
1XE7PlA+Bfb+ioeLjwT6CzCkPdPoa7hJXrJ6DwGc+DlxGOPfz/Q3NTbLCio9Ar58nhMnc3L7u+Xs
qS/WhBLDt2gpqkf+1StloQErunyIvALxz7Ha3kmcN/nRCSGbkEU80GejmLKYKCeoWl5uYoK9Lq/a
iSb1fJuQFIoh7u1T/I0ymSifhDb6Mqk5NO0UgMm63aDa8nAimfaORagRrXiTQWTj/EoGhpWRC3Ft
L5v3C6MOQm56MlfycufLwAx8/9jOVdRDmW8QlEKth3+D0qQ6l4BFMOgjs51Xsk6wGqfCO5w/SDaN
5JfhNooi3BuDtLARFKqjPhWzMXZnCXirywl+Oq6d5kNk2SBEe9jufTUjN07a8N01ZyoeyI+B7v+G
ua9hilfN7DirPiuOd65Etpa47hqCILF35n66ejgsq0IO/yATxFx7TntWMMBIbKrrnkh0qdeGNEy9
uG4CpDEmSMowKYdcAIzVwer92zUc9WbTvNKsYVQmfW0e/0BWH6zscrK5OEpgc/k5aDtpsruZGRG3
woCStObBkAmeT/r4jWC1EWfQXIiItAdIlEDwkedzBrDSvyupmdVRu9UV+EKeZ51wPKk1ZvLQT3KD
AKf1o+V2KD7HD87cEANasljfMTAMlsF+JgFiPXMW3STNE2yCsW57LMWxXunCfLUdD7JteBxW0qI+
1XZAq+Z+p4yW2svqOI51dvhtnmpeDepY3xwZkpEJa9FEqTLA2hpH7r45jgiElWtaBwMGuSCItlfQ
uDsIv16j7x0lLZkbsqcEPV+pxjk9So1hV5jvOjV9hninjv7MvdRYbTJQrYhGKov2bHAOXglcr8cZ
7sh5Rb5L3R2PTLXVuxdqteeXkCcyxSjLt1mfp7ZoyYinkKF95F+xaPA+vTgmwVpnSgZwG9PlWgTd
JOc9GeMQmp9zmkoW8w1U40TuuHLUMmBbwtc2iyNHnQtOKx5GXf46j+BG/dXP/rJOJE2ehRr4w27t
6lfJ4NFk46rsyjBcQtyNpF99D/iRHrtpDAxnb+WlLmKIq+vC5p1tCfbIUMvgiJyJW38W5JhkYXKh
Zm3MkBQgc8RLSUbjmsr04CmDPNoxiCgfIys+cAHwIvdTYoZOaDk7yTqSWMnZ1BaBiUYol6Wz7MgT
SNewEyMEj4aYL5UrrC5OobTct+qEbIeGiuy11PAdE1AuqwQaUDeZuUxUCQV7C2F2aSPXkVUhmza+
UohaZPfLqH6mNEs/QlH/fpcrLaHjRjUiUiKe1ASrXfJMeHHVLD58b51Y/IU5ci+JaipoECqGBkML
2BH9nz7MEiBNejNk35ISKek/oRM+PZ2KqXi1dJG/hm99vUIfJeQVnLhLvaeYpDcbUQWEHE98Z0gG
9tAYPw/h63bLyd2UxkueScvc/TCU+N8T/lAfOzEzhjGturXRhTFT2BtCyzxzMjt04TssFjN6njfF
5g8Fe4WGRiL7uTUBSfql9ega+ogpW8cZ3uaA9BGa3sC0A7YKIt8Di2b22vhC+7Kxiav+ynWBxkly
jxn0QjnLvZCI2iSNfhLOFkVItaZvW2zOifw9BTpoQNlj9+sxncoGcV8wZfwtzTsx2YD/O8MUErMl
SO0k+WPsIAWHfh8ozivJ7udqWrUXz4DrS6VkWh2D9wARlgKHiB2cefb3uuX2QBLq/5SxpIiXfrxr
jH4RlYl/EwX8HtvOoBX3OSVjG9w1QAUC0fWWKP81z/umSJM83vhWsksJCLX67zOlGG55lXlx0gzh
HUcuKzwxhSRBP2Ju+rgG4mC5GIll/hB5Foc9abCb3WiGeI6cBYfGCg4SRSloufK3yWa7yrnrHVs+
S5bV2/gpoXrjXtHAiK9pzsIuboB6u6qiMkktmlF521P9VNEU+ZlfcFofj1zPCYg5vtQkPGBVpOer
JPjMkGptELSG+zTw0siWCt4F0tKY+XyiunwkeXSpf0YWsyPRptdXwlDSob8lGrpRvsvCV11TnHZC
JHHCqB9FCLdFm9d/z3LenpeJs8QW1WMMPZ4cYpfiX2gSZKpzRGPHSd0w9Tahmf5qfCMVpibNg4c2
VYWiZQEuwWVuZvmUUH7w58mS+GWIe5674P++9NCSC9h4JcErJTycPJooxLX5HqZWbyJhYsJmq1LM
wYYmN60wKpFzFOYPUnTFnhWTzgcaEvkdbHRfwWQPekRj7QFxFPSVzb/xtZdbMv5oo3GJ7vGjn+Vc
V0LRh16qzyHEELubP9Cmbpix0OP6YATUzGXvcYsuzXSAteDRyYHvpReHHyW1enqM6sJHQau3ZY/r
+wg8ojDIFgReq2gRAvnqqNUL1/u88K4ad4NBlx2L/wXma5wGJjkejQtLQ/fz+v3XdoIw8xTubmFe
OKZL7piIEtUNbSoNMGjP2KTz81qjRwGJ4zsBqwntWQdXfC4BFAC74J4bVorZPQ0JsFNlb9zGaVDV
GuoSoxz8W97t+d004sd0s+jQl+1OS9mjY+WTXFpS1IBgQrYk7uy4oL1RxLmFMikEgJhsqN3ah/Fc
2MKVLzJToyCpbznI4k2h+HnlEHn1t74K6Df8VyfNmPIEylaQlEuNbhkpPFufJ+K6U6zJ+k4Pfk3m
iLnWRLLz/jSYeD2RWjmNsdXcfUO2JvW1OWeBj69iQtgYozGvMlOfx+44APzNyJJUIVXcmrZUni6H
8CB6bAHwPoD3dNh7biKu1J1+3dIYWMaYUgZZ7VdyQ5ddbhGMKejzPRhkv9TPmShCSHeVsGsnqGxG
2S/fBpgYibN5EiWEMFtZmur/SCrv3EsMNTDo+Z32DcOmfDMl0ndMwCR4LwrlC4MN/UXn8CWI7TjV
q0yu1P+LBt0bvQpDg5WN1ZFYhDAdJ7QXP/ucOhvQRx1K9+tbLLe876g8Q0WD6rtXhD+KJsCBh+kW
ucyIC9/E/SZMt15ybZWKVlYAciRWOaaeqEBISVCYxJcjYT1wMJRHqaOqTMPStXfjHDFWJRTNny+4
woopcqSLKx+1bZuAGA6oqkh8PfdzIbvsRIOtp/o32PI8j3ygbnzXnx/ZPJThA2wRqBo7iKdny3wc
m+CPMtjhjJIhc3BeD1i8fY8Tq/GHUGSAr480Niyprq9nen6/BxRpY/k1rYcXKUgwgQQWIZGNhX5g
WpOLxngSe5G54dDqTGXgmnFzb09r+3BEmFRINv7KCEY6SbF2OoC8+iY5nm3F9sgyasipkdKaNpMT
uzYueqzG+DAuwRTboaAC9rUB0tGS+N78fCc95wcIjhNqCSdnSn8ZfkKcOWBU5/0occ+/TZUxUy4r
33Es54z5kSz1OpztugN0B3mhkGLrBX4/gzBAm+Qpt5po9S6mkRxIx90NVCY0hTlz87QU7SjC6wdc
oRDvrbs+FzvHSHOJ1/VdVfy5O/YarC2I48PkvBD5YZ7EWGODcW0b5t6+AL2eNbS/MEo8EcY7EwJa
PML1LfNSpOCBY0zRNadLV31UNb1Poat3EhhlrQ33lvsQSGP2APCK+vkl0xKLAufUiMnlPZB1wnaD
0QSRawbn6JDe9MSTaCboLyfLDpSHZC1tmQEAvA+Wb3dIKvfnegiEcOHrNgVnHvgLH0q6/3MSpSAW
fK0v2+f7GMaC1R63T9tcTO/zXEiUlxfvAUsKewfwcyEaPFN6kj/W7X2DWO1sBLtqUIIWsMaLVCsW
3R8lCu6ZFhTBz0c45sxHy/UBX0NHhpxYwLJ8hbBqxOcWCje24mcsHewNqWzYx7NOdXhMxrQY1vRE
7OdRZamHrmh0/BpCpQ2hrxQ2ctyyjbMqBGALkCUFLCE5mKYFIo4IqFGty6PZ0MwGrwGQLvS/A1Zr
4hOIL/gSD1J5qWSbLHINcbBqm+xA/mHFUHLpiq0xl7c1sBfx4tLw7jdPlqZdUQ7gZvCEcLVlC8Sw
VYoVp5fl0gwZxeXuE6z/B7TEFTEAH2zXHVaPUys4lUFYvNmyb3WnXy4zRFzDaLQMHmTg5f5FDIPt
E2g3idjv6SKlIpyXo/OBq7Ew1TF51sq9VvFxPhjkZ2dB5Fo2f1qNMSx8q0cTUz4g5TRM0e99bHbk
pR8XDbT0kjgkiL4IsPNysrueNyiU4huRTIUXdQiRTLWP62RhdmBl/f1nb26ft6uMZ9lO5dVDz5AA
ZjsJw1LwPMT2+X6MonzOrZLIdy8kNfGXHYeNRdmjEkv1DAvtZGIx0n0EwFqmLyrCO+zW3UfhQ8oJ
PoJN1gzKo6lBeCiJ6xOdGi7hujHWvheNfENlWUEt8pLB9/AfDG0DARmiCzIq2yoqnb1MvbHZHr8r
TqvT2KwVNV5j3TiB8uOcFnw+uBA2Y3118rCksIZwiZioQTPBUe8Tdni4TZk8ND+1CTl2Ajjrs9tR
rKfba5G2zomN5+tdsq0oBT2bC4sxttR/G3PlbvUj/DaAodVhm3HHGCncfMu3OjpjLTl7om2cmMFN
9cavsluTPj3RAoHfHGMJjMnIXPXuFYRk0gWOA3gpqSilMnFjp0TYK2JG7sWBM9M6CSQKkC2hfxb0
XZMQAOmWTB45Pj2bezIH9vB9+m/vhuxcsDBY27oaOq4lAnBjYI7HvkEN/VxSBkuuiGZ50fmamliW
ervtcQeezGxcdyT5PGI+g4EwpCYZhdGLZQDVA8xulNZb28Zbf20Lhy5vjrTyVZ7V2+OQQjNLZdpU
xDs6L+e2JuEsIndQQJSNrJfiZ5xLCQ8vG2NOkv9z5qYt2Ic6eOvCqnWOQjGfAf/wewZazbZrVS5R
bx0tNr5DMh8eaNMvAlxZi0utWvEC0vCxXGGueEc7jqR6D+JuII50DrM3hbx/jfUUfQrnCViAaCxA
AXzWxPommS9JONQMMivEzFb52Sn4AFWzZEvoYKkfdBObiEGPGsRrWooG/PQc+PppQgfAG/bPoeEF
cXv8Jmh8+dMWPc7nFvx7pJgjt+M1orf7vUZbTpveka+q9WVQHk0rE6s23PoKrtBw9MrVaDePyjS6
TQ0d29bV8FX21ADmimsMple98RGjPrumHhQf2ldhMrfPPodwWkkbBFl8LlXw9rFC+D0z8JpIdSSc
Ptf+bi85ROMIt2JqRzc0wmRwNBHCGWzCHpAXwPOzs3xxlNf4RL3yfGbzgOfPkRMoMY7jt18n7xiB
uqzxkSueFM+CYgFz9SyaNpWLv3CvJjOlbW4LGoRpCrQ6M7SDn8rxG6fajoinOT5KdfWGpxKNJVjH
w/bccZHQDDFIx6+OPe8YLqjHHqzuZmP9D749JmQOVYa221zPJCN4ygw5uVaU0J9kRERiwOxIGaCZ
D4kItAokRzsbX1rqE3AuH2SJDkLDekA6DWPgdqmEQSPe/DGfuPIve9Mr0xFsm6luwqbteKfTFZSV
5A/4kUXeXhc22/mf0jF8ZtKrKf8HqDQPEtIWBpfMoINWs4UR9XXXnMn+7XnYczklwg0xPxSCI2/S
ktyY9ugyX7weAKK7VjnJ8ag45tChM44cypVEX+fm+q/7iPhkhLju7Cwxiw81S8usgvHQW2QIQ6QA
pwtXy53janbxU+QxHFdw00VcagPr3y0c5fydivuMhK7xNXRx92gbX9cK77xgpHnLzgYm4GGdA3jj
DwWqcm4W3iJiHbJ6hD0icISn5YtRjv/k8pHxysPDC2pH5wUrPY096nJg1VlyBHjpyUTBbViY9MAf
r9esgWY0AhBSvBFwvHGFDfvYnbnnU1XlLG27ddAc4G0/awwSxDWafCbEwpRmbx2ZwRP4VntK/3KZ
HY3tmODd5s4JUpnQ3kCC0LVfoX8WNZRArsPpWVCL00dIX028relav7ou8vJ/nk828xUhqngJCRN2
HdLygQzu2vvugYmifWti+EO+YlDwEKiYISeunu2h/G9rg9Qkbct7K/7SbeBatUEm/xxSjX6hUM6R
UE8J5zVMxOf81xjv6poY3eOKkuog1G9EthTPPKgHIAOUha49txiZPRF7D3E+BzwjTZQTuPlIKo7t
rmB+MEY7T4kC5tIXGQ4BwNdTi6XlFqWHGyl1G3KDRHPPLHFVmnRKVwJo1wpoEZedjk44aWE9/Ur2
/Cex3fbdLjZqGLuX6VrCPw5zhr1CEAJRylWZ2ltbyWzcOOeM54Tws5L70SQH0icMMThqmho2VpVG
e0Oky118psgvwmJ/0r8bTqDgC2iRdJt25xkCMfAAZyIU/65Pl1BYjSwQvd14i77L/nuV4ZEEEdot
LwxyldIoW0C8P6rLEYNei1WRqyPkcuIWlgHMoBL1aCo5UGw9ecZtxMxQO/j1PhNYeJRQxuXaFKoJ
N1JHrFjAewHfG5WTcroFZt+dxfFI6ejEY4eoe33Qnqbl3VnUbHRvJxFdRna9yvZvj0UkH+Hz1k04
mzcZC8YvDRDSeg7JPmtR0LuCsv6Z5Sm8pxPsjlc3NeCc6TTe96IRaQUV9WMHURd//M2flKIYEiU/
XljrZp8ekWZe+JtYqAi6iVqP4YMmA5sSBO9sP46vVv/D2slyVhCHV4ovE4V3qXABsCXt/incoMi0
wQV34i/9aWVI479c9oxIvGVtXqDg46vNHoOZib0dF8UY3JZfzy0NKqGoOD7z/09koMshNXNEuSc+
xdIb6Wf7ljn3aw0P4ikScRw2UAELEttGJSyAjYLxfi4eFCtPyIqyZQRXoIAmqd173iEcE7ou0nML
j5JPiVXHSWDAV89bHUbnshj9QiQLdwMnEqe2cTiPFERFnl7nrLvUQ1iZLij0V9EkerSc+CzILRQH
NcJ5XUbnvbQvBeuImgJNIWKLurUurjN/a7YTcp5hpy6JMpj98fCuy/Jr5oIylOy/YosRsEaz2TkC
KKI0GdC2ONS48Oa+YDyWEB48Qo1yUi1U9jzmcEQ2o+ywkI49kQumhvvHTUmOPtmBQntUtFwL+fME
Xb0s/xRzupc0tGiQTvxU4QFT/bIB6iy2V1zCJRR7vKKSrEqlR3bMLktkVb5fUQHNOgRR0GTU4xJL
hfTm3+/U4y2ejIFmJ93NMrIUc2/lD3SoadO/1pKtFJlNunJdv0zd/51UZkFBGi33RPfU/dRcTmwu
WlkbEt0MLR4C/7Az+NNy3Cm4aLqMewXKn6+43HbK3oGpcxBROeB2Pg6c9TZGbz8XsA8cquHr6CMH
vsZ1i6wz9X0yXUPji+fnC5ICHky2/OihThtodFiby7zQ0v/QTkVo5MCGVe3kQXjfHNLyA8rYqe/W
HQNQiZR1YwQ9HTvawOHBZSzqaCDRsM9DAf9/FfHOlLUOnGTNMFx4o/q/7XFWJnBOo0MYrVxbgjuE
2Qmg9CNfhvkJmksJNFBp6jCLm6pDPnIEBTwy8d9gbkbWkSBu+BLOnNL7h5jARWRQpSyB+AhJT+fY
HYqW3IlIU2WlN0frxsSbxn+hIpRidyVOWshDb1ng9V1X1h3NNOskFe/iGwabqAsVGsl79Cm37kzB
EpLxA9aVZjFzDTTX8FcapOu6lUVM7CJvrdy2bm9UgTvQjjQOnpyXZtNRsX/BACsSXWn8XyNYWB0e
5co7mHpx6VK3a/t22U+u8ljEMAZOd7FiI4jz1LfE/MXSxHTlP7ry+wInWMaV5IqWVKPQEo1kt8yU
lMC6gue/CVFyozpDxtvyQkOQHZVz3RNdNCDcF4gKqsM+cM4WI5W+e0kxHlt4jBA+PIDOufU8iseZ
2OLToR+QCNiVo6aPMTdYa9icXpxLISuf9jc4ReTQYT1mCIuM4siQJlPjfYBXbvU4/IVNqCZLlRBj
0h2BVBCj95FQIidyoyj7h0Upp/yAP1/WAhKI7py3PBsGCGtLe7FIMDzPDgFHj/bKH0HXrOYBfBNH
Y9EnPuyG1S1UHeE7MYNjRmM3hX7Rh+JR97OwCPoDVEIkWp0ILq8iQaPEd6U8dKZIW4Ezc8VX6pOM
Aa3B5l/kDwuFCsF1BBbHkfk+Ux9IDhSysOKx4C6gcwt6sfn98ceD90NMYahIy0T8AVYd8ESZqANf
ZFZ+82cImz1drcA5Ry3di8xHKgdzmx35pcXaiJNGTUgaLGA8HS3JXk+VyC5T2PUbQMkR84nT7AeQ
LoJbUkTY+E+ahKD9SsAoWWjzRSufJdubJGE0ehkcYtXS3WyCGm121J1/2cjRriOekkCwtH0HC4L7
y2d1ZJ7FbHdE535YmGN5FiGFxdVq3s6NgaBAJ6dPt6VpCH6QtLOsIijttakCsogn6BdvN6mWqVCP
W31t3hMwwHqJbmXsKVxM+oalPvvY26Ri0mxAwPJaViYyUwJMaJjuYiftv0Prtvmq358koUxa+xax
+VPvb5LNUj6Pkep1OJGOVe39sYK6+JRsx3egPRYO1i/ASc1Od1UZxZLXWnNx3hTZjXGBzEPl9mg/
Z671FHd1X/UKxrR7vQEOoteKq4ygni4Kwm86tIcZVB3F0kJ+E0W5LtxRnmPR/udSkwzXu7vqpWDN
9MrhkyNOnDZU69MYhjT9/rqFTcyxXJy5dUc1fvG99oFRvtNjQpQ4yOaIo8gqDfZwY4vf9yF06uEk
DfDUH2QrKzEg2jBASEZ1SCMXhCS2jJ+8WtW8d/8W+fslS06Du0Sr5OcGtg8lu4ZB8WuQ/56FMXnY
4LcP3spoyTrzd73HKHnY25/22BKkhT1X+WAx8xKiSrwD1K6/Hx1TOvvQGWnxQYI16xNYmMMzID+3
d8z5szhfxuFhGcUV/r9M9LI6aNEgOzV8WzEjlnZYJj9qmWdqbiPGxOlw0shEd6GFzapX1xEdEq5W
0XjJ+6L6BI5B0FvQoeeOyHq/G7VtlwCJI11WmUnhW9Qo5tCHYJs2F4bk2vQTBCre/bg84nRtVnxE
qDsKtosSFvDCI4JGagqs9pxlOdIZ44/Gn0twn11X7QkIrBTldRev4SBrN00TNIP8wdAh+Om93hW+
QUlFiJJPjDoLuhhEb5SCBuDaEQosl9vMmJRx6OqLrw0DoECbhI9XGk06Ln2UyPhrkBmi16Fjw5/g
o2mU+RUgNiJZEtBhAY6bligSlB+YQvqQe4pQveAM0dcMZnutW4jxxCOltdXZXnL4UUhOHkGcwowQ
GSIBISZxKGKlJWZxd9QWm7U6NKfujO4yci2/KPqttMFTXNhW0UHxgfrVKF7/2MYKUTHshqIiC/Fd
7KaOelSkjuioQBU0d5ct+NklNHfO4sAuXn/TfJgex+bDwc6cRol13jTXfFW46pyIZ1leeVE46zs2
7HTGRtBxUhJiKD5tXck8zP7knksnw/3feJYcbSbfJg1iyNLoVcSrjARwg7aPbvirRJxZ+dyrvlFc
DmOYRF6faGI9oBG57DzmYMD2W+9tFFItsgJShqzjMg6aC4BEjwjOaeICL5paZZz1gKlihu7b8fU6
NCv4gCpj0XP4hsSwjWO3No0pc5gAHJIfXvhviGRNqqQfA9ITIoDjhfAelgdevLgTC/g+vmcK1iQF
SMjsHZjTjnoUhqkgmxnIm+thRSlyQnPQPKjEuBd+ASPxFKfGJ0N/Uz0KVkY/AUObZAhEEfY+jtg+
tbInfdQhCHIdjMT72uzv6gxgdXlCbuvJSQaH/MTRon48RHMyanG3m0lraLF7uxg3z0NMW3wXUFeg
DTx5nN0uvoB4Si8/qmuC+zbkJn3eJg+RqdQBkrs5NzhuyVFDJ9CIfDCfvrkduOx/86PaiHroAcuo
UmoGCTqKcFOwaudXpejBYQzJJ5MehmYuglQG1hMHaTHrv8HrFWTOBSa4ax4Lty5yuJ7ahJ/6tyyN
6A/qj+BV1Nv1dq+/BX+llY++k//oyrdV/t/u9KYHr/Jg4LkcWYMmcAOhNIjrvjoRWaGohLsb7y/a
q4JrJX4ceXPhVPB3SNm60w8RvV7NTBsYeUqGKRfhncYkSYWuP6oC8zWnernkQxxhLobE4qdK9EuZ
0/nt6ulxkMUlU9Rt9gt+X5Fu/ackzaOUU4MgSroQatdyJDlLq/JLhKgo0Ftj6R0EYHDlHCT8ee9d
HAmVCqZLBTrBhAmqTTr4mPkeV9ZOHKgJoghtSvbyN5MVUL23DWNFxDVH4BLMGndsZE6SZpbE7pkU
NEaOHwO3xU5kmu/2rbcB1KjTP9CwkdYNMb54i7uXtylsRyoztFlW9PAFfBhmoosalJ383Pr8Huj2
uywwP6Xe9E5HKOjVJ0Dgus/BE+3G7jg5VH9FXZlWYvO8ujZXB35QsWeB3ijb70SEEJZyPFBbpT84
NrYoD+jV6jVL3wmtGxXeWwAR5QThrUf6Gu8+zgEUPa7Zpk17ocixC7uG+zZP9TWYNBZJtHfjpGhe
L8CqKN9stbe+gVvvmSY+M7RbYY/UhGS3R4OXbKMOC57Q3znGolIWNaMzRxOwi1TdzBvjyZ3J66k/
stkuNXKj+BfOFet2CUv8Lp1ehSAPgUrZUrEHdq85PeMDk0tOYnuR/Oda2S1D7nYXT+64AT9AQAbu
AB9FsztNhwze24bLPPHQfnJocL05BvgdEYhcNurdlYAPig+KQkW4X9raU4S8g+VBkBsgDkqIO4Cw
T6ePzQqWEGnkFAaZYv2VtXLcfX3ZaGcZB/8jmnywzuOD7KSvj0bFY9vIJDG8c5rlga4XNaQi3CxX
jd9Z4uwBofcP21Vq+ibS7cyKRFEtjyXs8xjYyk0fnzGpS9x/4ZW5mAzbGsfKyvajWz8w0tB5Lqy/
FYTP6DS6LYT9mj6bzy/n53jPhL+F/MBBERLq1uinmgdsteIjcZWZ6CxmFX91AMwWxwRsROHntWME
3Oo+D4bIaendaerwtxMkJ4ckaCl7FCQlZ5HfPy1IrKPYnaeNK1WM8c35grZfH6uMjlXHa9cpXN2x
JbiPEC0ew+atiTrc2Sy+Vy8isLZU0TBF3iF6oUuDW631EhjtJDNGfGJqftXToYOVHq+xAJsrB4Hu
RcI8cb8yUIpyVknXuOS1Z4Vr6GqaJ+a4j2Tu2VRhS+PONNF9z78z5Dwt4+4S+iexyGlqQC1SxeXu
pbmaqjkVhwdLSgaGoMsDfWvyEvzbpr1QG9bIgBUJ/FCFqPgC/jioQbg1f8NC9bKGS/a3f83X/eTK
bx2n29W3gT9pyxNGsRppw+CJ4uiNcJo/+ifhzYqgwCajyGAHRRkLX9zsmIYITuAS1JHnUSG5BM8U
yfJ6rJRdCR51QAvOAqQZ5tv60WLxIhn37CAlAyIqnfAkxpHHdohALjovD+5zYIqI2prqSOyYJnqn
TXc7pAW++GZG+JbIEDP0uFRmYNsB2jm4y2m88LpyBH4jQdAROSdcO+lFiBwZ4LeoguDfJI+m0OQ8
zfpKWp3w7vG8xbTGzMtsQdFX53l2gTFG7RKtjm+Z25OE7eU71/ECzmXpcybh3ykO/03HEWagfNMO
1RuTXjTde1UNF3GmqG2emnodbJlbYzG5zKi84ginLgK5XvPcutogJ2ksA4Z0FAzM7Jb71HUAue8S
M3q6Lu0EKVTgnlRhXkP0gDVZGB3u5xsDQSXHn4nIKh1R4KXzv1oHBYOVtUPhqHpmNZmzZGux87wp
GBcfY3KRbtIun1i5/lnooYvoViBpku6clJ3iiTkmaTc/cb/vL5i36TMdWmcTr0g2NRRgaPnVPoPK
o+LdULDa8JQqJtXVGG9DPGBqC2pf5Nvkq6hBOXmH13ssVUUYguiTAwe7OHp9ZQEyBrVlH1bE/IVJ
Y98UD5UTP/3i+wVWWM2sQ9YmSWtTy9FRtpijuhksI+UQQEuS2/s33solSg2mJxNtI5IA/4lGlb0H
PPzzFihI5HdMgu544G7wDcsIJZhQU6FpDaV3nhhCbk/7Yf8tqirCDd+CxTN4bIFpRwLdX0xk13YD
ZWxkuWwfWXqKiwLbcy+Iso+JS2letWSOaTiZYISZUFi9gOpdtj7NUmNeYB2qXf6130jf9ybwRBsc
e5ib2bFA8zRnI1gzllQEhXbqcTW0jj317v8TIDAGb5TJaxA7lZNYIMu/RxXADb2rNjnsF3IJYEed
c7cQAkPAF17pKiUEHekSu0iXnGZEJju31573p3FvrjQYGgX2Tcsj01/e1ul0QAI23RAUMHCNSsja
z3QV3L4x0gxlhzV2PA8A8xGRuIs7nSZeCk2nE/Zr9gBi1K89UBP4XsyuZPAOL7kTqCVGiE6VDPT5
tNjhENDuWLS2Poco1AsxaNz8ly9mI9fqPfdLq/O1R5pHq0hsOzSbItquc4g2IgRWrcUu/A5sV6QI
8zbrHe28bIevVFKoAqMYEN7YJkZehWfHolfrTyyHmydR1EUvw078emvv2Ht4G5fvUtRBQ2ylRhNS
yLDN7bVxXneTE23NGBtZT5yoxi0u+/pB2D9uOTKBj/2arBVY2eOhhXGb48ZYZZ9PddKW4hkx0WUI
uPUiVY9f7WIfKig217EKJwIMOcGuLEEkK7CCzIm6dxZvsURNhRrOaoYsjqa7U/SJzHtTgzT5OCrB
4cNbL/4Rv07u1SF+BceS+hksepexauzgnW0GXSmFr4QrLw0mFdQ+O+o3lJ/Z4hbAlw+LAbrCOs2V
AsWZYjUHeFiOSs2xci2LEBMxnkmhsi+ALWKAlmLO/HzahCUvvc/rKd7X+0yyash/IeWYY89Cirsy
vezsY1PGi8KG9SoyIaI6ItKT9YCtkOk3m0gQwjCmuyi+krFn82laFk50WDQWsLOE8rDGaJgpZqEL
p0wruHfKvuNiapBxu4xhFTHGNQrQVNgJjE+tJJmZD3JtZlSAGDr6cydfFgIRM01OR9MUbsl9oEIZ
+UxtdzN9saC4f2Tan1yKfJOE0TJ0F1huiyAZ0MoGpCFPd6FYBKg7JHpAubi1NKOaLd4BS4A12gcp
yUl4k5KziSX8DFFdm5fTuLNRWVhG5FoT72wS747PUw2S92aL0eKaeGE8cCOMUJrWzdq1Eg9J5yzC
ALh9t7DbaIcxzM+inwCSvU/pVIYaiIOtFrC09pUYEcK4J3asAnlN7qyrZP18x5qGkVdw39amUIwl
x5pXZupSekk26oy9eSxsdxsxbixqC3Pyrm3lu9LejJyKn2WBd3W4s3tP3JcDlNIa3tQahN3esOq5
lQ/0lmmcQpDFIINWDaz1vTfet2E0R2cNjDRlHwFIQEw3t84oJQ4RPHjeDAWj7ud/ypQiOOIb56PR
IczVKGOKOmoc+6RrXuInd/xkuJCti17AEMrUAL21S3d4yA2z3oeCUf2bZKBzO9b/VJnvaeFFrbyH
AVWHNCOCE1dMTIBynYtKqDwUD63F7OSDihW806tbE14wIrGTUR7QMzDkS2jXapAQ52TsOdCV/QFJ
5JsdWSONLCIvkm4qadCWERYeODuluCN03zzdJpsBlDGo3KcbEJfL8/e37FeT46HgrN6Cyq+x5FO3
H+1HC8TDf66lbCvDscY/R8+nwQeRWO0wJIYbpsEjcKUICmgnviW2cEjTBBSfhAFL/P9efxU02gmx
RIuVV3i37ru84uuiVxU89GQ5h2eFZFLZxOTskto/hmMEYH5EgbM48G0ccF+pgtLljxtjWCl9iS3l
T4GzCpGHdhwmeTnh+s35jWhzldT9PYO3sW2eIHtV6fsr9NrW+tjsi1RkWIeb5dAfV3w6aEtZTuCq
DZtoI4t9aSkYWr6oP0q9F8rixNjJDSuC5CxtpQQCH1iv3aE+IwQ64VpmIUVUsLv3xnD370dfb/TI
Rc6NRD1nEkJnUDxNvqRZ4xTMGM+Yf0jZ+4eEu7T++sdRX5i2T8xj2sLaQz8Ww0KA/kl/Xs7eJx4Q
q8NNrab+5AUiFKxBluuBAPpO2GcRMa1r6g5f/QKpQqQWeEDg/KCsxKNv4jO4q2lUQ6DxaCvM/fd9
6cDKDLthAphnx2zyCWy48r3qJI8km9lgxiYILkAImNCpGPPTPDOHcWCJXHLd+8w1Ce6wHA0YDXfJ
7QomSst2pG1Kd+qh+yfidKBZsEwYxw6cq2TxpEww3g8s14xWpGsmnBzcIN/A+gfOuq9jGq01Js2a
R8EJVtmbDlF2tcPUvzCR00c+ywRd7KpdhqlAMShj0SUfLdU6wsNkXwztZW5KKpWQvm7efKsyqfAU
U48brEwo42R8wMR6fIHjz2OLP3WBiKruldJzSjEv3lPPZ2BNsxey5J1Z3cUwDXaNiFcw+/CO5b9V
SbK1HLHcWirqUWbGpSXOKAKZaKmFdEbRx54M3oXjvRpFvwsdxx5FkONC8hbjwBp9AE9XUk56LRhN
jxqZ+rL9wESQFzqcPFki5x+mpemPI4TfdvO1J/h2mh3eoqJ4LVzaY2h5LxS8q9hNdjetDgdsrs63
Oo1mEt5AR6nEF871t2kQL+IaMA3HuBdqoaRlSrR3oYhoaloICuPJE4mBTBjWFKF/XeTkg0l4nyh+
CYStwHGFhGrZ3CMUsKS+v65+jBDh6Y0fBYYcLSuTA3BrN+IO4jsyXEit18JDXdUCsjO5dPrSE6OG
BLqETkGkqWqvZODlszAD2WOO1h0T6baQ8tELbIVUJapx/EQHi/iwy1ZLZ+TS3AOtAHENhim8a5as
2Dkakl7gOmXfHL4DJxyxVOVHJt3x2EVHC/svmlQ91Vs+GQUqovMzuWj7GPcHlfrge1f3hCttDE4I
kpCxRhcrbdebm9DEcid59A/5I/HXPMnz5Y9ZolQHnX7bpeoxIObyN0C6+6/k1WgnpJxDknAT/ZKO
ld9C0ktFAiySc4plKlLvcCKfiUNmI14t1EOFeiewE+afpqHyddgq17BazLrUQlBXJy4x51MgtDQO
qUhEkhvDFCFWp4/nO8bKuSqQABu3ol+KXNsAXMEzrlO+W25kL1XRie/DYr7klPwmYnJyq5JpMK5c
bDp7KC8pZS9ba3EbVJKUQPGoipafkuMR/xuJQV/sFrsHTvU1i+F9/MCZQ58rm696AIc9qXbvT59N
AwO1xhiKlW3uTlBCo6M6vqqL9xH7VcLqlNURjh+XMO0vPDLpM/fIZOZVcmXtSSNBxSjCHWmElMP3
dULswF7ZIBTu6w+/VUT4vDsqZrYeSzP70nh40o+FnkXQBFmjcraNuqU/qhtNVPsMAM9g7aAAyT1X
87qxhyhdqksiZuagYidE5y7yU0qe4y2DYaiMaTDI8fq+jOw6HZdrEBMmYO/lyFxHk0b9vphDk69d
7Eo7p7wW4+j/eu1DNOVklnLIx40vNFK4+Qb9cjF/I3udrg4vNJPzefML5irax0LJSPTY4Lmnc1j/
UL2MI/K52ghbtDDExYuUQUwcFN6hCPV+Sp5CenjqGo6qmAwCmLLMIdks0mg96budCxQzsKkEWpgv
Rt8wSQgrv+6mOXX5WJPIUS8W9jTzHfrVJ2x7xtRQhKtqeH1q7nzUHpiR3dM6sc/G7RP0iQiXlmMl
Xq7/Zzr5EG+tqeok3E40cgzIT0HitCpad79DdjtvjKrUhT5JoeMDQEh/E9xP6uZdu7zw/he6IGvJ
UvqZLS8KtF2bMthUWbi/S4GEEQvyjCD2JKOnLMlxstKgNZ6wLJ56EpmR7HRH/vZ+zZDuycJk6+8i
ifwlidQESxhKIUChF/rSedRB0VGGXjd+yHp458T48+6yu9Dz1UIVRvea9hZF2Sk7HMasUNxWgsCS
zAyLuNBHnSrfEeiUTSb4r+oezWguZqT/f1AmBRAO5wJ1x7CO37ipa9tzr8uL0h/oSvKGgF72OMTb
kGx7qi51xBuke52Nt0yy0TxnLNrA6Vj5faPLk5/NnZI8HK4bZFwadnxxlacmwaQIuTEu7r/gjrxP
KR4WjrDxxYL8E69Ywbk/12/4rrY+eEazAlm1J1hV3odz8KUO3iLrlSRRaVMYYvA4BsRsmcGVoDtY
0o2+uERRv4Av60PZn0obZKdp1xbWblsIJVEcgbBDBnKwwh53M0rV0977X3tBDiIh4tfTdnQrjTmH
tFY4M2h5MuvqD/zLbhIo0EqA0eOQFH9gG5XvPZtHSrzaPN8CTEbihjXeCMmkN9YfEkgeMZX/qFkU
GrkTFFvvW10fSErmAQyWyLyZlQtevcAX3y0EASrNAiKGPh0ZU+rPakLn0G1hxf83einyqwXLPWin
tF8C0plFvsNhChVvD3uVRFvkfQ/Um1TlKMU4q6mnn+ACrZy08NclizaaX7QeX7Hf8ZZVWejMhye+
w1JAfUK7x2CC04K+zr39LpVSb0tBgkDjBvnuoQLYffEeggAIlUdaCZR0e6yn7WwfNxRXgNH8U5jL
wMD7wXE6Fovs55AKrJNk7NA0zGZH8uX6eYU7eIsJP/k8Vg9oDtKA/aNtmzjKQ13NUOC1urx3z6F0
tm2wpg3vBrLhqI8FRlPjyiakIvP407YGrFA9eH8G0q1u7UiGAXhFqWF0Uf3ACUE8VHY3lsBbV3z4
9+BZhh632spH8YRjexU62O4IFMhsVc93fWuOsOnAuBYXVahfnng0MielxFQWFw3gzAjgDVmKaaIX
goLVo/Nwxs3X2Mb56BiY4vBdAz2dZXO4VkQWbBw53n2tmWmbZ9TGmm8NmQH0jBk1yAtiotkn12Cy
IAURmQFLFz/wyVBcaH1vD3lnGHVULkaC6Bfxt+sDI1pYcLGub3eLRMuVKc8mpKbY1B9vETBx4oo1
3U0GnqLT9LGKTyr0LfhtlkuVnzJSEaIzS/9Rhu28fpCC5uGZMcLebv+jBVvzP+dR2unCjS/hA6JC
VilRU0pDSvip2rW5nG+wbm/DH0U9QWoV5dzaMi4H6/e0G9sODK4o31WAR3wXU9QFDE5hEN4/Zwmh
1Frux3e/vPUSSQVOG3z64myYsl0KAtk6K4vZSXAkdHCtCJMS8lQVDINTPe7IiJH+73tRIaWI19xW
Go5zDFHC9MPHz3OSYmSYerZRYMwdB9QizfxCsHQrc5Mi/u18lGgQRbLNKHKTSXBYoxjoiCPrxnBP
QlyibzvGwgqsE0majXV3yGIEFca0bRshCdunMcqhkGs8ZRa99iY3KSq06C29xW7T6YgmpB8TuyGn
jIRdJTTh0hG1JY+ZNMf7jZaVvIXdH6GX8Fcdnc99UCQeEBM02LaID2xZmooog8MhbbfMOZH3yJtP
2xmjcgyyfppnru6YS3rqNH2mwhK+Un445qo88CCT15diQ65vUsOmUF0ZE4gNM8yLxibKdm9saER7
mMnqCYN7TbIIvs80bxNYt2YdTdNCmt9JhsU7Q0+18cMmZ/jmThJ2fPEtnEjMgwwb6CEuvFGsyCa4
qthl7KeplFBIJdUa43hKLwRQbnHMgJ4ie7QMZ+04WJXjgkJmdBgrxcBVTr6wRnCrgch4ZyMTol+O
ydr5r/xkPHuo/UdxWkVzFHUX9ZPQTqWIqi3prRuvSIfhK3AziygKkNLC8TRjuYTGd6ISWIZ9Nb5n
yAFcBTO2oDbgnq/wQzvUYoLeUN1l/bbNdRRi/ZPnjhWT8iL0sOjxPxBbtDthvSphJUq2kZvT+S5g
KuR6fGoN3XcUKVvs17Q+JE9zP7oygfDSMcgQDfzQcVQLz7Tbh2Nc0W88Ugot+fuN2WHwi65a/tfn
v8HsECDVBbpzu77wnepptkwoRZ/7uu5sCU0jSD9Y2SNoCN2LbcS072VUSq+M88cleinfK+BQyr2v
E1HuezmMmzdEEq5prNuTT91mF4Ckn6YyA/DbjaObpcwrXEsrWZyeLdkcaWHtS92g7706liIbCMZQ
JylRnv3ZEMFZaEDpJ5+fkJ40cIqbcTmfhvQW8hEqpKGeujXNVDxb6yXm6XN8uR1dSGC1vWKrXD3b
FHvdWe6wwJG9iFqgZcXI0RMA3NypXV1u+KlwvqOf5l5ey9rPm7BYUAuZhoDF5nZ494Txaa+d+E1Z
OtDFrqQ3zNvjYnUF14RU38vTKSpfWCnnSfk+972mN3VbiNK117fhQrTPwOi8M8ggos/PKzxCiqWx
WQGK2jeyC2NBvmUa/WwRgYMylf/Mg0Y1yjdk+uT/gPkxprGPgr3GANP3OTEMmk8blNA9yCpX153r
u2DtaNGZsLq49kqIh8CejVvgCRK4y1UFismWz1nmto6DUboQjD5HPVW8ZA0pzt415qaBVwVxTltw
R7soPxpVP8ePiZwjN/vYNp5LeZXwfGXu2h+jfebkxD/sBA+0JLVI7NS+tj/7iEfXye6MF60EKeyY
Pg0o+MJJkcokTsSbP6o8CtQqAvTZF9BP62b/KJLGeHX2IdhOrny50nEbNr2gO7/Ta4hnpS3QoDQb
WiD6IB//wobqReBUgaLXxiU4SA/8rM3yQyS/5nFNjqGCcViNamLAgFiQseMOkRSfHPzWaxkqJlnX
oxhmsIKN+TkorUnDwQtL7kfQYzJL02Z8DSxP2TrYprA844GAIWMXNQjZ0DHKaeLFmwMyy5BXriFC
UgFXeLw9B5H/rpophHfNKE9ATwd8m1eA0l7gro1J1NKHrTNzhytmoVBIxFD9rjRsl5BgRER1l/lq
b7pVN6Hlt/xxKzlIobxNSrsC3yqZXjSkSGkfS9K7pci9J6CIbKDUeOVvUwSL5jqeHlkAYWLZTQWv
g0SUa5DslQ2jQoIC1wo5vp8CI8VGFfXj0QRJVfWsSIWT4a6/vuQtqr5Rw9fAs1WHCzD7a8Sd7Oo2
SoFCJcNc9Acub9Na4L5WS4b4k3k22kuLcBKfe3OCMz2d4agIMODFdYTp0g/ayYco/5vlJMkH5VPj
b4masjZ52muV12QIcJdYEhXqDx36SHj2PcEYgo71CLrnS13t4DBknFeWM845A9bMO3cjRB85Cekt
lIw21yERlPiLyzigo+SAuaQJyIasFmhNc8DQIRjimYMw7NqOjOGmxbUatp3oEpERHEwSOvtS4UGQ
YCiNxJrlHugDjggV7uzdflnafWR6hK9Ogpt8BMhkEqAsKvKdt0nAwZ3nU/3Uil3lmJ6R56FoWxCw
vbyDFs6ce4P4/Jp5wCdGXQbKvAr+QqZkPYqSmA6qk0iTXHejTp43neeq95HJa4Rq8lSj/SLvSxfz
u37e824yqeyWyoz0WpjoF5kVO1kOgSdD/FXz0OMKq4oVD5IYV669hxnNqYCBtWk5sakHjeHKnAzq
7h/UpxkdTe9XFVUvd2Lk/RbjIwttwB8CF8hat8xepCmmnrqhqMURcwKCbaT25SGwQKSmjYUgAXoZ
ZkJvvn/tAYjNkTTu5NKTxdEZ6Ge8i2CN4Va5j8Kr449szmS2O/380aaqDozDsy8iZoQeovhqjTU7
APdmhzblzt+8SAMcHHvtTEeClwxGVSfy1zrm7ZkY6d0Z1VijgEMiInVJB0rFU90VKrRjLPqMKQP8
qm1bxZXwsKtfHmBbUBaQW9+N6ROJp0O5ZRLzWyxSZkv1DebFz4ltSHu6mZvQuTVJrOIOVx/fRvU9
4fzhF4BBSwjBgst/KXg0JXQE7CEpwHjQR3EIeIpwAkl71ZoaVJ041tElAJlXAnmR4t9ddN/HlQod
fbRmJ/BtJtMPs5A1/RIFOBvmt/qFg6AcJSBc/6jB49d31AETxVysXo/WW/X1BjKRCoe6eQUH5/H5
Fx8idSOR3oSB4mchX3FDb/MA8fQYQXYy94XzhmSen/FGVBkFt7ziaB5Mm6MVj3W4hs7GfRupd5vE
+AFPJeyt/p0sltetgG6+4uvEMpg6ekLDQfWJ2LLmGCakHlT+ACQd9dXJwuo4DCi74pnmnx1NRz00
JOsC6S2U20wBvU9CChBxaljmFyIUYp4AdIXA6k7BeLLUWiY6xjI2adWPRu/1WjVuw75CYt6466By
aiSkrZYg97ZtdoDMpktfK/+abcEEe0ksPWe571BmqBQ8Hju0w5xHIXIzzrIV4H6A8C7Kcr0fe3b9
X3BgPUgPl6GTjEB2VZ3SXoKraRNLfXlhbhqa8ox5hj81qRsSij2YF/fS5W4V3WDL0e0Or4a2/pls
6K2/5ecZKzLc6U6NIqQr4RGwQEp9gGb2KuStOuz1z2NMVqfM7bdsNUlw+spG/67o4Rk5NdqN6h+X
BnCfMnHo5knylL/PdvuN/Gf7mxTUCwU3LJ+SVutfxvUuG1zrRG6Y1XYBtrP/9SlPseX/KinMSmGA
dbrkrflDh87kRRIYlp9liqwoeApVbwnQ2r0EZf5d2/HFIVXw1shRTGZJEtDNvrVKwKFaNeWpmTeZ
5HQ+1GyPzxKjEaqBSAwg5BmBYnY+Z5rj8x7ks/9VMj+/gpSBYIfEFpcjLT6xtfy5Mdu9igQV3GEo
RgBDx+6XfhqmZvAZQ4uHIxwAESYCjjk686v0e8/WMGsDMl/wDK+BIlnJ7egO6gyCNnAVlRxEGdZt
6vbJf5cXRI7nlt9nK0f4dS3r9ZzWMVtxZ4cL6ZINIyNmD8TNBvDmwqav6U0vxNHSGPJvQMDRBJpd
DA2aqfShclONla/tlBFdRAhucEO7OxM/Q2F+sCsQsoqojF0vQt8sdTHtdhrXrtbXVmwzBhhyNCpM
DYKidp0WMeDJHTvqopq71TYFcT+deyhdxJnDHGH5AEO67ZAWGS+iQNTsGceLbkEOn/OxKW4eXFZ5
05bcm6+7vVT2dJSfUQeXOiWT54nqq730bnFeIcx8rSYWCLkj4DpCZgd8yP1FTMAfTowCscGCxu6f
0maJ7yIAGuPFIKVOJHRrDFfc93FrCG/5K0AwUUX6Xp3rPjEoWWQWUvRiRu0nR5ManukXNG5KagzM
WrcJDrZTRy9UEYomLxelFPwxFnlkbjzB2jreMLWqvIruXM7KjmTCv2LyA8rPLay4sPPA0JS5m8t8
4fGWHC15IQNgGyRZwtNk3WHTHbK5UxhdMI4jCC6xSoqwsYy3yIZMHl983WgvPKCkWll5MaxIK72a
lWVPdN6gDJAn+zcWjCH57+fgR8cGHazXZcGcyQim4Sv9fJyyXeRn+tka/CU5y6aDwxms7J1ChMoc
CZyMe5Rv/T0tcl4gmNjsmQoTjdCXU7e1gSwvLnq+TmFTZ5byCO8pO4anA4cMb2cHQoDDI+TvPlrP
3lNRnlvlfWY11hUhENfVavJ4x2fHfhcu4jibnbKaUdiHYLgXpI4dMc3TzgLje4FwqtXxoe9pOglW
VkPzVcG90VmAhUMtD7hJLSrr+Mtvjowg+7QbwbRcUVNhJkQmVzMlhkhtK5qPSRAdVrohnJnT3+/1
Gg49EcNf6SQnZH+CaDUxZVmpxfOM9IaXqlH9gHUTVzhmssuF9jFyXk3BA/WR9432ywHQ6xtDOzYK
Vd2APy7UWJLRxrX06JSlAYDVXiI1ZtUBWJRrQt1z36m10V0+bhFoFov9zajfb5nLLw/iBEmTAy5E
0dup0GCgrNZ4hIGEfmK1r5p4onNuK+G5wrfNR4fQh9CtL5gGB7YW3L+Z+IdzvWwG3Prb1J4rtpMK
skwTQ93LYXFdxQ3xVXD+RYTCDd/MK9FItCoRA/gXF1d3AqUAwpBlbGAqZtKbSenV4Kj1gxVFGrMo
VlMmUxEcGvvjtFolYO4ZqIeLBfqyw3z7+ktbOkpvKwVga4JZvT20u/S3xpdzxAN/1BqgVCy9FOxr
XJLN1yKCYhWdgPEE+19mhXgfhMTS7SKP7Xwh0KSCqnXgWQTE+PeW/jK6C7LiQZrW3DLZ/d5hBXGU
Wx8MK/qZQpziHMDo6tJpj8lJZTZdeFWeOK9cJIhM7UOar3iiko6fk8yQCH0EuJ7uGYX7It0WYxp9
8mNGd1gBjvYRMbZalb2AhOkeiNuie0v/Toi2WnRA2ISrgUjB10i/dE6j9hqvaxwfebpXSPE9UZSX
jlh8P/uiqsl8tvgZrOZkq4QFoaikwvXPUKj38w0qzNCC/hV9+EPAGI/50OcVnpTuRhBPzpIWVQEE
RJIDp453oYsvClmsIRlKfk2p7efU54JB/zPeM3pXWdykxF79GjVlIYwl4SjIZdbXkeM2soxyd9hU
5Q98Ca2qoaQaWUzaUJsalRfmhwlE0sJSTb8U5eNQyvzu+dixey4mfWrIzKWWfdqcZ3tNVCA3U/6/
poicPMC/tJt1L8Ntl3ynKpUC+rIgUX2QQr51xqw6POYdfH2EyahzhgVFlGNKO21p22Hjf6QSPlk+
fBt7y263VNSD4CSFR+FHA5s7yrSAuKpjylraU2/3GDOQV8efXiBiWDF4rX2XiPTGJ+gXjuzZgGvh
BYnIaJ2csXhkKrXy/KVChZkHexgsSRPDWb1hEEIojDEimXgZFZSz8LAE849PuR0T1VJ2iok4wGob
woNvs/oBqOwwCrllURF2vY/NtTVf4A1KT7ninNF115watYAYxTtdFg245rdbGffOVcKtKTOnDqKl
AIk4FeZOrpcUby5+XThchIo0NTuTIE1ddVi84kScv57HEt3dg5DAqJOEOLyX40QTkXgsycPrA0ji
U2Fe8KIeGQGrO/KcNdi51yj/LCk3oMcuM0fHUG6IzU6sBQdrDr6FzvlEhYKKTEY0s4c2UhuyXvdh
0aN3lewR6a6AxDCz86pVpu8GVvYC7YJJQ2CPZkE15EAKOZZuXyE/0Ivj8mPccejSdkn7t1SU/SWi
5B/FWtGVnOzKM/ex7qb9ClWDNUrXWgna/lEl3t7SL2FGeXkyDAtutQwWxf1KQgzETcMFFnT4ztEI
c0UHd5j6YpKQ13J0jjz9lPb2BaGmXj5K6usmh+WSUH4fY+KxNWJBPWMlFTlg8CVn1RsNEEMsMPB4
xRyOfe23Q+Q5qSmgbOnwTO9A1wAiMqei0fMO1q371eod3sWGhkSoRVuL/47IumGU5digIt/xeaeU
HqPiYBNbB2n/BIPhE/YoRf2D9UQBwXjQPF/FlOG0m0J0y7rp+zRKP8v5TLku+KkX8XZe5kAQeUJ0
/ZFMzU0Kg1mFyvbq5f/EHSrze2E4YYKoWZiCkGHrLNMfxqoShRAh01nMxV9SrjBuH19ytyenWd7t
Lwk6XYFq1KSg23FABSrGHzJhKoiVUXywgDJ6mmneYPZtVGcw/pzW+UnhRyJeyFKJijDlpDrOyxkQ
MmXL+iIlkt9ZhhpSA7vp7tFkNTfgAFysf290Xtw8aWb0tSHywhwteSaENdvSmAzcrZ8/QaoyLv80
F2ooBZU/glOSwPzZEyrqWgYbitlJkaXpgUjCIC+tMx2lUwimJx7nHdTb64PU3CSVG0K6vnQtDgGq
unxE9I5ztpbx8IyoFGwxYQt5CPz/uh6E73v40EZ1/sgazxiwgAL0R0eoy2ZH/5JZPeCNXdludVf6
GaRTmxO9HlWcWrc1OPKCnnoM//Wz41kj4ceU31cgoD0AcnJ+q0MpIiRRqGSGIowNECFn1nQe6UKu
c6kNLRXmOFRp8gJV2Dvr35yNx/lyxsMCfgH+PDOSqFC4PKM3KxaL0fK05B2PIH8MS17/2smmTLUw
lz+c5nHddXKqjLpIdsMcxbTH2D73loug41apDEgxFj+NimpDxbuoQEJQsvpoYZV00vImip/UsiGd
XymqemuB7Hro9wLZfKZMfyOzL1AkVq8lmZPvvx+o3t4m/emnnA3OQ8PJeWyI6zau5TPnJChFO8zq
Ito4BtU37pbV2tNaCIusH6c/IQgABBuAmxygJqGBZjRiKvl0PGMFCWXcsDJypfiMmLp+oNjnVi7l
YoHDJvBJgRoncAoPaFEz8bUGW/CDp9gJ8VVnR+wziX9I/a637QGNeyPkeFih4KKJGJ5tZPgtHVu9
dXxyTskes8GZaL+jzKLrHzf2QyZvyg6oukAvV7xfowsrle32zNLo1FvzIUJBR+9hH1gYA7+6Uv3F
qCTj85uTUm2bA0bKyE2W2ssb9qkpU7l6p5uabm5DGx00lKvUb1cNHxa8BxvvTmv5aObQK4maZu21
zp0AdOAvsnoSs9UlgXDxKm8wqED+HEDOCpYCmkS4ZTzpU03old91oUz0d+rXN1tOGghoz5e0k7de
wtgGqiAnIGugAssZMitVO5sxoIA8NJFhRNCukY6+UQXRjUMbup3O2ZD+ptHd6Do8vrgSoVD4Xerr
C7uyqq8C3jt5fIkvAszkyWDzv2oNnGnLMnAzmmXnVqvXbxgp0STgzAIY3/JdzX6UstfYyFXeEv0L
NZsJMdtLB7tVfiyxT+pfCGWepAEgggAqGVGHikpTo/0yJzWoc1J0sJjmMDvLMi63f09rs1O6oEgO
MycQYKTxpbDrawGOJO5GoKm++loeC0V08PC4wiTEIPKmHuorYcK6qa8HSscF5Gw22EoMF4dOX8Wm
lmLduxHG0bb82bfEu6hCW3jCrXxOugdSjDmnQV8LZ5egzra+LIfuKHD6dqX6vKRRVyrijLJmpJEe
yiUTyWonhSVteeFU2GYZ0+xOLwLZ22jCH+c3EGivACE+8rL4htzxuVOxFiWB+VWs2suDmIkv0mMu
8Tw+x+nP7JzraRwJpIdcqZaWN+ByzOUcKvfXES6G5n4zrJ8FlkUb51fHjGIwdj5rxYOD+8BLDldq
KaszNSff/4MvrIlDc307LcNVpLlcljiQ3DfjJSyIikShVKxb7x3g6p9i37BETjn9KqKNBhqZ7PNy
74N4L6TyurIQbZXoOAoTmAPSh/bXeR5CUCU3TWekMhJCRuUKnWmtfFjQzdbjzc3I17enww6RoJ61
pAdBcw5usl9lYbixufKH02XL1ig3f7SQp/MpU+N5SNTrdSr99wGQj4TkaXux1ujQFXTJgCeyBJVw
3zm6q/ErVNbZIIFQx+xddlI192E9LprjlnZtDpHbPnVcrJS2sJ0ddOzJBW3PHYES43+gEHpXi1hD
wryB7G0lwPoFKqjxW5ZunpbYNlxMc89xFgjUADFcmiRnvh0VBV6CUGkMVcB7CoJDLFP7Rd+0yQiw
vxTDS5nxI40eWGeKIQz01APqsZ9t4Ss7YlWHY+aSYK0z5g72BkHYxjI7WzUitr3cR1XHQf4kG0mP
ljFPca9z8s2iYEoBtBef771yOKPcvrOFrOpZ4U/MSTH8xO65ofDMUbcC9HFw4K0bTFEAU0ivu6xV
omEitL5gNiN88oBOpfgrtw6O4q3QGjD3+nHtAHf7DJINrjhUHU6ScqXYYoOY9SJ4+q8ElCUuYufj
C4Om+nZM/Px598EXwGX2qubMOvcuQ9B6Gnx4qwqvhAzBF0bzqBhj3405kENvlrNOkixP1knjnTHE
aNfj4XSwdl4z4GgFrOQwDIOj2dmN7aafv/BK8wLMNxdZgdZXrSQYctI6eGlMdJlu4+cLBHDjhLpR
TRqAN2AcInWKcuSY5B7NMaDZwG5H/cJcuNFGrhn9m2DnELVpZbOL7BkksfX9n7uNNalhOtn+ma5x
/XHh4Wo8BZxJ78188eAij9XG0rGQirYc81KvbHCM/nzCWeRX4epCmfGXoKWlNYrzNLI2oAhcdKU2
YMlVFboHB9V9JMtgWUu+fZ95OhxUUGGTf4ZZEN+xAGYzP5cwblZv0LwjBEYNKW0HjV5jygEEYIkz
oJTCsEIm+ZyvqLsFov/qU0w5Y2IFN911R7uQSI5J82FeBuQQlWkr85lCMCL4bf7wUDQcyucxDXrM
WevMJSvn4F5Glkwc76B52M+CA0n+V3P+5XUbyhjMRYp4hwVCnL2fCAFFYkpevaBzpNqIdc4mKdDl
kciN/fJAVI7m5/dkcTpoV1sc1d/DdsWUTqm+L19WNpFJGoI7MFKl63P68tg4e3eOQ2ByvsgNTcUk
nRaiBO7QAhTVY2MYKPNeCyHXg9a7qT9WYb6oMHgKjJarKnT1+i15HFi74iTh/d0gP4lzljHdNAxV
6Z8hVEQit0M/aqznZDBtktpurf9uB900mPUfzJdpuWgETbGRVFt33nytf78gjGsYifboZTcLKK8J
PuT7zzqE8AY/M8C8Oa2GLjAW0M2FuaohZvKLFTP1sqN8kEoMjV9wfrRuwnb484jRUR5P6dKiabFI
spSgkbL7YZxZ9NFePBuvxcjrvNv5GOqwXJ5PaLYgyqWe42Lpdvkalcjk+7LEtoZXqgcBD6MXoH01
/BAMb9FYjnKdYGyVZeQVhbXa7Ir6UO9DGYdL1S5pmFda8rBRTMR0j+lMVAxt7S7YLWIJv02/SF9e
v4JMPDMnsmvlBl92omJ8dXN4LHUi3AUaP9fUMComshlz9enA7UD1OZyeTVTqxM/SLVQ2WCd1AZvl
MlPvXJI921YkNe4y9mOULQDI9PV+sMEMIroULA6NnWoh/LWcfy2wb97buORCSYbFV3nNTfjA+y3o
ko0qCl3yXJQU0FI5P2V8R2ro4gvwQGDa1IJa8/DTtbL6P8IMhbk1sPcEgMc0vyIVz9yIv7XWWvEX
N69eURes5y54ZZ706SoL7M91U3a/zoGffB76WEctRwzOW/x5ysjzdy8epMGAKTMAj6KJ4kOJx1wS
d7OZTrG5/wBcq4sU+G0kCQ8UnXuIRk4a2Ioh0UQgfQa2W/zdpHwWOPlQ2DRRT7sYSFNbLcBy0POX
wmiDeI4rk3a9Aa9EPykzKy41j1BLVxEPDnHgExETcyu6E7MlgSQVqlOzO5KNJacyCau9CIxRCFNv
x7QAchZBod+uI3v6G6KSRBY1HI/MTQfeQ9Ajf7fbKoG89DBSCBvCwPQB8K6e6GLhaTWOuw7kyDXO
tgR/ARnGquRD2tqxiotNs0+M4OaEnB06t3Tfn2h0vtxfNx5kK5a2F09m4bKAnO/EoKCN8a3aMoOL
q9cAmOqfkgYmkw8mM7V9cQDAYNoCB/658zfEVjkUnd4aoJgLCAQDkN0wCaZG+z7khnWr/jxoHG0x
/LhJUYaJ5jGCQDXVtZV4Aro/eQAXhVNRkd1hjXhpn3orbJXCZtquoZudnxYjuwwXlYZ/ihK3ehVX
kxPAlTBQmCttPCMxKZOt0bmUEpko1PylOiQN1xiYOaqw1k0ISvji8Q3KPuXb8K6oYCwTWUrjQzgy
qO2zCkyVJjFmc0cNctY86HlGDa0XjaRgElmH5NZ7LUKO7GFHoZqcJZJpiy9wRTEr63dpl5Cz9ml8
6cZERENXtK9z8wzQMkk+J4e3zi9r9vpa0vlqXuvvYFeUsTrIYjUBSTIXTgEB+NHWxXpfSalr6ycI
D8klP3wU9uR0AxrdVsyvOxSHzxMCuTwDSdZR6cnXdOaO91pp8HzqV8dISPzLPsElzY+n/d7z7E2f
ImXjEpZxazPAPKaNM3GW7MalExGXGZoXmAMZ5DGgFW9T5yola74539qUNCpdJ9WHcCSpWRiUBMhH
aGqkeoSCvYhiwEdT7WWfkZRFzAegeKoWqVgpye6NgoxP3BLayFTVEibbiHK7BbV6A+ZmQoWWluGj
qWWhSz6BYgwevT/sFwrmFXhcet713rt300Almnzzg7MxJLysxRmHEnc1OdJeinidMvq+N6b83S/j
0xd6ub4hbJKWE6WEv+FDF5sfelv0akTRNTvGIBH0lT6BAzl1H3gWQgjIkyBoLohFqdCcio1MvbNA
yJzKICinWLBn3yRcWT/uR/IzlngFd/KmRlBJXfA4wjVQ1uGQwFwFbCKAPPkA05qMSXCUFRPna/nc
nIxjV6CQCAjl1t5uUVTGZjOMFfdocLUxoih4McOk7SQkwLiTCDXCbVHNkJEj/17U+0gMuJFaMJY5
HNeIJes8rWu3G8Ux5E9f+AuFZw7vf9hHZHrlHYz0NGWWrBonfRqd4wey46CaOGCSgWrkmjHXahGe
wV+E5h3+6EtvoOYnuhcz6UXS+iBfCy21MOoGQCKaEFrIP91+L36Bf5a+dKMFkZvvnGyf/Z0fhWGe
2Q70oPhohuFfrMgLVBFWU8/8Q+xnzILBL9YIbuhmrobDllrwIxlIhrTcjcthbVbFoOxSLtAp9OpU
8c2iQbKMAprUs5OTW9RdwY6DiCWh3ncr4H87dUPW6QnZaLgeE/gVGrsekO82n49Ni4YpnFhzpI9n
t3e+LESk30WLruuahN7X0k/ZkfNvTYOxYSTEuROglonsXuMFkUkd4k8ZR8WXCQyP13Wf+IS1FOlq
BCwHIOTh2neL/9e+sBVGO2lYbI24ULvEccuZwPrqluDlWXl0UuQt2j9asG0k7XoGPhKpts1/6On5
E8/XPXTchTllqc8thWQa3RurA+ehWIQuI9E/sA1Ap6hvLOjbLvhJ197PqsVS/6XwH5/p+nP4qjH1
2BurYz6THqPYFtE64+9qle3rPirDRsZVWbDlqyxvM8MqvyA1N7cy3ToDiy7lp+S4Db0SL4YUCJS/
4wM6P4bxNlPYHIgwI27k+K+2sdnLlbAlQFUOdp4fADOlnzPLQA5sUQeIEa7cSMMepZhBh/zjzATD
O2SM+SXskPTiSnSQv1uvqPvqKfmTkPe0scjWqbPx/eP1tDRY+pN8gLF+bcmxekI7OLLibw6umbHk
Fy3LsbCF1L2vyipXeBBJDWvskohDuxcHY7dSQY2D3HVQ3ihjbJXjrTmFKS6fT3JU3qapj2rlrAQO
VoR0fcZ1mlNnuCLK1bkLKa6bd0Xgkodkopm54Cc0qaHz1s744ndiJ+IMK6wnYnjoQ2khgsAfvY9c
QNZ6VNG6CEGsIEK3Vq2ksK+XsCrx468W29+7S+4cSlFnHPcGStu5YQGXrYF2oLz9lXJpS77UYL8n
PibuM1c2wGNowa6SwRcn6S+Xihfdgd3gX0HMdBL1kHiTlqDmccj8HjU7kkoxekJihzGgqaGL77po
nua8u9xzjIAQfnsOB+GHJvs3L+dv85OC1eqrGEIic49DCxgHlL0dBwz1XHwRDkj7yITyAo3RK7nG
wGTeDUjrxIrGhb/ucbDrlkf6OC6qcyuS3/00E8O1FykolZDft7lpecRnAvr0NUPGpY9DXXJjA63y
khfeQQmsdISNqLA1Q2MgweiIm11f90ZSbJyBWffyOaWwulDNjpXsMMrPDGABlC/jOJ1Cae6G4+dT
0ARebbo/v6Qy79nSQN3qx1GkS5Xh8xpGBlhGMKO/SLZricYxvIlUbLNTZva1Lbf+tH/z3kmJT/9o
KKhgfjyw6me4LQaQE78nKG+8ph6r9HDSZrNOWoIGy9NJ2NlC5Ugb3xroR7UcyFrvH05Lfg7D1PcA
w88fFdJIluhNlmoILavx0P28Hj9vRPICvfWeS/CPAfbUEJMUmX/DxwYTgwHdgQ443DdiqtQi210Z
Qd1rKhqeJD2P92ZBP5V0kvSTd4L8pRzhifzdgSzgbR2s5avTHTffAX4X44mN8OfGVZTjmBTDgfFg
Lzn4jXbkM7xvnfImRWtUJQ60AOwfEzv6T90eHI6EfLjN7QwMIYUZBJvsUa64oWkbo6/niStnbZKs
/7fEIkZoTKv2qwykyHIjRDfwSFpQfX0XA408MIEtSRqTIYjHYUszrWRcE5lZ5jmK1te/TfmSGBtG
ElW/Uc330M3zl6OmoKyUC6I9R2yZUe92Lbud2OvCtv+cA18R6vamLEJMiCI/bYzJH8a6RhhE7MDe
AS36ucS75jUXmeuXy8+nctMoFgrIhcVHZq0slYcpBLW0xVa+Nh264bqDXa6JTJ62HF0zjZg69fYG
wkHveCtCQsMfkjyDtidjCLdXnBF6mYrdb/1Wj0u315jASz4ijyXN7Y7v4RlBPzaE2tpiHhCjjBjT
w8ahd1VF1X8kbcePE6d9VDIHUFititXtCMiSELv8QV3Cnw4nKl4pbJAWoQw+i7V7Sr31NvmOQ16W
bBTHUVbBix/iP4gKTjaBdEiEX4dr9ziozFEiI98fObJflbF+mHDpE3+WSjWoEQRzHmHjqxzh8Pki
yR3e1IfI3Le14icCVYPalzLuoiW+w89CP0pNhRwx95VrWjidoDiEIPXMNWI30N9OG+nRts4stGYH
iy30V/IdJWRO7tI/o9h/EHqWi2tJM3AFtiAbVdNerwA7sKoDOBDWpUNL6GI2eSUrEYEMT7Lzrxce
H7qbOElLHh4trA1SUM7BRf1MqZvhx/ZYg5TmC3zoc1+CenyHOa49vHLW+5jbb1EPFoCMc36wntHe
V322Pw+LzdhlDf7W6Ae3Wg2EVhFHUYUxgvw3oOYb9pLA/bp6DlOGbNLKYo9V2yf3FqUNQRKpagGJ
lt9/be1+upJFm5Cr0PqRZJ+68bebCfzjszAMVRoQWoit0nMSVPQR+2rDr/BVr9TDBThEXeS6elMC
f63NjSjVf60mKFDv1dYP7bw/17NhGuO2lo++Y1LQWCfUwWdVz2FAsm/HyVN26TiXdt6KjmFBxTy5
++HAcwtxbOgNYYOpB0Z2REtrfc2D84btiFuymyYk3uLoB/AB6U374q66+n53cYcZlxJka0072eQo
lHrdNWBrIz2uhOeOC5rGNLCDL1e/ceqpu4KcxAxBHlBEpAqqe0kIZxRG+0Sar3lhI8ft+mwIk6La
+V5cZYralWA8mR7SZAldExg+ckBo0mKY6JAt/kcxS0UUD5BHPmKMIUxjn48ZnXQpG4b7s2fOFirF
2R3CiYj7SZtYA0g0VVu50kL0rrmux2ELDpifLFVUCd+lkNxxgBWtkAH2JjrkMaTxRnJpTOzfkrr2
cdo5pcL13lYlA8zVt0Oxhott4jQXltfhc6wsrKY0M/Y8pJymuBoMzM1wex/mah5e/rprV1j54DIy
/wfKVw1TD26qP5Iscv535CZ3DV6Hspublg4rAXYBtDRMhe6YLWUWwIrl+lNqDZ6EKLbkMqNEyU9E
HfLUeCp28OkcyUN0gI7N8TcZpQTm/hsjA9gYdqTeGtzD7Ky+Buu0PCwxsTSP3pyou70hvGpVae60
xK9mMWTCT1V3PnJNpMyxQl00FtVBzsd2tQG//i83PCQNVz283ZEVF6HRpaAZRZ58TZBLRN9Mcnfk
ktKCdyKI3Bqn+DZttZWYJCPYd8906s8+Jsrbn+RawbpABnwolCjI2d0s4KrTvQQ8610AXtdhGi4A
1MZNccIoHS+EcIgmUJAZT6Fvu8nUwWOuxp1MPMichsUADcMu4wegvdmrzMU7huv3BvRWB1HV0NNU
a3R8KL36V7nVnaR5Ed5Qm2JRdg6hBCGV6/tJfwvafMRoTKU6uxqIskz8q8qqtQjXfAG8VLwVPNKS
y76JSOqWurU8EwRT5VkQENHtpQq74lzoTreuScdl0+shaZ2qlI39HZOOjruARNBe9dVK0cogNkiu
TBKNjH23/mcTYNLkmteiKBMUtepfzSnw3ObtC/mRSp/p5q6P4F/sVhDXpwZVhllsSoAZkACZZz65
iwW9+7IZeh1zzExVTOdoE9I1V5LtIjCGXFBvsb9wecn9c8DqJZWDDKFDQppMH4JeUZ5CL0DqHtJw
br/OYosHxlDQNHN2butOPyhl6Gomz8NuW8aq3pMIu9s+7QmIxqOgPjv/+oO0C6kJLo37yHXQQ0Bw
lFwiETnPPXIJ/b+KnsdZuAi1UQOgcvffD/2tHM7/rnuTG2JjzfE9tLL43re/Hn4jqiZjX5TDCliF
IgQx//5yUQa8sVpIlwMbPQfrskDJFw9m7W1/qAUj5NKoarMrOePmJnaBgTJd0JM2fZ6sE5nrqo4l
XcTIuHOsniLjOA/eDFv2a9Yqv0i04BTGpG/ymsUlMoN4I0KdG1mjuqUqIAilVbUTpAZ1406+QRgv
U99j8281XscAH//8CepMOxW+/r3EzLeWYk4ax/ze3SL+nBq8ElAF3a497zgE5BKVTfZSdzt/XZuF
ypGnpQgduJt0Fp95sXPFcZUkoK48IWHjIkTeMkgAU1NZO1anzeBO01zKtXDflUbZ6I+m74vy6p3i
G9xi3bXPMj4zScBAcdT4FxPxgJSZk4fqFXHrasJo4PWWki0Syg9iDNonJSoSNHAV2YvzfAB7qboS
BgvtKImDkNSroGufRlLQ6vEZmBTnXmL5k2QXZj0ja7mNEOSTu1RhGItf2O9LT0mN6+R4bCcyf29m
2ph1VXAUbdOPpeA0wprIrprS/y6keGCjiCXyIJY1ZkYfLAgnE9pXX+W6Vr2jZZR3BKlyxvF3I61V
Xdy6d07HKHx6ThIojQLMk69A3u2EQw5b5Ml3/EjrA5/EogvIa23wHsFfblBtMI8/OhFMGx3LJ/lC
t+cJssme5B4rLpFMEaxS6RH3L+IV/eg40aZGGupr096vtvk0uE1bX0N84KdpCY/QiTVJ/X1JjE1A
ROdE0VjjbKeBHFG8FQBdHgOtHH6SVOtHwnbteTBEZHskLgWlkH9yyAIniMS2zc0Dap/mfeRdCVcv
vDyH6j7rJoAu6byiK0MjVKHvsp6t857ZVTCRwB5Tog1nB01buinJwNe5+dIsUjrnI7M4aV6Ta6ji
xkLLVN+o9TaY/ztfJTcIUgHxFbxjxAjWS0NTSxXiJc3eTm943lFG2n3pCc3/p5TLCvmKajQn7z8T
QWXQ5JhvgkwuBYj9NGbi8+/B55BlpaWwhlz//MdC4oJnO6GuaJUFHJ2SQsY9pttkgpLaOzA1p4zi
+7OrXOJm2wKpSEFl/O66uPAX9ZywfddYPJlm4QkGoJvw6CLqkVEu7ASetCHaXJ16t0cvKbS0t+91
saLJLG8ZV6ZjmE6ytBl01lrj/21uu90HD3KkJWItH7dRNiYYl8+Man9NbQSz786dbrjYWdVRhRLK
2wJ2LHPmvybt0yPRvanb23bhr0RYGQW6mWrFg1JIXkLp6cTljn5oAUX8Piobz4/qX/SrQWNAo2qg
8fSZeTDQTkljw8YP1X0BJg+mAl7egsKg1g5oER46+mYkAAiro2tpXIS9MMSjZwgj6sH61ST6Jhma
Htdjk0fOFGruHonrzfxfJUsTJwvWlaScrQzN5oTUyqlt1En84RtKdvgEdJOAkCf3V0lxPr4rPOqg
J5K0WbqMVT226h615MwCaNXLPTrmrmOVTzbw9mb++VdsBjCFd6AeUaYbrKfZWI1OHS9jO4q5MbsK
+ZzM4ARRulvh6MDYYPJP8PcinGEzinFVjvfMcZw2MRAXD/h7vHU23VBxxa/hw36qRR6Lo5jS+R4+
FTN44iI4BBlfuGaAZnSP9KPgN0hSUXv2hLAc66stxaSBmgnB8XQj80/b94tXJN1XT0aWy/Rc1QSR
I43NHZ0zcNTRKLRC/py1sgJ04uivzBa8o+dtR5/wC8FUNLiVYL4k3m04DhvnBe8fNa5cGfn43n9M
FEeuXoinsNbsOJyMQMSiJZ7UEFPRt2deUUcihkvgcRBo+52ikmVaBzYrqfHgXE6FEosaldPD7vW7
wBcvb8azYPOvOyc5lhO1afVkOFkCrvEO6NeaCMoq7FhOGjQ+Fq+RqHsACBZEEMJUx5M/WpjQ3UQp
ZQ0dzssdFvanD1VXHKJjm0OGHDg8aDt6tnGe7LGEpREGN4HJtQi7v44FxgNLDf3cCZ8OerxFug8Z
IBGUiGmmYJ9ES1LbilM/moziBVuZItcUVSK5l/6peQ5fjM8g8ZdH3L+emEiG+2Shix4JC+ifFSsr
O6oBlTn1fo6CE9+fTw4BuaGOb8XF3GR2kxOk+XFyGHEWIqDGXtXci+Eo3RQ1xmBu/teZnWfaec7a
GdoFFMMIwB5dMAOrUPGVFjOiWZcusoQn5Qo2NKC8H54LMzE7DAVqLrimdgV0D/OAZopx6vqFuNyK
xG+HfsY/ixzwgpkv/fYESz0WIFpDoj4BPYp+7a0qY5DwTI2TWAvZtDf4t+dtEn+PDUxxdJuFH49r
5F9C97WYfS867/8Ns+hRL/VI2H9hyJ6BTy2TX3G5/JxmE7oXnyWiSKbV7h4Wmt+2KgOMw0x58XTK
uozOYdbqI8wm3qQwlhubLQHmOkyRLDIUcPqdNe1LorDp8s6zijUqWvMuwFE5rAtVVch2Q98M6Ch/
5EZo1F6pVUjcXJfCGHBnai23MveAWPLM4uqKbSnbTDW+rtbKzs4gcFFTqxXocNnFtZCYbbX7z5Id
zs00OvYR+HoMzl17UUTxg8m5R14qxh0FEg3UFcH4XiXxJlOmLSzmEHa4U9PcYahvwEL+uDvEF0qM
KmhXwjej5IJUhTAzr2PqEa2ceDclYTGsWM+Sga6FMBffNRb/wxo0gWcPGQgZ3o52LeDF1IpRZ7Ju
u3VtgD1oANT8wpLwI0qF8yBuSSTR8dhZBQmQndfQyUxIprrF3ez+zjmPxtTc6m1T2swccZU7JtUu
1Z2o7JXX+H8J2Jmbve3WgGHyckBrQBHblE/yn26+whxyPH/Rq4F2Bq9nvKq81m7HPE3ykV2z4WEF
G5dwiOWBTjg0sq3ZKGoc/ujeHLU8UFpvp2ioABBq6KYALyJiXNB3w97RBD2qMxs29AY5rCnYaCfM
5RymMKhMFOchjE/OGgyyT40muvJ1YPQi7cc1O5RsZb9hI8edx10f7SMYiK72DMv73DyUh6GtHizG
fEmwK7ECvH8ZgNFR+eHtiPiWxolVjeLJ1pgsftUwPjJwtZmwoiGSQlycthwGIVJPe+dOdgddusk0
e8SXUl1hRltxnvSM4cLAGccMnbcnND40dhy75qCRygmqQunmPWFVxLgCioyEOnyHn7XqNcYdkFJe
UYOsw7ldwMfdc2QuDpVQUdRO9allXkVQAxOivpvnpCdDckgSnN9AbpaKABrbrBOa6dwdPqggAESw
HEV6oJyqIwhfwmnnaDz8GPjaqsH0X6vi3UJ9FK2Jt6xo5gHD30TJ1gYx4XsuvSnBD9shcfH07mqq
yKFv6Ry+NHDYArCeP0bYwQjOFY8f6IikKXKdYZOibZsf32Ksuqi+4HuZPWDAwgOucu8QAbV9hUVG
YiLnF4HhDkOi70/4Q+6H+vdvbPU/z13Sw0QvYjoWCWIsPoDggcLrq5udcn5j7md0CS+NkR4lMOxv
8/mN8I+WoZ+Fr+n3Zmab6SPb0PnXJuC9dotM9w6p43xtigq+Rsr8QZR+5O6SA7EcG3s8kJHTWmlI
up46YOvsOedNdOubNWBjVaslIqB57LZRLWQh2LKx1CUGpRfnfL9jSDi43uecZsVxbQr0nL7S4H0J
TJ7d2PrpwrbVr7ZE4rVOuU+DwGrZLcslcL5o1XGgvSBpMesx68kA3XMieWyMt6YxRCP6ISqKwoSo
3Pco/HgXnrKNS766YWOlKsEgMdc+wu4g8mipLyyzrBR2iFxwmY7H4upllDce/rR4IRhMu29zoc2n
LJ+PSyXdalF7aObZLqBbtXsAfX+uAlFMXLrm/AKyiZOzbn0M0E76FcDqg8f6AvGRYrdzQv7erUnX
a3dOxBOffddWgTdtU07QnAzoyS34mgX+uTedTG+CKdB2+iyQfK2iKX+lSDYsmhR9S4sfSNXcs5Ew
pZhnXpkXSTcjFYx5F7IM+9s2/Sdf74KX3nKLXwNMffhpwei5O2rDztO5v2qZsBwsGbPk7Aub+iz3
gwk4RIXJU9pkSt0Fzd2sWp0fZJSxtrKV585cdkhfo8RRXTuaIAFeUdAEUvLV0iwVGtQ9OO9KwQBF
JV64OmYSHl6r88eta9NQ4mqaTa0hk0+2rvn+7FcEYFRIfa+Nz1XiyONOtjAPlONTpCU0T16G6Iwg
JAgD++d9PDf7k1ClUKbZzrjiz54i3Z0mTwR7DlSblr9zJKgeAlQio8g9+0nvFDOXWGClReP32TQu
B9sBz54GLMGO0UDxOlVwOifeZkLG/TVFBllqPIgUs0+crmx3Ml9XQ/ZlOPFftbho3NXKRGzYCWiD
TRnh84JVZLUm0OpajIN0SYMRW14SbEHMW8YGQ9cgG64a/ZwV33zJjQGi7BZQRVTazIqChZSMyPxq
tHN5yHrTQRrvv+K0FiUsrnRDzqeNSp1vza9uxRoCwjWeL7YuJ1WAiLQ76E0uxbLHOX8u4MSk6Z4x
cBqhPLFhmbF+Q8eP7ECIQ7+uwE4GPK9UgnjQQuPxHzjf7WUxW7LkeppQAgQHrBeehrBADKI8B1W5
hhxV5O+NDCl8f0cAmZqqyBw2WY5IX/q8AbdhPi0cUDHHgkgSz+3NlsJdwT2mdiJhCkDgBFxu9chX
2XWEqFLiplc5nkcBnu2cFv/eIu5TlnAH1qyCVWpbVp7sm4ntWTnkRIqBdeoptiaGxym7izVvVpjY
0qH0LFmJBgvBZ6nqJSG6PlKhtIQ+C7hgsMEed0BzXw1CNGVFClXpk+FIrf7xMefeGIAYsBBGqpXn
UdUOG5M73kDAlOJL7tkpzcS7htzdmlvHc1DwA4FaclBpG6DKvMmeGXfjlSN8R//gqYTYA/3rix+G
e7Sqs+I0diJHWor8rgVQCMYuV/1b7MzQ/qgIYIFlpm5CrbwGR0YZvB7gfijaNxR3dPU4bUv3b7Px
Dp45PgrNVqUOHOqqNq8gUvOUfv9vgvNkb2Qapi15BvNh8MrBj1AH6Yh3ein8cgqOvmInkO3AqclF
uUetKOYo1yyekPiA25OpOlXeAUYLHiGz3Q1fPI00RS+oXFynLlfV9kdBE5g4ySfR5Odms0Us3Yjp
F8xQRTgiFJiKB1sI7Gv6eCrNBKTzryHkffRaahMFYSJfDDHC5e2tvDGxffkJAR52+2er4CvBlN5S
rVU9eLccK0QgZwXMdFNodHp8XgH/ggeW2pTYkUDnpa7V+GHkm9o+x1oIj+Z9saaBN1VotNj7C/A9
628TYNOZz47dO3TSBBUnYPB+01iDRS9XXhwT2xIBe8uW0CwD4A08GmzLlEL9qfuNryZA+JcMlLK5
lCT0/sA7Z+SFrcgn0ifC5oepbmiY+MkP2JYNhyGI4rk5AlaXPQ4GjBHSn0DVyMDyj2fddb3O0hm+
wGuAYxI5CRz20258pJbSUhevgDhnWHl4uQqLFhUM77K0pXYffDiXzlNdVLt1UU7r27JqJ12xejCD
BS3tczI6XMJL51B+unFVI78anEmNBuLfrPBhpbRLaVPUjlCai+1ao9MflWirxO+I37MmzJidJrcR
FQ6ZBdPdEX25BrqjG3AXTNE3GeS9/AvhrO8frkMMubN6Tod6kDs1Y6WdVIvvdzgdwyT2pmZwvQzG
LMeForZQI8ItFBlXYEREOPX6MJG6WNOmyZ9lMUg+VgqUx5xlFrs1bzMmR5SHE/QtWwsO3mhG6hf1
26jRHEejLll8Y3d1ddrnR5TKfobzHt6FD66IvMytN2YAllx1YNPyHJvCV77d2VXrk4DYmmnFn3Wz
Y0vw3rKZ8HZAZHhwiwO9T73LnSLOvljW69dmIapRVTWy1y7d0MiHwrXJ7e4YWo6LAO8ZsKeiwbai
6fD3dsxpAxdi/AUrf246GykGE0Tdm4pP8if8ryvnCTmOkrgS1/z8eo8rOe8tR6RumnrNqdNLeFYc
3+aQ1EjzRCsTb53JsYMBC51Z1byE35dqC2VY7ya7voeVgKlySnz0UOmwjZNClG37FUihzo2KNJXO
K1A9+r/EBIJufPtlRxAZGNEkz9TYUxITxIPzrGZ6+j/g7xmbcSZxn0O63ONb5T5x2IOdhEUmdlom
vpkY1H5Ca9NWTOsHavztt48iSOolhGwiq9tYB7G1T+K0mLO330V5IES8QAYblXISAg3KlbPB9M8Y
QpcFGG958fKgeC2W28t12huzWO+fOFEfSZB+MTb69K2khoSeWJyYG8IxEDIUkzWcbShEF2fodT87
WtcC2J3dD8RRUaEb3k5cRIj5KX6rBKoEevWOGowVtcawI6Jh6IeHEq5qBMyFRNsmqsfSv/ULCPKK
9Eu3o5WaTIHbeR8lKKHCEWyqKXb1Qf3glpPwJB1ipTZGcjPZ3LiQvx37o5jnOjdmjVb6vYCUyCkM
ufnACNXeVC28P3r+Lpvo1kLYyJwkScs2Fh3vn8Q63jOYyAadDzn/X90ODesPBHJMUG8O1quFIAaG
rbtG8/9csrLQ5AOpYfFLExOPtduoHOld10IAxaPwNhFE5gb7jOyMW2ld59eF5nyQ5jXBj6e5Vpal
d+qAzRP0S9JEg8EwxoUnfyi+PaGfqOdk1CKeYCexCJOdzIB+/2k1im4Q7JA5GHGqix7RUOylNXqG
Zcysbt2hPCPROTuO5YtfLJYfW3BkjLlpQcdQ75YE3qA3J/zWrYvjBnQkuJryKnOGCtW/1wv+9JOH
KztZrWI9pTLSb4NfUtWUzJNjibSs2FUvMLFljSGhxJieaf9LRbbdpvxdfJVai0CTVf3NZtFku24t
cb4CeV6s9fnJd2zWIK3jDTX+lnQ2VOMIlpnQc60f/i1qMNFqLFwwUcdG8ffQE0bh0jAlSAPM6BdD
YKyh8LQMhAQ5VsMb3qUcqMgDZhD/iEnpKGiKOFNI/Qzi0DYe88iHf9imry3R0UEy4p4SSb8pBT/J
c+LQhlWdqrkDinqZjENj5qvYS6XC1JsTK2pMEupT6z1u85GwefvjeKxmlMnUwoT8ztBXTsH0FFU2
6SuWuw29d6u+KMIp8eMl0bmopQuovoD+nmfYWJNLts373UguLyzhLiJhnJgInXhC30W1X4Lov1SJ
/0kqeNSI5jXKw6hqX1xp8zehyC82fNkeSunHgtYHYN3gEdnfaIYbO7GPWtXbOkyXJhAz9i9Bbq5e
K9BhcNuujlm9njCPQY/mwvODcDWKbr7yllA9IZzbeK79lQePA0iZAx6Bqe0Anugy61z/84wzv4YV
2Lm+ckhyeQxnZAvil1/ASGfU6xYV4ZbAc1jsPup/IcxcmT8e5/YbTwLly+Chi9Obi3iUUPVBdCxl
jd/HQaR7RhMKmu+KuyXZeVDNFgWx2NgUFYqVkViPey2CTjPr9NUHV94iAygJg9LOR1a1orlAprUo
ytZp9wvbQ84aKDsojWnFSe+P9lWt83K9AV6WA2r6b47NltBgf4N2LHmtXGCiXhz9ZGHKj42j/aZ4
eIwJGGCHT+4uA3GzUZvddQ0wgsXH+eg4IsUjrtzVDgT4OrNXPB3g5e+EdERsTTa5vxfa4FnqJJd3
LgDafuUoR8veOv1QJZzJVvlBeJiMJ6BuNkMEFjEnXjYbSjbdKptM/Kuw9lC1IaBFo5l1+ZITDRUU
E9We1KK+L7JDd7HhYwrWOLsY5bak+x3/4DLYg/5nWxQw4yFqoE9Ul1tHGYUDhOWHTE+DTB8F/5qC
m7v+vbPX1ac8w4cy5lmPgQm82QXLCHEzuIMwxzzbElzQwWxW2TbLMMJdTWNml8bbvrENBI4coeIZ
Oy95UK8htXw4FunuK/OxLGB84pYnA+IXrW2ty7kZ9+uFPGcC+YKLu3852TbKoDuVj8wn/WDccMLY
ewvZxqmj8KFrteWwbyCErD6FlEYv1Bc4mlETc7qV2WKlLNqSR9O2pmIVdxB5Tar9Gntg1zdWfK4K
1v+quLutC7w0Rmgh0jerPFhZK8IG+qyw43wJi+9MFr4YNrrXqxOz51/Ge4TLK6E5RoaHxDRylRQQ
GSuNusb84mc16caPiCG2izcVSrhX6OVoGvtenz/18PpgQ/p1P4RvSFKPpfK+Mo2+70MLKospVlvQ
du7nDfAe0+WHdLfDWIvONmIpDAqr0OlVZF1HRZhdHDiMjVyFbSNVkzZd9rg+KK68U6JLspVAxNkY
4Xmb7ikriJ2Qi6TzCQIOFs0ucdMPTEeeUJhgnaObTmX3q6btR9nDEO6QusFwq+jAtX5Y4r7tmwg9
NVmkUR6oiBUKpZJu89fBulhFfaAbsi5zbdixuHWHjD5Y2TBb1tds8UU+58HO6WALykfX/Pa4oZ5e
uNEHwFKdeKCy9jhxv5tILEsPopktQ+JM6NUA+ILCvwvRal06ZIrB4icouyYnsQ1JuYjgCBc9vlB5
9ZsqPP86BQosaK7TGFmIkuQmGOFxG5DfEcpsHoIWS8VSUuqHU4BUqKKiyP50WJ+cu+R6mraSQ9Sl
eYwCFeaBzBu54fzepKwfFTYv5inIu2vPKf39+3D45+5FegLk052ZruU9B04BUXxGVjfRf3RuGzcz
5dUypJzxeAzJS3BabrWp7bnrWmdqdZ33ys195PaiOqPm4St4nH4CliimfZ4+D8lyiZKvYT6UzE3m
ZsYxtSe21NddB4fkUXRoUhCqNKU748Cntm+U8cSqzR4FBsuW9N1yD/X3q9wrnk3DNhnsD7qbwKDI
0uSL3OabLeE1MOOtyU+WYH+w9oGgxw4XPjCh8T9gAMyixIo74BpeI9e4atkCQylGotWbmJUpk1W3
SeaJjKyLBHs/bY5YnjCw8Cc0IsAUzgEm3pzHvYPEJSJ4jFnu7eJKZVjr1jdiY+h+4rfFz40d2OHs
xlsQi2XXF32gT0aisrus/dFbGOsFSD3B0dvjm40iy1yGPqS+REWCU4KXoMLJijchXHrgYLs618/5
ozkLrORW0yMY6cX+z9Pchhzs1J443JB5AfdaLvt5H7VLVi3K6rCwFz6nJVYm4wcidXrZoI1VmXqn
5jo6cT102uuN72m7HEKVVGNfqk5DrcaC/t2yKA6/JgLsoFHhVJzPhCd4zAgOGb/EVPoTeDUGwL6b
M6GUUVtp7i4v3tOgAPs/TKtp1rglrCOUFihsxCWNm59zOoBV7XFpIvcjFMxxL/RdWVn3U/5DffdJ
/GVDiF55S8bNWGah4J30AgeB9rmMlmuDMhecnw9tV8UDqChZ8bOjcRlQRDCInT+2pilbk/Vg1Gdv
aCjxG42vWNIr0MyzvpFoZ6iEAHaW8WIpywuYptHuRk6GZsrZrFmawighRepcjoN076f0Oc+YXSDh
ihTs9aDDuMEMdP4uIB/hc4oq8ImRJubK1USVq81OqQadFeuFpk72HF1At5BCdv5INz61fPHLQHAp
9i6Juj2PhQJ6MBUKMWAKSN1yd5RRfHAaUKRnfMgLf2rgnbMHagZIDTmFzMBiSmv61iN7wlbYCZpT
FCoD1egYWDUZfG28S/1BONZdb2ovDKisIBrWp+NDua9WQFKG+xOL46wWfcIZrjmBT3fGfhfH1ubH
fzn0OzK427QI9U2Zl2xykB8z9KcnzYKImXYp85ZVF1NdvDp7y9IPDYADFbcEsJ49LitnnEq62JQI
POwUpNOUF1M+de3dGjRbz0ijz83QCEW0LblspmFZYXAK5MKti9/0nZzCm1kEC3bfSJXQPMNr6Sxb
qWWyajihiL+6m3hmQ7vQTBzQRd4AVa4OK5PGqbv13SZaa5j5sIK/oMRKXz7YlxPx4DcDgaZXXQj7
taKF1088btXMVl2VIsA3jnsObYnm9aQ5zG4GEm6xy9z/qu8xQDX9HsWUIx7Fj7+U8mQotcpeqYwg
j92ouvNDwcQkxfafhdzcW4fVNX8Nj4wxF9wUSESImbNHWkaUctu5IOX7wSiomzEd+e13OjjZQPD7
cOs5oBbjJtHM1PDIxk/pcWzreNRRwx5Gn/HCYeQdZIqgwLIR4GzouOkgbZq5xJ03SPlvFgrzpPa/
cpO2OujxCvyvJfBAEZoTewOgJ0m4qdgQ615ulU/8rOTzLD/ej9MESjUfUrz5ld0uA+ryRSTZl/z9
mj+O6fbbPdLwbakplUY/x9qa4op9Kux6Yn5c4C6mTpZyIBl7iQEQdYnsLdXNyylFAS+an4q6RH68
Oog7rG0PQE7mz43Io6iXmyT2b9yPBW24ZHJFanCT1tnFu9B833fBgn7v0Quos0bCzMor4WoRyyOs
VETK4QZIDIAvthsHOcx546UYERae2+VC/9i2W5hsd8ZDJx6kHKNhhhZgYE9Qj7vBu2U0nzvGRZ1m
bIZek/NcTJJCcTHP3mKKKlJgFYg9FKzIN+vPdd+iIHAEyxpboaOSPGGYfeJ/yfi1aHXSCq/GPNLo
HjmieE3LG89flMhLCHMw3PcTOnl06duxgh1vWr8rr943PDBdS2P72gSyANAOLaobRwksONg1i5zv
NmV1AVHPAS0OZv9e20zpeI4fWNtz/0ZC/8oobz5kf/hFE6rR8rMA17sosE8nr+09cYNmcOYvZGvu
UK3hT+xIJr0m3OAriQ1UXknYT7Jx1ICScaK51FlRGR15dDYoWSmpzP4XqznPzJV8YsgLOi/Ff8kr
rhVgs4hRHXLC4eE2Ghcs2dJXs1YO2z9/tR1MvCc5u1TzWtnRHasEJgCzyR4nb2mcd1YqQC/8giXR
Not+Yf9TwzeZPk7j5ldLHprKz3pF3rBDaftZaWCWh8JnxiEaTY9TKGJzRvdq7otpe+eIYaKcDA5c
9Mvf1e+zG9c+Iiq4L+Pomq7EAQym8sgc6XQxmKC/Rec1jkHj6blDTyYO9sCgBXFkAAti9EZcXhJb
/496uSGDYRS69XBABSYhE5uTiSJLp7arVtbiw6xPyNvM4sllENRAVdDHBy2YfmXBrRp190efpofP
rZFbnlvl9amsx4jC8ONoqyvh14XQ43VxoF7CEaaTGfkwG3XLJRtJWGlePkDD93arss9fFIaPEm8i
wP1lYirvRCL86vEK98Actbn7zhr5oXkqJbPsGZT6rxFFotUipMfp8H/xLCNFcohSxPp/Ch7qTy1w
EuGtc3rz5X9LhGdu2+uaCgVS9pKEhhpnCov4Ix7Ay7XjxThWq9pROpfPArhAhFS9X3Wtmxf4h9TU
K0NMpcGEu8C12QXN630Sa7JnAdcqobzTrQGxrNdqZn1sHiq5NFU0Er6RT4yaV5Hc5W582wMF5Vib
yLDBSkYitqWDUDEjAKuFpiekA4HVfpfQnh0oEF7+QPRlOW065odQyG4z9NyNxnI8G/JspHQxsZwg
/4GXjATwnvD+lfyeeyALm0Y+c/zdfTi08mDmlmLxFBy33S9CFUn1Tieb9sFUGLHR1yS25x+gFONb
u/5BUI/x0PaywEtX6Rf/TBY/60ZYujKOwH2clffLqbjkmRxgvyzmUH/7LDLYiIlIFu2yiSpMh+/h
xdNnqmRTUActqsxDnYAr0vumIZ4DZ/iew/UcgyD3Q/mxCUg+emXA2LJizo/JClrhbKANxCgf0lrC
EYHCdGFG1Xh7sEvUCGlJz/H6gchSUuC3+lmZKrTxNDmYcsSNuykdPBFT7gWuqd2L14eSdh4juchk
UCBl6vPjAmz9NXlx8xwScbnBSk7D+kdGNOpChqlcpwndouxASz7jTnwRNZCuDPQeM73dN42MGnqL
4CA/Exfmi38K/22IM4Zqsk0R9kWtXRLktvi8Pvx9JA5X9P/ZA7HkYKKhi1AeN3HeuBHhceunZ13H
BfD/W0o7ueByUi03qA91bG/IqH6WzSlKoRcIiHmAdW42UhR/Opot40hPHa7sCcllbJ8fsKzEEmEs
FeX80Fe7WLRKSO2GzUUDC50b/P49gNzlo2no271jMEI/6arPhYgLZqt5VNmasDoAfF5OWPYHd5tm
mjcOYsvAl0i5kQ8BSVc+gI9Fu+K8ow7C58xdX9fKhh+QGOdQ4nKyok6P15lrr9OyiE/yJc8Eswkm
Q5CHAiLn+IgggcubuRNNPtpHECeGQKgcZKVd9c1SrdZqd8lvqs7Sx2RY5UOoEZPkoSDHj51Mk0Zn
w8LgkITi+6w7Ij1Z7CQkDCKUuAy8v0Hb3E2+/qknouDt7JIPlaCJoB6+C4iqemvlLuT3IxRxrvX2
e/t8M+pA30STqEEc4WSrSVBn6VdCVO+F5bJMkou9xhjtggXhq9KJsdEmWS4AGiL6Fr70XgXaLta2
SKwMJJb8scimIE/7vGRr5qm1xNuM2ER12YEZsYBdXWdH4bqfVMLmfZGGVXKWYbjXH/04mfbyLVi0
19sINtOHvOrE6trQjXfyQx9d/Fq67+j7Hih5dtWP3mNFacT0W9HfpnM8b53x7n+2skWpxP+QMLEs
zHQYldXx+e5idl1OsdL90Nuo93TtaPqMt+kQmcLdLMJEGJ1LsU20nUid3pWkFL9h4DJca6swec/6
V056BqgG2KkzxfmuYx2/FOWkibMn4QPACZbsba3k/lx9ATrt8wSKS/fw75P/xV24iFiXMq0ieee0
NdzYkIFwd+Up09sHKyUpoIIWoac3Pgmgb6PbXQP8ueb4Bd+pcq0JVcXMzWf55c6QpYFRtVH+Yijn
eKPPn5+fEDtIziZtYAuhQSBeqwb2L7G8V8ToYp9iPCp9Eb9o5Nf6SIbWExxi+8B/mngz3VBn1QST
wqpecdbIhlDv12wg0UzCXZZiROh2ZGrowZipXYkpriim5xjwLDyciAzLxR1WqYeZzussiPSOe0Ut
u9WpC7yMv0oD7DMJ2PTWyUxlOfI5XSw0ULjwdEcm4YUNihWjPZ6GSSWY9zIkCca3+Q27oRciLv7+
nCDssIkUxbOVvCO5y9gpRQNOgaHYTAQMsOPBKI3519CK3aiHfpC0vtYaUmKvLkzJ5cRUwaLh1d1h
ApbsrknSY84hJBcdNrhS+pR8SmQ/XhGD3bibuQNQ5LWrzWajkTXsFCEULFciCHIxcdsLfzsd7el0
31GnX6276wL62MEazNNYruPrImQ8YmuvouTYh1kmnEGlETs648Gr/+FMPs6cTDNA2zJmOu5PQ99r
lGmf8tFleOBGdxwFNXgz5gVVlxYJMmm/OMYVjbtuL0gOtsxsQH/0gQAXwHicviQlY7j5eKDL2Vn1
53FCVz6Sjr5/mQkccKY0cPtXyZHWNNbtaVqq6PWrUfM/mCobs0sOOcGRHeTsjstrPpN9l/93cr9V
p4OOnu/wleEVP3M/mEMLfay9svhB0Lujk0+FQzvqHBHY6tY1FVLHG35wIoynBrD9dlg3Ww5S8Mr5
w05rtR2umZUa0Kpx0oYpoMPqnVDvoClGB2KGUQaWpG3XusVFHpXXjFKoRhfGL9g5GPm9NK59b/qF
8p2/jll373hV7FLGgP+Ug68oB1tboK+b0ndcCwdfp31mo8hkLITMhRj8J6z/f3wVkfve1RFLN2b0
oj+elDAs6d1RAotS3mSeLfWKTXa5nDBhxNqHJ9GRqwBpsh0vwBuuE4fHkHsZ6T7FfMwlJHQ1k8Xw
C+t+2gYibYFjksevJv58F6OY+ScFmpF7BMDMlTiwOuOML8jlWv9u9+xRWhr4XWajkqlMT/jffcA9
K9hRRQqrVHA5meWbqlxqyxB9/RlIL+HbBCtAXFnagLikvaTvgMlpRY/Qs58vvQWIq4nltvRJJbw3
Pq7JIJoOAZTR0nOS9ePeKYuaX4OXYotaE0HWTUQw+OzrX314/tw8HogsFrsRLYbpNfisSheVtaul
mB8eFPXETMOWDXCYALJdjrjDhTaJ63LdsTawwyG990oKYPMoWG7QZz0Ed4nIf2CFuHbor9jD0wxC
PqRgDhCOYLLzmh9+VChxuXEasphbEMyWBaVbaa4fYMetTyKzuSNtSc6NRsbuEw8bfKfdWjavl2fh
8P+DUcXeFqibo+eV6lB2EsonMqdM65kxt9jhkZwEC/BT34vEpngRX6QwwvjQ2SPPY7IoIBl42KMo
nAhbJZl40dM5Oy1VcULUOa4KRm2nW9nihwsoZzYqdmE0/PpuyHuiPMgukf9VhJu6TIQJ2+nfJeAl
Mr7VfTki2C9dD6lr8/3nsR0BFcAWrN7fMSbyiOZ6WH8kIsbWhB2IT6CzkFXFXpyvuaW7685AeNHZ
voA0w1t1NIcIAt7LnaEDFuRe3wzLPqlS5O2583L5NxuaYKKZbe8WQ70JgCZtHl3scmlFIyL8GYQ6
C0kpHkDNrqTLP9s+ssVAPft3OuJ7M3cvpptwM5k+Bzm3+e/+Lk/9ZV9Qoh46VyQCi04yzWDAiYx/
gL3PBZVu3elNIkg/ogLfuJSTMYHlzWZljDoFdOZP1PyBjAzPNkcT9jOY7BUA2YcVWxLGn5jGpU7J
QVtWpvsOD9WNO2dgXlclrY9thHmnnnriXhp0eYbeVrEo//zTblODMDIc9iy4xDlj6VlXqxml7vO+
Z5AC+a5cmwovFNcaH8m8wqaL57mNIqmnPEDv+2vvIei+K8KgmRoZ5bfy0KpXUieXSLb33HDC4shc
aoVxogS7snZsxtRPR3a/xpa6HdsSTdBrXku2veX8D9oXXi/1O9MJXM6sR4I4B9UQC7BfgyVxE1vs
UZ2RBW03DuOOTrRdrLJjN+uz2uy8aCeU1ufbmi82ZcYJ7RM+tNbEFM0B5x4OV6tdj4dWdwFbM/xa
F1yMMGV5+7Wl3HYNIotPew9HTSJo5SxoS97qJKD6gyTCTGvpvbof+7VAnek7Wz2dW5MPKI0lO65f
6wbMDs7OU36BcCu6Bl0pf+Dup9Y6XRdPfr04HvZjpUFGb2x0x+OmhaWUWtVafEl2Wo/sQdOl3q36
SJbVMwxbqJlfjvE6zPLDiO+Trpn5CTaEpIf8imbfzDKzBzcpuaHn2KdH+UMN7unsI2BTFl+WKSME
f2IRKp3Ng51U2fdVM29NBfl4rxua9Lu86FUAgJYVNEoYyWgxCGvw5ln+1/+ZJqMsmT1Qq7hm+RnU
4S0UdHhFVdxhbKUumqDWLDVw7E1chl8vCRvUOFIyXnjH8c25BkzDIm2n6/g2UsXs0ZnXhvD9qIvC
0WNj/mXlvFs97tbhlm51VatwE9LuLwhkgAsbakivdQEsRbOy0c1cvfYFhB+utRG1ZV6D64FZ9W41
/cTeGUABTKqCEV3s9iGFphLhia20EWJihuky8zTxdTxfsWRqeq8gpGJ3D9my63tDsUUTHv+luDPk
rMQesZySCtCe3WGdTnck4efhayMq8Ntrcxl2kcwkUtWA60kqP15nl3R20cdobHgpbF7Ovu75gGzb
t4YgYWBivlL92PN8PdoELEysQ+5O05AA4xwHtA1dosUTwNZSMKYZvWELT/f7UyyVurZk0vBK6SHC
0tRc9qp0eIMudhzlMscy2779HJiMRyiREnKuiL/QEKtQ9yQ2Hg6f46ViDRrbVhryCLmczC+xrq8C
yiFJjYYsbuHXtHUdTB07YSu7cb5GMZqKEKPxcC+pjMhpRXPIR+hWArNYf7iBMmgqzZaI6fNpbyeC
o+gquujyX23yO6md+C+92UzyNmps9kY8OShLu1uQRjzgY8c8rcX0GKzYwP3QV2GYO5gSKvtnl+0a
IIvxeCsM+8UqTlqQ9a1PhbYEKpLn9AVai/xfd44ARkRWo/XjdStw5KPoml6aw7tbHWLgeCl2uAu3
Xhl/Z7t5AaE5dhxZWedwZA5EfFHuBjqWvrgQspRTrXFFabJlwWGfO5Mb2tUw3EPDDBxJW9+hl9N0
HTee0JpKiRh+v7p05PUU0EJrAF9T35xAvQlqncLzxoe6Be+PxQvd93yfTzMgsm7DoDoVZj+aZGnh
EA8ie5Jiqw5bnyQslrrtcBR9m+Xqo/A7rqSY6vBWi+zW52KmXMmU+vNKl7jqkUlgPLFAfGSnKQj/
0YwbuFLf90A2pxNC0j3Y8YXqO4CUjl/b4PwSXm5wgoGCfDxHBK+9HIPl1974Ywpr5K6U/HsOrUxZ
Is5GD2IKbMtL+kBzdFAhruEluUeIIAcUskUJnPwWA3ursMszsSzro3k2vsPOM5+1i7FxahPjO3M1
e96jPSqQAdjl0rmFP7+NK/UnYbsj0v5nnlNPgflta4/9QpiCu2J4R/WTs83JVkpjzKx93OlwYQXV
HL0U5XD1ZD8An7hY5pVgLK+d01VNMr02AB0EThV5X4teqEAfpwsQlMT7PnqGWOLbmeb+xE8uWIxT
wvWg73Wb9V+jRQJ+WO8rdwkdsvFF2ImoOfjWcuTcWgFcqiqnpW8onO/egubyv1UQf5d13DmQSZk7
3QTFXG5m61jP+feRtyV3K/QohoT+i1HPe3GnYlkEdCrnqAHwFevcQWfWAaEOLA7k0CN34+jnKci1
GDTi2copCcysAqeXfeDl45cz81tFFItiMdPht2MxLbsxSvttLCBgQEwlaG92tESXzqF+J6FdaeLd
+8dZzlgdSp+j+FJFFG1CQB9F0BkXUfqQMnhBgg3+cknDbvvejszQlaCtCju8l0npZuewRAWmbiqU
WiMMSWwJ9C7gfBKbvPZIETS3qa2pbl3j4l10XIbjoCyc6KiqpVPHdqVTyhuRs3KCno+J7wzzRko6
pB8aIaFPFJ+4WaQi6CeQ8wzjdV1X4h6vcOcek6reIw5us7RukFbUow8xj6cMQTpqyMD31BeAKKwf
TWWRUc7A3j1Ln316DT9DRDx4nLzNPkUzqbEBORF59N7XDCVgwQvgV2JsX/KsPUSvEGWPf7fBo0VB
cTLw9vFDmAiT9fZRmZ9/9pCzbl9/Wz1L0/p+jsFbdF7D2Al17ZDqAR1hf6sTI8TgdLj/ZxyBzNoJ
xwxgq1In1taa3T9JLz7JuArzAGJ4gToirvRkqz18MhUXdEZVx3mwcsckjQ1026emTrX/4iI751NX
xmkaXvsim/Cp8RborERybIIShxrovhSA3z/MAkGUMLOa4coJcpRNOOZo6mGulNZQdsnF5DY/r/f0
WriUtVY/LZzPDaDzJ0VYDZi6HZYuw3+4SApih06aISZJIeAOHrEJvdC0ZI+TWaD4rDt602yaWoeb
io3liE2z6J4/MnWk2YlpLstuEc8p3iK9MkWPcZ3ff+JqVDnKIjtAuSz5PNJNm4RjAKeq/wQ1DatP
mH5058/mnVrXLwsPNmKOifwoAMTlzOXRRow/3EjEwiqhwgzgTQyZV4Bs8D/9UMjeS1tZwAA2R6Dw
TX5RpGUmHdkoqay8Vfy8HfZvyvFSGMcqddEY31wGbTPMcVtSOWFbjhq2UopJvP3mge2NMq69Q4bf
OSWzq4e7N3HPpUH4xnMIY/tJYJmNAerJlvzmTD15Q05xVjCa9WvUF6IgEDriTqwcgP8wfQkv1uio
dGxXFKBMTANgqXX4Sghp9sLXNMa/p8sDKXAZQHoBbCc4rLnP0nOFg1eyGEH/8WUfbeygUxQfn8Wb
Kz/KBQnmSkCUWTv1i0XCFprGKrn+Vrx91BQjfnFlrfOnqPoUGuzFp7LdYfjCQVyAfFkPx7+YrO5c
qbn2QmyHXmh0TS+vG71tix715czSvsvtZ35v3VJ/SrnOIwZVwsvpuQamNGgZZsjS1pCqidjN8odI
bHFtRzykvsU0eHbBDNV243vWLiUPbrysvBaUxVeLUggLGr6IJWp1JI5Z48p7Cdga1iCOFXtABIRQ
K0ZdeN1ic6z3nHICFBgtBlAnC1zM6YipgpMmxSn7GGj0M7TKdF3MzVNtSPGHjB5EOqokLr7r4sH0
x0WGDwViu2J1TWthretCPf1RCkuINgfWCNZp42MFqoW9H8TzuCq04BUFt5SnVMzXkj4CGXVmgXx7
62M0f+xV1vSO2cPrP+FElBjwPrarADpLy/kesZhQQH5DTvQzS7mtGm+0dErOInHjM9oZM5XszNkm
hw26mYytbvfLl3raT1MFX8iniI9O19XEa+P+xPdWABAnzn18oAWzEZQPA4FXGhnQq4G1lt8n8Mff
g6WUPAh1QoJ0FH2D9yKE3IK0iAG47G+uDKjM2czYbKn+chetSuiQ1VYpHpiSAZsJSIxdlmk4aS4E
LUuwEiwdshi0ebGkUQ43oypyMkEOfAZr/SYjYpWrl/wrfoDiJAaFQVaa+Xm+yOfVgoDorEaGErng
7ug74fSqVkus/i+7eGSio57X64TfR++PNyR1ncfk5L4FLHspjUO7p1DUzmepyfN5kEJcNCWwQGxi
90NAo+puvQMsxL3a7HhrNH7Q4fNeCioQMDVUgtoZPGu3jYdBrKZauSUNEW8/HiTmRTLnN8WGnFgk
1F8C1jzexRg6cQVc0aYAQ/37ch2Nh2A5rEhXk3iFVlU+hZ+R0q+pLmSlDWWmxPUfkceLRkGn2NPz
hXBFiHJKUcU1ISGyoGShERL5nt3My15X1h4eEsbJOT2jITOsgZg9H2tA/pjDsN8qKAwuJ2LBjHG8
uHwCTCAxMTMaiB0GCNPyuczxjGpH+JQJwyXL2macJ3eC/IeNrzMf/SF3GGSfGxOnn2uqwyqXtbkd
r2srqK41n9rpTSPdLO+UZZdM5NWBqAD7GXd1gg7Fuq9WaKf/qaABBT9zQ81qNHq5jWcgUhy/De9O
4DGhH2gkS1qzoye37apbmUCS1Xdm8+6Sx8jh82xg/2i7ZeYk2EqY+01E3VJJDIJMSMErC6poL0zT
OzYkiH3sVg1kpWGTalCm44umG4he1nolFUiErMnbF37MpATOwxCGNa1760ZDVsVMRl8DZM820qWv
MOle8XfBbL79lCyLgUJnDOqI3RMvCrVSMWrg7md7pYbz8bjHgcjCBbFwDB5MBG/1CN1FuZLl61E2
QqWtPCN8Km6OZTREOd/4AjX+V17eSmiEbBCKG9B9DjchylEA6upTnjmyDq/ubbB/uvzJn928KKPj
wJFkgN1kRJCmCx63T+2yDMNzcIUfrOXVtd0/ZgVgkQFHBIInvbJTHLfmn6/n6Z84LlnbX+KkUnnn
23EIt2oek9ELy1PWIqTP9AiD/u5bfRhItoXUH25DhzXbASpdNzXjzVEphzhFCpfGyR+lkOcvDyKf
SNlRw53yApy/9PTmx8ijcZ83UtQqkltehuUZgrlNqkQ1C62Vji2cHgSTnhPalSQCrde9QrL60zZo
X8HfjZ+FlFh2QDebuctc4sefBqenOF6Ouh755EQ5lH28rAhcMtF4EMYg3ZHsJJpIJldNRh+Ivdxk
acMbLlGc8wd8C3VclECgGnGEcN+94mRNdbKOVBV8lHVOCWdGAlZ5BYAKyvUdsH2BW7rUWEWlmdyw
YF8FbvADhYazgcfsM6QgdXrUDYCVCdvXTyjpEbSXIi40KAt0/ZSb55J6OA09iwEPobCSlFpg3hJ7
xn/wWPO6Qu63PNEBYX4Zd18+SSwQESK1sQOEZOzBrzOUx8oD9Hg7x2yuPrpiJemdrG+tySqKARRY
/O3rLII9bP4uZif5jvJv6BIZtU6D9bz3H9ftZ3iNIdyZWQvxTxbBjazE5+U7Y1arJgbZLgZ3p3Jo
oGjoBBShTBnHkR7ODRWlrFhqbJ5Vpbb3VgM6supc57rqbSynSK8ADv3YM6eryC7g2EjYZcTOzPvW
4NR/AzfmGfX0nfwNhNPQ+DiSow/+6KLL18SDEqIUH4zuNBL7D9GZDEHyNuF7sJkgTye7ZiTiU2rU
9mWSbqonaI/z28eq6CJLDEzAXuhumNBcNTG3tQKxDysga3UDoumzLCknhF6NUJiHt9ZtIV6p2KDx
2ZEGSaUObwju8IB7KbvsLYub+fQL4MTeJTXbY/jG96QQJKlqzr8URz8upj948iak1dsfsgvodSJM
73H81yNxhDJFXq9qJcHH7jabzyB70Ll8BfAXY4AralBDaNPt7qUAUd04gxRnL2t15nhOm/JuaYQq
Gq0phqtDJnApazqAF9x7U9OIwVMX2XUEsKk7XSeWXlgvpNgEdYX47MIWimv+YcIlJ09EmFozmSWn
Zus7MjD6S7BSTsBj/ADOwdmKLi01M/2k1UH6MJRiH2Z3DQwSBIQhz8HWAdTT9eC7ys3KjBUHPD7o
/ck0HLo7t/6xG3hvXxUneIxrUsg8YggISJSrmXNCOmILQL/kSOSaQEVGZGwwyX6Z00XOhTA5wy3X
fZzU9eph80h6ETJAeXkl01Jh3pcHEEn7PA23F756QWrH93f9s90TvmGvY6/FBUZ0eA2ESTBGzBIZ
UytsbMfNU+umpjU9bYJ628xI/3vm9kEte6AuijwBh86/bU4Can+c4auIs8R1RlTYeUJX3c+DbIjN
JKM06vX4/PgpCHvkLQbAdKRaYyr2PzWamIGm8naurZTitE03jjBVgEP9G5HRETwRGVME+OH/SAkc
cTGjny78ftBe2xftWJIzTVrchz5Vos23fTzcmOY+2LiJS42Q9VydMAYtiJcsIHZzLmUVlPwtPf6J
0Eoj7HQJeANV3NkupjiehiONlGRU/LyB0G7cuHDGuopmr789o8racjP2JA9yQomEePlXBS+FnKkm
dhrWCP0NlWaAGuexeUyX/3GtxpWveMg+oajV63uqitOih1aZYzG06HMCa0p/xJuP0fjQsTlNONCI
Tcvjpk6JsmYK2V60s9qrR9nekhfHKp0Rad9tJv0F2WGKk/OdREeKQChugtR829VND1ssCqTjgxiv
QKfHBFxlAKHF0Z0oMP8/gYOwkDU+HohXzc3xwYVIWWzTLd5z9cf3nGnJFYynKSlIlJRdHRynB/7s
WtgSiRMOPFTrNU615BOu/FU/bRlBenWkfSW9erQlDjq1h98hzXHVABzG6K7weh9Wy6KTeU48XHCg
wSmsAx8ynfy8RRatrtEmBPpzF5B/65jtoHF5OrdcDRny5gm5vGXZTgIYqPI2u+G/SjTgCQyjLEBT
iJmJwQQwAWCkyotcWs38xXCUbMtu+k8CY2V0XkZDPM6me565Y0ovNjduntwuhG1yjMC4UlGvFOnk
vgbiRCur0AgL8xjYpImV2eE4O5En6EXJEy/MUEND3OlzDApwmJ/r6Z7Z4esogDFG1eWIzsmxjiod
dl6yxT/ir8li4N51KZ0SqsIKAk3DsLZv6I0/CiDSjVQ61bFXFQJAmLLfwt9BDEdoY2/Kfau6TdYh
I7LXQM/L2hiIcWfEFyPq5QQNxGTBtALESkPNcsa8H8FYOFmnQp+kGqKdoeVQrKqvAAGtomISVqa2
ZJOfRpjRqZuI0FewkYKHLUocoYNO970wS9NVMCOVvGGtRRwdKSCfctiF1AhDkJczPG/RGUhjQCtf
lJOjjtPAkjZ+FDUw5I5uf67ltsG33yoLmLt9N3eJUIpheDoMua3PLvGN3nDx+NtTDRp3b7AYIyBj
iBeH41gp6kz4BzRffE1kOX0cnkgev8u21+qa5VZzazdIK85RkxJY4zToZOj6hVl4hs3xZ91fTZRj
XcGcfMqJmd2HeemJfplqo1I7pxFAsA59RGabePKRhsZDp+KxZo6oM020wEVHt8+aRZYTMAstSlBs
jdhmo12Lu4821b0Z/7A7hmPo1uYD2RUwh07RMIWNKC2Bsd/70JQYAqHOaHthVvmrtvULyBYI0uP1
JwYinFf2FF6N4Q0VOLCP0YT9sRgAOf6/821KwCJR8VnxylkdUbUAnp+870MTO3a0vphidpeQR8hB
qZiCJ/0O3QRsEJJwcKr+3QqZcynAk0DSfMvQ0+fV3d+gI8SPEnP1mW7hA9ZTCdxUoLbAzdM1Nzpg
fhzPfp73veNuhV9JZGi6xKHwC3+pgRooD0YwDs05ZQIae9O8EJJcBQFKu0CUq3Us0w8k1PZZu5d2
yV5odWkI8cHiLYtX0kaLUHqCjWc2MUzXNAa9q0oUUvyUUl53371mxrMrthxtkAmY+BV6T2RXBdUx
Fq6V8dH3iwuGagpGJ3RlSW3xsKJnIr43l/yWFl9G8XErByhFQ2gGjQaLzvkC3E0UMlylp7X3RzvH
bY87V7Bweofy7j3359I/bUCbSgSIMteflLOJMfGj3rUdHl7IqAP/P4v2AdNZDWrd126O+igXMYVm
qY5capZvrPvyPm5XMea/REnLhRqgzdt1LEGDaHPws1jIxC1q7vWR0eqwK9VvqOk7VmDhCYFqDq/C
gYqvmbxFFkVzO+JTJAC2+BSiK+wIr2+S0CK/aQ8kKKbizctqdLPDIL8bBnT8s1Su5JC64SpndGly
0PP3QG2ChWbQgKPjQ6qqNUzhI8ZPn0gqXn5FtHhkiwUw0Qmj/ItyO6CN0S23P1QITEEv2cP0LuKI
JXwkxVBpDOQVyPMg7xAMzIucghkhvJ6Logl8P/elIRzL/92mvl3NZ+5NCSudbJwAfSqN10BjzEYc
0oRCNrotuVd3VofbcDtMm2obV0GuTzQahu8AYRkmyEfvt8l/Xxw4easjgq8jXNq7kzBukVf8puC+
YJFTLX+eTVbQf74ai9eJC+F4bgva0U4dvHKxFLLpgnS8cylhl6LBoKqyZBOyqctH5/Aa2f6GUyyH
6ZsxkTzAeR8BKsR5GAWnvPiEUwlR4EMyL4C+lYMyfVh8/QZWp9yeYE26pGT3/VzmR3LmKuAFGFjG
7UQWMYKOK/YzKE5L5oT9eaTgGyB18ChBw62VCKkG/ysZsTlD2rpExZ9EBA0foB04928nQYZwQrPG
36r2fT2mSS4pnHG2sUFFKVdgIu0seibjwPnSu4B8g33hqpHLl8UW5wK2jN+36GFpCCh7dGU09v0Q
YNqjqJq7P/nS80ExQRnws8CvOiNUXVJX2WwdWII0Kfl3yHJwHDSAhnBOBoQHQzyFUIyWlzfh5dga
CsibkCrsJNqZ6H2FBe1PQZhBH6SnGRaDbKGW7plMAXPjvc1Fc0o4wz/Q3xkjoKf5KVS+4fdHYeZ5
yLDK+KToQirMRddqcYEhRHeK2eYaDvzmienlEL/1GlOKqcmJ3dDr7XEAdJFXnCYhBxoCQ/nWfzr9
5F24D+iTIGCf6ynL5dDy517y6zpP1xM2M3QaUiU98YOTPS4OOgxH7MdNAC1nJcklcKGpBvTJXIek
wNRsbAL4r2HjLN/zBctaKPxfjXUWQo5vMLCXUYqWpCT7dDBX9lHat/MXMQK7Lxhjvqc+pBa7NcT8
KqB822ut14T7+gOHZTrekQgdPuPRJyZPPgXDrq+i9q6MPc9TE6YYBMfpFfyuxHlw5GmVdKh4LYI7
acmNSzgQrcoMKDVUkxZH6i/wuQKNys4jK9Km+9Wwm/fmDHjA/Y1Y3ElqVrH6yQeaMjg8QxfupXfe
x+nKkMjL/i8E6yoDR6D04nJ1/0KEZbJS9yyaVgcEhKH8Kxqx8icsw67QAspXh40Dbiq02AIRBeFy
NGwGRalZ+4BLG1pi3RnlMp2lsc3BKATVnAstg3AM6abV8WrlpGPPmGzhGaNSO7/9YroHS/Bh+RLZ
LZKpS/1yR5cpBZW/KHyvXxWNnUmvx0nrpfkJ4mU3mCEntFlcwgqWdvOFlg1In2Ge3ZmwNTaFOeQU
AXGXWfYHKGW42/RQLQj09kxsMdXcnJ+OrqbpIS1aPym166xLVV33Vb6y9DyfDe6oozWBQdTYJCIX
aKfmRUOD3cScA6fdEXSNibFtusNliXYr1SXD7bd7gqLQypyiiQN9i1PLS0yqoAPobzkRBl251Zu1
3AgCTAXJToKnYziYihGL1MUkbulAM9XiDs+ZZBfZ+a81/cGaawY3vyb22k8T2IJXBrep/q8Dlsd6
QdzD1MRdJDFsKlFoV+nLzPXCaNXoDRfFEvU0exmpJsSGV391evFqXiNKTWP0ckXKdKUTNMwVgFj2
YH3uSYN0/rxVbsO8mPtJ1eXV8KlTn+4Axbq4HqmWFXPc9lCEjmhc5qYLERWk92U5x0n07eMAqtko
IO22gAN+L1WOP7HzlQ72B+qcCM4JpaITKZZQtBMwRlNIRljTs36nIMFZr5e/ev6ugQDDO9IW70y2
9ZX4LIcmYsvGXD2xywm7iLSkmZRDUHXe+RrrexUP5vTO1d70BrwAHm1wAz4CxatfVndHpKS6P6F5
Ml4iaZP43KRQBhhUKVlGdNtRvpSg/iAJ/UNOBUcRAuUysER3ZhgeiW6LxrATniTxJ28HoegbfAzC
P+O9/RGRojDuzViPb3QkgTP63KqUsoftDq/paH70BOtH8Pktx27jC2O1+/Yly86zltdIdtVj+dbF
pFUbG6q0l8lgnCQrVhjfIu0nXfbnWscpxOvGiAH01LMzXGOvY0hxoEEyyZH8iEQY2sDRzxC51A8H
OAy9ZMrYpodcjLCNGcfznBkFzNWN9NnglNC47Y29ZG1VbdqlaEXcM4kWjM+HDvoVPBBClXSMZa7U
MCUaVPnVl5TeSWON1y5pcxsKSloFaWEkuB1kswGKl9Sp0TMs2xvlHWHy+p4qhZFK2hj7R52/1Qn9
kgttgqFkXbFE4bZA40ZAu6LbBe8EwQGKUP+Jm8W8hZ4dsaS9976v8C/MzwBVKHtEEYU1uCqw0tR/
uDyKSelirum0964FHrOrzxXFTCeN/f3n4r3Z+NMOdL5fgU6pDVT+ACzkx0Y80atG9TOKm6lNL8O+
qMM2+b+EY3uUST1TMLGnpwzOo8qs9Q1wNstswauSnEYRwNu+cvMhMzKzscY/WBOocmONmFNCoIQP
D5K0T4Jq/eFkWufLJHSvaCeikdtDa7WCQ8EHcbbj4VOpQZTJPhnlGVRkYlL+w/Ni8zLfj95yxkzS
ebz5XqtOAihesWcopSgC5A6c6BIk09QoZ2RLN+uGip1N+YO3y3Cohjals87/QfAipx0eJ3HQmuNn
yo3dZqhe3n6sg5QzdZwRHrOujDB1tsVsTKYrl1jBj4m/8vhrolIqD1V/GMzdOrbztfOjXNBLGb6X
/XLxnDKMvlVsy4ERns4FU88lfyIz36CCHqodwCPrJsfpxQVUqRb9010Yk9Bd+qeVSM5zJPgqOMZP
d1iPkJTxAPmrtS70wuUv4oBC9+PWYlm6OtM0jPr7lX4uokjMi8qccjGFcOP/3gBkbDxFdcYOG9O7
eWAilXklHraPCZvOyfxnSMDynH9S+ZiHnOI5aTgqmfSit6yigYRP76xCbthALh3LM12cCUPXZSbk
9x372J8EIgAnx/SHCUjp+fzD9zpujyvVr2fqMCKFpVs4MnohDSEaBobeSoICue77ekLD88QVhdTz
ezfib8QQpQVb/+UWTWj38elUFRktnuvua2l71VVGEB60kFzH7SAuneCGKnorM22u+if+eLoq+32t
8IOn0TDd70uApvgUYZDeAsm9fKXkoQU8lwnDmnC1SczJLKZy2IC6H1fud5cNK6cufdNWWZ36aiUx
cG+6DKoAPSyyfgo2DhgbpfA94CN9TP1qIsMwgFgnfAebQshzNEUNvLM819ibapWcnLnl6JNpEapa
RyAnJRSbhgqSAu9wF/nLDbHsdj3kM7aF0wGnDymiSSsf5RCt/OqGWxBKMQmEZkU621H0Z1g8UeEw
rfO7MmYR6OKNs7P34N59YiNBczpebSRW1Ht0aRjEEKGFXmEOuxHitPA5I7Be8N/gmT4p6lsFgv/E
ze4lAct0Xa7q1XDiSrhYmw+zkrUtnDOJ4TFD384EMHjYWz9uxxh10y0Wdw90coyxw4r6qUiehJui
zumkUu+U041W4rrG3m+wt3XjgBEtzTNf4lu4o1r5hHcDryO8pA1znGFMQnbzaHQmY0FMWTUtN/Le
1WEEP82L7MSZQegd1tN3TjUjIkzNqgERzKk1CWIKJl+b/7p5lZAts7t+wYAA9f5RrK+IcEkKPClO
QvHWXWs/KIqPEZmuVUpatck9lmfVjxY9zlcvEuYvSYPbRsVjGDipCc7LSg5FjBTbUkMFLpuh5zAJ
l5ivRjc1RM4dCh6fEx47/38JnlCsrWmKAVXLwL27rbNpGmBvev9zOw+GospSe4vuYkO9SGt/KlhV
uYVdVgjKr3wLChj2MMXGn9DmOr8LBFgxbWHQ2w3gi03Ka8SjJauBM33p6HZs/8UupPf6Zy4hmKyx
/33XMtMNQJOT9PZqLLV6ZG4h5u+5GJyp77zR/6wfr30EqWs3jA6SbuqDtJktasprg6xDmTsfI01U
UKTh858zEhK5zHE1I55ycqB8Zh8/C6sEGEG5X7/FHZVWWeiiqPmcIBsgEp/infX8goJDRpXl4ZzI
GgN8pxvnOSk4YSN1rrmuB0v3z+PVCT7TfXJD9hTgdTGBNur92vckLsd4aD4177OopxFUm6X0jFJU
y6rZ8Bw/YWgPh9pth4gmQtBWDpwP/+bx75AhcDLLD29O7L6zw/B2o1EPNDFUdEDMHP7Sg6HHYI+H
7x+RQ39IajDb/JLS0RKFjIuFN+Fa6YQbzh8oGM/N/kNGWN6j4YYbg+5FBnbnet9gZt332Qf+QWJU
dhDiXFFbc3LqqB5eEgeKPNN4vPcp3y9+08yU3/gcyxVMGrtLC7s2XoXvK29PbRg/t3APdGy8P8Gv
pPj70gqCCb+4dIE/qYolEuUJl4ey6Ksw9uQpjKWk8FB+LHvSMou/bPlpoQhAv0baCczuIq+etQz0
EkVQDaav8Dd1uyHjgvhqzK7MbFSfc/nYLSlMciBHnTGdujWwz3LKozVDK1nNt1wHLJhOOtQT83hy
4YBnkXCtrXHIENtAR184hYQMvK6hVg4ShaO8mZ/SiXSV0MMEQkBKX3A6bUlHPHIgIggAHR3PkrCw
VTKikW9ZvBFKkcATerKIeaLACEAx0VWDfXUrfzKQOE/dk5NifM3mzhiZ/hecS5OXS0BpWaJFA2u9
kt+fHOHHx18TnbzzgPlaVIJC6g2KuBAZ2bJ4Mumdodk5KpZUhgVpwQl7hzXYtb6oADK9tOj2fOk/
2Q5JJWkaZtf6oVratgtFhw9rhpVYBnjtrPD3YHq0uo1M3y0c5p0mV/WCinso+HnLlwtrKxwx8Yic
tjpZmdmMagr58OfCdMqWSqCuaQJUnQ1NVH9NLGiA9DNtM85VgCBhNF1fXO0rpKD7TXIP8ji3ENSX
Y41CYhEzrUVATXdpyeneXyHhM0CHHxvYtF8dd+W19v+f/F71C7PYP0jUIggM1rjjjKP+z+x52dMd
/LivhqCmv4WK7TpE+hn8WH1x01S9prp+OqisLj5S1cVGTSZpQ05+iGEGttRmy8Pek7KseSs+022g
srUPpmWWH8Xv+dFY5o6SwQw4Bk+fxcnmdfIJtiEvX58PdFv3hqH0Brl/EqToBZUE/yGIwESp39/+
+PRmWGd+/Fd5g3sOKldSvwC4bH1zU1l++5KsdSXF+kvXszh+Q7VKDn2DgkUQ8Iv3qvesoBodS0Cw
xmJYTdLscKt6mKXITGzj9bO9xVl7mUjSzHSljcZd3YL8RyI02khsnYd5DxmjCCxbhRXqgjoZQv6E
CROtF3qH4z0NCEZhhR0wCD35nRlqsSrv/XOwD0AMqBNNGbP3hH8DF+RJ2ZmnGTuySEVcrxQ7b+Lh
65+gINETxZGW/F4WdwWKFNygCfjR/R62iov4tcqq8gdSN5sdbrlxuM3mAsmHWjvfP1AO+yjx0tof
iqmDquNG7d57KTRY8BBgupRE/pVUFlhW7XxqCPF9GIWbJ0XCSi88UGCe0UZs7EdLMo5a7XivMP4h
gHveKdRa9f0mt+1DaLdKT1YhovNXUQ0Y8zz29wIu4dk+eijkmxADSSfZJnEncMseRO2e4YIchZot
sCo9HbJFEY46AnynH+BCOB6O3qHi0nVdPlwfLYJ8J5GEMh8LFEKs8xDRreYpzNJZXcgckMPlqYhb
wpBe7dgIgFLu3G1O0Eha44ZwpEsvY0IHxHCbtlWdktr+rpT+jfBeq00ONUSA3hHJ8/acjCGZkkdZ
mcvj/BL81QDG1IxncnBJzS6NECzhgs5UTf4pVz1STXEWoNmIqY1ezvngwIHtnSerC88Oz6wRY5aK
nwwMPOSM0PwLxwCVqS6xy0JFScHbj8ImNu/FygXvzoh8uX5Y5DhtEbFU8LrczddP0AA4yTFm8Rog
xr4OGQvdiuQW4NEaJcikfiwKNtVs+aYuyItgeA8zxi4Qi/b8CjT0H9Iy45qtVruaElOfLTThc5CN
Tni6Go4uKAvztXRyASC0bpWnt3bPo7xT9o7TlOP7yBD94UnJEKbQHw3lcKo5SFv/0hYiaCuaT6pW
2NVK0yArmqeH1XD9vpQ9/5GTwo/Z9lYdKuXURm3MX0IrdAkoCwk2hwm8RU+GwK4TSRidc4xk3LE1
B6VOnONgVW1KqzY4O3bA1SlfzninRIFPwTt1N3j/TQx+OZmTJa6bSGYXreaX8Er/ODIz2hGy+yZH
axFjupH2fG9p7ozTelsvrKuTYCUUI3GJunKcOjPIphixBRoGUdV10joMEA19/xpCV3eSiBY3q8BL
mc0xhc/j/mK5i3ywDz/mnCpdaJK0yWHaWRFUpoeZNIWEdIFuiWH+dsK8simMB6brWjLyLWF2IR2G
RQC41Hh1ZVlf9BnbgS0nOjLfIXcWouyx/UWAMirLlftp6Dz6VU/0ZDuXQInVi8UAiV41YxA91VGY
Bh9LUFkqQihLIZ7dVAdz5z9EdjRV/ByeTwO5eT0eSYKjZeC143ooEgWjMCPyvoppo2bkoqyHcPt8
asBbsEhVBYG3ScctRhfoEFQcc+k21efkfKyQed5rHw6DLaAl346584x2cVVO0U6IsDgmL/C9hM6G
9kvQn7FQrgBj2ZWez+rumvKwr5Sx4A0JVtXpA93MyrsYaIpQVnX7UpFLNhOyermbjD12Pke2qoVY
wbBWwKERkRIdbPIFHMC4KGBYh5YhQI+bDA9iNWB4ClbDCvrMowmwD9JFtUW94gQTVHxZPVbrO0Oc
adkVk+JITN4e4J1B9wzIY/ryXpKbsigfwawZr9UmxUA9g7SudA4Zj9IxaUu4QJ6Zb7rNPIIJFoPy
W3dxHHmuNhdkIFlFpo+AdI50oEAQsEmIhZQ+KBCV/H1qVk9YojYuw8s446qw5CQ/eT96fyInvEw4
p8HNKhgYeAP7zRGzyN9P/mTVXMukD7EimGlDoBhMfrAD2hZ1LvMtRNIS+WrYo2HnZeH7El+50XPQ
sxswWuj2IGWW/YXeafjVsIGl7dUCOTRl0LBgQqjl0u4XAVJebg91cfvc5QCnkf+I/E24YG/wodaM
yR6rlBvzRyEJGZVp16PbVk4uF7jzsRO2DCHU9pXqprlXVNGGdZ20BF8AxMkpQFs/0cVKvEL16ip8
SlGf0vBtuse4r/JLeTCHMWrhEczpREu8lmWxW1FrCfVaGo5MnTIPEcdClu9Zx+o23muuULW+TkxE
Zdx5jV2ONeJkhC9bUpYTfYMi0rquST5LJF8J93mBzoP6UO3SzyC3GvA33zczD2Qg6zfnTgOi1Csy
gkgNncfWwDx/G1ITyu+u/ImMfwm/cQlgd1PRYqYta71godgJbaxJiJ+4uq4ft6PjO2Ib81k/Gb4t
+Hu80vj4hyeW7+EyyladsufHBv5O7bq6IiSwcX6p8XzhSEI3Z7vCRGuDyJAYXKD8PYp5AIJdJRL8
dXgW72YwZCyjsahQG9LEmVjicS5QCFJhyclqX364WDu9wkz3P8rlVAGKSFDl6odWi1mvI8SDTl8I
T0SNp4PW/RULuBqTSc++Kwm6Bs5iFTUhGsGptQqIwPFOXB3PCDfKNwZ3ZVyUgyoqPXnmbVin6Vo7
YynqVj+rZfYlDb6o1vC55OM/9Y+gEEL0zzlAl3Vn1SDmMCU04R7Q78elY5EVSK3XOWO6lU2WXaBV
dgzDlYaszvWM2DWF801y1vX9TIme6Sy8rN9c9oYfCUYse8W2PEgnGooZSlaUczZc8vqjGM6prSeq
9pHqnMFqasfvdBRSA7UxM3Q+YhZnwbBiXGYAhZPqMYFJZ526bWcFGI346IWmmm+0FSlOUQPIxikk
3/gH0SPcZBr3oMqmQfdn0N1qCRjb1ivhxdDJ7mS5xPosiCIFCwWXc5KdFJjbVQ4uQxPYJahbWsBH
nUtFQJzzUmBE89IYnkEYNzEJGrg8+i4f4r+s/9xuA5eayZgGdIOZM3BKtPPDKAEMS9REaPYNnIOJ
DsSFtwi4RiKM9VLoC9EspQ1CggPjIPIUMDikGLR6nMnQKJla8tNotJhd7BXw7zwGOidtGnUg15Dk
LvZN7e/sV+xNxnfQaSK8zoMiYs12/Ve93hQA5C3lliFG0SMaoI26RgxibpA9f4ypji6BOTotuhAV
hRJZDH+YvIIDVHfgK/O9KtCw++5IHeN1YhfE7AFW46bfqwZnRNgrzrGQV3zPvpxx5NVUU/7N7oPZ
UZ9Oqm4Hrxb9s1df7TsiCXNBsZsYPbfJZ6wQXRTz5unUbvYL8X3NzfZ22OQ9dX4t3ipLH/IL2olz
FWaDGXWYr3VQnyJyIIGsIWP4RKHoD8hWF4msbcu+p9vVa36cb7LZJkCGTY66BEPEdPM8ugvDdEct
dSoYPz3D1P/R8QAZfpUKP8Shv18Qvt74w9gxTW1jJkbIHdIflJE0PvPlpyUKXpNLLPfbqvQ7aKQr
jUcuAidL/QWCxNceMygiNcRHS5Pb7D31+RJp9pPW6GL+jRpcPq/9fmYlGDe9EMk1GZq+WlIlatxV
7vRINgzQDNMFel8OMiU3qQAkeJ7rfmnMegCK2TiS1PZfXC5uE9UbJGWUTPc1yd75RCCaaGniRPWR
Lu+marek3Bv5icT1j/CUyw78o3DfplLCIiEcIxQjjuEq0xOuMgQoqZ8a3iyMmILW6TBtMcy9tfSq
cDVtbM9LmMuKFj0GjCEpnEZkIBbFU3k4A/swPDJ0FvpPZyNJC4QM1twlNwMrpu2Jg/3u0r4sWio5
CGAgYyfQ1dk/8/IasapLZD4pC98WbS+KsEtUVYiSmJIxTuZNK8WOpWtQwY0IrKU19hgf5BAGMdt5
gesCQupYIXBCqyTLDIBAKpTedv2M1i4mOSe4DIiDA72mXwNMJHqeyWYpf8CsNxV6+uzgjkrdH86v
wonz52vZOA113LeTZ4ucCeE1ztBrTqRcAJDs48UNf0ANcYH/sBs4iH1qDWTvgmxytSFLtpaGG2dG
PALFV9h7gu7XJk46T566dL2dcmWY7aXERG3Nz+g7Ez6DaujV5Kn/HBVBRNSTqfonhhCXQYQPrpes
f43UeCu2adab2mhjdgTtu9zsYNx1fF4sVl4qZxYbGNE/+XUEJVTBnwo8EN1ukHWapd7xKYhA66cr
43Teu2C/F++21AW5ByHaYr707aS77L55K4m1i9T52Wch9Wu8uBL+bNXD+CRHXgs5E8actXx80SiE
vZ55wHMIm0Uqp1rvk9RCd8Rh4j3xm5iRo2efRye5R/zCRIkAnucrCp2RsMCZ7tktYkJO2GXwd32A
4RtByaLsBW9Sc+KIiJx5ZgzSoO4obHToFoRUDU8A2xiXeu7PL292fYYvIF4y0avuJK3vyFpVw0DC
sWB1s+yjjk1zg+1zoklBuqvX9E2F88ZW1mZjstvVfOWNbHjSBw795VsSmm+SBejkntMSlF6Ic7iY
MHZJexCmEb6Geku9d8fIUOiIZmFlsyvFvT1Vt4MyO08IE7qbQFc3eXVrw7gYGAKEMrbtqh8PkU/v
opYq4hhfHqQS1hln7a4gYxeiV6S3Q7lEklwrdciijb6bLtKfWa4B7JJpUYnQ0LXJXhBENev/idlM
uqw/t9EM8MpGP+gPbItx0gkv1LiH5Qtp/BcVnfYRnGaDBAHeBnWJ5lItm6VstKo5SSzHV2oeOkvx
C8rsVAYg+Po6We3RckLS7oKSrDL/KwIiwQtn05nf1RE5Q3AksLqZnRuT97bV3lWYJZe4vlldfmQz
tsJaS3klW9/dVlNZqvyyTJyIbw4RW4uqmte5wCkvxVaIut5jZwIMFmOi9ZXxpBhhGLtsCIc5K8Gm
n19PXQ10el+HSM2SKu9j0HDiGg8Q1adF23TFVWsOlQuUcqvcNuDvCKblE7QJrd6QQs8Jdm60eZjF
lPGZ56D8qQSen7neQ8Vz96Ilk8Yiidegl9rYBjaZhaxBnKAIiXEofwCCPJzbB5EqXA209a3t9v0k
vqIEKlI1cs3uf27hwL1mttZQcOJmroe6cCRHyO7qMT+lW6N3cXQrsHJnA2hW9bDP+MecUSZD6o0v
Mf3D5J3FcKod7lA2xte2/G0vVHomN2akFtdlqwMV6rORAY9nfY72g2PrESxYN4dTG+oS666q7+sG
FKp+brB9hrngEsunJjstxYSdR6vPsmKobnAL/sn8pAqimzWmsmMWqaZNXq+Y27qgdgVNvbcgHwYD
inj0dHe+5cMKbSPZVlv6aB+lBVDb1R2c9Ko0o9u4cvBmocA3cgj3RnglftbbHa6vOLQxaVR6Ifj9
NyqqgJy+GvKidIExJ8o6JzJr22MgTrZjjUrJPyCdSaO3W/pJTNgJKHoNM2SgeloSNpDfAe4WCWHx
H2xUVcOpy83Dllfz6TZqai1z+BdCo8qId7nNtRCT3ZXQQj3Ov7gyuV6oc1cSHvrVOR4AxXLLVI6b
a3EulJuWvOa7lEC/kqlWwRylJzSH6uxkcQcUn75O/gL/NbP3GHmLumWqOLHn7AJUR8ScVsjTjXaQ
VVFUqmQfRufbPhcIEAGEOJdKTtEW/rXPJfyvSQMTtzOhVXlwTnyBh0x+ZcD3XY933RwnkOQgJnBB
/77LhyFMMSXO3Ab/0uc3TnW+nvIPK/9tweBoQSB2K2fL9Kx1O7z4GQ4j4bSw9jyH24RaQN6K3o8w
ai0OvafrGD9s9VXWWBGNEZ23fWRk/nmXK/gv2BeSCXRHH4XHCyO3Xt1zdmMwhHNbJ6T5Aoe6dtcc
SXPwHj9n58pGM/0yqq2IhZ9s8ojOI2ISlcpGO1WAEcQeLb5TAIiDzO6U+gHKGn6CEQIvnQot0Wlp
vY8VVNsSIVPOkoJ5lleLlWCqIAOt95mQYi2dgpMPPVMM3iq8pjCx3ALG+xWCbBGv6wh8aP1hHS8J
RuwPIXrweOZiaKx4fsZWaJYaA49dZ8t7EsVaGPZ9SHJ6a4c2YyjJwLS8vnH+MvqF51lyKpQyJOXd
G0D3RqWvW9cGYEakvoBe/vnBUE0+PKfZuZJWJKe82FkKFFLQb83LAaJwPsf6toL1Rrxq+M6Cb6bf
H/1LQKsZ1mRI+gpvMMLmHePvTDRGl9kTwLP9Tg+ZImK01zR/jXvB/feCT6EOdA+Vw6GEUNYoavD1
V59woY1DIbAJEJ9a4tzjvEYFxYd8VEbgTCLJBseikV3Txfs4hlnGStIUIh8eH4gVN6gEdrAegJsx
1yYTUvSJYeR/yiFIn8/fmBsCQcz9a17hzxIFSkDUms2Zi5SpiAiRtjD66PLRifdWF8kavL7vczsP
xJECoZWvfk1q1Y9h48a12BzoXnw4//BGUAGKeRu0zOp7mFObVpa+KoAG0v36pNUv/ywTbYz1viDZ
NFVJUJKH7HXyPKLi75u07YN3X1LxNYkRJHVP8+Rzj23NyomC2lmjjg/OUPFPSdrc27xnQRMqcdHH
Y04hviT8s4uanCvLeB6Za8NvJNWXHTBVOR6iGgDYHO/fLHHRCV1etuMZ/1YK6dr2emd/TzNjmFxD
Ei4mD1QsgU9nyubYC1jq+RBOsNsNXbAODiVCEbc9kg7cmbhlomOJjAJKf8Gozo5x9FE8B3GuVzPS
JMgWX0LIhIRKUeALzRDMgJtOnpd4tzaoyb7hwfTzlIduDRTQAK96r5r9UMWXe+rZG2VvXJKcQgNC
yIXEKqnZp9Etqx5cmDgGorVwVHE9ArvFSHJQ9O2HWBMnEjnpxr8r7CwKcdU4eNLso1hitoiBVS1F
/XTOeXLPjCljMuhHYGKzmPcc7ibHjJizOsQqqUAC4U7LMFqeCzrtEuLUeKpwYI11OR7mnndc0ReH
Jaje9DgWk8UM7dxeD0QIeLwbchW2mQ8a3psb7Z/RJ5LJ/EjVuVmrVzdhN3kA38zoEURRaAmJsmnD
E7rLICjveE586apbDde2Qd2ONTt7xGRn1XvK5I209ndwZt0Osz4SocFeLjJfoG/lWR9fJ1CTY7wM
zeMgNV1oYboNcuSDhkfNdQn8PXj+ef02PeYf+Gjx/8AJD3KTnFYbrFAamnfWyiWDvaBdxLmsLwWi
J2SWZ6kUcXerN3Tf5Mzoqba8GRSsUhMlPxAVMkiqQHW3a3vUvxvBVmObG82awg4dmM3L2zxTzAph
rZOTRxAbyo2zNq4E1GSc9zaSv8Lf9XZZpuvqGl0jtyhwZiC8TxaPpYLTBxYWDUVHy+eJpgC0ZEQD
WD4kJ9wvF8YEQFOX5jVg8rhPrYf2vOez5dQev4L+rmL//h6CrebOZ6UPqUjkZEI3j2d9WXpZvFBX
kAZAlSPanSij7Dw0vVKaaoTJdefi0/G8h/Urdgaa6/FvaZYvKeHDMKgG3QVhOpH9GgAzSk0XpzCg
0cB3HtQfox6kCgplNEfPgOSQVJg1KPQwSErPiLYoSOyORv40n5D+SDJYvEZCAB1aDS7V7yIBqWPX
gpZdGo03G4Pv2MMNqm6ECeFflTi6t0245EXgxCLYC8FPXEfG1BdhPlfjYXyUS+rYqn3lLKBC4F0e
zk7wBS1QBRc7wgtSP9HoXLa2NUNBc9xv5X/Dsob9f2CNtahdFpr47RxUgOURb6K3JvgGqEgU7cun
9JppPgdgnNSKFH5BH/XNT6W6HClnSJhwaFbasFD1garY50JWS3clvM+2oxVdQsE34ofUpQR/7hBT
Vu6Oha6LGmzv5Xcb7bVgL9/UzI137rrLA9ldbDHL7geJt2SvUij8dHSLGATO1fZn+Np+5JqcSioG
OmckXkFwctFKScAWlmKNyKhB1LwZuFBcmthvOMfAo+fYRovT2xw1oMQhIH1v/c/Grj9HQkonCJTb
nJ6wBck89FGk6ibFzV7iLn8Bhl4P5h1XrBxZEGT22xVK3O+LapzJeJUiRqCkVOzHex9pvbGBMqA8
kRMdA+WkLQ1oTGp4Zi5cmh83+fsj5hGL6BspQnIyQ+2FXmQ6axHZB6f1ne/1yOfcJwsgGtqauwWs
ROSWjjib+zqqbXTWCiHO+MMC4g+WtjAMhgfXKUDc7qLczcnLqIf7jWivJrETbfRIn/o/keocRNrN
dt3vsRNDb8hpyBP00PP8Pk4JcgxGY8WOgEkFYD+lnslj0Akb04bjlmO7XRu7gMbvSs/v5/icYrJm
BEHF7ddmLj6onpEKJ1wt0zVpw0DFy4Gqxqqhejsnp5sK3pjw6zPvGIBCqSp/iIopKcdgMTy53CTq
A1W2/oDVaL6r8mqL1GzH5sSq5JveWYEvw2J05atsO34Qat+kfIGr0r61KROxMX17B29lZrqAlyel
XCHFUJ0eiZumY67i3Wy6EQpMxuERt+6KDXx9wTlBle1SLIMB0/Je5raHmnixuFxOj5ErW+UDw8nj
J8nNNwa8p9QdehVjd4EmNn7bayOQY0+6lHuzkgg15hUg4bOf32b1anHHGYOi7I4RrVut7rmufdfT
f7Yq7UwS314U/RWWib4WhrdiaCwuqNQlpYAfWWw7W+VEQRz5nHG3v6OqSbe/3Ax1cfScl0EmFsxK
PrwngGvecFw4Tv7png9+VL6EJB0Bgp0C4szs8zxnLRXx0Jb2argOiomJSgNGS0sL7JR4GZa86VPL
Pfl2Jp0tqNCoyA9vtX13CxvRcbP2qBGVRJFIYHDJkSU/Gr/H1E6zVTbAwDY09HN6yarL9yULc1/O
1fPV4rxbKeEJUpjKS1NDVPYN6V/1qdqFvmqGkjMd2j5T9YLXBT708DG9N9jwLkrrFokDXPZZhckR
xpZKqs6rXgklgiXTm7zQPlbtykKhUfpLlvNfGx50W1iX4ZSbgP02018ljDyZSszrUcmEUAfXuiJV
2ziL5mmniUaRRFfiqP7s4QU45ExEBHS/G9Mmqj5b1m/9qi4H5eWh+WZt7/LPyY4mKPuReto8dG/y
EdUaTjhZTmHP5KLdU65nEVZ/NDYk5B1TSqzqeVdA4ojVEGgTe0YcQ+LQJvQ56FxvLSH/4auSdZYz
7B/7A+8vOTngKhNdjOsdoMInADDUYdMtKF0ehImGX1vhLX0TC8Y6sYJwueJ5b7tA0x4K8mOdzC0H
MfM0g55wkylWeygwkN+qT4o3asQ0uIqa4hh5LvQCiObcbdTs0z37ZRHUIXL5GEjdcxLJR2pHdMc4
hojdHgfVT30X4HmNQp+vLFI/c7u9GbrG00/4wkJmaQY78azpSh3NUM2G+DsUtkyiD7xWrdQrS70M
/cV1rBVgjaZ+PIu6AJf/7SG8jO/4CgumuUIM5C5fS61JaDMFcGfYQM3LUHa+Padq0CHB6Au3nCLu
u67fnleRGyuNEFmC338j9yQpbiqs5SxxyD5QyByLPkeST7rINY8mySp8Px6n5I7h+LQt6LlhzTpL
k0j1tcFU13ojTtOoyUrHhAT1FpHL/6UQ2Ohhr/UEFARmr5UJL1m1p2wyxaFJP9L8tFQl08tzlY19
JcrjEW3WTATHaiQe2N2D5wDby+B2G4ncPmpcEaxyeg8yhMxBnnR4ER58nb7eCvwq9YPkphWjGYfR
rbbKId2b1xwc3d1qJrXaqvs9fJ1p6pzH8dWhsNp/zTEkbSJnvmR6GsQKjEDvgEy+vGHYbe2hjtcl
bv0T2JSODT83h1whLKiVFJQwMQU57vaki6pe2HurN6WuAS9udD8zsFxnL6JHKOljX8rm2mjcFgk+
Lai535QmH+ymRRjVtwfjLHZPHnQBHpFVqDYD54rzxhka5L4s2HrCi9LLUlZZkgmZ0Ph2SD4ArFDH
aV5Mm2ivA5S9CPWrS5MAth3qvHU+UEFujBBKhJsnq1AS2E8vywKvrof8jh9AWfYudS25eDMSHuDS
ZiPUovPaTJizapfE+1Hj0oNyjbVoc6etkM3zyxyDvolM75aX8DmYqBh74xJicj4Lgyuxwt36nGkR
BDicHbJcrbmKINTQ5pOjazVtpBS+4Am1EBQ9PJk18+8Eh4tUB83IKTzlSPf4iKR/B9UgujyYOwaJ
fSe7PAFe9fhS5+Ttu/BD6ZU7ldXOMJ5e9oVsiHPAdHZ7AX91Xfo/XsguB0CLztcsp1S60vj9Rw0M
KMMpwMORRAcCR7f1xBZu2x5WCjpPOFhhBavMDwFNCsFYqUfy+OBs3LRmEvn+RSFDUxY84OQdxAgx
qNf6FXR9XqK8N65EMuX+Rn/e0yP+p536Qqbrk0WWwfkMCNmJ5KVFwf2p93cDvjX2ZVeAVS+RgltR
QbFkFMEyJ2BhumOcCIbpnZxdnP/c4qGYPaCGlV7wBw4Fa3JXVkgn9jMFnTcc5Q7qr8DkUHJDd6pa
RuwP1CYhFfNhJHdgCyLeXewlx/rYrRYtJseLFM/Lu8H/ENstjVXAVEFbe6S4K0Q/WsIwFrGIJOVl
OKqeLtPgNZKAasa6Blnq5N0x6IchOwioJ8NjMUo4SiCA7YKZRa1+IHt6VOJUUBPuh2UrMFIwCjcg
+tvLGNAk9hNr1GfRNCukJKhW0ykPvtZ1WntxX/3alQGzxrnIkYpEtTP9iP+Py3Jlpzj38QqRdF7C
1LwGyUeoBvarOOdlxqBtUwHVQ5HylCtmRup9wZCuhw0fymL1laNuY7rt1TO6q1zNGyA4am47xoFT
vIHVG7IKAiM34BXrBGq/WL9SkbILvZhiSvf6g/2/VAAcvfPJriTgT2E7SGrMxCSK0XEJJSEzWglD
8Kh/nK9F6Qwm5KCOKBqFl8HS1+Ah5EgsbeCuO7hWIO4g8VsupkwNmZPmNZjJCSlNf080eek5yiq4
4nyuugiyX0g945gxJkUaqWIZ6j7zan5Zw1XxsKCqdDBcaHIzISxv5BbOcqSr+FtgiyfdR9TZ2Kp6
TvnyRGYrD1f7cWmXydaO7wMLAH7KVWF5w4FBoJ4K5lmJhjriZIxOqzRQWDYGcVF5Nj9aI8/B/YHv
czCyX3dFUsp6cLOvXh2Q57MTXAPGfqtvFkQ30d5bkHL+cq7wdxPvPTjycJWjGQ3rGOSRr/m5/jBF
crcA7jxl0kHN39A3HISKErjhRVgQ+WImcdyxQEG+8z2iffUowPSXpBfbKQdE+PNouXP7ucE+U6+D
H139g3EdVuV8I9TdG21JRSAaet81q8OD8y/ZhIj+tgeFfny8BhF62Cab+ANmjyqaESSDBUGtjnwV
NTUAe9FSCZMpCmu68AwXF0jx1rFaHS0uU8cIBLHF1Ex4tqwDv0sK+lhMuvDo5QT9/KGvkJPCu0vl
/vk+1h4jYsw4hlHmZJtPLdThZGX2w0VFGlxNS3uo0OhlBxs8jnV10EGKNKbINaPGXkWa3Y5Wc4st
SwMzKcQ09HvnPtl6wV21duT1wJ7WdJxYiQl3fMNpbDUPV44N7yCu0o2JXPdduxRHbHFZHrFz7qoa
mIYIp0Qir3OKLvzb4AxZxpiyyGoh6DL0y+re5h928iXDnTMJW9JhutTi6CnGJqi+KjeQstwz/RGA
aAqxRnWhpwU8+uRmIbcgE1T+Nrt2vXA1GHNsbbg7ErlIdQj+HkBJMkeEIew0K5PMzBTj2yfwEuFc
61VCydx/GsTqCo2LaEKdtZFwiSZlF5mNCCPtkI+wwmZXAz8flb08VE5mTr5BA1zPTOanNJVnSosl
nG6WCKdNHCkpkvvO0qh7RQiOo/QzFvaF43UKS03z9nsG1it8eaLGrLJDtq+o9taGopioPWPSA0Vu
zHnpgHaAeokcvnJMhawcjQlgF6zQXhXAi9dA/YUEljiNK/46eonmG6r+o2KLyEYWTCAPI9R8L+mo
P+CW6ajNMt5EWKxdy1dvoR0By7AAODfEta793U+0fGstpv/JFOSfGnlPQJYgH+U5W2W/RsUxWZLf
vGcsdXzjbzLECwJ5Kh7Bv+8UBp0gqC185mUnzSP2XEy+iwXWokuGGy3ZvUGODBRveAFFPFTxeDG8
uj+alJaHjAyKa6oUGMiN6AWIT2wwEC571ciYVfm3JMpaiSApTOhUBQufbW0TWsrTf2PWwVRILht1
ouSKKJsLe58Nl/ubSlMCCDxmQJWaG7/W1TeVaVTtrdHSQYZS6gn0wTkTuVMnq4t92etToNzu4ogU
h2ub3YcSJ7650r35cK7/tXrXt9sXqNhdeRa+u+K/huLJxmkkrYMOPyVTSjqTZuzQmXeX9wiKdue0
FVLQ9kt8rleuu/wC35rnEIp590SmtTKmuvf5qFguPZMWPDT8kZCJv6Aawn2qdbNcFGSNeMPCJOmz
NQldNvoxsUxVKWR0yRMwO9c5KBrEg74FPQ7iPgRlX8IytvC8zBhEaOpHCCTpGwwn2IxXz8o4JHqD
PQg7Qe/ovT4pJeD2OMMxg1T5fSBWJQym1EtB4b4vdlir8vbcqY9WmmvGizmoVF4FELhooILWbv1S
n5kdjGUa5wwatBmWO52PgSljMADEiAtWJ6mu4Z19OtgOq9EP9dP6cinsbKbalRm7Ji8KaiOC3+rg
y/p/PX9VUwOTPafZPRgwOTJzHvHETHRJH1rSMXsujQCyUhYu3/2g36P8kLgDnI8ln5XAvuBE8Amm
Rt0oQYVKs35FokPPjRz3dgvD5Q5wTz4V/IeolQkvMh9Cr6umPLPUEHT+qv1WqkWmsGgn6Yz5lZrP
KLJWhFeUlCCORvHeNYEHt31SClLPOWRhom3HtCD8lyB779m0RGSTSGMnFNGskkbRrKCZ3PQA1nIL
zpb44LY7cxjFyrA0TyHyhn3eBneTAG0bQDda5St7OJOqsJ/fY+0Cy2c6xBFaKeQJ7700W2YO+LJ+
QzXbQ/LipOLz/2zEP8m4o7PBpJU889PUb3XtisPUGxRZWsGnMF1ZoPuMZmsY7AmbnPHfShXlMTaW
5GQOHdAxZImwaDBDKc+PEq36nrZ3ymDy+7PqcllZtnGv36RvGnV3hBxLnpXd1O6BUY7p6/eafOOI
7IftApgyA8snvDqgxFgLfeB2kO56AoAMr2o/KiquH7PUYLjRZxUP5931Vg6CO9wyEbHVi9Tf5w8w
g71vVv95yvVpGv11t2E1BMfAsO6GU1KoAgQ4E9kaGuIsvSYGYeaYDXMEfSOrV8ydgKhE7SstXqpN
Cemu4c7Ee0NWgceSA3NMRf5ncNAl731Yz43GjAy5YAcYrJG5MGwAAmJdAzvZZ2HF3guIkFBYWVqa
LbazG987CzgRv01Nq+dIf4tfgDL7peZMMId71E60gVECFgXePprXn5+3AcIFC9QKfkVbj+N3uTXg
z2yohl+9Ja3qJWpAnk6sgfg1sQRC2DljPC9uL2ivy4TcwEV16rJ8jqTZoBn4q7aT/3sbjNGO4R9j
lKQW62yNxky268kztP29VOdcHRI+t2bbx+b3BmtgBQdHhQtbsvzCMj1ZrmKVTgLukGZt9kUkrKeW
MbtMKnmXG8XSJCOrbVAlYekPhB6aqx//P4u91LAWEHrJg1uiTb5Aho7R1RCUac5mHbx76WVKVOsD
etdPnerSj1wftE4R+UrTKK8bepTzEAnwNWs0WeFrjb7D4qz2kfJ7cHy5h4QJvpTujcI9Yu7fdl6a
U2imLRtXitpGFRIQYHVx12Wd57lmJSoJvNSJjgH4xgykgnT0GpgL9HSOPcsSYiROMMabIOGrU3X3
VKKcjqL7f1jA7LTub5bpEclc2MmZ9ZJAfaAWtSTesgAFs/l+cWcBDLq1geMBzM//KdkNmJqDsVWV
pI1nxscW+GPJbiKwxD9uQCyRaqTNLuMcAjvXJa9qVAtjcu8QP2p4yQ7o1ffRbnZD6MGh9eX9mK+l
2uqFXlrUsL+11p9w4nw4bDNR8uoTxvRJ3hu8AdfbNwhePA3GACVfW0S8nxaFNWBTVxxv/8BT/Jq5
b1xHIa1ZCNliLZZT35Itun2MwmoHtXQtLFa5yHv78NwtjV5WQGdchqHEGDuMbRn2bfOM1Jv691eg
yH2OLJ5za8TVU71zENhj7rdhpUAPwGeMA9mZvCfGURB62up3FbMuhwMcQleuFtAYRFMbCFodjwrq
2t3rKWBR3l25GZV9CmcmWSaJBG7U6Uxw+e2qjL3fyF/F2IbTrxh0Db1Jj0sM2Gy5rY0Rr0ONG+73
sS4w3D+e1LomBMFDpBBE3WCpeBhSxyWzR9Od4TYjmeQu9FWzdxRvtpj3182powtXXmZrWT9EdvdL
GeVYM4b4B8F3K4/cQDJrOZdLjcS5lpuIArR7GP9Ob6YZdoQhv41FGGFvJWr61el8mAA2UwVlsSnS
3ghzYoq3Cm2/cGA8KJLCh+g5XHSKWoYs+9kA2FyLoUunobcgAycXpdxqxQ9lSjzTmVdnMJq+5qOW
sHufa1xIY+x0YHYqm+o2L+bqxnsBVfaZ2a+EcOOSN5xDuTHXo4pmERGPFaQpwY//FB4nhizZ/pOS
sj+XuBZPP0OZ68hk7nf0lS4FQTn2eSl6tf6LMMD2mGaqLJpwe60pfBK205snv2nRftDlAKafmmy7
L9kC+oZRz83urBla5TrowSU+e6CDf5Q5xI2/AwWUBWT504PjZplRciE+1zK4dQa5R0mzHkkwBVNT
quSPxY//OXEXTDpXASJt/Er1oGfCwgHfsCOCkC6qWCmFm3Q0vi92yVhMCJSNhkiZcfr7FbV1XIm4
qFlFKcWkNv8bIbSDumJqEHHvLP5TcAD7V/1tRWSiZR7oHqFQe8pyCdBKWvbrPa/at2KNP+xN9+sX
eM1Tji8aAJKOLt8luI2kBgvhjLkGroCKu0tssSXOipH278hn7JzytUFkPPSE4W4eIMQ/ApbkyNog
vmFhBWSKcfJRNPp/r1wm07ToZ5Ahncuax99rY7DJQc7z3LiWAQtzB3yJtcsAxhMrplZ99HCApGXI
PtZqF/KWO/Jzd9SsS6AIFE2CYrA+EAFjffolevBhxidY9233foscw2ZmsNfuGXdaTT2z9aVBD5W3
uwWySQi7SG9YHlTaaU81qd2xz+3DadnmyWGTDlv+ytM28PQFfvWh+dozDdQ5jpPePKiynaAdw64N
Lwc0HMI5etZqr1MYSNTymW3im4lI8OKe40HeklMkMoUGVaDpz41f3lpNF7KscMAN9/ik1n8Lh0dq
+cQqsr5A6C+0oVDk/N48X2KABHEbaYc4bfb1u8RO+QHYsMQbeVS5Ef65yEkpdAKqfp80kynRORuS
VFAayMf6eox/eQBOkEXTN9VMWO6+1jPzurDmizQIDZD7k7YRJLLJFO6IzZFb/sB+DqxST+sODWIV
KuAFRwCnQnZwX9H7Y7W0I5F96pERSl1lSotIMDWpsNnxuWJsnsB5ex0e/6MB3iyuBPAfDVwJgA6/
1M0TbLvwhJgbmQKFkI+q8ZLUr5rzy+90y69Z+IX04cP+iSa9ArdVfIDR6LMYOZnQiEpTarSJnisV
1arY6yokQE3EhAYMDJFluwdbFfZiVNYwJgCTPEaMcLnVCikAUtwETjbi7Jf2MstPdWAGbpEmv877
rI3sXE+2CQMAFMTu+zthkxzqgN/ehM8MvmkhbUiAdIPEaDRRq0vRO12zsyO2bKYvrfFzLn0W4+ku
IkvP/Un+QuufO7l269M3OeKHZN9TTCH3LUY5S2xtSjGcn+7/NR+BdJ8WhvOLDD8CmYtWYYhPqHzm
IZjATeYpF4dKfLo2vL2LGxG42oGZgcxgdGuTHzdnTjVZyT+vJltbXfzTExYaugUxDMGejoxBx84g
VqStAjwAj5KnyLJ7dpsw0KVIICZtC2nRuF96W5I+/zcZ519W8cwlnMdFfXPKgossVDqa6cUKvSC2
FN2/WgGy3fPkeY+BQzUS3ZpUfhx8HK2k77C16SI8rRfPo5ia2I3fnM3Tu1o1QuY+7I83StwcehEN
ihXPv+0fhpWF03vPnmUTGraNUMn6C/ubbzi83dLB5TcsKB+tMW2XxjyNJXjtbTczCBAjLdrDNYa3
3EHkPJcWr2smdrlSjXkW9SDNQAngX1I+CL9hMI5AnroxmzWQECgDCWH6C/Gf504cIXqumH38cimz
x8QsBgX6qBWJtgS8ijvMOddO0g5aggBjNZk/ps5Sbk1gZhY/jrpprwqMJ1u02xt/UAEtw0W3TVHl
5cho5JVzCClVIq03LKy3cWGtxktQtu7XNWBq2PVXGNxOnkjXC4qx+1KYPCBzOTxyZS+MJdCiD8YE
nn0ebLeDMSbX8nkIv6ij9hjfio7Sk2qxOWDILycwqZ9PMyHRgoBvs6PJ0xHu4lJfW2EvTNUDiHE1
0FV2mI96BsTWLw3udxza7MIJWvNe3WOO6kYubAee0ahWo5Zjq0xoyrka/IH+KRZsYEUEJszHaEtn
yKpwxbIVhYeG1/zqvqrT/xlt1lxCpt2OozuDTuJPz7vWbZqQ9Cp/qF9czBtVsi3uqpwZ7ie+T05A
iwohJrwb/2wUKhq4UyL2vSE183RFsB2izVtATN8rpikziSrUjPRCl6mivmJUNqI1xnW4JUEpn4om
s+Ea5+aFOYwXUECUroWX0vEFZEDkf6uyQoWgPb/KVCUNquKoUgXsPGSsZBpGfaqgzAncaPQ4+PaG
oiBr52MhiDf8IJQuQ5FWa5zY1wD6Bvj+m/Ad44+azMVFyE3N9J03hldzdLuV4Tqe46kwGgrIKK2X
jSuoC4SrOz/aux6akvIL9PZsxQbXM6JzkLDQmGdt4Q4nsmjomE/EvP1l6579yElKBBKSuqyCNHOy
hoenpYNib70EyKzwHMwVVhYB3wgJPR8kBJwm64onf1mTTZ+z4MPuvLZBRCkBZqI1pb21yTyrURxA
/XYDTk6suTMf1K+sxXE8vf1H6HpZjZnvzYier05ccTNCeExceKUvfJPk1WQcd9lTX29eFaSMaG53
PvPgeAWNyvE7J/DgfAyb52KQMKTMuj/Nsi2jagyfx8M/N12gfmrXo1BaBzF1h3+5y/hnRZ1TMAF/
V6H3j+qxvZ2/qmvrm+YGjaCXp8QPiYLoGY/dUrFICN9bC9Jkt3vBhyL0vb3szSTPo53Cwaz+Uaut
DYdYmP8hiw9V3BZCYzj8A4RAznb+804JKPGE5GcoxBycIEtI1BA2l2TOnCx+TgYQgrysspDJjlKx
kO8WX+zLAFJQGn7+znqMJcezIDThLQz9VO7lLhLvwlAR+XgEf64T/8+cMprh2ZxmpKC+UgKaPCcB
h+6+5hbzk3KEcjZ9gI8S3PC3zJp1iOSMxMYX0gRpk85uVskP/dNW2MhaRt5qfkGI2yHnrUXonigZ
jmFNmhk6t0Bdwkzfq604wjocLOJ4qxFAE3YnJn8rXjfWbzV2/hi8noJmhvcN7Y1xlmQvTS54Wvyb
nF47MBDxbg9FrVg4+cQUNYmDPIH1c73igGi4gbYQQiJg3McMGDiSUAq3H8VXjfL3I1EhgsGXYM2+
Trm4McqHm2SJ4vZK4IilMsmUvqp1o1ksFo/hHQ/st5/CyiyN31nLNU2PhKHjSqpnANLNJg/emuBJ
onQwti3Ub+dhuEsYIMj1VocyrXsiMgJDqCGDNhosP9AC2H+e0e9XMgqqFAckkJGEei/D+pp5kJkD
uzQbJz/yLExFBt6SxvEsyp+IiNmaDVQXRK6dnaRkYQsoRPOUPLZwVMx9VWzpZgw/yIjXwETupCN4
cphniAlRqndXWTC3l3A60lL9uxeoPXY3Vea1FsGSFpumr8flGgUyAtu0IhPYYPSRIGnaGKJVq6Ng
LQSpPoTxERhif6ZCK5Q8hEvSvTgE0fA7wRN5zER9tn944QykTVman15fcd9wdT6fq1//S3oDaH53
xQIf2IqHnNf+pXXVPkAoUgQUX6tGGMAsvYpi1rIkTEOKXBikhnS8Q+0cR5OKyaC2s20sFN3czO0b
G8rLzkiwgXYc+SohWrR26w1gbaSsM+NMQYnbe+wYL8wDftLqsjnhW/FmlGpP7H33TwOGWKSSf8FY
XL51K81z6sXlkAnDJPg85fJkosttSIkXHaJ90Ak1/fZLoGmJpMe/rXdrrgR0zK+fb4UE/BYOMG3c
V/3TOreDI4sQ716cVAqxatmVu58AkgkuBB2f35apz6CnWOoe2Rij9mtBQVaMPRBaIzU5vqBUqK8r
TFhinW2TylBpHYlTiwo+dhybdSTJGjZmzxah6yFWXkFsAk4yD61qdqyjtJiHX3q+Px5x4M6NTTUZ
nZGMYZpnkbQAL3Vsz6AhA/r0UGTdFeuh9E2PM3bJbSd/9NH0dfzmDBDc3wBJKbFBWEYsE2zKM0gy
z3+OFfj3j8IwQkBG4W51WsGA+meRxJVZ58IORpj8uuSh/D+7Vye1tqBcmzQuku8kd4Xx73z9BWH/
SuDbSrMcHWqJiapn7IQGrYRGJ0cX5N1uctX0wncd9E1f+VBymCeuAPAUqSfcdKUY/jXnVWj9iw+h
iomasanR02ZeczeOX9grtxetnektcXwvUveY6zaIHEGBnvcjJYBKo+1V8wtyIeS6fd5j0klCJmEc
lG6/soc8dtGwuyhzatu22lCk2DqlzYkDZttOVZSL4hHfDFaY4Fn+nvF6jSF8IonQ3MTW1S4WjtL3
04f0TIFDzHum6CVv4rF0L1M3jTo8KcqzDI7eCUb1tUFCFPRexikW7wPUT2+XQCbf0Bo7sRx36jdk
MykGFp/ntq5MQgmU12H3HKNS146I7E0Mj2BsW6ie+mZdLFAzEfa4oXB0doJS10U0nxjIAGTUfZgo
i3NWIBXEQacU7XdkxgRhgTFbNQFGTwr6Jhh8y4rm/iEgxbPlXT5pJDu4fpi2CrjsgepkrcGqBP0H
fM+BFk3nBZrgzOczALNRv3bjNZ/QnlLvj2TDIa1Qq6oy4ZR+6cYIzeF20MhphtVlT3ZhuKf7zViy
lMTz9xhUDCFZi9b8n9RMfPhm1tQZtMh3cqEmVFFcQmvtTVA1eYFLSSyy/zvEBFkIyxPrB1lgZZbl
acJwi0ubaH+UkseQnpxzj7VxE5qrhRvxfCJBHiQOnglC4O41qDdACXsZgUkdA2paBGMnLubOQ1lv
h2cD4iAO8QVW+0ch21mRL9mp7sfq0Ob1vrVvXkESQ4UtVZiBSDqncdVH1vUlgJHskbHDjMVsgY1o
Tmfo4Se0coIe1PkJcyqbo/Yc1D5F7tioJAHr9jmvCbJGB2zVjRC5aLdmx94CDZG+dZMdiuQNQXSB
fvHR9VXePqlcIREL8l9rmIpBVwIE2xn5klgy2OYDHrpNppuoSWjYIupWTkiyAcjqb58FkCN/6ZaR
Eqm2NpEqInddqdNd2VDNNcd8V1u9zSTWD9nA5e0DsZyk6nQl+D4zyFO0PoIq1yV2oYHXNpm6zorc
jt0mXH4JU+3Lc//5SlLea410OCu4xlqr2FMiKjb0xfnWhOT/UpRvR1SoMEugO3jWfuQuYw0Fjx5u
EtAdq3RA/s6EOhnFfLzVlA9sOd69Z680jfOTywz/Ka6CMriUrHLzogSTMn12/UG9FBzqjN9tPcdK
Bx4+03w6+iI5rke4EAXon53dHOUkbt3Oj2Lw+hgUZYYeAv0m6mtcL18aHLUOrsZxlc5ElUJwRPAU
A6MaK+v+dDV4taK5RIWaI5lGtTyhq9W+X8xufBOeX6GxJX71mQmXejE6kLphqywu7T2dXTCKNHpn
icoVywdE8Io9Vgi30MDx0thFqBhfaDuFUTWKyXNHPJnQNtnVc6QmIyue8tLbWYIgBPHJioCaiPhF
x8ydIw7dldagpDnyex1rsJ0YOQJjocP+hJmha9NKSxU8w4chPd8Z72jllJSTM604VlR3QqBv9fOp
sLUo82zZ3H7ScwzB9Wh8hESnYh3Dxw/pymhDRSP4Ccj2DjKnDDUzVZHCwDnnyPZ3byNaHdg5i1Rn
w3DuVclASFX0G3R1+CN9lPEmvxj87vcr95Pe8ZnXLiyM1KWK2eKb7dqcypeOBn4pNuPfJN1n9EdJ
nUUGJnMp5BiJeY+O2Mg8lgVFayhICNa6PGZoCiQ+ULoMiPb4mNsW1/CZgwP2iwXRGm44WW/p0Ars
PlmmWBzrMTrfpI25B+0k9CrH4p4F29F0cBfWmyjIRr2EDk3R+vNJF4zDn9Zzd1o9EIR596TL/El/
hwRGuvHiL7S8iyFToKgyuTlk8h3Qs4mcGGJcJj+MtsoKfdQPbw9nyoYwDW9MPzNs72skoC5kUPKp
fwqVURzYepTQEiGZ15vGX/2DP0G+1Eq6LBJP7f8xlIHHo2XfGfCroxmIQ9UZoAEgHvusJxlBIAT8
Ar5xgx84fjG+0p+JMZdcjFp4TyrHqlEzCISqhLeL7RPH+XitvzsCQI+EDC2Qh829jqNBOM7+rJBD
XwGk8EIFMSG4tKLJU7EkB/Ex6rT+xcp4AjuHCpDOWrCkReq169axi2Lmd+M65mxRcTqjjtNzTJSp
HsMQSRUcj7ejBZkY9QONnrt/FWmLdk3TPClkEtEK2cHV3KklHBYP2+ljxkHa1Y83ZtC/sAtArkLG
lMFAK6vFx4SWo4J3iiNHw5pvFzXCTJVSfAQKLm2hRv1mx4DENpgXq3qr3NQQfaCNk1r+dwYib/oz
XuGhAAeUeZZ3GwPB5ImUkVqFy5lLsufeaoibF6Bz/K0I0TpFt+TJypU2k9jrFRpCvM+83VgoJ/Vc
nk8A76RjxQ/SXMd93Tf8y8RX9vxOS5q6p4EYUJyNwREUyD0+Jt3PMs/VSkXheXnpI/lbRN29HxDM
bFhPFHzbaVomU5pkv3kgu5/bCoS3KCZdkBThbbDN9RdZiIFNLutBj1oVxtJNRlPTR51vmRke89wX
hs5bq4O2MFmbulf12l9lLCnyuMXcSZ1sMDfLBBR3Wv6456mCku1zCFlWUlOZwTKjstv+zCb/Fq0h
6TSfXLR2myczEmT6jEXVpBAhosx0P/Ecnki5qKF3jUGkXktq5OI5ag5KUeANDE35cb7ZTAk/1v5V
Cxv4h2MlzLmL3SlxDaQpirjfPOLQXmM36EvGote0fGIX4M87aObbSfOvnuGBffAweMJwIY57zsMb
Y2kX7PfnS/9SQHEDXYATRHChmgGM3res13459mYVXuOhznJjhV+ufr2VhSKBB9ofA9N9m1Pu5nwF
kaP0EnYwOC3hJhTVia7t2h8Ioa9DKMxRzH3xd2y4Yijs8oDE3Ft5E3ZKUblNdMPzmKhzZsL1DLjS
4YNRKNi9omY260gyaezaE9M/mk2hh2NpF2GkkhTRoDSFbprcsVmcA+6v2NLhvPfqmNVUZQtAQvs4
1Z6r502FXqjZVr4LVeOm85R1jVN4nK+pD+7S6YIwFc4qs+Q0cMn5bSE255WmDRFjm0cx09LRgaw2
CoS5QOdLun7DWox1OXZnCHqIlBaTg3UMIlTTo/SG56iCEcfUmm6o9oTNYn0q5htiKEJC5o4VHAS/
zRP9pFz6Egd+bxlCp3wCvTsYaifLinEDBE47RKtNhN1ZezX0xxSBRGo9KOZrlCi/5F3b/QqL3JxJ
3+B5wPOec8Xk2fDxGO2/T/mpriU0UshegH/PSKSLVDU0YodTROl05+z5we5rU8uSMj05Ydp8nCs3
EvS3MyHmUHWu51OHP9guABK1e1K1YcEVelcgcIl+YefhkSYfKueR16HqGSWFh0tqdUkYJv1lHIWZ
D7PZUZRBK1rhyJBViLaZiV/i1r8pPSZQ14jVIuVFaHdJZZFoHjW7T+/66khsAJOEi3D4ujBeWK2E
p5oiNFw493OQ36uvgODnoluqL/9Ey4oM2ViQkluriDA0wnMHKSejxfeL+Dn+DosQ3KZmTKSJntL5
aO2k2OJo9BWLo4NbdGTIs9DPjiYhp3/w2vqizfEkNBnNVZ/wn5F3/qIYChcoJE8ryeNUDY4SK+rh
xBzAvl9B3EUYhku/nn0jjV/XPQEkE7MvrEElNsWvHIfjXv3NIXaFmVNs/89bMkvQc0hc5OL0FZFj
hE+Za5SaYJFRRgKyDZMcij8LV7O7aIfIZ9SXgKSDQhasnYNL8oF/da209kULSEiAefXG5JRVc6O1
QXWs4PPgw3IvBXs7R6qYUhp4Ki7LdFSEQpaS3qEvVEEl86rI4ad1Y80qHQLoXRbtXtd1hXieZpy5
8gxhIBepGSWd5dn5QB/3LY38hd6qye7MiVMABuUotvN1Iv9bruKkJe6ihDmDlBOFcm1fsAGXyxlT
YzDBlngaWpj6FakqYvE1w8oonyghiWwXHsVciXyFZZiYl+h0PDoWK9PhND2UOMckZdmPqoORe5us
Hz+iEGo7GhH9Tm5QwDbDHNSLDYOSaTdygYqxQIf59FTwJsWguzTWmQXtsONVbM8jZO7npp7sSFoS
lUamtiAIUB4PlG3ESMXwswSnGlpU9giNBb5cebZjUVSKcUiGeJjoBfNuMCe7bvAVI4b6PRv2p/Wt
JmVvg+XDkF2Z8QYIhsQKJ3b8SWsMfGdn/LGLdgeuOCyygg7Z7l3CnUrfNNbPyYZ+C/9jnFphsCzG
YftchhR1sOEzrWIr/dpL3UD2U0IEIPmj5T+t7qJU3ZzfJUur7OBW5654jUw5gJ1ZL14qFR+zdHsL
DpBWyI6Kv4eZ0ig6xpJvj6m6L7/SGsdum5Y2kLDfuvdyagQWfGIY7OjVlHHfRDEt9nysAhlF0Rie
TvZJE6/HrwStbf7OaBia7WkQqLWYKgpS0lB21QrH/ezr1zIboAZ0zHj1ufraSjLnyyBDqrKUAXZl
xixW2Z4bsIl4Ol5xA8YleVaoq/yLGmh7rRl0LiwFeTc+PFbZeSwg/r+94Ut3m2EVNtZhBW9dWl9H
+kLIaEx/X1F209Yeo8ifNrG59JW75oZB6Wm0Q9FpDix9wXx06+GBOVPwysA4/grj9RHmo7EEyoKp
YMEQtJFI/Z9uIpOISEFvvljaHqVv6reAduDjMv8NBvygaMAMtqqNizEaZnf57L0jHstO17XPTo+I
oa2547G6uyVoZOfykU6OHjxNuXGPed0QkyYmpT15zrHxa1p0PHe3lGLJ788mTH9hBPoWxK+UOmNV
IOwIXup8/Pf49JkP3nshYhVHAM4lUtm/LmVnS2h6THH7+IIepf4kPuG65L1WoZh1lZD2KibGaUxW
uTRAcE9FGj3jCYxZ8EwbV5wqJLDz7aQpoLS5ROriA5OQdfAIaj4x04FB9bjFyy0h8Wl9bZWpbBgP
kiFeo8c2AnQQjcVIJAYDaxgkcwqG/dOxrBLs04H7fo1dEVJUkwW6pSXp8IvxhUALEGNhjiEdE4Ha
KFFqJWbgd0QFTpdtVOUrjumd6XnhxPnVRmLEXD0c9i8TdW/f/7vesesg97qvGJI4xeGdOMx//OlY
x/zmxtHQ7CdUwLyZ6T71oQ1OmIqFY59aVWpAge3f3By7WsJWeODluLh7X9E+GOEjYTkMuP79BrGZ
iyQsbTMywx6TynSlba0h/cEQxhEUeSwusO11kDrZB1lucrrIhDVy4zvpbLPuqILztZlvLc85+WXl
+IKYzXSPUe9v3g4zFUcAZ5GXb13vjgeyVrbn2hjCPSge8Yskeb9I867KvR2WDanEZ9B6WhdHFKS9
0pTZbCWq2EhtM7XI97Eh/3dFlCXoxkDtYrbps/uWBuITlFjOxv4+w63bDQ9a4mAbQ/fwIv746eA1
YTMxhm1lZkN5f2By6dt4dQacyvD/ZqMnaNC/Jyyq+oI66t+C65p9FiEbs8cQ6tRUOnUv73X6XWY6
xkLYcOly73tRnAjoBQG2fQ0ktiLrI27N9TqIIdYOumDawYeLrc360FgAE0nvrkf77LcW9r0S+31o
lIR8r0E8AECwfzkh2nUsgcmc+eB22+ApM4qmRmENjR/u2Ex2e+r2I5M95/8Y+TsEdFBG3ternt/R
gDwrE0tDLrj29lrwrJYTC7Ke0YyWcAfwqgJejoxcqZbDbBvjdIjozuROj7Ph/D1/sVQnmJnTZCqr
BXWEjKsDeYTePy5kA/W+PMdhQrrWxgNgUfBOcioFrVPjoCcP3ZqkCSSz+jAQ2q1rCZIj7rK1JaI2
AIf+VD5QPXAGFUFmv9qDT9GJSgdXB3VnPStuEEa+6rCfVRreLIbmOQFFZ4Xc+VrqIcT6qgF65Z1l
AmeC30znNtOy77mHgDfEc/w1nk4pi4yQ+JxXSaQloZU0xzsuNJ2u7cY8KkkglWJC7EvDvLMfGdo4
QWyZLESQj6tBwg7RE87RKcg/xTReuPymvm1voWRRMrTxUoiAccJZccKnSiZ828wlK/GSbPvSrxeE
GxeDdKgiI4U/WF8Ccy5CV1zKu8ukP1+PA87vzTyxfNKRjxRch8ze0BEkfiFazQGOBFfZatq/uGju
KnHO0cAJOEVthlopG8sN2sI5cI+BgiyRTzzSsLYwJkrw2TBKK/ksb5tz0xahiIrnZrZrfyx4/A3r
nSDqzbAb820GT3g9OBoLYlSPUYBoeddt7vV/egThuY60giXAqbodXBMgZehS5MCcwruNPHAtGMXl
SVPwhKvVpuMm0br9IRQP+LhDXe0RMu0EsprpsN9g4X0pEcXJ/zDZ95PGeHWHXhSCaEz6jW6ruYfY
saZwCZnNxlKJzOCM8gUTVMrT/Kbn5QnMP3LpvECisisQ3Wexy11ag7GydS3DwegSHClXUFLO4whQ
8BYGYL1+hWNVR/m6z/9FEx3UFutqOwCD1nhb5TBQY22dxOFJoU9/BV57ifCeRpE5Thyk9gof7wq0
siLaXKKrlIeqIlnX54WFEtVPAu/pmaiBq490gYgHzifNDZFThZ3UJCGS6sjN38ueggFVQNKlJxIu
rfAh6J3+HWzJvBLu4mtquhqlXIWyP1/AR4r2zg9oqOMByZq6PM2ObspGxwb6bYoyscct7FhTAydh
Jm9Uh+VmebDckk/SIwNk1t1ZAZ1DnkvekM77cPPiKZduy2Xt9ijseRC2iBJIYsMxXed1XP5CLbFg
Yw8rwagopUXfvZU9A9sBWJ33YuU5zX6hC61hShp5rp4ydDJs0H2OGwUv2/lOW73u5T8AqYn3YpqG
EeWmw9iBT7TWrYEbScPYoaSvp1dk1jwRcD4RsMwA+Sf+yM3PGI4GPfHcIw0Xyhbk99fQPCCXsTUz
yOTv3t9ngkq+2wVqh7UPk8HYBSn65exrP+gPddrtVpb+gbfEy1JywW6nv74f/+8Whpkt9AmGTv31
SZ5EyMGeMDEmr8RXtR7JG8LUTAKkn80Hd7B9fP2/c6BEOnBDKQln2D1+0jkH+zrp1dprP/JbzAmP
MuGhEhkmkHmoSJWK4+XdPMyf0hTYReWj50yTZm/TbrhqXrTW25HvR6aFL8Q/iS0KXZ+sl3fjLsfV
VCweKrHkEs53KX08KNypmU1DOyWf0QWvKp4YCCwI7J1wm1xkaB6AaeoYdNm8t41HzKULstZcd1nU
D7qZVT3JOlMfQw4gJtNLphx1lZB2n0x7Gjy+zqd4yoIqHfg3XQVUEVrmiSwpifInNWRkra27c+JL
N8xebJw1nw0E7fdUtdJX85nIylUiAve7DsbPcm0LCRKWcdZeEhkMGJ2W3ckW8YSxuDa/VoGBXJyS
FGjgPRQF3yXj8+JgoP9T21loKRfYJ5U4C/Bug5QcHH1ybewiLx6Rrd2BHiQZn8eJxjKsYG/RlFdP
MZaHDYi7gPUCH4AkvQrGzCxW8gHU5zdT8nJ3LW+N4AuXEEZITNFEPNOJeZrQg6UL4l5sYcH5Ml4y
Bb/fDj9bJf0eVhehpCM1mbQ54opqhujAEy7EbN38M8VMvqIKPK03zwXLFd85J8Pw7yG6nwKL1rDO
xj0p0MbF3vxN4lh2jcWVluOCoVpffRNWrqNusPqXNnY43oPRPwU9WX+oFJ/jC6WDEtbjQ4jcAcEM
GUfDok9JHlulYw/6c8Z0eMrFUaw73RxLjV6fr+rgWrpK7ysTsfw7R7fPCH9w/UYNLSWxdl9qgoXI
cVI6Wf/EJMt9ul1WcwdFb52m6QY+K7kSUmYIDG/VnB8KTYoO+Nz90LF09tUpBbBC1FyNu2/Cgo7/
Ko9papZshgN+TjTCJkqW0JWdbaiokQv2NnrV5tNhfKFN7uFD35xqIDxu3g1Q2PKQ1sOJPcCE2Yt7
bmXMg/HmEG4Yuc6u2FhAsTcWJE8TufnTzV1/ZtyePSy+cRAUHWWg3lNsmKLmknSdc+KNXYb4vQtK
k7ggfuyUSr/9ly8F572BW+qbcK3LfgkRDUFk/AZrI/BeA0rqaXw85Ef4MkfV/3F0OhDB/2v9iD0q
eMlAs3p1Ugfw7FCUSm5onAa5JHfL5tx1VHQIKXfS8RkShykhRV6bL1np47jFsB8+0i6JArWYsDZd
0b/Qu5YMhT+AMeEGM8Vu1jWcBSt0mnYizAJqeFiCmsu/U1CTsso3Uqc2oSLGIj8RxHMVd1liIUmB
ofVlnQu/CCfG6gEpWIxWB8Dp2rnD69IC+mRkqaiB5LKWZ1BCJ8Sx3liL6nmF5/ob4M4nvWJCoPHF
I7nmphH3eboULqEU3LW9NowLs6U9dMe82KfnTzDTh/Mu91WkaqEIpKOtv0/AgME0/lXoHqBosHgl
EqSe9lxZzxJyUTC8C+CaARnFeHigiq7rd6LqwBQr6Mt4T/EWIgJu00w3EHmNN8zo1sMUwHwkVu3i
OmXdCauUWYGj1MVpUt3xgpdjYY/sKJwNkjch8nXWBTd4A1fMUIkXjk9eCXQgWZXt0m0rClU3zIuz
tWtoPQF0Fw8pAqc9TmIW8ukYhFq2kNwunnZQhyT91Aw0bhhOWl2fJM+QiS5eyxEXwsVWYEAowHCJ
4Dsp6bxYdcLW7m+R3LFCeIkDpouwDUuz9Iq3rKn4WGa+5NOmdFM8GvXmdA5o/1leayuNYiu+id9T
sflzAZHMxAKu6zdAlJywbMvVzcBP0OfeDQuf7VlLZtuDW+hiqSc77PzpY3y1+U97LQeBkaG40JLf
8NIt2raMJVXNtD0L8JxPVxnj0+7xIU09D1DSnu++HJbV7EA15nY/9lUgILv8Xz2noNEI2TAGkziN
EAFeT/k8T/Kdavd4n2rvCHuekTuQv2nyqyBmG1/tx3CjAdGgkGI/WGWTiF+w7SaFQ9ZSBkgeMtUU
QVrLAnw1H/J/NyTaEvHi/uJy1L7eru84GHlw+BC1ndeEv0V6ooy6Pj6zoXdTUKZxeu2z07IUtSJV
z2Bx79xHIRqcGpGoz5J8zDzR5npsqPtVraWJdhfolj0ZLbvQzJbo4ZJ8k4jn/h+loj3uFbOlY2so
901aILkMhN+yjkhR4F8y4l3dATfHB5ja7VJl6lZNUAYeE+Y86QNZ6uBe//EHRzRO8BAmDyTbwRDI
VrwGx5WsZWPdAEm9wsHUwD9lYhOFjkAhWGByb7Gpr7Hbq4mTb8duxjerBOqJ5ojz6MeNeFaN49WP
pKhvWDWpxiBm47+hjiAHSY2QnKuaoR6bMxfdBZ0zHslf3mszOiMhAUjCtrsUUNpmim0nOpxo4qd2
mbL/lWSN7cEpzXWVRzvgMtv0bpQc4CXwCb8OvKxCE930JNRbRthVBi20mxp3H2JefRDbwHdbivdY
SLKKxMrhXfSD+qxZx1FrVGr9E/15muwrK3zrMqCdtjMEAliJC0H+kH1QRaLuRJGG5+E/XMqXGC+p
3iiQB7/40dTea2WnmAYK3DeOWI23eW66uRXVPQi3A+NFeSLHf6n2oJXNL/D0uRME8ajQjQf1afK6
vHddqwDfUQctEQGgHPHLoPq9sjlEBFSTffOGeMtSA6WtXKoqY4TZYo4zR8CEZ+dUi6rcMl2dvc4B
QNcwbyd2rXLnsE/EoZH0gHGkVLFb0LefAKCbKgrBiFguMo1Pe2hZ0wK0IS9Xz+6Ui1k9kLR5HQJX
qMuDJPvOuPmCEAd/Gea3W90+Ux/iY+xjz68Bd+3J5JxsjDPzKibFfhSwhtShQz3Dpjva6SHfCrQs
tTGVNH17HWgDaW6xlLiE12ogRG9JXFo9FjyUihNMKCc7panWIOnaKTqGnFxuG+MFF4SRt6HhzE3W
tiPjxxIBVVPcbikDNM3wjQ63QbESNBE8YDP350gtauCJZBKV879BEqQJQnrnHLYZM4xPRL/CH+wf
FInmedIQ4G/iGMt/URcEWWyfn0HNAAip/dNr5/isy9g0Qu6OH/4Rwyki9/1hwgBANTH2vMNNoXJa
auPofkFING9DrmGYU9Fqki0pF3AoXAkL5Ca0/DQ44/U255eM5nOsSLk+lGDr6tAPmYR2tU2jswVf
HBvLWqESlp5Q/SDIA3ux25tY5e6uAXhirYmLWpUEJszZAS39DTaoipq35UTpdbodbELn4Sv0Zubz
eC9atfm66meyjm2K+jlo1z0gsYyszeV75Qk7xeNcErrCbZ+p9NpYaz2c7HhAoitRk9HwgOR5jeKt
1xH3PsvYKywxU8omQnXp1/rWG7q7mFEqGvL8IQD086bhXs94NnVWDiFZzgs4sNP5V9VnCOdxc70V
0ZzpkG1cTy6OWewQaPYwwna+Weu81lmTYmp0cRzN4G4oXurN8ECOzgVdezmlkAEBbAztph66tyvA
fvo2db2IL/onnzUblR33EzYimwx+TvuMyY32hJL0rrMQfi3wkaC80JwjtJqVy70f2v+4gFIs7D82
/qsgk6gtwZHmkCFlYGYn+22JjPwN36mg8si2EEgmJAEGLSX5OeDsyQOISw3aX9wTSqyMixDxD0db
+ZLiNFFYBI+w402FgLHqv6vsH8UxMUnY4fVVwvHCib51ueuID21Q3WWKKMFspPw7G4xsstlgASQZ
O4pJgQfOZoe/s3wLiQxeIEHgI8W7PufUY4pT44FZGAjOed+a2neiXts3cpY3R7H7AkYcVm1mpSeQ
EG5N3ribUhS7AwrrEj5FUewCRSAaX1rwpswu83yMxxVZ7F9s2atQAy3kokau91XDnglu/sw3Dgmk
hY5nQI3MoMQ7zsfWPLXSkt/xBXoggeK1qeCwYDXnqj6Frm9k7uHfNMQvVaFMWh6vd2gDuKtNGo89
vwak0Gtqn7HOLuGmmK19+x93fKOu3WytoDSyKeqAVnjOepo41DVCkoWAtYlKEacH6+T6j16dv/ZX
ZpWUmMRYpxta5/NZ/atKYPSOYhb4QYmkQ1z+Bzb0l0BCZTVUlqblTMjvlbrY74YgLF41EyXM8Wru
D2doW1aE1AtyT2kqvLBN1hBhN2xCQMJDo8a9w4FqXNhuZQT998OHhWFhw76OEXEGndm34Ht6KZDU
5LnJneYWFyy4hMSBfkTlicMBsCduN/g2jyQ0ejhFFsok/nWYHI0JsZzg2ZXYEZrqgC9QK/SJJzAu
eiMLnvO9hegu8stNzV12c24qjKt5OB6H68OT9c7lFufsAJ1YTdo7yRkNJcGYnwhuUWogaTAs4p/y
aIj8wCduO825Od+l+h7u+7/yZ8yiUhKbXYThKSw7avZFxFAhqDft1fLgi2tgTqwexIWiKnhr+WE0
to22z5PStLF/9QOY+0G5qGUDQV8XB2RanDVsdT+3wWQTC6e5o6p2bzKjV5/aXsHMriS5NRdA+Gbk
0qm/ivxNGNcQ4ahIOGSWjjOSw7R+X+PE8RfzeEhlmMD5FW4vAvMbQH0cSFK6cSm+ivGJze/67mf0
RfHmt1GTrHe0pkVrGhwx6RQurv2Zh9YtXHz+0OgsvxyrqMUkem+wpo1DNWzsCp2dL77Kknf09O9h
rgOuwfDQTe72nGZMCdf1RShbAKdgVuRBsdgW/hbu2vZnu3ZMn+8HDu/1KK99k1+RGQRgf11srUVR
5ua4TYNCwKcmR/r20DX5CJ2OsqQW5deblbY1ZSLusw4GIxt6cKupvLRTVUhQ393kjAM9gt/DcwaV
QoRAr9Lckmkk4Kh508oSwmvHeQWPpPil6gwHLUWkUpfDfx7DI37GH6au0hvWxHOap9EUc1SUoIB6
OcHGYD2b8ExkgOMb41WfWRKjh9mhXChn7kjycKmzlXeu4fe+4xpfuOi28eKG7kVIxuWZUp4gFLYF
KOMDbKsuXK26ofnXb6+I2Tntw2dTrhO3uBiDemNwVkE8CnJUPt+9jBGi78HDWY2ciZg1riWF8RMw
odZEAL7vA4Xcmi4kO3f20bQVCZf5JjKSQodZNzDUrFuxKmBRAs75whxqxf4DosaBiPviJpgxmR5Y
JIA2SxwQH+Q1cFG4rMn1OjMvS2JUjPVMbVmukQ+NN1cMb1MXMbAVozoLc0ikDzfGi1hXFEwogvd4
FgLJ7RsekuzA7jp9XCLiSsmXn0paS4EOULrmqQjYQ8fCJER0yslr6/4l9apEkH6n3rfGeLnrJDFM
KKOAZlpjQwffheq/8yg67ZDe0VLLCyvsE61AR0++VqrW4fx0nFIdoG//prH0boJGZccESs5FRr10
wQRv8SvM3IGXWk3R8s3xVdHoYaEO2kverPfuV2Xjg955JVfVwJLr228W0pbH2hF33vc+AtBhHvlO
d2iupncdF7FZodvdFIkGYph62R2WAXqP5AQ1Al1pKuPbF3/iHOo87W6tiFve/JvIaSVoEj8z4VB0
bsTGBS+/T9wHhMOPH0ZRLwvVNfg9H5xtmQaexsU6gd4cRSN9ZDmM0rXNDNmjYf3yyETk3kNycaoD
aYdCqZF2gCJqFUjku7xg0zMdwuLArkgeesgUZ+3We2t1OwnujufTEAJFUa9vo5MCC+VPWBti4rc7
ZsW58RGWubiiR98PdatlM0UJlgo8/Q9neURwugewA+7qWOOhsoRmuBR2xMoQccadXV0d2Ydn67Mb
6fx82xZp+ot0UpCUQPZfkxr2JLwF3dLI52xp4JUehWEA6XB9K7XjB7nfCDwijXScxPcFH+BkUflA
9Lxxp0zM3Uho9gIVabwB8bQ9rFzCNgiJxZcJLKfZ2Lhim08390b2zPCDNfji2UzBJWH9gMUWz0ot
2v5aN5jqydGuAPpXfAPMUbR7owRWGM9TCFsZlkqmSFAM/yHfIy1TfvJC14SsyMuyvRrSW/M55HjJ
HmlrWurpJJ25g3Aoyf84MBf3I0k//a9TY1s9XdetF3fDhO5M5ksrqWrVfWIzxIhsDAS1GIFJyQ2O
opu+GjWcvE1CtADeHyOmkru7tqR2FGzmTp5kMKGSsKqtEArWDbk+fkRfWCfhsJ+arf35PTNePumA
YMB6eHvHDFxG5m1HQA067Oj/enHJxso5gD/WSdRq2ceohP6S4peRVL40Qwy357w6San5nqAFSppP
PKG9M+Kbz3fOTmQQPxBO84YFg78lrpOMeAbsC6JYVAtvPd/zZFbdiWtzNTO1zxXuP/A+jZ+LUGVy
g3DygJ+yOPvi7xdLzPFiWpNQ9HOdo/2nHluBeWr+2NDX50/4qyW6i/QS2q8U62UUJFxBoxFurBZG
2VwMRuSRNVxChw5C/rQ3REji7ggqShX8aljqDjH0guCJxsjK4X3wy3I/FyxkrpAqEQiETX9rR25d
gitmvP3DIvDBoOdJB3pbCr/XYwo+xxF65PA0mpIHj3ZQu1108p3rrbJfM5wBfFHSMvL/4KM1gzmr
DtmO1K6jTcxto41OlyL0abI+OO9BwOYjWkgS4MTebAZ2G2Azcf+IVjU1KYnn83hRNkz+X4Mwid3T
hw4EttapAkXUr8CMWCc3d4XOesi7Xmm/dkBb1B5ujpXvfaCoxh7ePuQM63wcoTFj7gZtWQjDzaMs
RwBCH9o59+ntC2/5I3oJFTCHVTkSnXw/KH4vkqVhjerzYHdT9XLY+R3b3cmvMxdoOwPhXHS3dyph
/tJxk3nE6HrqIuLgP7QeYU9gdPmRmGrKcjIoMlXR+YO9QY5beBzJxGNOHarVAzNcbFqeJSJM7boa
E3qxhn3weIIq5U5IYwNT0dQ+EeXAE/jtJCQz/t9UN+EQoG1q6yoy2BZlK4ssLtzvdh+VHOH11cjb
TYstUDqyOZgIGg6QUFeOK3boJKi4hQ0UU5a9doKyHE8qBliLtoizgwaC9nXtayRjsR2yL0+AKS3r
IXx5k3EFeW+jKGndvEkqRVVpN41TX9fkFPAcbJLHgavqX3CG/mtsdu6/twjNjAPL9T/wrBYPDPPo
fMNeRhGD5JttRIxTbtV3sV4Y3KHFiqEukeuIbIElbwu7R5KhlnyDTr3jMbzOJVADc4ePPmmXleP7
PEre1WNfXPcFNZKMtsygcB/wsxdB48dMZAvp2if/INh8VulOAIIY1J2bxB6IaFOKdlKFNtQ9Qc7z
4n6m+wzTskOPtgbAahrNu0Jbn2mj2pNdJU3i6eovKZO5HYsOOPi+3gYDC38XOxHVvWNbRVHeZQyV
hacbofez3SgTwK598PK79wph7coXgMsz2JrZBPlikbjelXdwsumHFNprkNpzidN5RtX+7QsMCcb7
HyylCbWY8H5p65Ji7z6/Vcqpi+MGDE9+sur6OcDklQ2aQ6qnS4zqJNCoKOpG7EtRA5+R5llQfwIv
f/WbWhjHdVvsd0M0m94GH7x1R4BLyHmkG7FRMOXhIR1CDdrHsb/DrXQTJ8AiMMWm4FUa0VnT+ZW8
WEgjSdRJHrPBm3npWFqJwu/5iNBQOiuF3wLj+VphipGUxTmsbSwXI6nWCXMcKRthn8a5D7W8K7UP
08xJ2WddVNhlatqa/O+69UEMGLpiil8LYLS8xJfsXQ34pkluT9lSrXNAHASygcHbKQMrRiYp9mEB
9PWLJ1VB5AoLkABrhvLaNd1hMV8KS26w9XeGL6BTqqgEjkx2sTC9pXARdszerhOvFwJaT6HiE1Nm
IVAks1YRA3wqQh7TcdgVwuMcEmwCG0jipl9lUGJc9lnIlwDHz2xYoYsh+S4AtcQqSwVkkMDtgatt
QCqev1W4r0eQpKjatq8ZUfpsHVbmZwNnkzuxJjam4ldowDUB4GwZTGtWNVLEl6pWH6MqX3UTpB0i
6HL02C8SX0VKWpUk58IvtdfhBeD1YbSOgtRVrLJPzftSoxWtAoySPk4Eh1/RXcN6sO25bjR0xPVN
HEMlFsJvdTwrCe8SW7z2rCdUlGGLa4smSGIsXY47W0++NzfU9muAzEQcTn0KIFhwg4vtrFoKfnAQ
n2uqDTDG7uu9vuZV+WQk8JKxfeKuoRz7gA1hG/UfyzMt1FKa9oeaXdFZOtAHO+PB/2F4BL1vY+By
4HHTS5JE5nxwhwkCqB2VV3+9+yiO17cf9xov4rtdKp1RuhEjOkox2Nv5hQl/ASIimgXWtG4FBQwO
9VaZBtHG9rdfZDnAxVLCZ1caTgLcRDGp4GSN9Zk9nZQLogwQKfS3FOaY1FFXfgaGKenyAkMYX+Fn
cPyquWLY2rOJsWUqc0FlVe9+oSqILVA/xeu2fv3kdc8nUbkKlFG5RAOVlgsIlgdfoPWl14SW5G8q
M2u9WaL9Ue1HJ8xlsPdGRLnu0HQ+tbg48pznvY1XO+6FdPIYFLrPzp+4XpNJXAGiS+tiofW+pUAi
GZPxkiMB1Gu92zguKeWdakzxctgnLd8T7SeyDSTfPdrpFB9ga/U5drN0z3ORTn6LueG8ryREWnZj
UCI+aNbTx7iPjytNP7FrxvXreJV/4iuiYFsgcFKUtph0d87eNvLN9I/UeVQIQWaygljqddbjL3t3
SMx1027n9rhi3mPQUpIKLUhBeGoGCWURWi80dlB67XOq0RLb1BKuyLGNnrQYdF6pg7oXjQR/QCzx
xV1x2ni2I7+XWfDf7Hl1guHEp4w0bISSR+6FSdubOl30wLyVkr/A6zmwwaWFAoLqgbe2IDm6PTE7
shIkuC+6U1WUAESIB9ozra7Hph08AJ68+UeNJGMQc3WVZVVMe4XmkqEhvGnU9Qm4UtLFxJblNj48
HvSLElhvoNO27+qL5EWDghi6l0AmELn/wGS0wi+E1d7kNrQR8SDcOfyoBx47tJKUd5qlatAYHs+E
/xCNg5hdOwRIsv+G1ieFMPnxQBTbUgl87lbyHeCmOoZNnStFCXjeILj3Zyd9xC2qpdTrDgc+Wdlx
PlQT2NMGJb3Qhiqdvizvy61sfCg6vkIhgq3fiTzc0IUO7FObKvbfxyPumZOIK0l/ODIElxKd8FPD
cPMvrG0bjge+lYkpL9zs/tHg2Vi+siDG3KZnWTJvbIIXEcV6dWE5erHCHK61Pv1mKfDMLv5kvK/t
E++Q0B+QzZF1YGicDRiOfAp5jTTzxjLry+WWwcQuJyyxcYgZLNpygigczogHQEr0u7RGMif2mUAC
6f8WEGc0enmJB7Jy+zNezgLFuY2SHrATp5iiMF67DzZP1PSs7A9NGowjtP6rMRpcfVbRu3MeTO/q
TmCGY9oSF4IQK7sevovFUrbX/6M6jGiT02NIrH3p1rNKWJHrWJynoi6CT9FugGbQnPcGiXIWyDWh
w6GeduTAEUkIYswFK5BswIgj+zSZuk6ju71U5l7uYFbKwwskxibbAxflsJNk/OrmwqXKg9pEm2F6
Cx4I8srHYwai+r0POt4hMR1S+SLf5eDijMY3+1whdS73E3LwPaLMyQfU6QCmm1tOYl81YBlhr9SW
YY6NwBE037oRgRXQ3bPyQ3R5EcKmLY1IkFRy6Ua0Bzsv5tksc29WsYCVz7UJYYgaQNl4eY/fjfIA
CNor0nbIJiMxS5TYcSDODcWABN4aVqp42za14ai1onZn37qe3M64VJCxeZUcl2zpS2JSeeO2T7D0
aXn1NjS0zjy7rBqObhg3BUyKcUGoex7oDoDETNFJEiMYKDmY23FAHHNAr/PtHefhKf9Q8Q74+rGl
WnHdv1P4/aEZ+Bi/0ZoQFtqkfQWDfd0adV8b/DMAOeNxNTfcGjko9MNMpllKN4xFeXSrdBDA3GMV
oOgtGo8hFT+7WHT8mIa6Y7YMDnieCsYCGA1sdtCaHglAB7NZIKJ5slC7asb/AP6qsU9oGveEGxl9
B5Ao4om3P0ykJrJOimaFxD5Q8bYCVciuw99Y4hC8PiSjLh6aGDZRgnH2Fz4J49po1m6SQCG2Ud6B
KOr2yY2sChHzcyljiUUPGLaswwkynO23thBibe2NUo9QMEVWPKhqbqTofR7ap9OLjaSpdFGbVt74
i0pGlUqKqma9ZsK4WnmbfnsVjzA30SAbUitgUY1JR9gb8y2EAe0bJCHvnUlyL1Hpzlfv/rQgDGbo
ZIw4nGP32XLwr7auZUy0IOb1gzo/f1TnUM5CMMPrGT8/X522OT+hka4ZJnzBfUUm/zUBJ/T9xudC
bN0epwqCqaQne8HjhYKHNh7W0TmEJ//7T1xWpJscmi69AiJLcI2lIwr5qmHPZyVcdNae7jfO+zK6
7KiQI033uGDkwfN+8HTjnH9Dyi4oiJBFkDHhidiDInnKuKkDqka6debmP2hifBBqhBMpTIwWAnhC
3GBr4jJTluTQ7kjFltwl/XvN9/AdZlWoswLaEAiWTfm+HWVvYoYUS4E7mC4jFseG0hUiXtm1Qsem
KX9zcNdPPnEXmpePnTTIduYhHbKNdzzzrbfE4v023/2uf2uytLXyXSCIa4+2BXZrd3UXoW1xD5tN
fNaAnzJzAV+X2Okk4Ds1hPJV+dlUCgkSR2SdsGmOd6BiFMLbfD3bPn/XKOhdQ2RtGTb80pjlJU4C
WkHknJHZyjtQM1kXjow7MJuD5Cejo1Ae4Lr1iJLwdWj5LUHmnQPFlpVGGS+oUKb7XokaWSDtnDMX
oUSGFBYyHezfjWL+aey2ICQ8aujGjCJSkdvYlJT1aKlnug9XV8r2OoO3qYvf0Pgy7lopJNbAhJFH
pR5/VvH2fe1nuTBYo4+1v04o7o4U3HW/waccAdIe6ym0BSWuaqiopX6mfBlY3g1LajFUkEuHIK67
owbKMFNkHc78jbGdD34WRgw+c8ycZXIAayxQsrxasw+zneXOGiZ3DU3JLx+gAMPDe9v9pvI3hnvN
i/1RjuQ43JvrzeGaes16F2t1Wg0zvmGjWoM9j6I/TBoMRQDLfDhxWW46RJcZOdJ22Wvyx24udM3n
tfUUTr3yIRvocJo2OlfFiKOA8rvqiX3JhI/pyvioNr34YnepLkj3/Ymq3nnAI+FX0B/7/dQS2C23
/kziJ/HvIUoi5qgdjidfcGTAeJyWd5zm51SXCAGJOnI96yB9987P11p1CL2GpaOBmrkdMPbQu3/O
L7HpUxat4c0zen1N4wLza1rmIMmSHmYJdOnUu63J2g+p+VU94s6eus2leXMe9J1Uqo8q5FGopLeh
THRy7yGUgqwwUbjB8ESVo7eWxCjDUspzRAjY/ufg8fcbC4KSh8tZ6BnIP562kcMA15wDJ4+zQc5g
rDmISTHUB1ErUEiH8kr3CNuUr3YLz4pWCOl5hVBuQsF4hfEyXM5dG8wli4gFg3xCow6+tFe9gTuC
1xb4wM/O/vaBiCJGLKP+7Ab3sEFKRKkNtAlBd83m3C2uCl7Z3TofZ8yVVSlz59WGD1NcYQM0WWpR
mZQQqfQwD/ogDnyJuPk970i+9YBYLtYOwO92IF4Nwm02oIr3xJd//IjvspEB7oz35A1qKQkepygy
6+4QEioRfG1ust339qkn77E96aqObqXYxs5ho9hI8qwbifCcDhrm0031cRi9jLiHEpsIogyP7USY
8vlBbcgHQiO7qAD1cGR2jtCQL1xC0wljacmnHYVU7OH/BYKpPMRVWCMNEoMHvgCWWdWBQru1kw68
0EOXo2ApcsdaVuHRqqB/4T8gBoRSSZNewb8iUdiuGcIluAWllopmbNehjpzL3x45Vm9QtigF8MnO
igCEJ0FPuzIWnEBopfpgAgYH4NDbpZVGcZVCUt8laQljF5dNxdz16vgdS4nEwQ6N6caR4fyXJvZw
SH+LtTBO9es2lGhNtJYVcfcZTf8nmBOUdzxPKLU+ET3GuqidaGc5LmJ++LV0PnYYZjem078J4BNl
H3w7cV3IsIopBS0jfp5lbvUbzoIJrB41C+Ye7KK45MifFytd57XRQ1fu5jlDC5ci0rXYHU+/lbBh
/FV+IE01/nZQ9v2iScFyng3CqcDfOoknkOvKLf7v+dz9XwXEQfoyO9iUqw7a0je9B1GzbvEFHlkL
fB+hCVW5/KiCECrBr/gp/+HhqKAeD8UOKU8SvGWsyWCibyPa2bkcxQDRNCw+fb7MXvZHXUFiFpo9
C8VmFF/f7NzYrvg0Kc2LOr3fUN6s8VqmUMYAUHN2Di55wT/NmW8jZmf+88Pa3OTNqiC9UAKrKUpb
mRlGqzVn2t/y6ubngQrgxW+mY/nYXl+X5xQ+5g0lYkvSzqQJrAi7VEjEEZ1zBe+MGp8i9dk1UkDr
lpuR2lUriLM70jlhWyM02LSozlyrhWTjcc2JYQ7finV0eqorR3zEYtVTlae67ebj2QVrdAeA9ILX
/UyQnjmv8veYPmKwyhDT4+K0fLn9/RgcWyFG7XoOMQcbaskfD/cFSbgBKFdb5te5Zjkirv3zv+Z4
KuWNRKV1dNkcFU1BPjcUDAoXQl6UafIWIHdW6TXg7R5tVC1DSBdqB3m0t6m9pi0z8Wa4M8w5niZp
xXpwrTRl/UioknrBXowpszQ/yNTjfYTcmk+2IfQd8O21njtPEYQsn80d0aNiKd8tJSkZF1K/Kh2q
8XViRW8fEKFSfn1M41y+gp8OWNOmMl+7SGwOINbJZnMgPDt11Dz+Nc2FRnOiFHaagWvyM9FX+rsy
TqPfkcLk8tch6YUa9sLJSneYn1PInxLVNsoIKWzDNJ+T7wkLWY8LqX9fee4hedNn9kJ7LsQiUgRx
HxMX9lLMT0NopK887n76hAfrkUHCuKvypQHD3G67TQ7AXbzNtEz0Wbi1sIGUZ1JDd31j6dqizXFH
T4VdVaOT4BxXIUwr3mE2oUOA2+wjm2P5NItMqeoDcT5d19rEG8PkAX1W1DbmvcvIwoQ3TUtx4gma
dUk/5cNxBMFwvEM4jVFtysnhxSq7n3cT3rcWEubtMVADlxKpVqCWMY3f/FRg+RVdbMHq4JuHGLly
PQHcLuSDe76ifF63YBq6DsigEX6RUiWPBssIO25GT4cTeHfegipNGPXCsujB2VKP/CnD6xKLZhnx
lx3lLMZiNkDFOLTObcQ2OWC0lOApYHt1fgCsKCKFNtbuQwPd8SBZevsL8H+0gJucKUTnrbjAWZn9
9fMJNicMSQjFIx05VcpMTVI+GWafFvH6BxbpSYD2rh//98QHKgJmApz3KmtqiFBnn8pjIicpApR1
/U/RumXClLUofMxKhfPnT4tWLt/pZ+MT9urCXQTeysXz/c+9Uq11Kzf7D9WgrG7NQ8DMHyM2LL2Z
+6SpAiwmKDaLGfTR02F1rqiuQAsII3pZpe8M7pOevfTbzJMfpt2nXKTAoGzESr2cUL3LgpDIFDv7
n4wzduaFPP6/m+MAcntVP66sP2Rh+hQjtPLqyoFkZWTM5pudvBRZnIoIxpw6mYZ1bjxUFY3o5ADL
Dvu1S7dq7BI34QeO0VCAqiAKFk5WhsW6W6kRWVOTJrvnQsZqgmZKQoBTxFfl2v4B79d4stxZCQwD
OLEe0sFMxBB/PY62oMPm3UZoyilmJTnJji+NdH0zwQAyywTvETgX23sIjQItNpvdX9jlfECbaj4E
IY7oWB1nMlO9JdO/eSi7QQeiuV8ozuph6wtHhpsSQgvTaKae9uCfc/RphDefQ+7fB/69TGSKgHFd
BHTsWO7HG9zYc09l4zZuh6o1X+1RJnPdP8He6W4jECzcZZuSkKenF0gLI7NTDiKyV9UeRFaYwZjM
iyVIlrkr4dVjfqNsCMtPc6JmOMyg+QZZAN+8B9avgN8rJR1gvfTMLCFxIXbCb5k5Um2IVIFltYHj
yKh2kFhg4RKqpbsgXYZ73CqxhswwksOF5mNW906F+DsIdNx05c1oSoOhIQHf+xOjPDqmiTFDNRoi
txlDeMFlg3sAezuL1e24hKlMc2VDzh/E5DmZcbxgOLg7CIlHHpV3w+Xf69QGgVm4G+xqG4R9c/Mt
vtNbaCH725bEBee2ztUwCZP8MBxv3bcOrb7XtRLp2XfW1x8UHdWs/cKo5TR/jO1DWiSNb5oaiQ2Q
P40MntGg6Ed+JAJXp1MpqhqdnxlSfUgyg4QsaCsLTUp/d+xBGx/P7a0iMD7F0hRhI5FyM8oRoVZ4
1lqk9PMWqYfnAtCsLDl7MiAnV9EJrrbRunoyJlSYIya4/2VWu0QDLVAwrvMC+PRtkTVaQ3WD9aai
ezbEEpIEU9wYfvNMGi19Z9+JyRUuIXQoLs2qXF1nUTlQ6mOZyzt1MmtPX8MfOJ6VMiFb0O6NPk+n
B3Dg5DnRiI0HyHDLNbX5tGFMLcdHm8+Hj42YwpK2Um4rK85Y8ButItosMfg5BvrN39WLbu7A0wY/
5jZ5f8GAIuJsXPY6uqJ5EhFiQm7nUT4eDDsx2rK5J9z+CwYn+ayPQtwyfNTtu7yHx+zEZuiY4NOG
x5fVaL+zuXkCCej2MQp/WLK8z9btcFPZsoww02BPMDoqeckUNCQuJyb2JZjwx9GK6f1w5UK9d29R
E+fWnsgWJOOuPP2NSkuSJq/DrqZWn9NJWtDheECsWckkuCvnkYPQZclJz0ZhAXHm9CIdQYV8hdks
N9N6qouGUkRuYO6yACiXGkuzK7KcSSBEsrFwDV3TdzCbEZ88EChBBpGygxu2JpOc9yyqqjbP+cl7
hgIC/+KYaeSTDKM2aUPnFlicfyg2Xi7t9xl4qoGkDwosbm72VCMZpdmgdvQuhpZkWc99iAl656hs
BfLZ0Tl64mTcEhI6tSRmRDwJnlOp1zBErLDzcybbJjaaRJF8W3uPnKAB+WrXmoZ9EQvBoL2pZwmc
lAKt0J3gC+oMLDAj6jdWQ5JUlnFscqhFQyQ8zkHo8e3Z7umr9JvoUMZzcA85TkDguObvFdZYhCtl
zpm6hUnBVQdwPKj+1VuJljgbDoMVdCvuCRaxQax0ky7SXtIATdY8e4T1adtjZCJXxUAmv1N7rMP/
SuOb58U/GsvfIFsR8YyIj45MEphsOLy+kk/qQR2u7C/R0S8XWZo6HRWJ7f/QEglv+P0adEMzxt3b
vnQZ9WV1AQqy9AG2su8wZdU103Gbg8O7pF5YMsAqKQve9rAxDXOn2RzfTiDHV2qoGcgBNdgnCqmE
CIhfH7mM9Ro06rhr4z8CkVBXQlLjD/6qcNFlvuVEW9HTOEwhixVmXBiUB3E926LwrZoooSspw/4T
uyfWVoMP70g76eUPLCW0XSMoWXcyNjweCaNY/e8IJ8I2iTBuVCqC8en+J1zCfdYFGn1WsISBBGiN
lS3ZCRkP/ojkib/vOIs6wp67JaKhA65xtA+ElvYo5xCaGj5/L29s0/9YWvyr8AF6JUVJGPRwqicn
ViHzb5EUahq+3b1RiJ5lv/ljARwbgMxjVzz/HunenhTgoDA5oP1M6CgH4ff6458zBVaGsQRIcqb7
KDpOWzt2LYnqCq9eeYaW8CIfTxzfE5UcCNrxQWwJEfbvtHG9x9ogwywnNobdEu2FXQ4KmrT6ZXyt
NcAE3DEetBC9Su3vQeZkgc7jPHbRC12PyG9eds6pt7q/FFjgLvDFUquco6YEDJK06a8TLV/dhonF
KlWD1CHCVp60v7buV5jBr/XW7ndBNKCwd7YsrAx19awWufiyC+G2ZhzlNKpabza9hxIoNPH9n7tY
HeXrPalX31j7v7TMyhhaxfl9PafI3zYHpUG6nx7WuUzuQGyCE6VjAdN4KrSAR+gKx/9PxEW2ZH+A
OvJ5r46Hiu73CCI1roqXHAqQpm9DhIghF5wm7GJ/rSEfoknI6J9TDbXHCtNT+aQZhfV+m6eo3qNO
cqmdMPvPbMmNY1NdRSP6eFIo5pZzcn+Xtfm0n5+mfvZMqoMnSXxxcx2Tm22HWFv5iejQ1YSSrgI6
CggKOFWJDxHpmjEkZgyLfVU+YgcNq9OpbKsB8TvyR9N/2yhzTii2ZjNblzBY1JZWiCs2XHT4rS9F
HcIYvll5/Vo3zQY0mhn3KcBjFoLD8P3xr2Gjmglm7oQUllQk0lQfRZ9+E2Rch4A5yjSloiN4yLkD
KfVlFMGHLO99gokFvsVEKmVS/4SYFhcHNga/2hxuwRuK+r3XPVegF2pMlEQ/xH64H65xjcp2yHHK
u0cNVYSNCqvq69o7VpuBRkpmiCjOiebXU1EOinbTS+9kzohhhPQcxW9E3USWzZhX/ThTSRBvSbdA
83ZAFtm1gfXultWvl7CNBZOY0ORC570Gl2Pl3NoNOcm5h+Ynm/222sU0bVXftlKF9Kjiqinz4NcF
XTin3AAJfiBiVlzSQ4T06Y20dwZToDgYqyAyjkSig+nwlu/0L6UPd/WWbjNo9lzpk8DnJVDyIOta
Z41oHiXazm/Ek/AoXqTtuI8dIUWbhmsWEmF+znTwcdprlLrkhiY+rYgBsFcJAf5YgMCA6cCEts/+
7+V92EcsrgJuMvzgBV7cZNM6/kb6OfHHz3BaA4sPfah+dwo7f/NtJyPqvQxMse8PMXDuthg1Jgow
bDNXngGZaPWsFz7XCJAyLjqtoHjnLsSQsn7fsD2coUo5aaUwrV/mTm5fWROzXv/DvqELJg0S1ReO
r+vmMAPo3LiX3Dp0Ie+yAROYDlvowxwaaKcyCWp2I+G6n+94UtZs5co030AQfppcRWGI0Zj0Gbm+
GxifdWbVNbCSHkZkQpptqEuNoO3Tb/0RTEBdENleHAaH/mDHksCQumshNMWI0qW9aUIGS5xAtvtk
QjItLyshNxHKjpDgQYSZAtDJeurd/lQOdhrUj5P5OfKbBPzUqN6bMXBSvdU8pPcJf1Ek4sBeMx1D
dAUN2sJ3S3/v5kc43+qHEKa9LrvyB0hjxHzWSzICHeAG4jkKtk8i0x9X5Rk5JHZFl+ff4Chvfwcx
tm0/z6n3cvBWgaCAlIufSsrG19e8Os4sk8WuqL7tnlw9K1qamccovNTBLpeaAUYDatCKm3SyqdZp
c75yGkcu7a+xvqla1lDRNPnega0Dsvj28xtGUha4UWRwAMu3CbLFZ3AUhA8DWZ2seJZR5xfYmfxR
2HmVGF6avCOgmxlA3Oc9vuzPhASh9xlK+fZ3xAHJUrqrxdLk3Rium00x+8eDJ3jXSlJS611nwFv6
VKV+yBtEqQh6mT3UA5tTQEEWrWNT+jf56bpISgOMHzmG/wXBer6GP1J2Mi6gH4mvCFCcXvpbF547
mnXG8Zt+R3y1s7RTOWiNBdaJ0q0o9ssdIMDDigwtxM9tN+5cLfdoTzmFH0sDL23MWsZFGkItZF0a
sRP4eXG7ctIKlnwU5jkoxwKiQaGKME+B6w8YuNwltFoB6X6q8Xfut5XKRTAnevC86Q3g6zMvgdVx
9mNabcSltxtW0Y9H7xcbijNpnhW4dFJN9433qT3xCiUyxGEBpvaVJPfjxgbPPXNpKuu6AGXMHaIT
rFPrk51vwUea6jpEizmzfOtgLa5Kurcf0Y2dkrKNTl6/anUynMgCe5ug61NZ1749vgLkvo5GOK7+
t5Y7g2kM0evDxDJMnNXBA6X37pm3CypNu1y+sfnxe5TJSbAwM0avNfr2VQuLej7WuFYz3hXQ31Cz
stQi6mTBojBNWj66q/S4aLT4JaWcjQ+Bhe9cDao62Mi2clHvY5PN7ynU4CZbYHBed3VOlCMJb1OX
1v8T3VydulqhT58IssUnAJ/TBiKW06XL03yb9Y9PjBBfoYkKukispjmlz30/KfNDvgnClOPvSCps
QfqEW4AUIgEZJ6zzKujX/uhcKjoTVsZQ0iM0TQ+gfjnUQDtbMLkfGHu3H53JrsCv+/l9BRd3JDfK
xIZbh1JYVWtCfVPunG98ktzITd0FBpwbHYAkHlXPY0LcdTlEfxnrt3IvSUw3YZgYItObSP0shDsJ
REn67T19rL1EZZSDZfZoeicAAcfICFM13/iNHH8cIPck7tZktjALvT2dlzjw+xT+0g+HCH4sFmzY
cbQIYBx8jETDXczuNHudRi2tjWKuSKtB7MOiMSNjPspmY88bObfxdvcf6JrFDnIDKNPEsXbg2Nwj
qnIp1r8bZDzGCfHjPHoEwi5aIcpzVnbyh45OfyMpL5EhMyYEKLiADvC0Wb1yDdZf9/b34aOy8ptA
jyrQnO1RaYQTBSr+qprxnME+BsC2nRWHG8V3BZKvc0t9mtpdwrt2f4FBfWKzW8FJ4qglRKaZA2xN
E1Mdml4zp5fwZ/H7MIm8r2SyU/Ximd29EVW8QTbhCiJ5OkARxGaJ2lx26Uki1MGn0u/S5iarVx6k
dDsp+0B3/PV58L6Xj+/hSwHDsjOp8Lwggh4uyqQe96CBqu2hizvRLeNShlDEW7GDZEePi3fGNNQn
/Rq1FONYod21jZ/x0XC4/azcwR95qWscTKrCxSl4qk0D0FwrPu2NZZKK4YjByl7k9cgYesGihviM
L1kaEcpnWqYQ1OqFcvSyXhwj572mxfQnqQRqssNVaSLoVCHZvAfi5i/SdkuC25cq9+5oLdOGBttZ
nzcb5mmexP2y/EymJ0Fy4Xs1W/nFNLM4oG3xWcXaBQ8DmfjbNhtx8vyNAwEnzpIol9D9+TUEjPOA
Yitlorq7IkggepY5f92R5uzo8+KWP7mYJZFxznLBROCgeKDTwxVTs5n8xabe4b+pBZ8tun42uSKu
f2rakoOlZ19+vCez2dayTluO8+7uF/6Q0zF8UK1G9V5imKjGa0Ml/KthVNXaOgN886sTrpdHrrf9
fWyhQtcl37QwmwmovMuNkaHd5rEmGWg+kEnic1h2jPuDVLCN2nWNPMKUQ53N7fzV0mCl1mTRQOfo
q3qUpVBskSoOJDrtgvk7VD3Xzlf9D0Bl5eL43/R7lAmAEa8SeMmvlZDtQL5a5VkXJavjGukqH3WS
ICkLgX+/M2YrjnX8DT2CCHb1lj1xYX1jHgW9w9fFsiqQCfSw+WDkjerdY/TEtslTxZoI7UctLplO
KUmNeFtQE5GlUs03JOsHWW1xJH1dBvzZs3jD1eQOAzrQ6Qm+R26K9UWtEAL0OFm9u4yJ4PEzRkpm
f5Mi5HHhL04thEL79/UOHwybiJvyjtDaH9yP2U8GFtQpKU0TgBfSxJtghRQyMhC67mBum14IgeSH
bmv/6AmLSFDhdHc7rkSQ0kB1f7yP6EDBUmiYxYkE3ZGAEeUdLhdMwDVxB+ak3FZSYwHteRgLDPvy
VzNO8QkNLBdSzfxCwBFenhC77SDz8IbyCxGBlVPwRYUltz6TtdoK6poyIllq8NHz9KFI5BYmtZUp
MToYsWlLXwGH9wu1xdPh4oUAh0AJvofiVqEHSDuQkhcctq3gDANQI9Ud67Y2AOCKkph6X8aSeyl1
Y6Bb7YZ0ZnxdUyQVQG9NShdjEYvE4ZwK4IEnQD7yonBnuInJylfkIPZ0+QV/T/IUG4qxzrFV9p0y
w+8Ll6ppgVGfTzCmhTozZBvyqtnt+zNDdM7USh2xdGBVTTeO0w1O6gTZvMAKfiGYh32YXo7ZnOOm
JBveeZYc+XvSHXFGA2Hq5fmCBG6IQ3ZZ/P0LqvWW4hlQQIypJnr2/Ym+De37iVVmL4CutJVrYXaW
wqkMxh6t10O+VvBvWchXe3WG0jZlImjGjlg8UmtD6U905bJx55V4o170d/siXL+szAUSW/9LkPPt
C9BzZi9+eQONji08hvNVOiYI64kdy1qBUGQh/nzj2u1xNED+1eiuJOuXxE49kB8Ge06ms08+cV36
kQugy8Yw7tZWThnT6tyramkH21PLDLztY8u/vOmC5p0yGPEDMS/ZBvFt2VYJyclNg9KCJX41za9n
BTTvrLu2sHHcCD8k+M+hxNLC3bxChblJfq3bCXIAePvzZ4QOsCZ3a8MLBIWvgxU4k3E73X82312/
MWS/fb6lENNWGF1t+EH74BS8zVzrXVgzD1t7Y/zDW2dF7WDVV2Vd8joPtFsfJBq2cvX2O2cdcjgM
Qm3BH8yO2/GjNjP4LwCc6Ix+v4ICNHbmpu0cq4QADuP9/tkG9mFxWIOUt3RFh6lBhzwu0yjZBcoz
7bW4GEXkXc8he/+/FK9jrYLG+95khQR15jQxoIYCoVxdKHQJZrVqHqx6sXOI99UU16VLqrW2DQ1J
YxB6JvPIBZRMruJSBtgGD2m+YyygCidD5JzWliUKtmoTHSv9xYZ314LGCmBIcAkE0vi4D0g4rjGc
mgZgbFDDxJ2wMLvpafaLNkkQfMoNUIGFUAx+gzvOxHvOnefAnI/dDmJOPTJdf0MJwrnJZuBTCYYI
VwhrDL5SHXyPgsiXEae9YTEA6wJjVI1JmyFJK9wJ3Dj0qiCNZywtl3R0fZgeTl+FQ12FUV3hpEIR
VxTJBwI+0urVEOJ9cKxt3aFzMhJUp2GG8rAJBkSeNVJjpzbLHFftmGs2Ws2AI2/bMhkzh8XfAbsU
fqYFnCP33O29YD4z5EFWioGD0Pnc6/W2PI5IqMK4wHjF7++Ig9NSHTYVWbcnBAfpAnVn1wp0ZlOq
HxQnh4EBqefzjG9sgzTCg2iQBg9a4SrFZCA5UvTExlRUoUJCcbWXP+D1pyb1mfAaiIUmcFb7PSlK
sd1bM8xuqIpkQMF/XL0VNlEr+AKHh92EFJPeWCDpFxquUEEPqYBuexAQSsh7qinb+CRY/d9z9hdq
NGvgjJ9X1f8qFNzhL8Ok1jHrlwPS2JLq0HHhPjRNOXj30U3XINk3FhZ+TYJeNPGGfxSoKLFoAkJ5
9WMUR02buR+ns/GVHJ8v7x8x8jR/E9X6wYnd3RycWQAWEDMFzr0h0fuQQe4jCiKzINi65PHRxZ50
TPY6NBD+dnU4DGfv2YObZIN3SpwiBUPFRMWEFmR/GDcgzA8lgCdSTj91tVSRUwjx7fQGELHsq+dY
Kv0BymVBhv+KjstjIvw8y8FDBycXg4iKLCxUPKuvX9HYAYD9xMaJMZdYpPTBMi9dLTf80mOEewzg
gSvzY7Qq7ebhPwLOfD8JAFFO6UhZrhz29xbm7LSuhjbNby62xm+ulaDsUeAxi5iM2U+dFpm6dSY9
gGLEnA+e1j85toepNI4uev9x7z7XatcBitAGqFpQ40oZU1cCZTwXghdP4MM6cxjCGldZKnweBc2z
+5ei5/iSIdrEdKUUB0quCiF3ocuXQj/w0J97V3JE33EdaqtgP20ZKq0q1k1yR6aPmAz7owAg3szO
GinAROyaFVwz67DSQ3lHbkTfb/6UINxbhKKCcUdeP5O6wodWvbN6VwoiNX0xvHigpzasolc4Mh5p
MtFdJJrXux2RSTca9Jx7AIgAblOtBGmurc3fwrZfoHaMEFcaDWuVc1ro441Besea4m/pnkLh6U4x
rF7XRyO5TIQ3jDy6PBXr8pZ9dzs3nkQ/f/33KjK7CsGgmU5z/j/LP7OK7kyv0AUJFqqOT67vzfDb
1FK9wDw3Vllvv0e7hnjtWDVixv4Xhdg/vd3yD2aPFFCayaWYkDSMGSvtWP/9n7kXBLHNyRuy1zz3
nrRZDYKcGy4iHXT1a24Jye/ogEKsj6v/Sg1h6t5Tki2QXSOrUNrOQVlR99a91jTY51iWah0Qmx2p
V0X2vDZpUP9//Y/hxUZiynv2Km5rKizRp+GUwsh/Wsc28N7bsgwhHd3B5LOHI0Mg3qEqZ2X2Yrl7
ICgPRFwYigGaaSvyQiRnluXuIlz10Jv8h/Qef5WgJlpzrsLWmyJzCYYT+kNVetdIKGzqILAenI1k
Lkn9asNEsSkKXQyG2xiZkLDUYOb+gxa5wPiLjIXvxCnE20oCVNgHQ168Mlh6AhLtNU1BocaxRU6W
BwusErbFX98eJwaM09DuCSaXnr+1PXqAL6Luc+lxXRY6kyYk+REekRrOg2t6Inz4IzJVCbqmC/7Z
XFBto772rxO8F9rRwImcOg3T7c2JNQs3C8RXn12Td+QortcLGJtkHmLYVnlMLtH5bzaoeAzoVZE9
mkCdq7q/SXLSrGjdFJb1aBq++VKE+RNCvyjUdRAn6R3ttk+BobHcX6tK47Sve+b8SrIX3ScXWjhX
BQr3c48y62/42nAk4kszcCkuBT53307IyLx9XRkiARVrGyJi1w5iSWwWmh58Bs/wmLFnj3HnMhwu
yiCJAVu+53WCx1ZmD1cs4gKqcgEmc3Y8YpmOQaHt7BVp1K5E5ktX5m4X6PvjbNA4u7e/5NjxVHAy
NLT50uCsvPQckRAJ9GDKYgyFqwuImJY7Q+GK2mFw3VnG0FHA/ID6AyDm/qqZqHYxMaX96KZr+ydp
mBmSw5E49MvZkFkA6X30lkI0Ckp+azWrIKOsxUokeQgxHpucODqfTYyXFtzjigXsn4W2ZO8fnBA0
/JfTOqyK035JUhM1XK8TBavC/Ghiw00pnRDPbMLLrkHYNyo7UHFZaPD/ReA2kcR3LkcDDTuKG15P
mmBkl2q5xqyE1sVLOCoyMm54ZOQM25/05RlgZfeZ19JHULpkIpLw0s5fBkXpQAoGQAI9sGZE/wWg
SbVhUyq09nkU1m/B4rW1Q/dTWfAzuoG4PnxclhLdkKpIASMaofElaxNm7H1lRYvswvkVxA31chq6
0GaVH0ujdkBzhdgEHtG+BVjoft4btdAcbTLcbVm0BI/UELjp6UrEYtX20/gga/rjDZHV3foRiPsZ
9zglIqMfboMQrHPCLMiaYKuDM/LFV1J0in3rhX4WvppOmJxq/DEd1crkk7dK5hWqwZPTAJatf1XV
jTVp0py6LW/5/mi9SXQFBm3H+zhJXc0TmG7aVHFKScPhZN6PPLvxMkCPvithbEGOOlYbikvqOyGK
KOPvZr0EU7SDejnUpulZNecYzehVgowh8z6kW20b9b4n2PAZa35ZUbCBvWMU28lyKC2R1Xy5911I
sihGiBXs3XeSEdZwukp3LfU6w3gq5itsrUt6hmMGS6qdreJwuDJ/zcyZNQqzwTFGj+/MlyfyxnmC
M+w466cAcGR+mti6CdMocjYVc2We3eA41hF6r8WZ+PaKT5RG2WzsN9M8T1yZ80n+QJ23JQeab6eg
tA7CZfWtWcE9aBjETimrI/MWO7uxg1wxm0X/vtegX4fzR+RgxvzzkLsa/ngif8zJ5SrXEiXEBOwa
LojCXvEm2s3y0ErwrKYz5frKtkW4C+aQCqjwCHeWwz/9Guhgs0uYfbdNVW4Oz1UIpWzGqa5UcWL3
5UBTBxYAiyZfNAZ+BqLYcG/poN7fXlSRp9LQfrWcphYSV75MB05fQtXUWVFvgqeJLTJIPDG9cU6Z
sibP9mDlcAtnStnwLDNbNtVEuKIdk5evHEnWTBiUQqPSEsrAGJp6zgyP5v/GEXTjuef8dT0Cx2p3
G1DEKGQko753917F9LKv6k/djDOmrETbcjXfGYKrQneZIJ5jUTbBoDU9MIkfvTpLbuh3F88F9Vu1
iGMlmIlcsx3poxd8uw9yf065nTtkodBPKEpnwGv/ByjU/8aWZN8NaBEXpMkmaYm6pvKDBwGB6yiQ
ShAb25PFWA0Y5h3MMgxdiUW2/FD9pqBNB0yJ6260sC3rhYtMRQVAdZqk8ASZbXgIX8z0nK7Qdidv
Y9nhxUMHhaIJypppDfb2kurGpYI5sGgZF1S6jN5V5WMdEQ7sYtTTj999sdkNoqTvXI0osfx/OtxM
07A7HvViM4p+j/bdPibiCEcGUrFj6sE8T4VuhJ+717ZQiFieT3GdLES+zR2G7d6Gn8YV9AjCpSPE
ql5wvmp7tNgPbCv3Zgw7b2yL6Eb1ucyRGD9edqt0dLRAYZy2ERBUgAjuu2/hrY+mYHmDTPde0+GA
j6RaGhyAgT87hw/ddzG4yoiNr8w8ajk6M4k+25OIAr6r37ol+4BE3ZzUeJRdoPLDPCU6Tv+buBy7
UCnhKZgmk/HbManT9DsEWtQ63NL0S/bM7gmMOZriUa/t0vUBELGS0yG9cEFMHqFksVfI/pmcyuJN
KH7F4+JmdI/swdS0UAxFNU3spsmHl3yUqUtXo+OQCV7CiB62/5DrEUMN+Zvs58tK0HxOiAQGE91k
KGCPmnLVK5GBSF7qogNnP0Uh/gp5Zq6cW+hz8Hzo6YDUyrBr+8WzMGtg68n2hUCl4Be/wmrAVtEo
6L0+n0WyAw9ZnLSNsq9PBa33TnJu8HqhC1b4B19H8BW3YMgEZ1bJz9LPCe+Fyq4G5zgV/DY4B8OY
fyhQF7fAsHKOoqWmY95CdFS47sZueYJwBl1hLn1cUj6g/cHCvTtBM/C+zE+97QnuOb7whAVeAx2D
KV6kGZl8DT8kOUmxUoFo9uyGljTpvfQhjwuUlVQctHmO90R4lgaWLWgjNukBhfOOfYZguHA3mdTq
l48qFBXikuQh8C8K8hcAbYbdfQbmFD8lVUoA+iV85hWhXF4jsf8mVfAF/HbXnxe3SF3iNoiQov8N
Utmvv7P4MyGG09AiYb2NbXlFh/1cXYFVgyOtZkWNpQqPq4L4OCtBr+AbH6TMKxk3de3VvDL7CVdY
feSXrwBJXa4zVhk1wUzuDrTmzm6ft+Q+l0Lx0dULHwy6q2JOCn/Z2nEr8n/bDXxd+HZEHLzXRCEN
o4LONTgmHltQfO39/xESx4NSf0U/7vdyNty+IQDCPY7N+yL/fUHAHoL+SzUoDArwSbjh11DZfTUT
NL/EpElsVC0EypWDMTUYB+vHeWpzafh0gwbnvWV6vNTyn8VF4NHQLNSfPmvgp94k0A6w0zt/fxdS
PAv89FsdeVfdKCJXz1QwKSemqyRkgThPBxpgnInGN775OLpuvA+9+pKW/XGV0GiOXJPVOOWuWpo1
rHoh2le/Jkjpq1dVSMbZCa4BzqaePLx/TFoA0wWi/aqw9kq9eqV2zKfr11oCML4OUgi00fCaAQkW
Yc8VeXtkPI67v+v6kG8oMd03DgVUelr9V51J4h9E+94w5fuCiQwmnjvCNB/B8IlIAYu7eoJBdfmb
o38w6c10mC/vM86a59oLSZGdHibPfl/ogJVvpkybJqANXsw6WfmN5oKaUjynTzmQmPB7F0FSsJYD
zSeV0AZCzpFNeQQawIHTiLGZ7Hc3Juxv5sm5/9V6BjaYq5YZT3u4LvQAouyGvFnbf5F+2QjCN1Z6
NYwOcBjc9OwP8A1dE6ZFP/kvnjpgTnRH5Ob8a2Zue5/t4KhqjwnpaFJwpCv6UPV3SEWtvLXwnqeP
7UxAGf+TQDVrk4UGmN/cvi/BidOtnjVR4825dPJPshIZyAxtrK+Q90wmeYZK7IbOTYtJuRyR4AiH
S+HJSJE3RyA+KxwjursO5On+Je7OSQo4IjhjFlQ/o02tU0lY0t84OeprOQmqcbyiwDNU94Bt34sw
+4e0fiZ1FJEO7RGyz6/4vptZcU3blb74HtkmsIrN3t4CCY0pzb0du3NdF1/JUEyu3Vm0WZuBZi+i
pQNrdyLRLVddfgA63OQvW7lNEn39q7qd4hX6nW87FB924yqSnMTaSek2QZQ2guslBE0/XpjyMVTe
ncrLdj6CzOu2kKDTvNiNi/fY5VS/LYJd4s4EnpCh7Rw1rLShGsUV59UAK5J898r4ijbNySG/U5vP
brBqVNi9pbQVWgvpjcWKsjaAvMygyKN30bjbJDJxZV0xXmQSzFA2xbAGykypJiotEgEOEnZOGxcH
bJ8su89Ln+QQJG3XwCHnT3ZAq6fFolBBgBvvEafZAo+wtWAmztXQWzdfNMbFETlF7ZWu/e6CWLIm
YbilbWqNKlwnqym1l2Y7qNeAA1uJgRr/+AsZVrfJakDenp1EGTqAE6YcgpkgE7KVEdkcPrv2c7co
k45jiwizqHItP/xdWI9IBiT36t4U/1GK1c7nW9aQjjPNCyLDiQBvBbiQX1yKedOigzVkJsxfbf24
VpAzUgCXLmSKDWO5Z3z4oyqMPOa6HiomS0FijRtuxL37fUKRH8dzuL7jue3icm7lF5YQ0G9dPY5J
ac3vqrdhW9BjnFwMG+Cdm/GapiCywqZ5YyAwO8eAS5Tw4A3HLHZW/+5IroAbPKLKHAEyfw0guBgx
Y/rdF7UjFnV1vx0t0Ikhf5EWzbIdcpmqfr0ol9DKCoAcOWe1cbmLc9tYKpAad/VDrn73kLOw0fd/
9IbU6ixIyzR8km5/ZHQSEVNzC21YQIrZ0Bixwpm3/kxsVq+SSoqW/n2aPzlLr10XqLNh6wHEUlXs
PZ56JGahMyhzf79aQC6y4XfaMJKhvnale3JjdghixN9sj1JLbT0H7NVDhus2ICt1tyaehKRmgasL
gwqzUBFsGpcd53n+Y3oIwNrwo6vveUgdmVLrRWco6pt4R8PTGy/5fSJzkUaXId1zS/0WTUXaLSUa
sS/n3nzua6csGJzPcPGk8zrLbEo2x4i/NmLRUjgSEjrQiiTjqG5+2+2KHtxNy4nVi/yranXEObOD
+/vM/SPdeObVxQ0zWDiSJbYd9FPXvoOCICP8BM2rC0E4dny5XKTU/tNLyz4aAi2XUxHJej5SgDya
mCXcT5P0zn76Jbgy5VhMN/J/2MMRc40cIrho2TgDwm7IQWyA636teUPaBbZ9slYAKcctq30O2LWV
2OfDuly8wJNxB4EJKxpsu6xWRHTg93NGr2OwiMuOVC4/GsKJIJeGJ6p12iDq/vFPVjP1PWIV7MEW
T4jfkc5JHnnMjpVTAqmkgo54QZ2ytlJEueZboivsitXYP7ZgFWRAMLL6F1VCKA+co6jsM0Spot+e
tFAv4LQTkxTdx3gjXCpE5b9onHV/GiG1oLMJYYKHh+Ytn23PYnYjpEYV+TwH1LoVuUL5Wtc3O9DO
Cr3FsflwL6aF3lrl7gnKZ8N8uT2ZpjJvUTRmwx0XwAQxl2KwGDY4fBBYNRLNcn1qQkHkcdUdvfNR
5PhF+xeHwjduIFJuF5yCxWcVxLhr7AW4/OZZYUSu1AaiAZ16IODhYsFhDSINV1l9tof3hblWuMu5
C5KKwC5H6dRlIPYWt2eRvaYh9A1zF+kbSD26ts3IYz2wy00J6vW8AkoNh02lXMLWz+yPV2KQ1xEq
3xIuqjlAuNiDvrb/diwwqBBDeezMpz53Zebbq4ItFpldirnRvJOcJPGnuaDCMdMitTCOpWfLWK6c
JyL7bdu47xthEptyBV84GSO/FJvhDPr6rOxYDrXn2DtNlbgeVCgANgafxCCaYtq11EuRGaxnG+bK
zZL/EqcntwJyykxr20zjtkuBHdd48nogwVhKGcU79+hGY6cDJpVplq69OYZfad14p/kIIx3cm4Gm
wmAZqcYr95zHiHbeHFix5cIPwM/t6SudERdJnIRV4/UAYlksNQO1vDSVGtE0hLKAHSZ8Ne0X8irG
yrUCQn7rozwHcKsp7Qq4bAPm47OplqHisz1LXMUD5KiSGm2g5sdwtCwXnRRqbLDEYdhp1Iiby/xN
VSDMhE696Mwf5HwHgpmsHZ34Z/iRl6I6/VU/uyKX2vioR/3wemE0b/3kDaYxSiIjzJ5AlzkXlh6S
VMCrKMyO8NXXhsJ7+OhvEyLKl7cOad5FiwujHNVlXcLT1Q2eryJpMO8QtWHkQlQchPBrthhFzt/4
VxDe8BhFoX2AfOnozDZFAhvPHO0ag4hszBgTrxz4jr+t6LmDPTkqURU2HvJ8csnvhk2dQ6dRvq/c
Z+YINDfAYmbBXLzWHNhnfnhNJKNZvGRRbzMFjJRQuVUn0Y7i4ckHIj+AtP0tINkTWj46EnTL98oT
qWaLht8rGfetI+WV3/17SCdK8jaDzLhSEPrKb1YyT15d+uVCLqRAYsWxswr2/rl6LXfrRU7H7Jqc
l07hJiV7sneTmVbBDYJ2g65F5iZ4CsoIpcEnt2hhwfsvn//6gANUnEKPVDoIna6t+SQFMLN+oxoC
Kek3YgbbOzQ7LfYuOyzGU4WP31ZHIZ4Jvvm808ZJOyXEqrG/YfjFFwLZor0LAJi2O9DWUWcLSuq+
UJ5bmuacczVLfE4EIagQDOhEC/VYojIgTyZelO/ImjE7AJVauqFW+NUTHYCw0kzmu4ocVV1cEbJK
N40Naup8uEIqXuBAS+cM+jKVnRqN3Ct4jw3doR0iikD6m8UCd1p9etLmMCCGLjbqv0LLSswNqnYG
k6ryoKpx7Rl2HmeKHCOvxzOXSx4rIGhEpgFgVA9jfrgXFWJpvs9cFT2GCupaR4rXNiAXR56k/3Gx
0Q5L3SKNEftcWYL0y1Yiinjr+UK7KJjIym6wT9mxNN5l9II0HUdTkIyRFZ/wGnz4hIPxed7w52+P
GUdxuPUaSNKxlf/SA+AsgpFg7d/FVRxzkpUbT4zTtZNNQIdm+UFHufOBP+f0GvRzvlxPUyuCoLls
2Nou4kOQXU+f2Of+6ozrQ1W4Anm5H1c02HuMHUtY682krOrO+cVQfw6GeL9kBRMEnNchVVJYbv73
QL5h9+ktz2sZhl7Mv2oUU0VOBWEL+H9Cysm0YBxYWB9Gw/XDgabBDSV0zo2/ZxBTKw2stzo46gmk
rD61t4iAwVvEvqNlRihF1pRJ5UdVN2Ea4/lA7LXNMr/bjAZosod87bVRr2PLKoZfLm8BbuareboF
0FawsRR3ve5QgHTUiP1JSLuIKXNwly7RYMp0y79pr6GPjDX/5J7k2uSM/fIzXKa/S/9GWMXf/2q/
TbHKvYrXupEpfW8UUnS9RnxiUegUZhfnP+pZkJp+tptIMP7/gZmGPBBTx4W0mIohTM4/eRkVf/i0
0adHwNAV/mZqrwWfbXggdMKROeLhc7EUvBW7S7NMyYfDmW1UM6ZdWl4dmerROeimuEfr4rfgcDp3
PuFvo0olP0/wvONedB9zOIw9GujDfU4HYjoJM3vFKWTWG1FWkM2tg+MwqHh0zak9oln2UbLtRuV5
NhK+zrIbV45I4vPRvv5Izs4EnQgd9t4uFshrkUFTbDxjkuVFY0zi7kjnq2W9TDxVz/n7tt8nNAQZ
ISiNwSpQjblCEWGVPchTUpaqePJhluLIMfBNCENuO1qVZXNXI8ZD3uepbffvHk1xP6e5PhwFVa8e
h42NqOhXjyjySHVi468j0tuSGHt1xImGriiy+aBV/nl2pJMicyVyL/8xRSTqz/41afdQgb0K6x7l
0MeD5cZt8wFj0GuwY6rzKwSUYxu+Hqgy893iWUfnqXYDJgZn4i9pyOHcWw4mcH/Mij9FKZBkUIUf
SXOsoy60ZRjZeXs0P04827p+njiX8mAD5MZKSp6GAR2sbA8za0fLpaIYrBYQLSTVYsnKzUQ8AnkW
eVQQo66DREpJN7oWZKtv74WbEuaFuDgD5R/GIQtiEIKzdCr2uLQ4As0Aj2Z/LDjZQfeDAmneaPlR
IB1LsYfNMBKhn+M0jOyt4PP8oTNNoQE28CYQR9F62VJM788gmdgraF4TeOwcTxSQ+GQGtBe3es8l
M8dieuhqV7nIJzOes+BJUsXgdTfa2lJgR6LnInD8+KVA3MDrmCqIlC6NsymDHSE8jkfKpcPYplWt
0P+h0/wa0wpGTu4sJmG/9zB94P4y8bUzTR7Vbe3JBGL+6DigFLeJZV3QgEp8kGPK6sZBS9j7RX5I
Cx0wAgbTXD08cAlKq7JYvt4UYyrdVd58CpVY0D7psL6aRzrSL1TTDVGYsiRMe1NugkxdQ5Yb/GPH
DYRurZoedM2gAp+sR4QW4eCeGF1p/R7NUGG6KzyarCLEGnNL/Hrdy3pZcOwYz+683r0S/QbSVXfa
o3JT1o0GuZXNkAGd1maPlQSwiWH8OgB781hnS7ulbmezzzVDm5gtNVNgjCv+gz6o3+K0c8MPS0Xw
qGasqGYY+JnOb95ssDR1o8CjL2I+s3PmalEN+r4TkPpDq4K22k0xZKJ2GMmMZfBOIKSINcWmwWsl
RBR4dHaRAsoXiBiJ3IkZBO1p0xuysD625KFoW4kyfy2ALmn6I0AqrJrmXw+2SO8x0jA9vFayw0Iq
LmlwSTCRttFAaiIagjcXxOClBY7te4b7jf5NPMviD8VQlL4oB3wLoOgmNj3QNif26tljn5nnv6H3
a8bkclPsHD9fG4qMDPrWnNCl2WFG3ZM0LPqqWYI2FEkT5yVpqsu3FPTKHWHz05AU7FmXW5Kz6D40
TSgFs/3/oYkJKLhQYMTIQrgDO5txdqQ+p65wLTIkE+CCDTgvTh3AQb3+JtC/nKRevr3ZkyxE2G3e
eh7/Yl/zYzlmfigkHp7VgHnTz1nw2Ylexah5MBXj9dJABNWloYXamT+Da4IeLj9xoOnLDzPshOBq
/xZQiaaVEe7C8GY4sQwNS+pJr7OWkeL9oBEoM68FvIX0609kIKDXHuM1YZMdpxPmllWYLHHyzUur
s1w4wvcFnEBIIJWWNNPwI5NO41sxObaeMthsk1cRBzGAFZ+KCb0ojFFO03a8mYa4gsdP0TWbi6m6
QaXZPoksFBAjTQBxe/Olk3N+pklKiOxB2c34nUq2qDM3YgrVg5EIldx040xlXSOpKZ81Oi55SMui
pK9XDcgvUcLLXToD9ARQ/1ShunDwfQ1PQfTYn9cTik4jGK2+ORdmgeqFOCYIOaF5sMk765qUb9/7
Qxjms+obJKGpkk0n4svbDeIDK3Ws7A6hfmFc4V3/MjFip4kMnKzGvV8rKYZDsxUPOTTULdz4Cswx
/DP9vlh1nvY+v2FGvNOmnF+QTFpoqbAQPE7gdKaHvDoan/x6N8rUdCzPkqtI88umlTP2sodohtnX
yyuX9I9B/GrULVs+JkYjuhup/2P2NJqs5nTTqb6ZIxTrlrEHsiMNTG0b0WcwiSqCa+bybU/uC0IO
XmPUmJ0Z3hvFFeOzVXUG7z1dho3qfQS22HQqBibFeGxAWU+kXdRMtlAiyDF1+qAnX440CHNimXyH
aUqOwWPbTwPa4pIoNFnZkDj6kNRnT+Q57jDY9DCIn8efS0Gy4IUGTI7FGtgSel3KlfRaeFKSLbDJ
77PQZrYHE9Fdj6rs4u4aVszNCDrV2RgWzNGka1jq6+ga0fyrB8FJwZ+ctcLAqTSW2lG6eQ1yhCVH
5WegBVfc4gZK1BrTn43IRoQNVb6avLWZ94uPQ1wa9+iaFVUtO/rpHi/M168AItSj4rY6bBUldLMQ
VVjsWhClGGpJ9fEpdjzEpozZST7rZ/45gezYv2O558KWsnFkjKJ5JteBTxQIbQZBby6XI0djlqa6
Au0AVVgsaFG5oFpkyPMoJVYDM/a/07hTEGLHjHqdOdA9oNN0kHD0uh54PJ+i/XYeSFhomZWScvoy
3DDSx1M8RXmllTuEJGlUHXhMfy/sqoANdD5jdxuaZpp5xn3IvJMIJe0Nq9+l1SAbPUdaj2+Yf19i
vyCmtoKzD/HM1VqMLQ1GyRtwXIa76jCB6JUjoAomoFTz+pmWrvCCxZIsSXBIqEosV3LPvUdqazRl
i//BZGcV3uxtepA8238Q1DUddednDoXHL5B4ZcNNS+fLe9t4IOvguoqeARKtxbN+EjTFzB9TkrWV
EWfNjTrhTgYrUnQxQNUgUxQDd1F5yHp5/LdUjVUK66lYy5QKMerodD9H0hRH/JwoXFdjIjUz/nEl
CZqAFIZl6pFeZPe9dum06fNvU9pb7jShoKD4sgrIZWZ/ZdWFnDCYKN1EKMfOv4MayrG8IU7UsakP
xQ7PRrpSvhMBKHQtL7JsuNWZop83bGYxN5dKSrjIrsJhIlS3VXFDBhEPRgO8jdu0srFYA3hRkmE+
MxDSBnRF4Mlf2wBJFdYjjLQBQRkbz6/yfPSHCjw68ld7VB0nyF5Gl0UJCBQ7x7FEZ8OSc82eGb39
FIFotLw7YvDDq6B/bJorzYOFO3JXwtSyQ+GY8Z8Ve7RMZurDoQaM5Zo50hvKfk4u0LqrNDRZFMO0
KYQKbIimGNQmT+FBZOH/SFqDdtIm4Jhde//ypROW5ukJjbCoVenzwOjbEM1BqKth46IIm7xHHb7d
Woy4cJp9VQe2saBi950ufkA8ZlCCDypIi+fqdu53njOYsaLfU2Rg7tWQml12RXedKYDBKiVn8RR0
29KTBpYOP+dKIoAzGhYDI57SDlXlH6iAlIaiYCdVBDbdW2PXJpDIYpyEendWxmJVYWOftxflAk0Z
kvi9eTLVkmKtgVI5T1QWZ/ynKWJyV8MxM6+QHb2yDo/pHU3jZTwGTre1Yybg8ljUrVygZmKbSeWQ
rhbkAUDuB+I7pSClSkAj7UO5g8mRyYR4JIo9pSUqXbY+b/FJYqCtltZlV8E2r5/ZZrvYoMkW3Yhf
o+qPIbseq5LuG6/CiVMeWXfCv/9bfn4I0tu4bagZgoPzst5OCnhnM0hI1s376WzTaTNHeyrnZedp
0nVsvX0BYx+BAiAuYVarJ2FqR58FRlFF0MFZfH0pnC8KAVEY+Bt+FM0BMFt79CudpWe0IdiOFkAb
1n+Hg3TCZQIDNxONplOpg01h2oLlxB7F6HCwc16dEgiEfDzZTBTpVEAbq7PvYUM0EWpiPM3MMbcS
oLjP2rb20XlAnUSFQUbK11GnhBxDojhua0/lDVHGJpq0oaI8PhZV9QSk6uUu6R4a5YJ2Ol7kZmIQ
YQNEgHSTgIXR7d+kDl05pPqt1rJDfxGBj4gqzXGllashK0+JRjWUBvogc3enO9y25zG+j17mZxD4
qblab11tf8XfjTqpTgtbtH5rlX1gkhmbq2p10deLYTopfxvxezMO6uzooRr3lQfrRDPDPu37g2Dl
SMfG5kWT8d+/2EKOX6jxk4yl5aAbujkSaVgZyI/mUpZxQBui86s/rvTFv6rXbCvN9po0fnLLsBlb
w/JjPgoS0tkZDj7bxDV9BDjpXXqzZlS2Oz1pfyu5QTLuBgwBVk/BB8gihtsQNuIIPylQifcI3UZj
ycHpCfbKPDmtBalVhCti1dqrqS4RyrVisrakGIMb2a+4RwqTRBBlC0nSXEucva20Cpw7EeSN8ZIp
BDHrSvD/E9izLvhokUlzX5T8Q55XPZGmDa4vzwCDrcFnOfiv7VcmZB9RfRxEJ/Z0pJfHtdNu872s
lHG6zQCrcmrbdUorqO/s2KiGGcPGl321ZeU2kvlRAlgzc5TdUTQdPpfjGNvB2CKxZ54ypx9ddqJI
I1IGY9dqSz6jfddmWkK3qOB+y9pgUYfHSqgSLU6Y2ibTOCWpr0RQRUt9Duu/SzBeIKvL6Bvpk3Lp
e5hBb8q7siDrlN/5hj3qIoXQT2eRP1ro+h+Nll1S6ZtRD+EtmDl7RSa4C6n2iF3/Y2ERbueZ2agk
D0iWeM7CSzDBJhiIF4sy82pZJJXRtVSQh8Rmgj4GRJXuf65kPUDlsgTSr22A4y8kxBKZqqCfI+oj
63mPJ4eZ0oZxv4SYLI/whkoRXIVLCWDPKLg7U33DqRmgjdNyVC15w4HaB7I1MKPMWL53NaDSu9Yq
vndv/0UiAftl8pu6ww12BhPQtYaZXbsyg7vXhE8AcJ4QhOBgHHaKCWRstqUWRSjmAceAKpERpe15
9rtRFwXWeyXXUJ7Q9C3XFU/hTzQ1rYm+LFvcumF9hKIJ4wtINPPWmmHoEFo3ILQdlH/KjoSe3oEH
qQSBCMKh+4RCowoeYO50Ut1D7cNbwx22Lyrx/5mt2Fdkqbiq6e1Rnv+3BxpWQtVP8OQy0bBk4Q7t
+19sBuPNX+6ng5GPxnMDiUaXWjxybbegXsSMU2ayVGXIwBoqjZiplMEl9f4u/se5aQ9417CDGdKo
b8A7xS9eiZAbUJtZBqPN2mQ280EBblOh96qAHp8GxLPUqUAlCIr2qOwsBQ17rIeUBaMc8KkUJlWd
t5DTTRW34aJP+uZVxgaSgQId8aF7weK9MHoNWEZzOx4QfMCQXdgzBKi8HHKnwoNf8hnQEi9QhblO
vPePR5MpXyOc12ZY9jdgt6k4dnJWiZRa6jx7SyK6OvdZlEjCZkQBaXc0JEb5n6RTnMsDKIyc2QlP
/X852SvOtQtuLu8QS1VNZBFMNrGBmPTqGDugqnYN5cHB5BfF9kBs+ELK60TCR2a/fCXBqytsHm2b
5ccL3rO2GDIecdkN80qKP6mCKswdPHwFl6kTcAMLVPtiqRg4t/iJxTyb0p+ePCUJKhA3FyZQviif
b65qM463JVznUlG/t08AIW7asps2q9sDmfA0VUPsnfMTLcEFgyKDyg91dzCU4S/ZPvOYE6DV7M5/
oxGIThT2w2erQilJxKvAf566yWe6GOjMMSZegp4b4W5gnOip7ZkqmT8tXDCSdpQsh1yUJ16ntS7X
gk3OUFdR06+0Xkf981pw6U58m9VCaymLyHSziOM2wjt5LtBlJ/5MCMNT/4btQJ7WNR7Zd3tpmPIg
w0vPp9l36NptxaUzqk+nYUxyRIAlY0fthFIWStcporCzROyAAZNSsM3r09CSDgKJpU59BDcfCkl6
e0if14GCgPh6w6W8Punq1GqY45USSLAIF+DGxnvuAd0mbOmJjB1DjKXXDY1n1X6FHIokqg5sr9EE
UEb+mAsaQFfHDThb5LHQtXwMtbzi+GbLWDSNpiipIvMvDhzNPe817cwX8PTsSude3kspnpbrwtQR
W0r+tzNUEaZrzujkAAeyJCh8cSzcBoo33/AI0x+/spTwUUVn6pTpHUGDHF7ATtouOZ5+O4+gNNvx
bXET6XCiGi1sDU6gA8svOuzGPHHqtfJt4+RB9bix+FJwIyz3R967m0niw+Wt9TwL5/1O3m0sPyHi
S8VqkCS102GNKY1hWAUdPjKPb0eFAi21EWTojVbCB9HKjbaE/wIJGv7AB1S9621ZMmAL8ScfcZ2l
JX8TsWnMDhQNBfuKInaLzaom2ualwK2OF7EOFH9YnSZBIh9+pVXOy/jmkbthbsGJi7K4bxP5fgn7
b9hP/d4LZtitsz0cirYM63TqEIt0N3yiuvQvT5jCwEhy8Lxu7po5LnNNyV+q5zDXdgNh9sD76Fp1
xNPbk4N08mcbfqU+HeoiuF57zHW2C++zV1wr7LSQ5eYt3nK0uDEqkc12WGcw2stpNhzbidaMr5PT
3ci527ReMwUjmyHNthPbd8QC+SQ2up6dgJHGGXgtP2FrNghs/GZf+zxhUxo/6Kf2uK0FT5g8k9+O
AMUMabPphiQkv4vTRy5Lh+/kJhM5/S3ipC7vfcdNMn6tXxqcMQeSmR+y2hkq74Nwn9MjKvYSmB+E
uqa4g3pJuuqncy+hFHo8DvwFyRjlpR/BrhLgIMxvB6iGehnHh2mUtoABhQjLsLbkAMkEDIOo97kA
m09hDf3eGc/lPch1u4Josyv6MVfgA3lwS74gbzqrLNDj75iq7qR5V1gbO2kfPkAVk0OdAgRiFEQc
AGBIhPayFHwD0pvdn2EDSZNqMvFqOdjgZ+HJUZVQ64CwVpXqVCC+VBodqQKIs+vDdOFwNoDOQ6O6
yxMQl+cSnJZHQI0eWhcg4wX0Er+izHiYe0wH9LcDbXwdtQpeJVPePhf7Pa8SwuNgZyKVgbnVBKZ9
RnzeHqop1u2bPAtbqvFP8Zid1TEdSvR8z1dwjy43/dxGpf4MZLeMELcRCSuyEEU/oWwdNzLaZJmL
j9LkN1vnqryqLCoBbyuvCcq/vWmKIGYEs4m+BiSb75S/7Cgx3z0HnxvVZYijHtSeuQtL8En2Q75e
U2NPHTOl9qj55ORK5/5LUI9R0fsfzXR4aQUyl17klCqK8N+GYjJz+hzatKmwbgm/B6bmKBunT1yT
aTtQPiFWVOXB71CtiZHTMEEP8i3m7J5c0CcdUsVSShejiT3scCrT+d9aIkx/zZRfB/y5S9QnVBPJ
wn6Rj0FKW8duji79v82CIA5/haTcXhLZACyk7V2c+VmxzgZzSUN20R/Mc071whBq2hubFMWLija9
8Y2ygVCPiogeGvW/GIzGQI3wJ40DY9t6SGL0FShoFPap6rWl3WZ8GZwhfQ6SUtp3xY9l/kw+J2aW
fZkytuBmSURpewVsioWr9QEEW6Hpqhwo+/pQrc6niXsABToyK4IKNXAcWi1Ze7r86Mntnho/NeyU
6flMJmH9LgxIqNFQwYL06uYLvFcxp+oNsiAGV4ZLhGHU1Gjl09f/TEu/ZM3OM1QFWKfb6KIKVR6L
rmrqfnhukn56PL8H7Ouily5zzMBlg85v+OO1e8AIOLLMbCQM00xccWlQ6H5MwjbuAw2YQ9EcJz7U
0EuCoVcEtxRUPscr7gJmHHXeDtqO1F6AxrrIjOs04It0o/63p9zD23Ew+XDY1CpuNUxVDyCCoNj0
k/vkaAJCin5r7KY0O4lumjXIvErBHBeILkF3y1GUgtHHZYPBlvW8gJDfEC38VbOtsN0Acr/zNJP4
bJ/CeLHCRNmGTq1vOxjMXaBkmq43CkAOugoECMRMIu6ljGNRkWYDBfJ4xUiRB75cbXLXyMd4MjQe
EtNKux3mt3wDJQNx9V5tK9AY5dTjM+gpGuj2uuM1UKiY+Rw38cUS+jimU6K9Y0Qonx96lsRifzBQ
O21MRDGuPQniLJXvxmriG1MN4i3lmpjRiVMEEpwzqHG1wWaMSOs8tPaNHHogeNU53Rbbcz8Dhx5k
o9jkmR0jP3qR8NUu9wxQpvzLrlp+VOo8wMq2WCvgnlJHtqkqqr5ax+m0PTIDvOhN22fq/D9XyrMY
RZrLL9l3oyfXFbhA0+9gD0XjDrYeiWdR+Vzmh+92FyZ0nblCfBgdqslgSZ4rO+ZJqkGE7LVcISUW
CgYKK2MDOA+7qFaTctAsGtwF5Dk+weXwHzkUi1HnA6lJ5Z1yjYGyfkZalQ4cM80kg4Wpqez27aBj
+jl3eU9lUccIwbB+rdol2oi01jfOrxXwCfgPaAoqtU6HBLaWSIzqYCxi25UShHwXPBpQFLpyLIpC
JTlKBfVt+9KSGbPCAV3Cekjbnkwmu3cez/2afIyp+Dcuegdr1jaewCl8ihjnjWo9fmrJjQptEOxv
EXyg75ray//LhYwtB1QEpcQ4VAxEyzaHrVRd/P+Xro/ZXWYk4pZFZstEk9SP2qs4UHsnBt4+NmkM
Fa/luwKM1jT1bbJ8dDQsciv7F9kyI7mB2ck6HxleLnl2RKvYnozDzyUWURGSFtsUg875g/JzRXJ+
tAbwU0OmWiL+ur+VnfisZ5Xa40vUk1FvvayWLNZWtoFJ72DHmZyzcMCvzQQUZ0lSem8o75WBV9fu
jtdstABU7Q3Byo6sICWkYnTEUI22VNtQxqb5RB/4jKEbN3gprYwpwg8rubkvnieike4zr8SYCePZ
WV2lH4nqhQqhZ1Puu2/QYaGp5S5VAcqdXT2r3MX3dz87fbeEKoJfa7yWPsOF9tqFViTAvvlmt9Pl
ojv24OW+UpfwR/dc/rTWA1UGYtDGS/FsMIwNWcF96ucnNhqg8xG8NprnUdUzyFktYJvYfstCwZbY
aCevP0bwPRuIy1CydIsYRSkWK++pGX9aaq2F6akHMF3gAXkyBYhiI+rvOLn1gOaitFZL7FGseQsU
j9IRMvLBS509eUQqOk4js4kQdnXTXiBOlomLEZXcpNhVBFt6xtwQjJwdZNabORV5ZtWAQ7VL6j28
G3DDPR4kYoMfd5Rp5fF7S28eo9UNqjiSSBNSIJtZVqYsTcvV4Y5n8P7ZSa/u06XDpYfgKHuNzNWW
2EnovcuRy8HTq6xKepTi1ZYsZI2QyB5bE+hQUdpoUxaWyuDZPR2o052/GS9HfoxcKFTsIopqEFxM
8SMtdUz39uhQaAcBXcrhVaflkHqIeas8KO929WvhlsoJFFDDUWPrq8I6uuGrkcYgGFITkJsEePPn
5Pak/8KJ5e92ASSK/Z7WoUuIcyxzI5lOkk4bAJwMQLIheOuos5G0DDFJVRKdzSTYUw2p9qLDH4QD
ME+DuxwSh01Sx5cx1uPGyVbYxZ1U1s4ICAr+1jC5sqzFXr1WSqHggMbS7ekBgndxbDsjh7m/pNio
uwYWHHkVJKzWFf9DiCost/dhjfDp6EVWCIgbQvg9AM088sA9xPgCb3NqSoiUSLAIjiKE1ussVkve
UBbCQYjKXHwmHk0zJ07V2NgAij/P0BWS+JYYG9P5rOA3A6yuwCnzFBfhYLlx361iUS3gctlhx0Wy
dVwMK4CjJUtIWnQDS5OwtSZsfE/lL4UaQsXVHvCB6X7VIPyBHZMmaxjnVUI6ZZ9ajqzbKyAOCotQ
Lw0QvXVPESfqHB3ivV8Wy8LQM1E0DjP4Hzr+/us0O4I3gKvKs6uO+dgWyQnEZdOrIbvhc/nUHEGV
FABplpO/iPYklSWFC2S6LFA9eRBwKwgQ0BNqJJIMjwBzYSSC84uYchdoNzCYsjQZU9GcnrcgGwsN
2azed6vPibcbktouXx9jIyBC7uMopUO418KW3yAhoeuHyQRbxSKWsnpiszzOtSErHK0lQo2g6N7E
zT4P51G3A/TuQ9VHw3m2DLyPgeBtT8WKBkJxou8Q2aJsu6Mena8JDwOJsF4Fh2ZF3s5AWizlyDdP
sGPnCZUgw9RAcX4azNzXdterKp5YL/2TR1dYV5vGyuS9WaOgoOVPujP0k/cB0Uuv3zmqjqoaxvqP
foR3f0lhQK1Q+TcdMnHNZAnn4rPESxKsciRHRDeWrmDbhHo2j1ZTZkDDzZE7vr5SlK7dTxOMKdvO
ruiRIao830IVckYa+Y//bUTgjUXMmWZ0fE/09SszfjAbTnAZv7ut7d3LBSfYIDgxsNQAAFyMlgyX
rXCYs+2mZAoZvFxEQstYuX0K3Qu6S/pAlpAUm8lPqXFkc0NxW0+++aOsOHGDlzFBeyL5hjKU35FF
ekplfDtK6aatjhhFrCt8asb8ouiSK73/nOI0ILjZGTA36kwWDvXyk2mLTnKuMTG8/CYgZQLrz+fE
+ljVkxT1golVWVwD+IvxeHPOPffvU92mZONRp8xYi8qrukxskpgkknmrmOCpAeaPPQLnLFHLz4+O
/3IzzazRvoxB6AgRdZs5FHhNreDYNr/41mEPbVROAytLoBBjsWHjBl0f1yPlOmdS90h6R4FBoxDb
P7MB/Z3xCngVE8742ChJEkl++CddurC0ZwSEBuz+frxO2Dn3EswNaVdnMEo8TA0wptl2ciOUQ67D
Zc0Pp0yFZe+vn0lEpq0YdKIrQeBsB+ZF0OC4nxZ+G11eywClDyXJhgu9ESLXzkAbhT3Biq4Pm3U6
6a2Ro1Zy/sSlAQ6ejoF8pNytNPt2CDLJTJX0Gpan17uoj52I6VoQZDpjZ7P5QZ4vVDurY0zetAhu
kOF9YVumCQkAdweQn41W70mALy6xIsUjiCG73NNM6/9hgJmnWtckyK9g82L+nQpR8bPv499ZREso
HqpWoRbBA9lU9pIYT8oVO30BDRD71HqOplaO4EZuCr7nG/28MVQtshWwTmcH2WWEYNH8E9MorBFc
Ot82c5NHGbJD3zltcCjbPjjnRBM1aoFqwHlSg/YhoKdlfcEq1KMPNvKL7dj2GMJE6SoESO8Mo3Bn
lDePvIxjdnhHtFbipzz3ICZYXhRhDpQ215eycygTd0DwOXqK/HgXBEN/nG6E0iLXrnD12rJBYyK0
xNUDZVARxEzq7TFiorkRM4b4EmmZskPfJVtK6bEdT/Dmp3m2ZQlpniZ9y4NDBjVwVzfKkGsUN4zf
wUoxpXsoBk9MCx7b/DNbkZ08xLiQ1jzP0f/iDxzXHL8vHMt6lkM547R1J5n03oBR74UcyIjFEXPy
jkr1lklSdUDy12Pgfq7hJ5OeISrO0bIfPfuKyLNrpskJNQRBVEs337kLOqmdkeckArgb2US1tfMW
JDkAegMaJ/C9y18HWiIamrHiX7Enwvl2UOB4k6TgJ8L1VWn1Bh9k2f2XI+w/DdixhRBPsT33S+Ne
WEJW2/pIg/AaQ+QGADAUTM6SgBQBR0EkttERWnDcKqo+2p3zhFxQvuBnY03JKtFBNTOzhoX6Ev4F
ZyIfTMhgOmlnJcg8bhlmVScX+/KlM3Wx4SX32yGlGneQmaPK+ETyJk1StBVd6KaXU9Ks1AFKYQEV
UQsUm0gknlK6Z6m28cf5cmj8SwgTOFfghPJ1k9urE+CHVKLA7FeJ/i/WuERvINtUVs5QP3tQ3W9u
0zl0Uy3SjKzq5vn3qJCp8AENk4FdCPrCtiiXfrepkvHjubTiSPERmrxnwi/tZvc3/9YA09uJdtSs
fr/e+xESjSH2g/z3AhECs3RMx6zq609oeYsitx+/riZu2DiCT/VMmGYybW2HBqrI6OueT9tvI0v4
E3mm5+9fsDHawAjvZK/oPink1E3gLci+1Ggr62ZQjo8fLvb/1p2hhYC5VZzPM8yAkK0YJRI5GecB
/oEi16AFKyIw4IcqOtgnUyD1WRqDKm8x3mjG5L5HpUvjULpyl2XRch7zEs++nEJHOjQ6ClIOgiew
Xw6pk4qrenvxbjrucFU57Ploj840u4xf8QEMBJbxcM2mFWhs5mgUJNCb56Rf1vBgu+0LW/BWLjTz
Advgdnd3wzyZHMW+FiK34RcCylqs1KXGOgJ5KX0gEFBC8GdqptfDMrDNIcFBHbFROACNPYHdM7pR
bPq1oJXdId31nd2K4f2bpT6Pgqwi+N0ccWptgVPBXsrIZLvL895YH6TXafMB7pMg5aIRkYxWVKgU
SVlz5UkaPHllvGKvl3waaxjNb8FvS9SQ1U8HYUbe0aFyL5X+uJKHcTHWOrGPcCcsjHviIxmrnZ6w
rnYQYEbWX//iiukiHDWx20fYtfTDtz4I+98gtsCzzv//8vIfKKkSpas1wEcB6nRhHVJFj/1Gj9+s
dbbvQTB3/qjkjKUq220FUBhCQ+KqPW8dVmqjyUDSHU9CzYQvKgt6DV16wUFXt3Q+j8KRs6hwVwj1
VYkrtCtqJAknlPWsl2srUd26cT6wPw0LCqWV3nzlVSwwOuhICzcvTo5RDZm2259FvtU44ylJcdOP
lgldqvxRntM35Dr3/dN+2JSghTqKUjI9bOdAJujp8lb2rbY+F5vQ1xvMX/k4CHT2+j5bZKjVvqz7
itjhQ7Qjerg4581VIjM0GdzywOt4rOIxZCwauaWi/zkHXDFn4xa8Ft1j1A7kF1UrZhkL1OplFwkl
UbzIKdn7HnxM8ywOMukd2QJWQCvL98OdNhHJzeZGsz8kHtu8gY6KFELY7H6VYp4Ron3yc5a3sbj2
IFv6nxVrhI9eUJ6KgtgSQoIo+wJFDfqXoBifdsTcjnYbuknDqShZtiCX+9olFTjoxKKXPutFu2Qa
MqO7WEOTBCUHBDJNpgrZuKLwnqY2uC6ofe4py5haSSMuW2atzw9N4V7mNtR85aaf93eKtWVyliz5
GDRhHPVSuf6AgcPZj2uIGTMy2CA5d9f84K/lMiZs8MaNbFFA0BmvyD+OG2F3XDFcC5p11n8l024Z
MWJfx9rzrYw8UxW32oD1/JOKnolNB3rI46EL/P651i0M2UI5Vmp1dteaLnt2rxneTef5gaPJQ5/r
EAmh2p0iSz7kIva2+b7PsEGLU2cAQGyxbxFt6SP3HPhPem62wXqUW/la7U0uxyVpiSLhxwtqsn3P
7YFZ9/e3wBYg2/UjqS8YDpGykiKgAGFGL8uAsN4K62jXkNOJtFbcDjgk2kbou9EhPPMA2Q2I05qU
rFlRuksPKSiOwm6THUzf+cKbJjY6n89gkzU681wZ2Yjr5t7Ayy1tn85G/cqK1/HqxHTLzZmWoDHD
1ctR01HMu5oWb9PGkT3k4CCsXHDV7ify1ea4vJIYNu5Km+orBRKuQp4doWYsg5TWkbLIN/d0UhMc
7uWdRP+jh2XRU9zVTPoK584TJ/Sw0M4nO+yV7JqU0vjsIWI9xsir4xrEURoISBy8ePIk72fTkiA6
VIqah3Mcca7TBuKlZ7kHqJFcj+5qwQvuEKoh6KIBbDLdYH8wWsVPD8ZK+dTDOrbhXbcjwPLNpP4H
Rx0bc4mDWQRMHatpN441fvbCP4K/n0eZhUE2J6wFAGDebaBAHxKg7kb7gaEJ6ci2BrnfVTAsOypU
Nw4NnCobpNIAJlYK6qIefUktK0waLKEZ9/RwZWHjkEk86sVnGNpi80fnoP2/4MYmlOu12DMIyHcM
XUPjmZVCoCKBRABr23OYJ3+EwzVTVsWKbT9TBr4Mz8KthE/0roM6765dsJhnbnxLhgiF1PrBU00g
FCKABINfGeoI7ghG9Tn0YvxR4rJUPn+tTzeD7Hw5nw4Zbn+sedicSHGyv3FRITQ/WB2goYgyjVgx
LcHbrten7pt8J40Rn6ZTQjKb6VsA6fmEAZZlc5N4le0YQ5f2dizSco40wQPE4vF8ELI/TFeTHZSH
dPvJwDfBrBY2J9CD7F2Ko3qGfL57LZUMl5uFAI05vAFMUfWXntscGANpeGUbKJq/hn+pt3FJ7RC4
veLh+xAKdM8x2m65NL7Xc+WLLeaggid9h1xf3uTO99laXMTsEnG+B7v8BoXI4bDIO1KaDumegbJx
Koinb4YYxxV24eqKxMOSx9b5VHsXfnjLEVoKXKnU+mGVbluoy36VYjfe+dphYfFZEpFS0dUMym3g
rL3ZfqBjfgHbgTIPbYJq6PGUHVUhtd0nwjaLQ9woSiSZsNMCZpKInZKEvJJzWf9MF+Qe3/4rdB/V
n6KqIMHqZ5WfVNG8M1sms2CC5+24JZGruCkPLXs3femIiIqj3XJ+jU0J627TJ/UUFJy0xv83T2yZ
DX+dBxvbuacN+hfaqneVNGUTuezdqrOgMONCR3aPGlXAQCL4NTc+bov9o16rB9ZuLtdCvPp/dskl
/o+r5OCFXkpy8jKwvFmg6cwn9FnvmRuDicWHmSEJ4a0WU+59RQpHegLeb+c81ge+QLuuzeZ99KNa
8BW3JKfPpA/gua53DBnNZ8PvXe9tOg7KLRvp//jlrAEFoPdhavIFDsDfjawKXhfablquH4/UxkpD
lInNuaTTLaoVKUVSGKbPzYtqjLkmnqrayKii1XaIDuUD2zqenXsUzRVAtM537JO26UmnxEaLmgLH
Y6FXaQr7QP8pNRa2/1UxwV7IGgJITwbKUz720e9isQ0nTa44ttOpi0FdOnmQMzr2yFNwhxVqhZbv
DnWXVp2Kljh0+joSrzPwPHgOb/jsxrDIgDXh5RmSPq7XCS9nM/8jZ6RLg/Q7K6IJ8xgvDM3nPyYM
Ys4CuLUxqCfs1n692QUVR3AaJa4eSCsQkx/9aDzuKFZJ7zFI4n+FMh9Uyj9LMBstBRef1uDJIBhx
LkWKVLh3dxLZfnm8sUqiJbYtb1onWfTX54Zrg1BPH2+CzgMpeZvv/v+Faqg5c0pzC9kwBvm7/4N5
3eJWvrdf0RqrtlDEK8+hlW0Ig4/I7soa3Zd7VN9/cvsXZov7j6A6FUgQLq2gcPDMrIz98C3IWQMl
+U0STWUU1P5CiGeRFHnp+S6Ya6BL86JFxyr8NfOhrijAFs8z8ppoRRsZApOKFrJqTtr0lWXMwnt5
33C3eX2eWTrALsWbGFV76NP1x1AyXOPymobDEjuVU0XL9HoiMrqrNKL+hltg/dXHCrjNT0cVI1RI
KAtCetzNEwWbaddPM30yIQPsVWtexWHTcRTZuC2DNCvs3B1tLQcwOpmSki+tKSsRyaLJAnsKMsqw
Tf1z/R9vxbPM+fPsFT5SnD+HL+FsPxyVrrlsPQQ75VJlfhoPLuFarxVCSiSUSPKV+zNe9Q+DSi0C
jl+Svw5cd3oflYqJOhKDiMqtCUEZXJ0POHxE4qfY93seyXuUWkhRYu9bUA5kWsyn1WQTyHsga15/
iuYOMZoqD/5BExgZcyjXsfKhHkpqQHw1qQFhzPEqdLyJlXva6TwIwUObMi4dJ8RNrnlD5CdlQc9q
b5CdcKhBLzpu1sVBloUtkQAEaCmt4duVnUq0x7ndGhjysKPm+iQd4mxrFu+/Dj0WEyoM3e88C6SA
hFvCRh4AfNipbOHwfNfc05vr/huNQqoHKWwVEXsz8EHsMuu92uOc+j/gWK+Kz5e/wsHfZWaEXQ04
xbk/3+7w1qOWlVY3JOEK8YN+TiXrqCUgegQkaoip0G4ygaxVMEbDw2EmwoO/S3DA6k0WZUmNRxlg
QT0inwlwJenZs+AaRX19/f+AVQ8oMrCCmVzC4HiFsyQ+jzd5aalGGGXfKI6KzxkMSPZoxJd+myy+
4INgB9xAguYCbawe1Am6JWreQBsEzF6JembtJHzV2tmHf0qbQx/xm/eny+9Xf5d5bew2tCOq4n7z
UiyJjDqcScCfy6v2KmXlscZq1UHAf+CIMtJpN5rV8X3J3rOwIBIO3J+JoXM+mbgCCCovZfpLQuCp
A2m728PdGt+cQX7w0STjIaR1r5yFHVUP01JUeEXp9YJyIUDZuKygx9lfZNymtdKSavFzaBxH7zru
Uc/R0XPUfkiialBAJ3Xt6L7edhqhGcDwHgNufENUvmh+0C8EG1xgc0JRIuFj9sotSnuKaqxvgKi7
+OCGp3fxSDNAEDQ7WQ2NbxyMgdtU4Vgrue2aSvBqWMCKVMCkMDe02TRU8d5N0Jrp2fNRXhkFjC/e
DQnYg3B+yC4Fq2nfD2sGRWwnAEkCdQi4AVfeYSgUhe8b+47hVWtsXH5n5g+ZnWo9a/DMDOO8jw83
GbBZ+xn51Y+wKXtP+KmaarbBlOOZivrsVVHNbe4WlD7IZ0Q8xmfxscSbpyjcxi2944pwzeTKOTY9
XJETC1X9m5tsynDra3HFEKruxO+XvPWxtKBei5EerEp/GD1ylg53y/0w8JtiDloJmu7CeSc+phwI
xqFrWjjHk/PIV+T39nXwa+wH1FQBPDcKouS+GmWbAyJShuewEJ3GXZdhNd8pudo8A99Z39ieYpMC
YajYdHtN4FcSEhUoIlpwM25Gh+MxVuhBTZ+0rG0Z+TLwWLwLJqCu2jYgHzOmvVbir5BD7fN6YI5+
jcx1jFWDPDB9Wbh6fJ+LhYu7kNOuDqBzvcca98l23egI5ZjDE5HdH/R0qHaNhbzNVP6VS6SE3M8x
y183KhXa/rUNtMiv4RG1PVGu7fNN7aJ8QqunWfb2iJDYlIySaCqzf8lj5H8fr0zDryKJFT/azY6Q
jqKH7ik6jbxr/avWcmssL2WgqRkI+YbwyXmOZTs6dU4ekhGxH9+y49rxEmZQGBwg9gU1qegy/kJ4
p0tPC/Q6I4Gj3MTGZehCgQkD96pX1KhIitrMJJB+ZustVo8tHzbklHmxnCVCJQ+zHcp0xiLpsHg8
AVHsr+GIWflL+hOQkwj7NRG24k4Qu82eSre4bluUlYwYxkDTEh97rqFolpPxrkGAogmiW3M/tt/r
uInKk4U4SZmimKC4k7ikOzAaXUCabLCfrVf2xEZILSpeMzgm1zHQPCJq9wIgyLUlLC5WEIXsC9S7
IDg/wmvH1rRMuyLyNiHqoF7c2YSaeDpbVpWFpnevuUsAVBRQosHSRCwEILDaFtoGeFroL3+PNiBn
dR8KY3gc868u28CHsIs5OpuadxIh3hGKImgi2J6FDyEJMV6SQDRVqt1mYHM2sL8jbqD61LEdwPm/
nZT4cc8jJPthxuLiqZZIWzciz4zusextE4fj7u8pgjyaxA+f38wwPIADcmETlhM+7s9gWh3WWNeH
Bh5md+bpLnGSR7QMLfjK1H9HtRbNh77V6LYOnMMGyolpHA/OfRT6jcphgr5ueBddlUyw+A1FrMyf
Iv1i2JsrAlKPAe11qZZUdBIWGNAZOv4BeOmueaOX+Zdce04I9QmROq1VCxDi+ETjXuqkIaIh/L/p
loZw/6lywtdKQUHzH/4jYWW/VafnqcxO1BeavMB5sKMer9Pu0DDX2io8K6W3zCUiW1SmUSaU611J
FpIicD2pbL3Q+NRfcKQMXm9IghD3dWVWQuUwFSDhMoqsLxnQGxu5ge+WoEoTC8d2k0FtBEJRHCdM
qxcnz+0vTXt+oxai7zx9QAmzUhZdANgllsTYBfQIgdDd8F3254M0nlfjy+Xr5slh6zW00pzlnVAs
QzSPau40NP1QZLDhKxbifJ18g7GwvTMV4RKSknXWRN49+vAGskepTwDRx3GUZawv49OwegPgNn0y
Ahxu253sprT3pMf+fWi9HQbmFnzvuuOH3B81LymZ2Tdl+arBMPRazFU7vsEqq73KVouE+WMY1EsR
CL754V59z7/NdStmteFQRpxB03tNSG6i+W6G5tP7auec0+ASxxzv3j8FH8d+F3xWnxhkQpfAJPbN
/2gmTI+pfVbT8UpyvAMeZchUbBcIXp+WWdoDErxURT52f4GkBY7nPXm6gOgGhLuEU5P1jlJOgHad
6vmzmMns+8K3OLYnqnbGzbfZ3ZXs7uwjmqqtyIdv89fpvJiLgQkxhCnAgtaKGXHTEFu4ex/vOnJ3
NleW0Heb274htre8Dxy7CRyG6GLlYEQV98VT0EeypC/YvPYDnOk5XuBhMoONuMl5wtC7dq1ghact
ql8mdiRZzzaGVyJ2WeWnVFstN93wP5vUqju0FgfIVn8YgBQA6lyTI6MZET6vrZCO+KIRjMNEOMHD
JMNPgmQl9AieqcPn78exYWFzSvhJg56VxY1jKImf0zPckhTL5DZocCFtCuCHTGaCbYB/O9/u0GvA
D8Ga94CGtHpza+8SRRjWSOm4xttPBX04Cm9jkjvpDvyHnTY5NsCEgBQ/LCpDXUJJLZYFPNETjUKR
syIAnm4XXiqDDikXsHoJdI069VOEeDyCpZhUllt4VWb5HDJ+kZZOoVNfYdd4uKBkp+9y2U6DTWje
NFeXMniiXHUa7JHqJ/14WYWZ3PERlf1/Hu3JNCrU7k+HE7Pb/6YUyt87JC2/Khz5tB43Qfi1C0au
HjT3E2yhjByNALbgPyWutXZ/OIuEnXh6D8hnN0tQR6nPo2HTqQKwvm5uuz7AD63DedrYqMt4Kewz
WUnG7C4ov1kH+lGFVpZa44XiqfERGYWmHOzZkGc+7Lm2CbFQio27bHuojMqAJlxolaBaExaMD4Vh
hZeL5zDgCEJ5szBkIOwxqL12aE6XbnaT6Z7KKWi8dH4SgS7VPVBXlxO5TdU6QYlBowh5pT/HhK81
CCKEGkr8+VvJUWt8GjQndX9T5D1iIHCsWVWRBmcdQOCNFMGszG4telYmEjG/N+D6EkE+ShABkqiX
JHM/FNDKyKWdAo6T+LiDnmkYiG5iUgtw1qEyTX2q+WFOPaBmYIlt9+dT8dIyV6SHoLEhLekJRHV3
ltANIDunfh/DGWlf0ihjLca2M8xAW4a1lRYfPDsFVWSPWmw5cys63J24K1AjQVHRF3HjUTarVAXD
8sYt5NoPLTzjCmwxkV3ZRR1T7gPL7NLIUF3w8xRQu4hz+ZEnB3fUs0igLWb6CZJddEAWLjvdqiqF
4mRQTRpx/9Ur2ZedkbjHTkzOAJt89tzI4epLwsqhirccZVcW+CKNgt8NpSxUKZSdhIzTRioZS/cX
s1hCBFb116ciUYJ1ich9yYmt6p+vh3GLk09epBY2hLlJeTlngX8QDLtXx37LgyO1ykmEZ7q6ywG7
YHbvVE0eh5vwj5ToKOZMvAAKfu0kx44UteuQjS+PeKzJ5D+pJTHyX3qUyq1mhQkVHCut4EmAoLRY
Zp6xGOqyPjMo5T36Enxn8LeazZFgV1Ka4HxagrT6Er30R7vxbBcCiEEXz7LWICC5VDSKsdHfhFV1
/hj840T+FgAKk4A7gEj3A+vJj6oRAM2NpCJbdrSaqptYhipM3L5Jp0joCI8e1cVTUUZQs8RoM0Zs
2OilIJCPQnFpK72UEtMxN5TiGSFd85orh8r/BITh0Qb7eYJRyb0wRu8/1u9RE2Qs5hZfFtmix4Yb
iAyidcW2qRBpqVxUxCaTSLT3MG6uKvpWj5QiOuLMnFE1Hc9cNBqtHB9vH3NsjCPBnMVqvQJcklrM
v2gGQIoKzdqPMd4FUDTc41cSkq0glMVsH8zaxKX0LTABVUjw8iQtzIdCImS+z8GsutBl8erzqZIx
me2dTIFa7S24c9eUccC4O8kA1ufV4OqghOjwwebJoGYuoWAlim4LNfrXmDRSP6FSCF/6yquCnmep
V12lj0PkRwwiLcIDN5FHc2t7N73xHWtPYLk2Izb8XGSe4QrxukyvQl96wY/J3/EUgqWuQCEOgs43
UtrTeEApnc6n/FGHs6QBomKBGr93EnfxBSlVIGiGOO05DSOfSpLPR2qUrJeKzhgEYEXfqx44qHaq
M6m6Jyr2k0vay/1gVY0qVLkeyWJLioQ45jyjw1X6nHQk+veRcaoe1HgUZo/PRKYhIO+npTPSiFit
w9uPTnjoW4LXp3uDJA8OmB6cEfb0BoBxUNaXGtJn5xRPV25esscppvEmjkdW9611pZTuGvMnERqb
IJh0mwBUzklIiIXoNmRlyXLTdAgCM2Aq7W0yW5Dhpqdax8D19+F05AKXp+HKssJhur79fhJHXD99
4XUCa2loL+8P20w0EMOwNm21IZhECj1SpmGsNVv6KC90x79wh1vnV70mSwoHSccxWQ/RBUmm5prR
QtfhnqxJIBiibQXo7yMEKykiwDxTnX4Ij70ggJtKSoJjoRrVrpoIJsjJgqDIx+y9MiHpV9p9Ss9y
onmzZMDykfaY1VUeEa9jLTHFP02sHIHBXyKydZDeHCO2C9ou3WwNwhDL8VOTkmvIR13BpJkRlmKB
r7H2HyvX+tMIB2ykSLzMEl1Y7+ebXNbPWN0kQFldI33QfhZmkHp/JYJV0s3LL1+8M8qd+2UkgMHL
uuUwSAcB40OypVaOg4zXDaa//LSZOz+RCUZEqAB5lGjsD14gVaWzuP08L37RR8qfBFSoRoj1ljWO
XOgsmojXw+mxy4ggJTYtCh0v36NVFsWqcmqaQu8xQ4Tz0ttJygdT7sG1rztfxZQqof/5AtfiJ8GC
IL0LJ3JB6ksEKC5RpYh5YFITSrctpvf7kOjeAv/O/403dj54Ptmh2wjMfmAPZxbarWsejK1mk7HB
jePekwmhSAjyiAlsIEmQ1jBpGweoKGFDF4ZcQzJpUFyVqI3o4ilet+6g3ip1tz0Tv6RNqHX0E+PL
dkwlmZiJ/Ee9xtFRv0YDlf67ASXYaRdRoD14hHwE/TLRUJ7GvrhL4JCsx2UJiXZs2VwhbtjFkOq5
4Mku63Mkf8gWL3bgPZLO5vlaU5gxsNdapaJ/+4X365uOTlDto6LUyZhJ6c3e2/aaevRV9cp6DY9T
zJXnzCA8zoOgWgHUriHP/p3P2hnxRLHHPr51Boni6fENwG0AGjuaEwbBMVitBxMzrjBAF+ZtFFyo
uwWPBg3oAeWKkTYTPRoGZK4h6AdnAcJD3ngsGP++vBzyCL2fZdG1xaWIHoXnzkBwsX7/9GmWOLld
43scIEucz0B6XC4m21LzFVxbD3KjwJQzSpgMtRyd9dY+EA0P5Ark7zr0IiVPtQ7Rw087oheZGk5S
Ta8KC+JAb0EI+lCidCT7n6CWZ1+/0sSb+RFGo93IYk/pIYSRK1lscJYTvDR+mbHP7jEn1f3kaUJb
VVzF3QZWHsRSkq40+ZM+x9LfclzviodVti/BExa6ykOmvNWlgm+wTYwJRwy/LPnY3F/xS2b6nDvF
IuzrekHmDmMap9q5tOLX6nW8y3HAqrbXDl7Dztupx7YeMrCrhNbeqdIo2nOkpAwYj+MUMFkZhowO
et7TCiWwQGhvZYdW7iQjVVsiw3O8tRC8t3FQH9mkPFy6Y4KLi7DNgo84N7JRxfH7orf7iPcM2Tgn
sbnr2HTPj7VTQxDMy5YK/tTH8rsmrsN8AAZvFOhatzztE3iUoehhHJCHTjD6njWnb1oyTL1qhnm0
R7azNrkxabUFRfp6qWNAeeyEaFzB8Ml1miYGPK0/HtTKDXeRjKNPAs9flOS56ZfGYWZ0q8V70XeK
ShSNhacpLDFn8UCK9QzyPfQQp23dF/dW5g2l4tg6TWnR9paGYXCVcBRcR914K3LYXxleeyxHWZ84
EL4NKvZwRA2/v6tVMHWqYxZLF0Sn5b0aSPf3wjnAh3Fty9AZr2hpoA4a8CInztfxWfChQVte5VMI
Jwv284F7lheJZRrBaZtooBD3uVNOP3CB6/RxOOkDb+ce6oz9MJd+/6fWEtObJ6vLyM7r2Fgqcx2x
DMCfyDLAfr+S78NVEQ4w2/ImlO7GhVzY28+0wYAucTgPLnZGjlXgWHkwT4PozXiU/B7ZlT11HvIk
eUJLu8qClXKloh+qa0KoBM2cUCwtfHgLBoaujNfsTzeXrMuY6ki/rnGfWnHisL4QvtSP9++COC2U
YqqWy72D/wxpzlxHW1rs39idJ+JMrtC8Ag6rVvgMgraTdCadqHG5UylqClmMBnJfvNU/7T4Bup49
Gk/58qmtJBmKR8LUfw3ATviMsb02wGC/B6rfBtPPnVTf4krum+qQxm9iN2OsTzW8CdCj2KO4EAXG
sOCmNReBbpZcBGDdyMC5jeeYYrE+gMCXm2mv8VVDq8OKXUm5o6HmEiARaDcZvnVwuwx5xBPKz5tg
/6T63+fBu9YatJN667B/io35AiquqJtFNXCfy+Rfb0mxJtuDEkZyTF+/Nvxn70SKHgtGu95NrHtc
768DAIySKWweyiE9bRyVWAGRQGyJvvALG6BOphCdLPWLC6vwzTi/dmqGmdQU9vtWZ0eyRhNsnAq9
P+HELZysa6uNe+1h1LsMuTvn/dnu70kT7o8uPN1/8B0QfvaZJMR65R8NKjBN03QPzUbooNrm+cgn
WiFNhPktcPikyl1aKLx96QzMjWKxNb6Dhvr2SqmuDKCti9Dv9/cmPo8PewgxmLt8HwRTpczGVm9X
BKyhy1jt/NC9TOqVzMAxeKbgnQoOocJWCcA8fPScRhV7C4HGlfJQ4NKXo/1Ms8FHs6Q5if42aBp4
hNMmekq3yb66A4qJipv5TK2YtmNvW9AS4OLqEwe5m4MLu420NS573gjH+34BFT4eDMeUrsWEM6Fj
3SGAd5EAWiq9Q8FWqMxaIFOkS5Bxv1z2xRWSyYttoDwU/yNo6NjrDfKQ2KtZgH5pscpjC2YtrgRj
FiSip0JGZDrqD0esASzXdjpasEcoK9BtspF3ECHjgvovcyMA4UZAcUUdnmdGhqAWP3/2BwY/ossV
hKpELF2bHONgDB6Paw7S+8qY5iCMjlaaU7aCVwoH+k37NcbFqNOl0yXM1zfO0P1XVCAu8uYh6i1O
bu5G8zUMt44nJlJQ4sQbbYD1D4awmZbIIQII2XlHKgKySc/rgXjQyED3IQb7N++oWw1ami7JNqo7
LAmWva9LZeZx1C3FA2d2gPpkWgd62NoPzONbpg8sJW9TKuIOTKnb3/Vc2p77aDxBtjI5W5U3YeSi
kJl+067vFR8rO3MLdoxVt74BqYGBXZgi/zjV5MBJxVlw1pmm93AhaIWv6vAnat8rO4OTco/vWo5+
9G2v8Kcl/dYFb42+kwAfh3GY3vO3g06+zvvmH6FAXwL+LSpSXecswc4WLZzBgPI454VccqMxWHJs
RAauCg1i1RDqWJXqC3yfe1mSmjhqwOURPdJ71b/YRlVrt8Ad0URGYTIqdA6eEZqq7LCqqm1Q48Zi
es4rkVU3hd7YTxp1ZCyloI+1rsGVhTJJ3EWA41UICf6RxmRxglWU52LDraE4edhSku08sR4+ZGe5
CrAcpikD1zem2CobfiDNLZzZXc0Ky4grA5N9Xbyib44TyXNoT+0WQQTtNazCTY/KCmAeBtCo3ttH
sOeMoDEr4GDCaN491GoIZyxni0+crIHL6YVWiRHBFegBVADzxCKuuqB+crZdGS2XmwgXZhzW9BQA
b/ZuN8LCN6sTmw/Eia1rq6W3ZjW1CvYgzX98RfuDoA5Cb8kNWVfEB0H+zwSfXEC0Qc1mjdNTCG5R
8VAOCkxjmRGmhLQZz/5VwLOOTZOQP3D4tb2nTv0/2le+185yHoUZmUUF1HFp+LxM6LOYv3eDQN3o
lcDkAPApwHWS1LcWanUGgDQkK3H/VNznrlZM5VZRjxgyaZ4og/DDBqs3XyJiDjWy9V/zkoG3JFEu
Wjlo9hXl4zvLbdVPtxwI8fAfE2C7BkGGFXNGqMzQgXeZgDkGAma8UrdnqwCkxUj3v3H73XMwSuEv
7PNSop6Ei7mk+1jeuiSt9wEjC8tujkWoEcHRUZrpqNECfShwM1UX3iaOOmINzwqpfYKayr++0NXy
aXB204nyNRxgJ4DmpTeHTOuIE77j6ZS9ogB/tegsWS7Ob5NB5tfeUi9ttVllzCQNr+qihiWXSwvm
u836YXcAD0ucTAoeTrX0OzthoMfjJEwfxOgHUYr7Oy9AE56sv0Hcmsrv0cR6PmYYL8VG7HnhWpDp
NbQwW6+xyR62LifmRzMcq8Takz+IPKI99dxUk6xTpmWXNs/3tYJmW8AH09C7lLjMJN0+tNmLYSY/
NBTxB7obNuQx5QDHuDP4f27pBYXgVNRSy2l3oEEKgp2uax5Y7imToS6ETs01bCZFHe3c/ux3Gmth
7DODMcCH0bFnxumuUSAQbpsEnXz0NSVoUSPw0dp4teK0dI5W9/TP7i1LpN59uhG5+47EZMtT1vu4
70+E60fU/EiTqjQz3G5UWZJKS7ulPoeEznPvqmvfFDHuvbiKXodaJrDn5F9rWEvCqw/Hh95mid6B
QItu5zP87N30tggEkDEq49z7GRguWSHv1rJJ/iC/lSu8X9mmikOmKDouX8KH2taFURXhkA1aNlDj
1WXCIRcUZOcV8K5wHqy/NO8H/M1F5rCrUqwZChcTpn8dN7wcYBlDJpvmO1RpItaSQc90dU83jUu0
Rr+DX1P2MArwHD0hi3MTjMs8QK9e+fGCXIvU0JGjS0Bgx+W0VST7T3MGzImXtEuzwNreFKHPewCF
6SugELy0ZWLhBGaQWHjzCLe1AuKWhIwB20b/anZcMsDzzMPMLFxDvy7fs/VwNGRZqVFKA2zmDn2+
SHpugvNg5k3JdN7HOkenUWjY8XgkgloQx8XycKlRJzNNywwozRNk1BgADtRcEnOoElIVNvA8vPZc
z2KIuRq6s5eZIpUTd81NdY6SnzM4D8XSNkQ2uweF09C3Cfy+SbBlEXQa0nTY9FCzEZa9v4Jqt6cK
V1KRZVDD6LvvQxMXOXUNPrtvoS4aG7TfuFi7nh2lFz1tZz3l0ocvDdx8h0EbJs3n7IW7JEnY43T3
hvEETpCfgqnHRHQvFeiSaCXjz2s3IsOEr3EWXWx7M4Ahw3L9z0sy9WOwTHULi+QKxMe0mIDrhxo+
NZXxF3eJxOQ5uMA0XU3upzhEnW7sHuoK5dft7vSVCoePl65566r/I1iqao94pOjT+N/PAzGGrX1+
CiyDmE7iZQsiinBR6QLaC6AB3//h5vDI9p0VB39R6cV48jtEd8dc4FyDgfRjLkahx2+MYdDGN8tD
D4MH5z07EWVXyGrdbGmXpjYCsdfsFQhk/32FITDqfgUjRwZcovoLvjBq2zTCb/dZb9WlYcTQRlTu
iY9l93+oWnwGmFK9eQlqqisb8c4U5BYbkgSsZQclna1b2aiOaDbrcuvWx9cfXJE6k+p1CX3+q5c3
nkwSqCfpePvxwHJVeU7O5LIMb4TRC3bbYZbBBMVDyLwy7YRHSDtD/1zVgw1gIRYSuU3ipdhhk/dP
lrtatJed86/i3ypxmdKMMg6JYJ92k0QI/0wJJOkUooNadyOXaQzVK+gwh8htguj7Sc7D5izYujZB
XCr8OW23uTiUNVfVPKYOAYcpoou1VUP1IjKHai+WIuJkmil80w1WGRyarvl52ZSOtBT9DqYIdOhW
xkCTD3Z5RUHoSknnq+Mju8tZUfdwoEMFoyyazkHXtTXifHLBd24uZ5VKlCNiAnGtJXWLazZrzze3
ZWCZBn3OMR+ya8hLROnF/pjx5f+W86NAAAY/CIXr5y31A93aFAzNf3mNaW2iUSd2VqrjtvZ747mH
kYazygqCInuwLScpgjyeXD6gwpp2E8Y5YJKOAlX1JMpLgob5020lTChloE9/V8a6VsZczLvIr6QY
1pDEiaxkvRobxsKc8kqTuBq1LnSVtY+zPaoJM4+t5nwRpFITSc6LRwQBikDwYCEvs6RQO4La/743
9e9smlpZGuTsl+tgFNqzGKpor0i4YA6Yss/K7n1SygPQCJCwk1bNnV8I2MqXsB4Vg26t6KUBUU7m
/4poSiBtmZPkSnwl3MiL40eIJSK5g6IpROorZaOjIjgY6U34APojGJifGb3452VYeud6RFjEMogs
lSPtcPHrtERkFyNFMrEXQcIoh/35V+8bgekR/asc+PBSsaeAbq3SFKkieyJcwN5jZS4086h725BX
eNC1hVohi0ptypu7i/Z8afMVhhmdoJm471LaYgZR2x2YoKu01JKP16iDtwgOiCb3RBpIuQvIK6ny
SUvNVTDrdwfWWAyGtABefeaHGNzF+5mL+CRCs+HpuZekpStW2DkstD4RUdIwXaAwKxLgiJJB+DtM
sXYeBVLP5DAUTT/LlxjaPkV7ats/VZaXe7IaHzesZXo8XfEhWvzIObQdodIt3P+8FoD/sceIcAts
gA0pIU3omjMjvVrM7/pQaoCQhioNu7Nfho9Cb4ak6tqtY+ZriazC870UdwPQgLcI2H7GYTM7Xz01
0EpsoCukcVFRmrxQfa5h3GE7eBq82pyrnCEixve0zNAfyJgcpwirOn9o2kBoqJnMkX1QaDyh6iJJ
T5E5vi25vh3iOkegtvB5oqSp52Q+20pRPtfsmAuHBCrTOeJtuPbZfxbOzF0BZHfo1cTE4DEqdrrv
JTl0743M62ceKX8YEl30hyBB4Ik+Ilcv3V4woOoQZgbxVV/yvOZZ0vEcS6YY4Z89tywkfB3UKt7o
Ju75YP+WYaYNDtJYaMX+q9o/cQUERN1HGbSDC+O7UpTsQIKYdcHxcq6rPuVvFq8dnUSE543MSSWj
X2+pbRTXvARatsU/jOzn6RdZAg4Y2189cl5IkN/QimguFxdJWfaj0iwD9Pc8qCujJeOHaDA9bbEI
yJsRYZQ95FpVl5h+yhAMC8q7lKakp6B1zm/I1yaAthcRJBiwPtXGJdHj8E6rbKyBJbyijXu3upvC
AFJcvjh8TRTeHRHU/MrEJz49n1qAXgM1q2jXrsUsUoc1DJ2C5Crb+O4Xe9eZtW4Ef836ZoZaSndn
wt6iWpmv65/8t0RWI+vLzIKe+q5EeTHusz3ZJ+35UXbqBWBCJgGQWLGGwjpV5CaZmFKwKmoLfCJK
YDfW8T3axg65LeSTGIfycgpIZVaHCJbvMuWz63BA3OJPMxAaFKTV65VUi3hFlxtHQXLCJCbKVCoN
p7fVTiv/jzohY/UzMYEYdkryQ/b7ZFfFEc8lPU49mKkwl7QtR/jWsp7jITCU3xpMqnxQy3jotGw/
RP2V/vQg1wM/8LhIv1MwVnF8a+k7QT4m9M2iRWwi7XfOWWc0PX9oc14Ochkr6KR1Ag+QDL2lR6br
54Lqc+XE04nk/lUgqACPTgOPNtir7ypMZjQa+k0U37X29ZaufNAVjXqU1kKg8gIlF6kD/Q5qcubc
RQ2o4fs/1MPRzxUAgAHcNPmZTEkxQGLmOl3EpPy2Ads50jzl8xP+qQc3NMyveo0f/oV02s0hgcNK
DqHfk0bOGnMr6Q77AVEEDAPIxkfWNm4pIJk7PYOKMPcpy4x/ZKhhE6i2lCVHSQs2pin6aQmKw0mP
pB6nRS3BmFdN8N2jLUsW9e+96uasrCO2Jll+NBkO5DnN3NB8iJTN3YDcrNlSxWAXtiwYsZZMdrRo
zgTvf5EK3fdQfAZFUBHoXW5ceDzHRcuwPtNZkmunAFi36UOJVo8ZDXnYcoa5a/QTPslIt5247EAU
/2bi7I9E2XQVgmKvNz2HAHuq+CRvZ5OIia9GdW+MwyiJMqX1SV32yzMkQOJwqteFL7xW2RPcdAcZ
kxqgvjw6SlJEq4LsKiYk0IP2LZbMJZVv/+6d3EuLd9wiDk1rQfuXGtZ+S24sI5XlZZtYlQ4TN9XD
oiv9nNUy9RtYE/L1jnAsDWBwY3KpDCZBVTl2uMNQAvXJL+IvQcaIB4Se8ahrJ8Ir/rIb9HbHaVQR
n8vDlW3OJzZT5ySxBVeO4sVaToKMMVI19JmLIJf0MfhD36mbuXxYT4y2CwJAvXqNKTH71H5MXROf
o6duduUUYMK8HYU9afGn80GlUV2KfmM6Jt73qDiKDJxJ/vg3LicQBiEQBFksww9k5XhCLTtHtsa7
GDwAfGmChK5+TeTnlpbEx+npYSgg1ije1T/hY3pKMvPIXGbewJj/TUhXkxHVZoa1/tBtqDcpZz7x
qJTB+rtUphV+Z55+arZT1/xKZCwZ3F73SM2GaTshdYuSku072yjdDhULx7L7VeduO08DoFGSDSqf
LhWhPBaVhkVkWnunp+UVsBDdrfUiBHVQcycXJaGd4X3xbyAYMc2TEIn0Nvqg8HaO1syPY1I2YrhP
f9cNx19RHPe61coX/4b+xsyOAoeVMMD+hNlboBJla2wUgDxMetWKMxeKE8LmGSXwR82cRyVwSrMX
Vd+ROd26NUGR+hgyYvEWMnDonZopGJPOIcj/iIfHRI96v6OBXz0BFkuWk30YohzuupcpsZ5icsOI
9KAkBdd6qGTNVIs4ZXfcE2NAIsWroZAOLUTa/ogc8eiMX9TqaU1qhJAfeJmR8E5oWGyGeB5gKwmk
9ojQjeFOA7lfB0uF57XMs7lKdPoRIfVNP/ZyJJFTWKelXYfKjMAw8mLkgII7G/iju7nr2z4DXS3q
bcYQCti0hIuMm/qmE+SxVEoAWzVsf+nVazVuGfG8JDoaPwUfmg61SJz002UT9acB6xLxO57MuaRu
B1p4O5g9mb39Z2XnYIqZhv7qi46AWG0nJIf1QIPvRGyvJYoXPL3aqjzyAICxLkc5cdj74hSScS4k
oPDxd4C7jPE/0+sq3+81zGLcrAuDxPbVNHA1tZ/EQKhWeFiGG2e4ruRikpJRUcqEc64xNSz6R1Wt
2ebSidT9tkWaQ0TQiaSynB3UWbcIZyRf98OLkJ1Tsb+McQ6fbLblBlC66Vl+L0XD5oHsFhq8nyUa
NWST6qW/5bl0VX81cwgYmzgQH2ejl/3V2zhwWlMcaBSUpVN7braLFxso3JgeW3xlGGGvZxfOUiO4
kaERn5Kg46WJXTTFH1AbGMBySsVCshCxSkWtDcvSUvkZ3dCEPweMlh4EpcUWGFCkp8tDf5LE41fi
Rzw91Ec+gLqEbVXCX4FO3OlndN75Lyhq00yqLmuXb+VmmFaQDvxWAsOqkoBR2JIu7Spc7uxlEdfq
pTeROmLVjIok2D1Y0CEo+XjmIe7G64PPQATvxtMaqgXIe91HCUXDV39mNYNUhRKE2JtgQzD+We5f
quJiXBXnFRTyD3BSzyxFAa7VRpMRHa1taoHxMmIMRvBslAyG5n24dozw/c1IuR4mkoCKEvrqnjrZ
5qwrW9AyaWAyXDC7e+t0JuIK/2pVt1/8aKKVQY/VyVhf6Azy6P2S3Vd2ryZE014cbz1k6k6oaAPb
ekz2ltpwV8iUdNZk3Jrgx4flvUrdnfrRNk8KGhDuWadEfZm+HMwGeRXDXVrMY3a1Mpiz5VIN2grU
i8WzlIcIFNFSrB72I9+PSKl7iWo8vvV7GcydwJ+s9235IzfNbJP7LfwUGaefCEgU7xE7ECF8bi9Z
gOnuw63o3a5z80h4UVhtShBWREoBZyYflAc1KUeQUNvsz2HeyatSvq55dKW9BHXpsHkzbNbHohdU
Jk5QcUocjDkfDXaoz72dYabPd3u3d1NeGotdgEwDptiKpbMP240g4CwvjnPTevn3wuiAexzQzVEZ
Q7uft95cLVyAVCLdn0Jg8NjnbQhQvwHDbXp1F1RjGVR5CucxHo6L7JtNd0j8uxV1eUWREZdPIk/A
lapt0/YvNJLaC4YtACSCaqwtznbw/ahi4BWNPexYaJOKJqS9yLwqGTS5L/4AAyWXSw8kB0Bjq9tS
VOJZeLIJVydbiZasInH3w4dgQjh52vOwo5zDuUbMKrWGGWWTIdYeQoYu92O7LDo1Ukg0KDZa1HYZ
23zA7pp8T1SWhVxEceb/pziJ26Yzn2cLxD2f51qy47FkHqfbaMFSh483j1GIJf1QaVzCX151oa5c
ldw1VRTBKORWGbE2L7EUUUZHlWbpf20U/NaL8252xUOVlGEvsUtSr3Bb/zslxJAxlA/gFUkI/UUj
yXVEP0XK8NUURyC1OvmQknKgHTohKcIz1b4fPvC2kRyvo+1DF9gJS3dapV36B5rlF+QJsqN61KWt
T1rMFFnIMr+Uz5t10m/aEfS9ftDxHC4kvQJ4L4353EuQuar9+/nzBYGkgKEDF120sLh/3N2266lN
u7bz6j/aNlgnpwk0brHsDSQz7o8mnJhvpAhj9HnHGaWf6a/IeSQlrGurcUw8rwqgsFHaTV1bBFJr
j9WWjeMFrHHbitoA2r1J3V+qDroKmCCXv/mCMzM1InRMu43j+nR4YF1LZfrHrv6+RNhyteoVNEo2
udk9qY3sBTHOmEXNHvf01wPShQK+LzdpZ+NP82GYz0S1vTOZLPVmQzICHhKmXAZFtJO4Fe5QutyF
20LFPS8PmX4tTARhpSn2QtYQGJIGigB/YqggAuPP7HaujmH9IwwbazarKH4JntIvyvq3hhaGYig2
UywNJRPkoqGuDlVgYbGbThx3ZtXIWmXZddpe715326K4et0U/AYESk5FQ5jYze6mBBgId/O75YQX
/wbiuQ2PrbIuxA7g+dL2cK+76eW0b62UlMDklHc0YBQ5E8f7YR6GaxK2te9W3RjnD8p+clJaL5BV
lqT8JI3k37+Y9GR7ZbH8i88qFrtGVHBk2XIOY5TdGhyNcMg/Ruxr293D9H3H7GcJK+BI/6AsmHUD
NYOTQTskQGvMarY6BFmjw9hg9Ym9cn6NPi4Z8cnphL3HOHjiiV6qcZ5UwbvNFuYGYq66GCfG9UkO
A+XsCnTwU+QM/WXUgYLgDYW0IVYZxaNqFcuUhjxct0OOgnfzOsn4BAyWWs5yO7IRG3pSJzpSxyN0
8B87HU8m98LDsClD86N3c6N0B6wk8k5jwYoriSo3OLPnbrVhEV5W05MTIFxgF5lq1gXAaplmHqLv
wvaFngkAdbywmJvLxAWsctGRc1wxXhFJgZyaeJJBDezjamNGhCZsZ5RXy0rRuYWCqXmlLVa69fwz
KiKOWuKkEQqlFllALFawpfvfIeaE1dYCh2JOtOlU3FdhzhNzfjG8hYtmEnJnkCUOmgUk2ZRcWZg9
7N+dTZ0se9YF6QXTG02MqDfC73v1Buc7BudXem3nYRK/1jPt4OP7mc0Xh6ZiUiMZZ+tEpdz+ltaP
DULiQk21WN/FCDR5YZFiGFa/xHHieQUPT4tol4SEhcevJ8880w2fpRIjlvQWdA8D/0t6Qf418F/K
LImJ/80bSn5w+HBPPWCiI0De8xCz0qUmsE7yKEpr2vxYCX5FmumIu/yRMD/GJlRQrrvst73ohhVa
bhoSktiXCMUG2ARuMsqh2XaJLo9kVVIcSQQ/Zqp7ij178mN2Tocfy63EG55WdD8miXsLyEk7d9x6
t6iciy8Ilr8tUHRurxH6XjRrP3RPlP4uDvmof18JZXOEJ03RZJ/UnRaRWa3VtNVjdnDc1n+Ngiua
eKmILpOmaWA8KKXTKxrvzMgQzz3hM+IWpMz2sZkLoqoUwl8AWgB+xRkNY75UyfsauFKSYwnyHYF8
14vcw4H5pDITrjpN6AeI1gJeWxxRI93Y/GRnznFMqv8ZMIysdC01o2Lmh5QZmOf7VTC3iAT+1G0O
8P1EeI+A3CcjGusEI01oaqLjFVAYxBjnXb1zeUuv2KIww9xhca+yw3mNSOLXPo0fHMBc9HOHntop
9tRgw2rO4CHgv9u+erkRH63UAW5heTccuk9wA6Yg1UIlBCDCCAzslPd4hh7YeaXzibqP5a3IOxwc
NEb601BY4V/dyq+AeVo3rMrjBg9hX8BjdHoVprXOApILONJTOG4zE3kmv6UQoIgQxiP515q6Fmv6
oc3SHJKGlreF+JfDBCRkZTjRvFxXbLmnayfOgS1FoKdEgHzktpnMKuyu/DTWhaL5V9t7y/WubhnS
jPPbaqwsr+2dI91Vtc5gGmP/wmO4kOIFxmMcEZJLy7EyJ6y4IXOUHV9CoLORcktMvp5oluk8kdMM
BSrI8Fq3JSA1XXv598/k1KOqMGSV7JfGIR1YEQOr3H7o1KUE9IzPtjTbUdzx6gvHVSte2TPXANYH
/PW6SWUAvApQzBjH4IiljouhWLimeqIUfs6fUrqDU/DP4/aZxy+uKNvhcuixZUMsvWbxbLu3ZVYk
YWpi050HRbj+HoTqDZFclf92dMjo8uUOoBPqQ3tNDjMMTO8h/yJBgOacxMzaKhfOlgjFBZUOfplv
0jNa2AN0NaKR8SURdg5Vucrp0MGvlDCKzGELbtR/sijBhEEHNQOdNsW1zXT6vKQtBssZn8nfVOM+
1zgbxrfmi2cvDuf1hsNx33Meq36b7UMveCOw53jCtJOEOOCQbycyXY/C+sX3qHmDKNcs3uqIbchr
5zaS+SUo7SYUKTrKnwxE1ZPDyKTQgKfGXscGwN5HlrYLfHL6mjkbHfFZvBf+o+CNFsJFCBZMvXGJ
FwO7Jy6VsjgA3EWnwsmmCdPOLrHMF5/X4TNUqPM5pOEyc7au57JxkNqm/zyiIqinG3HCE6TZiICm
U0G82UDRjkwjVFvN7d4wlin49DuotqU8JLzNP4s1PBbmDoyNP3oVJG8oBZ0kc9nSwkCjGUGPorgH
Uwfb3wuW2hQNFFiGhJSLD9WT4+87d2brouESDFVXb8afb1+O6Cq8JELhV7B6cFJHP2f3ROmPWomZ
FCEYTnQpdp3mMxtw0gVSZSYj9UMB63I1TcQtYhFK5xFph5XJqLAe35W1hWGPSKZ/RBNvkzPNd0ny
epJKdsXQYkvFJU9cEpXdXthMzaqpT3Gu06jNy9IB1qJf0WLDbKoKVInkFWcogXfSKrwynxQTOXg3
Uf8u6eRAF7YS7s4VxrZ6ck0Nec0A2EQDN21HKO8t5rAaCWxy+TfblRFgX7BTz9sFj5Fl0SAYI5z8
26sMupgGfgEfz9e3053Qt26YS00PzZWirTk5f4VzAk6BXK+C8GcdKwtSvDW+reIJfVWdMzNx20eA
KFT1Imt7a8eZSJVkv1oqKwWAgAsBzy68mYjO2x19AQTOzV3ncwIaV711gp9xTiDr5wftmQlZvE1A
d7bJ26zXDSsM2Ho+8YIGzt5qs6shp2wYmfZrbO9dPa9wzBYguzDwJKBGl3rs6d2p1r6ASdftBKyb
fy9qxAvojSzx4LWrJ2KVCn2A12D94POK56y5DZizG5rW+dKYQqizig85SMcFaBw2dfCbKgd7sigi
Fsb3+LT0uXMUXpwqp+l9irB4Q89JW3I5qlgIOjzZ9/VEH+hMpnJ+5ZVaLvrStYe1Sa+yXMejwxY5
ymmn6h7cJG/T+9fHKWvmzKhZgcBDDvCQ2JhAOMN8Db7YZn/Rvmy7erjhA5D6H6Fds0jLrn1ZqD1i
cqYOtsQz9gKI7Nr9+XHEISuvlQhEPAi8Wp5sS45jRQ7LhFb5FSiIbqwVIOZjnFo+t+YHaiYLdj2d
+t7GoqDn7kO7vyAHVQmg6B0NMLsAWxmMBJoB0rGbKtaKuKC8Ark0+e46JzukgPrKh1IZcJFPymDu
9drFNBGLyX6Nrn/cbhtZv+N1PR5sNlTwCxnwm+E7uByUkc4ej4Rui2cKkebTDOESbKNZrQ7CkMFm
jH6cE1SYDoBMcnDZlY9yC7kip7NL9epHLZ7iI82LcaHfoGD2jHYX6FBVBeOdVXOzpRNzyKVAA26d
8jq9Zyzu8oUQgORwSHsJvOFgzrDpBN8ePb757VfwHZJAK7mjLNS0sOosc+2vLQjxjf71uo9W8NQ8
4ls5vyxNyl8Wpp5AKnoc2/yMxPkcgCkQnTuwJKLV3cvfDDSpf0SG6ukJpaXyvXjkJFB//DcFdJBi
2mPo0e77Q14Dvx94OFAekLrubZUIhIMlcXjP0CxZvjd2T1ewg4/ANi6eIu1LeW+q63VxEWXW8bql
Qbg1T6upnabglg5yfa9pDg1S75PSNi7u0Sk5Fl5A/DblJdYUWocNU6JUtMLczpIJo2+aBIxQ1IRh
IfrMsR6WgLHB8+6+cQhpbfXSn6M7XqYOA+fBMSirWH9wj73z3Sy66ofY7phiMNrdtt17CTmn4H1a
nWCfep+V/abYcGvZCmibCrjyeYFXn0AgBAW7R3/kP/Vop0P/RgsqPa4xJatRGxZOfUUCWjYtCzql
Z4DDNHepskbCufORSBVfcOuxNp/yMZbvBICQShKPliSCgpiQsk48UMaf1LAnCMYQt3FdYWnclNC5
hu7ZTH9+yHrudWOq96XVIk2QvkyHgp52OWYaQJaeZVNcrgFTXfG5C/Unhtg/7Hims/PKtGxojrIw
IdiBAu3s0glvnNPu9jvKLE+og+C1Sf9/LPRpYNAjtsyT2MXyZ4V5sbfQeAjl4ijhRxRGJVOcWXAi
XoWmTbtepp7DUlpg0h0Zu0RAp1XK0hZ6e/aAU2zKMyur8ibBu7NHgHMj4s8gaIrhV2fF6q51/Ip0
GOIqoRBDfWwE7uhMYeiD0RZPeLHd9MoXlar4LqMlfkRY+sRR7ofBfFd45vjFRCzjNY9ahdP5zNAJ
X30em5ptKnBTCCd1XvO4veBhXobyNDtTcRIxDEVTfmyO2NFbvc802dEWmOHVAzcPOO5JxrtV0BxP
HX3udkQojmXMX4GHnstlthcQqflNaaldR7js70eVhyMhiU6dbgeUTWIVQH0xaonV6Z5NkELD3Nst
mxRSs/L30YThy2blEntEgYjXB7x8gbXiUvE86uOas6HRAUVOvKV5y49XIHwfobsHacgOCp5dDRPD
YjGyFjRiEZUgRM7C9gaeZ1lWRsLJPwnHG3EThVfGTHZH+m8FHXSUFagZ/IHAq8MwYZY3KggHTnRz
rdG4eXJfY/3N6AbSnYl2M29jDMSWF/9EFZxOOXf4dwvyTKEjrz9kxn0UY8LSfYiytCx6r301SqY7
Jx/BkJGaWeL0ss89rPfIggQDfHm65pDmwwT9YtggGIvCYarCD3ZEFHiSe2j6u0oolQGza49dV8JC
rbmgP2b5HdWOChZDIlzO9m2HAAP83KRYXgSnFJyjfhoy5NXCyoTo9nlIIHH/gezdtTRBQfMCT1tJ
nqTuViW/02dGr/gwkPcsEqaaesvA0PSUshWHiM9cbbz6Kt0c1feJSJ1jY2ZUvbyYfRw4MHus0p0i
6wN++iJVDFeM4OYqXtI+14bIXOLvWm5JxMp6LqKG+WnBzXPX3v1oPEQTrvsCOwq3kdtmA7Dppwsv
rPg3Xu1f08k0nDlO1f79RcuRV9fN8evOf7wgfVfkzHJN5zbeciicsz2RtDgnrKRQM+xbM1kVrzU3
dLStBOQexnCEp9ghIG6E1A1rOGo3yVU5pKNRLI26PKZQk4pvnGerYj/2E0OQ+V0LInENZHJJ48zs
RK1lWnWa8mvsEk5QMD2HVxdDHKX9dJJjuBeQ9ACAmvL7pFc8G4uzgJE+5jJDpQzYnEZKFN2r/js+
VttIJev8Q3y585tosSMUtZkJNGcdncmXYj3nPOBcMvqOaKniQHX6Cj5DgLesYF1bCj4Y6qZRR9/N
QIp6nLFapnS2HU5vtnhzWSjM32LpAnTYODDFiTZF+akTCP/Tp9Dikfus644nBadbWhqXXAEU7om5
/nR5Pe29E3SrkkA5iUlBeBieSusoNJPJSQMnbdDV91hKsVyv7v+oM6Cnxh1hVxUktuQRZ0gaesAL
lv/t8VGAPC/laK47dvNVw8WB9+52jiVQmczIGEC19HUMtDYRk4+fu5O+l+C++T5w5tb7Guid5os1
vDmB2XOhAUOGw+I1PhbH4lTUO9BwhnrKcC5uqWAexppZLPdEttFgmfcqMnt8a2uWPENExSGUOWeZ
ifIJxTs8/Rx6OVBZIHCd2JcWKpu5U+ygZcvPA829rgTa3C9aqe3+Kki953jzcmmmNxFd5YaTJYUO
t2nIljzutD+kQFIpooFR5HB5zcNXBs5lNngre3kf0eIbYMKmY5DRI/uw8rUJZfBXNhRqzuJtLkAi
PymwCHEZAoJ6t0JSSd7R3yll0tffjBBNyfTGrpbt+CP29IitHpFzk/EolnO1qo4U1oEOJnE5c21w
BS+0qlwd4rDHnHQ6/PsaG5MfBYjHpgfE51KWAA8ANJQygk6Lso7JWlu8ydhoiM1j6WHbKhLLqeIh
cPqlvoYBBt9fyoEUPVWSH4UyJaDwUrp1nt3YU8/zz/Yzl8UOdJA7+lUjRix8FYuC6OYgc5Gx3ak/
r2Xa8WF8kMbXRG9f0CVA//yPXm5EaEElkZEnCb9yLmYjNTWhVaE6JwMlJBJshtJxglkJRG8kfWo7
5Rg62bK4FzyAmE8UF/nBmVOPW2bUE7e6wyrXf8kHDnxtCmlFBCETw6LGfnWC3jp8nt5woT45BOAZ
6BPE8BVPn45On/eDwh0V0kSSI+N05NqeZFrICILRNeQjvKRbnluTtP9QwMDmjo1zZbBnW02EE/1E
GMhxwsONIEeQqkQitmNSd85DbgWfuCFwIJn4drE7prZIaSiI3jiggBtK5Bx6r6jXjs9M97yQE4ry
VhptAvS4VISALCaue6I5g3em0XhYOYxl78I5ikTC0rvldANIZFHI3+fVvBIQjVjQLpn1yI+6+rf1
mwI3gwLpy5ly4ufAckoX8XV3oIDxHV5CnmQRsbXZDVpVJYQ4uA/PgO/7/xiwCRrpMl0N8gXTGQH3
EkmUDtQRWlJIRj96pRdo9/iHRl1kYFY3szyOYe22AnYIaCp7AgOzCfhcwqVPOdorwY8psPRmd4sB
JawdA+js7/7HMPZWcvvkIuPTz00Ovdc8FbW+C8llfp1pKzyNF1lLTt7jG+RRThK21iRLLI7V3LLX
exop5puZ9HoylEcoGKS3NJLnPZuA9UkQGN+HcUObC8oKpQ3u1S+vhgIp7GfjyaPhgnhM0k45lmOL
baxpcMIfnXCLVGTQvysejIx7SIzdvHHXZ8cGMI/rLg+Pp3EFiaDAyPnGxBsPL3GuX+Ydj6tmvbUr
g1NFm/YaBCdpmi3p4ID+Ps9kO9VyLZ4cVfWi4PXvaHXoS1G7PhXxztPxM8Q4PdC8PYcXuZIpUhqF
0NG7a4fXS3Dzb3pPfo2g9W/X7mhfg9XtMwbLbujh9Nc0WbaGnMd+hQHw0w/6PWUevhPHEkvEB3Mj
oqVs1T8HIe6yukyxALo1JANpW3uo5RUNtoTUTN70XUR6TrRGCidpAORY4kJX4Row73SEsZNbMqCq
HNLmX+xLDT2ETUawo57Hcs6zLwPiUomqGI0QFiR7T+9XNveOVs8HywZRJO7C+Nlv28XyyCXlNwU/
KYxi6a0POkF+wneTyRt+E+oIst5anER6xGofX0aIuJXLB400qIu1knJtQbK8dPmoEYEEJYCgy2Jl
Dqk7ZSnFu1jvwQukF+6uSs76V7ACugqxWSyxUDgeckR7GOu9Sv3msFP2A6u4Q/qNSY4rSV+kLi50
yYiQIeeR85xIVuy7CPagiY0SsvrUOvwtQZ85pYmj6eR/QSWwWJ7gz3yi+LgTBic9jlJz0H5T8+64
rNi1CQK5wWj1eJzl7IyeTO7ZRMZKK78pk8OOdi7Zs9+AAPXp1zMsTRcXP4wEUIeYD8uCZ9SB6M9d
6QA/I4UBLhmtbfsqJ8lxbssG/WiEWD41HncTDTSYsmjvarzYTXANiWU/QmN+hLoaYlA1JBO1zRFl
V3dZjoBXx/n/IJ3Zboc+4491Bs/82UYzusu4pp3s1vaNojPwtGTtU5bkuQEQ+doDLiEQSd9I6VSE
Hf3TXkKXE4w/b7hIT4vk0I8eb51tzvXR6Bk07MC64YphAYT2wTv2RxgeBYZF5HKyNuB3RS8M0/gQ
ynsy8dny5rwYUW61TghL2mvRj+wIAi+KLLdk81nKtUpi2Pqq+idn3cWjmXq2KS4fSeqoAm3ZX8rx
WggGMvLk3dugGiRLT0SdKNf8OdCfS7EW1Y+dCjJ47rmdXy5BA73gk/aPXY1A50jQcFY1zVd9RFmg
gzFgzlU1aL3BlJYk2+bPB24oyx1c42kL2BlRVKmq0bMHXX3VcjUYYDyd2G+Nbwidbvgr429zPFx7
oS2FZdYbv99gGAFe/Ceq0x5X0XcvTR4/enrbV80XzL3LTd1+tzHKCzMFcIl8IpQWYYYSvKPLTgH2
oZAzR1AXdF/TvM46SB0dwJZsMddhUHSVPfHzLnJesc/4EpFDZ9gcRAm1bQMn0i0HpmOLs+Jt35Zq
jYiDCa2swT+0vSxS+zuj3vG8kti2CxzLZOy+WyVhSL3DyZSdI0EIWypingG61LjpoDG9hVAYsQbU
87DWdW37D70dsujubPmYjbhHsCenv4us9O8qjVW+bFOTTF/R2viLTUGU8cBjTO2vtH+by8v4kJHa
6uCuaXPuUW4rkKS98/Z+i0WKvyiea3uRn21CAn0Q3qiSzMTxu6s4yAAvpBNKIhs7P+iCqVHeHtPO
CaNJZLkl75sQxpZawpPaEL6NPcENrmImyrNF4Zt6pLe/ltT8crn3IeFlt9LKDihDaaReE3hYoABY
Ht/yQPKFv0+mj1J8x8e2b/y1zQWZ5cU9W/LQZLraCSCApELex/dPmRg9Jg/wSrDWUWbw+bf4qFtF
ar8NuTK4Cc//F1Qv8YNJPs8mE5H1I6/dIi1LxvDiH8qDCHsU8pRYZzSf7RlWf3uqF9sUnDns/LSO
FO3ibmmjefjL5mzcxsK143O4PIjnFo9Pns96tsHfupbhPh5dhlvkUx6sHCnlqGOV7wzPwo0/E3RC
dQ6aqox5ew46T/HT1KnGin8odREsVlgsu/hrt2JgcT8+0dvSGRO9WBBwGUpEbMuqik/3W1yjDYE3
nbUeZTJfekd/YiDItM7gFRG49jRxZOPPll/poLqknmdO3KVJ9Ft0cxuUiBxvfzs6HklHYGBqmZip
hRsaT0TeR1zBXlxmxL43AsfjPGFNexzcgsFa+6/9ukooyE30eOQptD4YLj/NcAf/bB6GulYtRvli
RRl6bq17FymbPzB2MOB0hfvYJx69ES7E/s9YSjYu1YBhZ9V5I3JzAiq5qepXhyC98qg1uf63b3cf
1OgL9cxjNiTFWztsm0N6kamZ1AtL0A9XcHTGjvcG+JzsL5FYUnZnLfQ6psxU1xfzT+AwogBdvrLO
a3tm7gq0od7o9ggcuaASpeois5sUe8UGdPe1841DzuoNg9rojz0z1zuj6krtVLTbnDXX7usrKE1U
3tILcDtj53T7vt3ZA5b1qrEPs6MDqhyjyirNNRe+MN8RnWJZMw7WwkOZIsaxQGOtwaxZOxESmKMQ
PzzfVBjiwcdc0v9KmAMfFewwOXW2jFbQrnCPCgezTH+GSkqiLRb9zS2MnWZJiNrLLS6xggPeMUOg
cgrMz3fupv+Nzwb55vYB5oRWQiaJaE8Q+Iy2NjVgwvijCyzbMrrUhWcUrZzUNEFDomGj+mTNv0Oi
OM+z4EXb3CwiAzH5sBLReReSeA7ghTmEiah50zcRO7AMDE6shK7cuyE6odDChI8SOko5OtfdyGwx
GIs4c7ZHZSSSBGanUcmhqI0CHT3J1n0ePHJHbw/93iqDYB08BSZ4ODlp5UIfH8e2by+P/6gXESnA
ZqZEbwtSbRgZixCQqMc2lilyU40ClW1xx7m1SZWTH07fnoEvVDJEhhv4zlb1/d7a2c10pbHOGoIA
Po98ez/JUx+1hFalR5Y3p/zMbOTIBfWTlU4Q48SsNoV24nD9BepVJTCUU+xE36ytiQd6K521IGyK
d6ijz4rV+5P6Cynxhn9HIjtJwmMCAY5LqRLDOKkXlfOGh4o/f8u7e69gjhbsZsntKus0L7mqQIo+
o6K0PbNKWvmwS6qSTyCvOrESilrp/mM2hGcxmgCuvSITd0nL/2G5w/l6KN81wlAUA3wUgFMpNF7x
3G08COSNU2UmxnD3zz/i0urXRf/Bvjnv6Ly2jTiz45LhQMDtr18rMELV7S92/EV7dP8310cwZLPa
DV050utIWquWzpT0ax+mEK7sv50RTbPegzOHsBv/1JFPJZSaDesWomp+tE8ecO3JlWoBdfSYBPYO
b/VweyQ3SVvv99SHduB8qTGct/TNEn2x1jX2VFKj7I3pdu3JyYjigGnyYIj7aKoSqfBcyJDHD4g6
FOjFrrM6IpwMUOe+4NgF7Qz/aOf5uchJ3bXop0mH7976K5ceI+THHVm6LtImQ9fAiJnYFfj7Q7s1
yLRAsxp9OPkEUPEgw+QbPxxZ16s0Z56ivF0j5EORjEZbZdYksArjEns2ug7qiEnpg9pzCJq02N57
2+aircu+AcjRzlS8IBceHKCQmvvxIRlyY8hndkeWa2aVOSlsfzbC/7vsQcYY+C37n1o5tLNMlno4
pffDY1NMaZu1FgW587FCwmzsXIwrQsWYAm2iaqHUpx1RmtcSCZcKHoZ/+5hNOq/bjEbc2x2Ikmhp
BWziwtLfaiOnZVT37Hn5U/de/V6a+UmNBJcPvWsZl/qXEvcDgUy86eWml/BUckr77V87DjzPgopw
MIvUgZ6Sv5uTa0T5drwP49qPYLWTKvz+QxAESh0oS8z/LIOaFAes950oIQhBHXGZ0uuWMBb2J6n2
5HCYWT+TSW+jSDU0DjLse1a31rT4MCQzRRHuUrHnVIfCA+frFVGnqvqle+6sx8/Y/GFM+4a+BOLd
vMfk+Pb31rwzezqc+W+tfMjnjIPhUimV2nO0GwJpd27XqlqSHfDb2c9pRa8sVpLdzlIM0QR1dWlS
e6QKX06g6i7X5ciL+bG6VFjPBijY/ctUIwcwZ7XE1wGD+9tMRxF9gwgmqXBilf5PJK7RAxb8xCHB
AFVhRxnjlV8bjI44SbnOHJPLp2K/lnvmKbE9qN1A6tBfIddqQGvwmRFx5BA3xvL7KXbjDiLYXraP
tjgI+56Bll/XbFytcP5/8LNadR+kV9WEedxV1ondkUNNdzJPl/wJu8crdexwdiEjmzmPOJ0RgDic
4KJsNNH6vP8oa5XZVNxZNYhO/4XL6GohXYjZro7LNNaI3J8DTI4KQV1O4BnhEUH9MlyodRgTIa42
WYnWAbABO8hBRFDRBML5SWFG6zalkg3y1kvEKopzktNEMHu/htvOomgnQ0dgdxGo2GXxm2IAS3jv
WSBLZ5lVBvKD42bTci13jz7vfBqcQHglZhx/WQNFoaoHJy+DVfPhSaReT96mjQ4cuYZpH4cO3HwC
Tt97zDr4vMCvQ9kdhK/Y+vGzfPDnxLqlYj7oDvwd4zt+vhBKflhXxYTijjYp+zpjMTBlzY8aPuxq
BZX4i4kzfqqjc50f1UwLdNYh0l5okhXlSslbNQuouJTfqPuT2Bqw2PXPWAx0arhYOKTgJKatRBGw
KXUyTXmGhXgFxrCX+Aoob842iQ+eb24symuq3mBug4q/9L6tcn0s4AiU9pD6BaupAHNsJQz0RJtw
m75Xxu74b59++Vy81fR0gCXo9/Bi1vW8JrMYfTJhMlaBa7LE80d2X8lMtAhrdqUAsaT97/j/34oH
6GwziEpCLJwGL8aM99SJwxLbFGHClaVbtIouYNHbwr2tnjkhP2UOc5y+4BCxxQSoesTdvjOE+mvJ
uhPkv878gYOD+SEj2u0g6xuG0yl/VNuG3H0laAIzKlScs2zQriA3UMsU/JilBmBSDAqSGLwsfPTc
g2JlWq+SdZmYU4/lCc9voKKotFLbrLGFeq1Ylg1yEXBevnfV9SLLaMxiyRCdDIkigA5x4gJOHn4H
cL2G/R6fwigf0PUWCN2tF96DpfdpAcIKTr3s0DHgTKslEaaQiALG23MAZ+QKASjCLWi7WSnaRx3m
qM03xVGt8RTvI6V826rHtuacDuO1hbM1rroVqdyC1VV2NPoFiGnDeYnkdtckXyWWnax27rzym+2B
rMhAiswb/rmHCjplQDK1WZUD5Lw4Dxy/1RHiK+F0saBT00HKYY/Yf3JgzcjyOL2u4M52NqkEBkjC
PWRkHoK3gHsZp5ZjLMxSNnTq9apcT+c+haLx/vG9dUeuCUj0mlbTbN1C1K6JsllsU/VRgPvUPJUy
Wb6F86GOBqlFUAKvqBLD88k+osDP4cW4jUte2labva1qLZRF0KxK5bEwEs+Ln04uwVjdmnmbYkoU
ye8aeMym9r9qAuMcjAmO0JFhHpl9VyYIRKu9rKhxOHSh/79ezVFkmBdFErAm6j+AqbmYT/JYDAtY
5D4KG/wl3zb5K/xfAHdHgChiQD58qPO/O71BChkfpFsS5pcDI6WgGucEticgjhge4J/Xbba1YNZl
7YJ2K+HVn0Ud8VlzgQTL8XBrPAfWKCWd2IegEhfAu26CjTpaQ1fZ+Q1x+NqxNdkAifuVEziqscxn
q3wbtqdTV7GONuVR9d+z9hkM1LXEUVLcMA7hPDwYJgGH9pROofeKRUhGhTGr2e28rL3oSqrf7WuT
4rSl5GpUSKTfrNZG/AJwoCCZLtRvz/uoPgsj40iePXIMkFXUY43uSGsO8QqlfpTdBqptqXeX+G+m
PdsyasV/+tXnd9o1+Lc8WYHJF5byCtUTuMJ8vJfsUYxUrPtN4D36rbqgiVrvHmXA9wkOdJHSm3sh
zFS2GRodcIEXVWrRqbpP8pb0IexvrPFExEWoH8+4JjHT1hjw05OFu7Nu5AfDP5g2ah71tjP/hSyC
6BHGFHlkOKu47pFPneC/nh3vMAlPZ2Dh4bnzGl/vC++Vta9xfVGasraPOs2wVcYm+V+4B1fPtFzV
qws6MoaHBcFLuBrITGdNljE36uGzVeYH+49E3EzTtZks6UyAds18+aurTC9GvgBZBLjYQFTS5QeJ
n2GE2UtGhHYH/rLCW+LbmbpKFzRzBflJvSRzcGpZXDVxXLziQhOmGPuUP7Gv1hTm4QO47VU1A7qC
mI/hWP1LcattwPYsMTGxj4k66CPB3rLLOo4cS3NIbRPBqZyLK4AlUXG6WHZRTd5B4zo0gOLulViO
72dBQr9kbW2WEf0Xq93pcB+XSFGznTknI6BG0YKaau0wCGJemBEjyvKgjA6NmPLUpWMhSRYanL4D
ry+E6RQuFsy+H8T8GVunz+/Hq8d5QurujMn1PyR7zK8kBzvpDusuFf/F4l92Sa6ui7HXANQtnVrR
3s0E/9OoaOq15nxOPsAf9u+5ocHHCqZWJiU7hoCvPbXBgFMEfKJIwyefNPY+cscagTJ29ZE6/1+E
vgFr+LtYILA356vesBHXtiApoOEQ/HIXcXqtoW6zwSqm2gmze3UORgc9iGg69jDxQiNXnqY1Z+ja
G4uCv14DnIG3BrRrkVQbYpeU/vr/yp247C+ieeGjtJYAQ2YKlhnNra6PeKVLSBrFRilnlLH4lXJh
Ab9lv+y94xZLji13UKkeWs7/20CDY9u1641HXa3Z1WLOgSdJFSd9t7OfEgSNjCDLtxkZDkZvFUG4
lqa7RmOszQGT5WfpcXP7zZV2kf84XQh5LPR8aKUT0w5VcuBlsHdpvhXewbsfBdPVwmDVe/5ahBpU
Ntv4Hf65BY7JWGAgvx8sxkLcH+ChkKwgFqQSZmPwBkhMwR01frICmSnxjddmFHxFVWL9mLZFhiTq
BE4pzYILuUdPCbqdmZ49lKNMjJA4OEXmXC6eIXkO5g5YGBnVB3jORDHFks/tdTUCR3anmwxBp20I
CYzP3403J5Nnrf53UipV9vUv7cko0q+5K8HShX5CyTVcis376rsYUK9pZLRamzSknifRn1OyEOXt
YYwx5UunNNFcZLmC149KwcbuTe5zWZJtmAlKY2OBZeOFT0w4KdFH7KLv1lyxXo7wgnbf8k0kEuJf
RlsWzMKPnA5Z+wbTmIOsND+avy0GQm+de8CM7pX5AoRYgzdCMYfBwf6CiPpua3r48i4hkA7gt2mE
6ba0qpCY71M8C5erxQlEKOIRHzXItwho8AwBdRKjN9IFnf7O6gyfq1ej13iTzQyycYf1OHb94J0Z
CvrPwY/NQeDWLCQZjeLU/u+k3TqKq8dePFuMA0OiPxbl/BXo+XNn7em3C3BZettbmlbf5p+z8oWp
YQUSEma6ANwg31ioKN0oKPOIAJXq8L0WpicOI49RobvpEtLXY55dY5QkFtFelDc72tTmlJmYsBDT
Yq5PP3g+4hGhPmT+6N/t7zIKNUerRtTvz/snJId/zx2W/3ue8yG3unBdxsd157srJK0OXGX20ClK
a+FvSYG5lobw/jhUwSb0tC30rvb7DBOFMnpIO5fuwM1sZYv6Xk3gMwI9TUUGLRv9Y+chuozRVV1B
PDyyuTOx8lV40U0xUQf5nr8wKsSWNgNufACJ6JmgsNKa05vV1LRDXkOswNHiOCw9HYl0BJLe2o9S
dBu+f6jOhn9XJLR37cj3/VFBdOuQMoRZRM9q7wnEgtMy+1Ftqexc7MiBwRayMtVTFvbUerV1ZTdr
1r9tW5z/N9YOC4oK5DlQp681lZDN4+m/T+O9r4wM4SoQudJtDZ9bq9edRK1n865YkA8K6udRVDE4
ceqWA7VEHJ4QFiAChULbfbne0E09nGlbPTf8SIG2AiXyciliKR3de649wG2mkUATzCNuGyriUM3b
uEgqDHHJpefE1/XZzWo1aBG3LXLdwuLOITV2QQOZphxiV4bN7CcBFE9KhN7IRa9VL9cW2sZhKerE
3gJhDCaszNB+faeii9zd4N+4FRq8EApm8QWVpUcRHNQPYk1rjh2XhHURFeHKh6ZvJpxldCtA1UJk
JQ2ujbvg0ugAobDNz3dmiEuGW/qD1iUTzy6hoSdQ7lFuN9GGfOSAm9bAlG6OoSUUJS8ncEce8ibO
w8EUDX5UhJwAbNYuup2LbXg9OpQ4aqSpD2grUVPDE3IQ7WQ4vTWLHYF4CGExurrWKQKvcuit3sVv
4TF7tWVyw1oZ2A4o2k1pKVsgTFkahGes+t6Oc7xRakQWH1iCD6k/KdhQyGJg5DhqbXInUa5RrVAP
Mii+k3E9Fg/Hr8it8EJHNvNiLvk1AdnqdDBEwNgWpPh+hgVRLhp1TDHzKgriyyiqb2T2t4qmW7N8
0uethFQ7BzFc/AqrxxtoV6BG5LYlzWezuSddJut9n0Wlf2TQNm8Hg4YtSJfO32wBiCWB3DFyYG+y
vbYKnI6aC/DqIIYB4anpNgbb0Zt60Qg4eEf5XRejWqVBNPveBVW9cZWM6js3bu7bStj/rgX8uNMR
sP+qiKr2YAW3EL2N7cL0hezq2vXFARSqfA2CaOWPbo5ZVaFbLcxSNWkzUAwRzBL8SK88xSk86OTj
XecoOuo+Z3O687uFmmWWTOZcBtb5y6c8mx1vAEXZ0eks3R+LcTu9KBx8osUzfi0RhEQel6L2tPl9
W10v0YyIwZOeY1CBy1Q65P2OBEAw7hi/THK/RaXoWRNpazeUxE7CpM1GsKnbbcSlxzJqJNg4yAZo
CtQUvXN7cwq9elLrbspVqlpn16gRXJrfjTFGuvxOFWFgk1FtVl6FFXC49gvI5jSNhzswVyf+HCPh
8Lalp4dgMWsrCzD4vQ8NMYJBG6FzoOMj5sSdTXHte75SXODDO6W6EAweWOOu8X6pUdqYnq63t76g
9vfzEoAVmeNk0CEx6Vi7i/F/l2R2A++pim5g5R/kneHBomRSCzWjMrlr+e8qypM8nO9+8eOFtOqw
+WbYDmTwZvVU3on+sOwKiUuMVrzXlKMdNkVRcGg0UlFwP89ugFxiKehat6JyjazPPsRlFbL52Ixp
fZIJWjYHHWArF0DtorEMMReQPrDSlqqryZBz2VZ9k2qLDxKRlgshjZFKSOEVk7igedCu4FntxiWO
UUNFpSo+bYDWFp0OdtrrRfU5RsR+024HrMD+AHu1f+w8wc9IBNPCRSwyb7PgB4AIwNwtvqHIYV4b
OPAPAWlabwHhPCzynzwDXrriYFW5Q54q+d8/It6qxjuLOJJSl/COgn8cq3BiaP1S7QxiIKGGSrIH
MunUlIdNwDhwfxpHLNNiYwRRjEuyBLk6LU6baVXYRiQjiJU6q9v7M96yWyrTjavg2s0Z9DZvxwMT
O1KU9hvUMFmi5lEzqqAyxOsdWRwZx8ioNFDE2Auq+yHnMrGwYN7LD1DlbLpdXkaYWzDWEJrM1Y1i
hS9thRDILgpR5cGhCE0gbkI203C85nyxhEgAzhaBw9PDW4XEM5SPC7GZDflr/Lo3PgBiBbluhozV
KUQNvnVGWJ5hJSHWcuDbovWJCnHztV7Us6kp2imq1ocr5fdsuZwXfu74X+KRf9UFNox51Kgm060O
vDtQpE37PdSjd6NRKw1ZVPEn+fZpNyQ3dCSpo1LkRHYobyDYgMF9unvUOOtn5BHHeMqrAujaM+s7
RGLvfycWeZJOZ63rolT6+lW7skGlpNi0lGNuEr8R7rVsbBd2J0Qo+W7uPkqUtf1xliej4TTM5W/y
w1Hsnd3IhMSW/9f7Q8QaG0XMlJGv0Ew1GpqJWT4B5j5aahUQZ0lwDVTct6PjQxzhmKQut+BA9T0u
o0zhAGxvK2j9Ys4Nz6soiJYXvFPy9uwsgRoKIZEUuRL55+UjPud6yfgcflvBHbo2VgTaoP0JoFQt
I2py5hysmFYjzLITN0OmBQKeoAUxMRzbX+1lC+mYiOl6CDlRFfB1On4ONT9VzAD+JYrvdjTSK7Dt
3CBcRTH0L7QQV/pYdvuSIjbB+NB6o4OwlAi+XalHrlt3Cm7aSGdaNG+qULgMH96bPpnvSrZXdON3
4+XgYEH+G8kNrORTkxzmGqRh4O55FBfkCBBaz9rENZdYpwPkzFMkTExJHZjOl1ofRoJQrDxbp3tZ
Q7LBReKQlAjG9FTsqtTG+wnLF/T+bz1MClr7De9qjk13BwYmnkixDpmYrWdv3k/UNfRqS6uHF7Ll
DZNKovIMVBwddAQnCejropFBlUAg6kGtNVVpnh/CoTSan1s0X4PG5PuIaCFCLz/Lhgg9lhsfiThX
ZhEVmHz7vFuNa63ztG4lvab2Zh0b+Ly1yaCj8i4IXnGkJ0GSmVt9WmdolA6z7YtVqY1F/G3lb9RC
7lZTWeIom37PSnng45WOMwivqSDVEYvKOt8K9opPDa5gfJAI0+u9CJNxiGRnSNScHQOnlwuM0E9k
QJ5LHxluE9cnOIig0xzpSxapK6YWTRow0rwoqHj4h4RkAErzbUuovbRfE9uycYOZMHbq5g/sq9/z
GPycFO/xgvGRRwKaTmEkl+x66ZYQQct1HAEZotb8yTqw2pnee9p75gxAeMUjWCVtDonwa1L13Bpz
Yx2OFdevq0Ewh2LXoe2gTFKtBiNM2KS9DFxgIfKfBZnhZUiVLUHRDgAja/tpnzc3oLGpKMImjvr7
/qxQoGeZOUuYNXsNOWSrtzc47oYskIbesFXKMp+Aa5NSYlZpBBBW8s7xrU477Oi3FlPZJ5XmV8ul
yygFy6Be1LczbPuLEbyuPqHO8hq4qjFOfCbbxmLpes/BD7z6BFX+VH2V0bdEZNd7IDkGLuKYjgvW
sCIrwBWwbDS2vnofVQyaIAp2wZ8vInoNHq0y85YSA8baUz6C7VC7k4LCza0PTCwxWGZOg+4ne9mq
Z7khMrhuWdfgb9xM0i49jZYTMNqEiwaK3WXkeCor8q3YIPyxwzy0cqv3KvQMZpHYCTSblK4QNPQb
uvg/dRhwLyrdKHYYbxZhdLj88eLFEaXlTHHk9H3lH+FjkP9eGljI5PfxJw0hEC6iv1x7qo3oA2OG
squc2hhblbHGIBpl0LNmNGyqz6zYEWcUVPAl6nGfpu5nHTUA32+aJw4EoQ+5iEX0Q8WmSBjhxQXO
4aeGmA0VzDKdfWoQzb0/E5jayR5Bvgk0cpNxYhkYa1orEOHuKiHU04Z1C5Vt4w58EFw8ZFRkha1i
kPcE1dNrzetdW1WpY92QbWNTN9kl8tornCb2i5vV0JXDPNgJVHBgYaVGOCjIt8cE0o2gXVSc7klt
zc4lysGMGW2ltIlnlqInvsNzTqoHSFqwHW9ruuKm1MP+78jdujMcr2v0ibBQvHwOOaoYiG6Ajmzj
/clbal5uSzFe0wTXbVWmMfr6HDoFvI0Ewhh3EMWQ/qbhoaZAtklCS61Xsf+bSB4Kwea43UXR1P0H
z4lI5RVX1VvGr0Egc8dql97PUO7a59WCnnbv06lNIm8my2xnQnl8sUP2prpM1vhMGMw8cevhGGXW
pOeeobiv+vTzT5RGJAD+D7UPxrgzEQfhvaAcs511cJ3gwhbFBxa0s+6HM8tHuEkW1jJX2tavvzKG
NaVlv7kRqZGvS7IXkX5eT9h9hTfY+RWHjtB8V8EzWpYhmGXf/j9gNUQYCPmgvXqaa+Cv3NKJxFW5
hFPitlaoskUxSAQiJJjsyzCnd/ChKB2HkQVUbFNp88aE38S2bxvgeCiQZW9YIshpBm3ooMyru7UA
QR0DUttfdTQplwbHoXffL7CeKrw8mqj+N5EBy/fLmgb5pUAn0ypTqKMbEP860wOQIw0D/J/lcM1B
JckuW3THGeTV8bybjknUJhT04g7rWzfbiXo9DuyFT+gl0vuC+I2KiYjnNSYSKrmaakpcPY1rxKCH
lv2qNMzI4Q0Nw3qtaLpm2jsAhtvTSAftfwlM3YiZqajEKQ2R+c9u0G00BxoRIDNRU/iR6421BQ5X
M4fBBE/v+EW+zSa2UQYuABqYH8f1MxxknFyto6DRRuehDqiKy1qNI96nAdGjsu0u7ZKdnoku9zSP
+O9kaEEfdjjZlvZt+abD2YSd/2Z7dJewkaBR5FfUMiJtW7ZeMuYFlop5/L8dCAcMfDbKik+DAGT0
T9dbrImseQ+DH+zcLFqbah2JdvnycUc6WabUDUgKIFIAoK5RuAdFs5OSn0Cf/jIHXJlJnrYaEXZg
09oGaB+9fPcbngBpn9EGs9SKheXPraqGYzEPaziZ2uUJuKymWWBzkDKW/R8GqtXupGLqnSVBA28W
t4rvolXE8Ys0p7QLmG9iK04qpp3TOBR+W2Ky8wrjqk3KnN+ex1gf4RllXhxfU24dDzb12vAHnR/a
s517K8wNV9ARiRdVTnCtQ44fsb4hAmubavLUU24EUAkLpBFXvMda7bJqJhWvDCmSk0qDmDgcTYXL
w5Klz9aDXN0VPEdfHU2KShoafi7f9rkZnHbitw1QdOSdBe+p0sYynXaDT+u7D7KPnXjxdsLKxQcP
A9f290JjQ9oOaMbIJF75yM7pK4HYq9yYU7pfnBruvKl5isIJk6fvr6rewBqTznl3Z8uRNHHH8QPk
wTGbOd0M729Uihv6xagurKrk5kjdEDmm0hfzdtk/oUNwzex3rDOXV9NKWj5J8Yik2XDbfaw9oZJX
l1/DUrMZUmxhupnvpbFref9Ms7vvxtRchkHSJ3auyo9SpfuPoKmSZC6EAOSM9IwUvP3R6N4MD4Nk
gGxf9R36wtMPwyeJdoJkj7KB+6BVU7+9eZYdcU8gDRJxd9j/S/m9nWxKuH3ED8arDgw3OgX88xyT
xrkDAxHndeo2qADW/z3rH1NolHC7rM6Vik6ddRn4ZfrxZOoha9idm70lXpgrserapgY6GXoPDq+k
nXhPuVJ6D9xYAxROMcyB8XRz6p6sOAL/ApidLi0lOUHzCNelieWbGFJIhXt/b2URgNyY8+nkGOn9
UyPoVIulSKyNDOZ2/V3jtXi4cF0g7oKirLL4bYTrcR5da1WpMoxT4s97h2E3/pIqxJlmkU8fcpRD
qZsjli15yw0DdcJNdClpRzGVgx2aRcOjqpJ5xiI3QcP0PeqeaXl0GrPxnPfDP8xxd86UIfBFZSji
HgdUNZeR8OjMI6lJtoAni5+1Ra94pIl2GpZJkDPlvKpUI4N8oouV+R95HgX1afUkxFx3AKLnj6Hh
9zvW7jMVc4VaDdCGpW8cNY5rP5Jf7FH0tB3cLHPyNcW28UV2XoT3f4tps7ckZ/NhAG7k3WZ0ChBR
TeIfPG0gSfv4bsT/W8fduMX4/CFT6PjXvPtKkfVQM6/BcpuJPiHzHWuBTyqnSaDS+RRBFjFadnKy
5Q/s1Xw9ER5xBcB1RStwE8EVh76sWvFDQacXIUwmTWYbqmZ+j1Uf6RQPzUf5MS5xDbKjSZHq3CrH
ge9FqocjzTqq1CQRDzOQYMCI8t0NUB5vpSHIpLGAYVmIjHjD8XocgIe03xU36u7RsSQKWFC6yWRU
eUuZF5fxDV/IxAAOIEqAwKBe507VxmAkiq6QDT9GY94t7BqrZIsR1LTh6z0cPAnvpV0Bzu1t7rbP
GrKKyz0Kol6r9esgXUfGlkL7RvlnBJe3rdSddHQmKNuKnsKr13YrF8L/7gyCY5N0d8Urb1Eu25W1
BQv7XaYEYkhlr5mhZejwuS5EqaGoIglieBzrQeX8svTita3wX83x3B8Kd6n1unfPdYp1DsDp8xqS
+ThPaYchpvZ7AsgumsMjO7/Hy5vNCTfmrLsIzNvi6W87ENoscGCQefQO8/57qP575BCT8ecN2Cd9
3X451M2NPA9brbxM8aplL3uu3wwWQ129U/z2axLlRxi54MoRu393xfUXuujOdvsjwMEEkCPbr8cd
5VKB295SkBgfM/lgQWc3JyEkiHVFDyp2VoGSYGI1+kqpVaKD46KU33CEIs7YFXX1vKadAYNLL0M7
qAI6v2WR9il9kbQZKTXYdctKrDQaCyG92eYyRQrSCuk6aYkIJLflbhgdE/m4yXYQsifY9Mzb/oli
KLYRFkQ3vtCc2bwS6vizWuj/rPUdYfVU3iMA/Jyn7kVum5fDuVCBKJPuPxWquKvt0PsTFz+F80Ct
/IDnZijWSPemEAD6H+q7aFCiSM2vHMJIupr98dtYYfiElmB3y0THBFhl6849Zyo3iRurnIiw5qXT
KQ7M/doskTwp31kay7aeNw9AKIEMN8753z03CQRaPYOPEH8Nkc+VkOdHjIb78Kq1Lvna7q8BpGFJ
Tmjt24Rmt5kTH+ocpGt3Hq4cEI8Mr7Pjq7Hhn3pl6DI9wtx7q0tN1mEew2e5qYoN5MI7obpLlhkz
c2nRvroBC33Mb/jbxE0dchPQqrStu/7E0meLbSQak80KqUk+8j2eobVI6f2W0PFDuugaV2kzBXqW
9Wu2tgOXRJyWaNj3Ow5guIFmPpvS9Oah1ZkbWGvnucwCrlrPNA8G+EAy//RAk/EZQTb3v27qG0nh
6F4LEy+FySELPTrEcAnoqXN5jMRQcjBuoddJaNHxqddrtXipS8ohwlWSR8lDc/0NkhFnLH0Yg68n
9Vf9NjT6zJ9awc7d/dGXKlxn0ZOf87ZkpzuXQLXPkJrbJOIkSDHUoUjS8UW9JDRuyKSWGC6tHY/r
vKhhWOIiFF4enxAh6hc6F3STMXIr5bT6UznFdmfu/Msh85tmn0bqnp+XiJWQ5ab5PH5TBDQ2SHzO
k6/CpD7WE6ZQDNscIvBK9kLPPbn44LXMVGoHPn/rRSTRryLTe1Osch7TwYXFKLo7i1uaS8ro5TlN
XBOCDNX+1o8MKEeu+nvJyfeRo8QReYTp3IZWSOc4Yod8JQv17k404mpeOuH2xTFDLWcE6JUCMsT4
sKTDOYxQfVfagANDDhJlA9SuqXt2mKb6KOLt63491IxrD8wsbHQTq/RJRURbpVCht6nTBFt60O5k
0rCqaK/n3ho7R9UFm89PIITiYx7AU76vddw1SiTf+8zCI4sBIhpRAshGYfgOg9M8isw6v5XtM+VP
s0PYaEhMxxFsU7gqFmbiTb8J8MXQU7WBGD2FiCEf3nVFmlTCLU1b2vZNEUHPfBGDjcerfmDkMrDI
XQE2cI0U5Wwi3/63ZBJ/pVELM0oNE6Mbl5yQxC92THrtsdCaCa7KnUy4vCnK3RmfFj5xodH2UQRG
vMyt+4t3tVQ5sS5hny+izDoFX1iUqrWdwfT7FvqyWuhq2rfWYIoB4I+egeAANbaqUZs8Kbs9tcL6
hwlFrKRdOZ7krEdgfaIn2XZO12EWRsHqDlVZjZmUvpH7nV1SY+GRCVRCKjmSpKhqmZ7PmWBiQlx2
j1QNE4f+pWUwCjR/hFgVBdp2sqMRtRvVXSx2qJNPbJ9Rj4XEpUnynFn8OtGPHCDcJVx5NM96LQ2j
aQ/AKLJTXLFoXr8AQaA+MC0AuTAhnGi7MgcxDXPthmOEGs4Oox8rZqJO8qwRI1Nz/AyVFfs8NPmF
znAaG4K9mI+15qoZhYWZNKka1Q+VRyozJDfErbRlA7vTm/1adGFPSsB7hi9Al1iw5/qgI0R0AVtk
Rqm7DPoxidHg0lmUmsjepHyq1Z356214iAl2KjZ9OJTrGtPojjTO2e5I7S8r3qigtPaoCJv/RhYb
aQGH8NzE9a0QFIITLmNpQv/wudqb07tRTHnSnRu8MJB2BHwrvvZxd8UuyK6yGgXc3337fCJ//ygB
ABYrlq3dz+Ktvq261Yx++l/YlVd2crqEVg/qC8OggAZvy9XvJTOsNz7pfUA5oBjsd4HRiH4hN5qR
pcuI0l8o9mStzIsuSiFjorBNzNGzd6xJ9z59LY0nkhs14E6f2OS6nZH1bSYDLDW1bZxC6iANhbDa
Mq4MD6w+L1lDSBdViGJFdM0T2XzGbxGI3Fy2wao/jpN2LszEu47NaraDPERrr/sHXGV6phk9IN19
slhI2EBaMdI5JnMAQUZzUP7AlejR6pCvMmfx9Lna6hl2xVs4Z3rp178xVGwBNbZJKXednx0ZJXN2
StjF4MUf5Ksd+Xw7BJzEE93xRpkcRP4fqdoXcVOOJIWr9/Bqn8c4COiTmqo/j8Jxo2l3xV503+Lt
PKVEtEJg3C1yk0qYxsS+TuU8Ob6ENcMUggMZ/wH6Y/1UQL5BS6HVG94c2jlOK8ZrUl7imooSSVgx
WwIxlE0PtDMxUmfTNFFXKWcRdqmQ5Ijt049NtCvC68xGNzCkaAgxEzDbd9RMajeXDIg08qyEsLqj
wMdha1eJUPMhpq8Wu3rXIsewEMDfMr5PE5c5y9EEwwNSj6sVOlGmiWPWl1A3o8ZMO6G/xVVyRIzr
dYZ43HJfCorFYTfC38B0fju8WbtH31KPlNyhAjXIpjunfuBTAXrfRYF5UOsdk5jHv/4Jn5oxkx82
GKwfDfFyo2C9BbHeUcbzjiY2u6NVs0+Fo2oWDl6fnYGo4xMBw83o/8RF0ETNzugC/1p0ZNNP0G7k
IHQeNNrWLdZPmV+hKgVR2C3pTf/SLocz7QigkBJCP0pQ4ByaMBMIjA71URp/uFML5itDywQvwQ8G
Q8iVssmol0+rAy7ET2/xR3aM90PqW+aSsmRHYCrAwIyCALTbhgJZXLBT7Tds8TK4E0krOA3QvkyV
SANm1b22cAsSN5kuFGSqlZtUnPB4xrhJmph1Bu3H8CxUZWXExuUXdnZKaDhe87GW7yj/KKi3P9Nc
S5fBsyBuaKpCH9SNeEYNJm7I9x1okL8Cs/XmgWV8g0yt/o7aq4mi8DkJ5Kk04vQ/lV6UlbdjJl75
vphVrs/DD4EpEooO3lpKX+OwLs1yys6pIVyJIwwEvMhLZhnbqGbcBYY8Ej9TamdtwoHOymhpEb1x
j/uovvG8ozxDkapebhusEVaMX2QJxlD5LY+7XiFG7FlDhUD3zgvmtrLu/Cb4ozyvXDzhW1XGgar7
7Fe8wrZczwL4VNE+xIMR+jyBzHhxJolOsMdLyeDe7HO7SShrJbLY3nZ9RG7ep7x0LCTTwYvYow7/
ABUAIzuIE3/rHmTjHvg/CwsOEx5SqwRaX5SB5WDX9pMLgpg6uKhPtek613+mSAT6jj+nfarusA1J
F9t4Y9YoKTcJCBLz6L53Aie4belKvnIg+lHwdchIdgp8EuwM1gcFKIew8F4RWzEXXf9g6zNDqEtA
VFAzQHVG97Ii30QrpfUa/dIgVf8dS5HKkkFCR0pjZ49yb31GBwr2R8wthYzYAn6OG2+ZUr1ZAV/Y
c/zSvSOrtYK8KAiehFg/JmpPxlTh3r2KcEgIaaRzTip/gCCqCDbZZvnbFLHpOh15iuX2O04JEPxt
8ARerIqW4219phzgiGNnq+1An1IbQrOFUcwiQtbWU/BTTvHA4lMEL68JTd6HGuiBzEfei95PtLNC
b80jMcNZ3bfLoPP7wMdYN7mGdzKmjknDs197uIhHj8hNVNZemcEpGc9yFvJXleAxciKST5/P7riS
UXC3XWzMB5C+jJQ/jdbYP3sTad4foVwLeTAiIYtkscxKS3IVqMqxuBmJaFDsZ17PIbXWhUKjN/hd
n/8qPwVpu13TD4MngJBehB0sO74UgeM2wzJdtgeR4sMw+AR2B2bTaixvjLwHhayocM1QJ3xUEuqi
rVyX/uA1TUqCeR6+5utOgt0rFjAdND9NHqEYRFccj+AsUM3TFjizWbbDHENeudqSF8XgY/Frb99G
k7R/S38vLM0OF1PTM2VurqUs+nEJ8XuJn43TSDzCFXO/4LiTSFGdIfdQOl48td7RjPjwE93FPYKM
665L8+5pwfe8I4m6S3zJnz/3kvfwJ0YxnnKH0OejWB/0kBjhW/vAIQ3n6hTuuNN7OfdPmwf4c9Fa
aJ6Wsa0XzbNHeNFx+xXDvkmMkzTJAb4FgDlD1BoCTovW4kTikQTueOgc1AeSiZfjtERrK8ZknseC
FvpNtLoVZmr7QpdLslpH2x8DyGB1boOIBivZlJOwOr1qXVm7sxL74z/Mzl6Ny6vYDyXd7yG1wt33
CdKCe0w3WkoU0Gy/+AMImvccnuc7PE8iDSTI91+mV8NLdhYjgvJ21t4oiBDPvl92gcl2t7wMgHpf
ELzsm2x5/ZP7BuHkmiUslKp7IiKqczWRzu9+nUsynXx01zr1sFcCJI+YmxqvRsS8ntpZ1h6K5CAY
LZcZaW3Xl26LXp0vAvC/5XgLhIeARy9EO2y+K2Gy8r0UPi9xMCOi/dH+U+wNg5sjppKJGsqvjCWM
o8Ngx48fzGcinpjWMl76Yd2lforObT1v0iGngFC1iY46SqwGaYj12gwfAACgaTaniLsCpDbG54f7
MaBv4zJqf7rDh5mjPzvqv63w54ACBY8VndTOiUu7qimAQ3WuDQT9QczswF7uTVdg/jUP6GYgET5G
28TIvXksiQXecodF+hJRTPzacUL6jrQ+Vvv+yAqY7a29xYQE72h25sIbVIljnM9VCJdULGPOpRlf
WPI1bacxa/4xEO4uUJlOWX7Mr17TMjhTb2gcEBdIHnHhE+SjT1A11HT8zOgJrm3bEtUNHgdqTKeq
YEm8GEcaDi4G6Zmbon39G9KuoXl7S56KzWW1RbBJ2OI4YzMBKLKlWaHy2ierUg765x+2Ih8pEJ4h
tKDoHsee2O+xgputOY26rubgGv2LCThCw4SYeylaReMTu3D/LyLNuyX3upV3wASxIf7xa+WHAN/+
z2Or5qJjTXXFxV7PIYd8QIRpg1bkMiBUaJUxJ/L9dKgrDcf53Q2xsVShwFAgAmgwOMQRyicCkp0T
jXfOCK4oVKhxe1aRF7m2FExQzD12zvrRnh5g9RVql8GrhkfDqzYfMCgLVZzuiVq2ZrVL/MV4hAu2
9EH2qIFaokqHS8MQzZirqoHelOcL79v5DZ7FtsGKcGcXqC6YaaoXDqm7lKj8CgaqGUdhyaZ6YY6m
Du+2lOfcZ6/ZEGcmA1Omc27SSOxDH68eKWxbFjiPGM8b5i1sqiN/b9moZaChITmsBNOIOJ5WWH/D
IewbJ+ocAXAXEiFWWY/ha8DbiivIwq3QNC7s7jt5MKtmqwpYKqWaUxYs0Hd0gf/YqOixh2VR2lUT
O9NmnjldHGij99rsw10z+nPPIbYh8SgLNtGrz1pSD5yKj/PuGnHFaWGa7G3LXDT2F7gv+kbfjatt
4Bnr+bjKnc4OyxmuTWUBLGaE+evigjajiuR62KqbZonTgvse7YbvjpynxPmNJpHOQ9sjW1Ilcqsd
jxczD6Zy0PFpTfBa2AYg4gtuRbwqu6jXZSAxLEbopKgdGf1fr20LYVh9kHQ0Zv0266I9LssGZHPK
uu/bn6MztwMe4QfBQKPMh12OVttvBZgNZSBiOPvuUjIDU2C/7/7P/0aJYRjNC0XOS20V1zNxCq6H
MeOme+9FnByKYKbF+BD/4dUsl61ZQA0v3/2+vVTO/ULAK45eOvKxUrbaOQgkbFvBfvX+hZ+GwVbO
vM58R2I1AW8CrIAYCoG0SI+ogfX9gdEMYidM6tF2vLAyoM8n+z9XeBoeW1jnWJhtLOJQZQoSBv+o
yT4pAT6Z9AxU8o5N2uSZsOqB8nUdu4vl6pBMyix1+cglqlbt+tISAwBAyfpb6gmOnQlVxTH9y0MI
+PrIuSF7X8GcCvcqfJQKe1ykUkeu/NVvhVPjd+VeshQQxpy3J4BrKCyn9Syx9+obvy5c3ajgaeZk
xdoLg4hyImw74lD7ytwhcLy+6fNIeVkSUoNYEAegWLqV+/iJW7VzrGxd29zGyZd6Veo1ZYUq8f8E
zixzinJGRRrTL7+whNfG7wGcUla6OPfnLIZd8Qled/3gfoQ+nLrjDr5iSq61gvkDHqERQLArmxvN
lFs4KjtBYSdQKpwcGli1Ss/jvRFtlwCYmPHtGMuJuJQRmM/MAyLup+lwj1jOSCI0o43oHBUW69xc
2biWOjCgXFay+X4AvB+iPiultTwbpCCIMQpZo38sEtJD9vvVilx0WoX7EuywysJtQj76jMWVFahv
ZRRdXg0aHgW6UX1i1skLz2DlkjCytXhnXn0CTT4ODMWa1gYQstYHkb99MMs6h+MFlb7ypuJryClC
2SeV8Nab/83ZfzsNt8DqUhNK+zdJggd7jecq4No2JdIHQFtTNxMm6VlFkMnI7Kh/0hbnkYfQ6KKx
9KVmBW1p7bltzByQFCxF+WEqj7ncG/MVbXjuCMJFHkUpfQKDwuOkXwwbKBMVbsYeu1LtMr+O94L+
LL0/29UORHKFbM0YChwXZreecM+kIXKhyXeCPAcGD0Hvjv+RVbSqh5V0faFzae/N0T8rNVZyTvJe
KgXVYuEnQJrrA8CrylozDewZUcXFg8YLAfy6p3rf7s3o4KBKvpTVLtHaEM1sDVYwId8UrxjuJ4B+
FdDqOLC0+y4OPca7/WAlMM7X0m1LOmYZUjYeuZjlwJKxnxP7z4h3/zM2e3pF3ZQmIMWgJ1vjYDJr
Cj0H86zVTtECpBIjGFVlHpuex7Ld12gc5CiGF96kPgc39KMSLm9bxEglWvaPmaPXhWaoEZOXv5px
h/VL/CAIv8yGSpxvMxDHECLICMV2qC7m/dxRRmUCJmEF4BFoQG1iiiLfy8ZI8ZB3oXJ0Xe4p53c5
Doqo+BB1W7x4Op5F4p5AeLLcnUpIB7hJhps9NQYv3SrViosWs/AaBf+TzJA8X/z+O5SL3vjkOVBC
9rYxSQaU/q6u8l02gTuX07k+5w4O+ORhM9DQ4x3/nN9i1Lq6ZLbcfw4cH8IQ5BNJ/XU2BRH6Esxn
3l7GZlfjhiYMzYriv3k9Ol7uQzAKPqsyqNjOdIiIj9Iw97S5HW8eQREsyjDjZVcVWcIboaROPgqh
b0B1wqjRtLmMwK9qR6WxukKvCVAvMdrHwaXL6Uuz13EKmSnH7KJ6I7Wv69G0HwoVbJ4RnIsqc8JY
65oQZ9+U9zqPtARzujWIYK40rGSpiFAiLoAsM8dC+KU0q65p1iX9fSa0jdoX/a5v03bDk5WvjdiN
dqJOFfeGCFTagwsFLyji3mYFXozMGgkhQURNraAuPxDe4ZCRsDMM+SQIx8BoKPf/r+p6ynLVKIvY
JFh1N/yd6+7j8i5rPj9Vppi0V+HOlYFmMmpJqQLL+uSf33Zeor4/GtBTo4Upr5mvxaQvjn61tjXF
5zZ0pZ36RQVYh53Qss+LhKCcNz7FPuv48yte4ALnKSH0PtW+GquUTwjDAW8Q3btnT5fwV8gPGHHU
19XADBFbda/UbRVGgoVPlD/Dkqpr4LqlY08biCGFKujxHmdqr7W1kULBq5eiUDff3xmqvhaOEhy0
yK7fJ+xTxq3pxCMrdX7PeguBJJx60MDNIt/M4l/JsWS3TmFkSboqEH4CRZsVARz67i6rDOHfd51Z
Ob96rkTh/IcUCA1o7c4yGcP7umP3ehbLuZtf2/Yu9Fm2URmcAAe2gf3ThzKKEWojnKeRhBxaTvD7
FAD+WOvFx7YOrJGJx7taJSYwBhpR/vI6oIF/Ta+mzhpu0G0abggShRgjI/R083tB4UyownDm53YL
th7TPoEZggpX3QK9e9RBDmDrBt5rf3Jm8qkBvC0YOkIFifteqJdBdCU9WToAwmhALNPbGdF5pTP0
12g8yQVPvSM+IlOrKc6WW95kLkupmTXRA73ZwH/qCwj3QR/bn9gTMbTuxnA9lsUiq1HeYOf43LT4
NxLJzOQjHvt3cRxfuEgSMeLP8P8Ywvj1uyIrCD1r2lB+N/dJr8N9a4LnyL+rGAZB5Y6+eNyb9jNl
mTsQPsp3e2mOGW5JCA0NNUskMUtz7qIziVQ3u3NDqBSfdIOYt1i8ZG98f3WVROBqkjoGKiuGr/CJ
pwh58twltueE/vIgkNecHVhDFQ5LYNlYqxLSMOHDSFESWJS2beP4citssKAd3IkFWW0yVFjd76CJ
ww8rKlbW/+XkMgm6t+4Vi/DC1Qv8aYcWg58RDYyXmHNcbcjrZHwf3jhwwO7NE/pbCKRaBOESKO/P
1XFFLDzqnk2CWyHJ8Oegvl5beHJ47l/L4RNcg49ksdKKTwpNPW7qvgfG7UDUaaz8LCw8Cjwep58T
MIBumPOWs4vzyQWWmz4/ImGomfu7T4riqZGkfmH3RTA0REOF4Lt3Y9EEZw+ccR5xfES+dLzGr7k3
UExVwP4d5lUHfbhC5bifEppF6pJ6uVdc8DaK1MhvITJo2bmpGnHrvV3h7Z0eAH4iBGWOeDlD4c6R
bUvvXXwNbmTdWWdjkJrp2LmnLNpsCy8ReerSidjffYDeddBUx0BiB3IlHfb/aisX0zCx/9jZUF0U
sIyGtGq8dl7E0iBqyVbdi3uoY1MOOSTfQkZypMKqUV3mCrlyUA+6z5cVQWnOvL9uPukMZnQAtQri
UH+fzPyqKTm3+ejXaQh9D//wPw40XRA4ST8ZU6MXjfJrlVR88TY4jzB8PUXec2qnLrbvuf0BhoqX
yJ4tz55VLZOiM8PjhIAiu/tnkkHpoFEibQlXztukbPmuo4YNNrcLhn2yTVhr6nKGE3FvPLJIlfkg
EmLGw05MDj0ppZPGxCcBcEbsMgMWXxHTsObMkdacZmqM0QCcDKe3zlAnj8sjqhQQkuDUL0gz28Ye
j6G9BVvp0As/MOrRAOdyuzVeX/q38MyytFO60Sd+bcVhnAe6OmE4wFVjMts5l/Od/kyvPuxIdIuv
duahTBH/dpVSLPzlXmEWwcL+VtiFWh/acxOOFqKfcCLGFzMt1/hqPuN5yyWaEPCU0uHJIt+arsg5
aD5Z3CW1fTaY+togiCs0i0CHTlTWKe6W+c/c8ykHGafg4pqGmx7C7NyKpknsujivUsNq0Ol8ay22
+nXjltaH7fHnw+MZDd9jFHxz9vVFMDzlaOQwO9dxZtZ50rLP6XMgDUOk+dEo+mlZoSIok1QCjkgp
VKcdp1dxfYywuAtPRh8To8KOryDrCUHlfcHpmWoGHcvPILfLhkeDBnVXJ6iBTXP4kNo5jprTqNlE
YpfdPvMYILIuptpR3I5PWh42cjSP3n50Z5niwmY/WVfYyEJZ0X/pcthMZZE+Sb1sHy5fTIU2IEWX
bEAfdf/wLo/F5CEn+HGlMlu+azlvJVvKswtlcxQTPLimsegOwx2PDeT1fY5G49OATpzfDXJKKl0g
ejzXIRW9PlyR86OfFAfRELcSl9HTCK3Fm6Jw/ltkxu2XdxZeZIqwnHXC1RI0TGUdZuGa/Sc8VVwB
Pz0q9s8gGT60bAZTBuOQGj8ZgqbW5HEq8MJ5K85tThgzqOwgL5+p0KHCDvW/JINcp/tuISaN51xb
UtwI6zsVfPnnTVVsDyC9/hP+YWwgJsT51PM43/GfLOkIr7G1KCLtkv6F4J3FYCPK3eZRycPYGycK
9bAn8/7smyZrE7I32SOxy+jpK1tVeMOcTnqqg0AEfoXvyC5BEMlJ1cEpHAJgVmioiQdHyLFR+AUK
HQpjVnOzNEQk4G10lDc9/PLRdcmsZUVN6ThOAqDeqT6YfQ8mOZBhzk5FSn1eTpVQPWdV9yaqENwp
UC7xe+aw16tjoMbScZS/RQRLEPkod0hcsRDXB4CXQjMIgsMyXCZjW2DVEiCIM1Gnv8VotjanpGPu
vMHncypgvemI70SkUJMAatAY7hgtnTYkoqrZ6pnozvFq1ZDNGIiO16lqhsXtbEs1ESqYgfdY9TRY
/UE3YIzgcpQA/Vr1DIWZzJYqHCJedttgclGPPNocK2yOPnOShGO7EwdAa7rI5gUdBCx4J09ZTD3y
cth37P0BYayQHFxFRvpRitrzq2CIaCZgB9/MA5yoOzvpFsMCUKR9DJrhpPlbx12jv9TFu6hyUfzm
65ifwZR0koBvfdOoxEH1FSJHhyJJ3fCa6DKGWvwLRXcKZW0goXXSO4lhOGOHK4W6mnG9S4HNFEyw
oRPmlbhMp1noMM6ZJGgt/LBfiL7ZBZG8/mDTm+kZBB/3jAR7PpCWG0KKlExGgfxeGSRDbw1h7lMd
0ZZUeOso4TzQt9LljRGGKrfWd26AFbtwEw8BkWSq2xOhlvwj0lGBoR0kdE7qHPigxAK1B8K8ddaN
Wcp3TTf3ayzYD2vCca+GHguHfRCy+6F5VKuB0cFkY/s4LwgKRSvPqOa9UR9Eaca67jsN+9Rb2L79
XENWB9auUbN014Yi742swrRcz8m+d/KakJDinaU/UAaGgHDoXnsB0fqGFFqxGALLx1KWQM8yzma3
nBDDLCMrlbB0R5687tRTHiDBAwBJMHpAMLeyqRhuLbr18CHP8ro5H8J4Tp8gxT6twN4P2IZPlcNb
gSggrtCXNg7bTzbU8c+8lwh+lXyzCaNicFNImjSrE+wayC4u/dLLiOkZNT0Imsh1F34NhwjX4KFY
L3v60nVvcbexC6sl0F38Yz0lwiQTlpR0gJJskZXwkrdmwG/G7PBmtqxS9WioAPKB5YawpThr8tVQ
XQCOKVZ+LCzHSTRz1NO2EHBYj+303rAX6pEXrIGxl/EfY/vJ1pmG/3Db0a37shW2F4Nj0o0ErAw6
sE079KMjZOFlBiJGMbHR4asWYS+5tHN1bHRAVq0ocLg+zEthFB3n3XDgM7rkGjn15OTB81C+tJkU
M6QxLuWzegGu/Q97Bn5+FrJr1Q08o9E80BUdyIti4F2mNg3pX0aRMv1v5Q3lRcZyAdxAdV8WFLRT
ilTplYs1PGyS3OtnujsFtikTmQYSBG4/iswRRAcabk9IxpXSdCys35IX+7O7U7BQVzK3fCG64Ntw
uXGZ49/cvv18bgvNBGmcWA2ao8izjZcbgUt70m4xozNma6hy46tFTh0WvRwjuize1h/PPGezu/ZP
H4fjO4PQd3IkSnT/dM8xul7OpaNhqGbQd9evv/u+OLZyTiAIhtNBa2PfYM6Hu+hAe0uoC6VPr/WC
pDvbnjGG6bg0NVv9O4jHdfHH0d5CbhWsVfoMFU2++Bx4LG+YVQRWKvV/MMkNwxuVQ3BKmbqI77ki
wAoVJ76N6aU+koBUS2Rgu0vXIw+L/tU1swIQU2P63GBmDHULX5eJ9qNHYD8PJirn5v9YiG/LqRHs
d6RUgpXrDT/zZZzjtpAfnfjCaPEL5x3sfIGXNuP2VGL9afhdkNGglafYX/ETH8xCziPABLd+sjEC
80AEZhKK9ipIWC7dJEEtVeYBEUj0IepJYuF3lzokqrlxT6pjFwJYHl0oojERB0ltEtp2ZUROjAuv
MZI+7IPZVeQXjRouv94HJSN+s6kxvGa+zuqkoSRslBY8GuDG7DcGJMPIfS5Rv5lgt9O2ALuT1AFK
jFIPsThJG4PzRTFFXgjXJYnWbvIQbhTHFXluD+vKPvIuEYx9ADT++3G+42MgY7XKwSEOyFhXEf+d
32YGYgYr5LnjD+rLmTUltV5WcWqEOnhvPfsTRsi9tjIZeJsUEjlHwzclNw7MqbJG9j4kmcnhaOrc
AdqvVRUr/lY0SV/HZMLlhlTgZOXhCH90d+vZ/TjndE8DEM97egQ2kgvIiCGe+4sgoPzWhNN/JnTJ
3fEnKH7F0G6meLdvRQxbMbOvzViCUA/4RXPuA4bmVBYWXxJgfNxuajvgWzhge5hVLMdcU0W0XTFE
Bt64KNUdZ1mfw+9VRMWXlB29+JfdfKryalttldK9L3XE1DPRvvCBoXGbXYTHNX+2ES2KbY5SC8Y0
AFTch2n/l3G6v0koScAmFuskQ7WkyCFbZOtz9fL3SkD1vByli63yRAekdgsUeFQu76wWIqAbQ8mi
XA17nUO37oqwkMM+HfMT2oJg3CQqApTp4aS6UsY0aWc/UZIUFJg2rOH+7klBL0eenV8T8ekdyG4Y
RsSLg5ipFJQYnoySpq7uLyuPzjDMz/OQ/TexjEyxb16Ul41nLGxADzeFxI7NHvZ6Yc4nN6Dx+f24
qOwpxFUEEBf0xTW7b17g9ekqPR32L3pGbI9eiYFQayLE/75tPZkI0salvZDWXBHxe8PODjdw8V/7
ooryM7CBWSb3iaIuJiDR6JBDWLjGoSNfegDbPHekln5nhMsUslutdLbL714RrqUhRKkVgTCh06Lv
Fu+geOYT8HtJkcB88vDdlby8vWoqj+pAWiQRSIHtU4GIqQKvtjnWP0tCLKsOHBsxdWFt8AEqDy8w
EUXkaed2xzPujSg1ULvZuusBvbR4IL8ss0kJNVgcHUXUS4VXdX0il5bBedt19yfSvcdZVd6FvzH+
ZF70brTTmgKJyz4DcBGJwZWbM+R+GqeOr4IdTmAQBLi4R3qVLFNdmDso0TyiiHQ858k49f1Ks3r1
E/doiJfGuVWHJc+33BNE+lAAspjjRiwSlJkoZA91I3K1exwcMjPFU6rNazaifSy/zyqs1BQ7cy79
U/sLjE5LZNHUzRVkkAB5x8Rwz2JRDi/zP3LQ1efONlJRJOPT0/KlDjXxaa3XkBQXsJvqbA2XXnTt
ZwbQzBOkAFDv9E8be7QS4vPtdEjSJDTb0OBOejY3bK0xL+lPTkxXD2kFgmE2iM5WI2oCajb2ycfN
J8kebupzE9hIqcHD7UFTrbs4gCvzqXMb3zOlNCvRtiJgUp+XRQm63+dHSh0Npqf+UWWdhhjXY0tL
r/gMXhnCXn2Sw/ys4XG9viwm3asGZ1m9N98aql47NyRp5bh1reekMwx9HStQ29knizMh0sY2pkng
HAR+Jh1c5sfm95+uwBCyIyMorfaaGmjuY9BzIIuZm60mLWo4T8FoKSLtCInaStI5G8B0JC/3L0r1
dwHSGSoCBvsKtgWCUbYjBbW9tM85MLaP+1zgMhGe1mE6lkWirAZ4eGtwdqKnaSrdGw63KLdaYus9
n4kOKQW2kqnN7HQnbJKBBwLtdjlBlhKaggSjdFIztYkSVs5tSMhxM8FeS/aJwbkQx5BVN9icc6DH
ZyhUlUTiU5HWCbojj3+/s7Hw2+ThiIO1AC+yjeU7uBMLcKzpEWp9zgARRyf7jv71zXyFAsRsp909
nIRnWkR8XS/P2NvVcgQYrgbH8Yyn5IUoEPOKBc7Qhd5FvgPo+setH0dJN6x09+MDWgb9H2E4l9mk
sCzYxcExcjyKTF21tGmHHlDey0L3qIoNumqrE/f1ZMXj6N7daty2c0sPAoHsI2sNvh5Lc7kVsl6r
hlOTY/6Mq1tRCsxePLvsq0kW8MXlZwuu75E5+Bmy8+9bmatO2RjEHq55+hxKkZpfnEkp6Vamrnaj
5FCde5+gMfrXUYsqJ/fb9RrXSueQXrzEEUm+6XJrvW3HPK5Ms9VVVObJkDNR3Akshbv1BrWeXUmn
VwROdf/7ycCQYaZcxSU0Bjgie2rSYKwIclX0qynlyDkDhAFjDhuI99yh3B9tkkDarMBzAvX0O9dy
uqWju8rXLEJyLxV+y6P2Gr71pyFi+wzWWgVvFEKJdNMNuDrH94gK1yI67TP6z+g99RsHpsxpTNsZ
OH2/+WGWR6pEOcfK0DMvLxc/Sosn95x2N9CAITqp164WgxH40Y4z2jGNibaPg4mMY6E2EXoGMEXz
OxcEPjqo33opHlAAnw/WmOP4dk7X17FGQSdZjr+0RuFX/1Pz/QGmsrNksrsE5K7E+7oJKpE+pLzH
Tqwhq02E5TeTxKCEctbLj+A+Pw7zNA1XLnuhe8omHLf/SDBLNOMIOfrE9P9vqRUV5ipY5uD/2QUL
9277QPSrtOWO34oXIw7nB5wHTeRQqww38F9oGr0BCXx6M22NiGGC9YUela9SCurCtBe6lS8NHjfo
fn8PaJ19RxUjDS/xPbxC75UdbNdeF4lIgYuJ/8Q/GDfKwraE3QsbWMqnxl4mf2FVcf1ZSdrUg0Cx
66Wpzq6O343Qwh5kdfxlRrQKrwcjMYD1mDTnsnMeKlbj/TsFApw8SdQ3lyz4VqXo6WACooKR7VDR
TS3WBq4s817QyoMvddeM+gxHjSkgux5AzHMC7TRnWxOFTtseEuQcy6rXyVNuKWRujMfcLa9knSRd
xGDGnvFS71GWo/sbderLJ4+aKMuUFY0NTE2hYcQ9OVmwuQzMcSbTwLc2uYZ239xYAjp9M4hgqgnc
MkEvLQRAu3XrjQ/QIQnU41Ae10ChA2dw5+qOhu/QZBPdTb/gfMkAG/gpsyGSrC9Kh8hrPx2qjEyu
WcsoyQvH5DApkv3sS1bedCSBFdlrl8TM2uQAksYDHSITDgqeY/lQYEQ/QrXPIvXtUdpJtPjbuBlY
VvP6+HsqeZdabTFyL3T1Lx+HFZ1MwCKIRwwxkNxZyn1EZ+bbql96rlJH16piqXqKwjXjSX0yVWG4
8xDXxHn+1r9LHb8e2PXRXAlSHEp66XxTcggfho4C43yS4kQtEQbiYlSil2zZPRuwU1Qyl+Fr9G2X
xTaSmTTu2TN6BagA+5OkMq4ZlwVQ4rXAXZLOKnAdYAch3G4NhDf9fmfWM+A5EqJa/W/QtoyVU0FZ
DKo8XiOrUm22inwEZ8sUEzTwlXKOGfnFtBCOx3I83FPLkSJPR1kxvfIZprHI1rLituDEYTxQlePb
0+ydkqy3QQ4RyLHb++H0olGyBpT+yBYIBg/LMBrr1LL4EdF6GGGeCpJ58+ozYtThbTjX5thHjCLF
1EFwQIVxpceF1aT0eqm5W+5vDNrHu5+P/gu4DiM5E+GWnxqhIMsxsM05FPeDivcsB7M2g3c1g0uY
5iV4z91WJJiUkzfOSKrmbjkJFRNjbzlrfaWlOxFaNF/gSrhMt6q9L6nqOzxMn1w9Q/njTatn+/Lc
q+zFmO1uv/tRB2ybXzEBmNQyYkObn+auSz5i4yu0Y3qGBU+d/OpguDTnKzafCLbVqptM/ZPv1YmY
Nxxw//Etu7ETFc4htJlw3kmQYc7cdrNhhtY53fORPACGQkJ/YMbQf+HO2qaxILTrUpJ1KEGmyx/W
64szELmkGtw71iQLEI+yCs4S6E2FY8yRFxrU6Oea4urOGBtOY0OFioUQzpJpRiLa6I3V1bA/fOxM
AbHo7RPqxuLIWx2UEQE9ZcCDiCWaQHtcs7Y+fkYqVNOzZ32EKUm/ZPOa7tyF3LWT4el0MMlMsV0b
8rFmlGS1oZBVvF63yGrR15Q/NCyodziPk56JbzpuaF5yxKhUcP2PMVR4fxByWfvQmYoO7kXD1ueg
bn29FW+mvN6FN5/PuDdCBHRGYXzTzY8p+BRCHvZ7gWQKk8K4u86bX+OyF+9vfOgDrqWLo9MyN24w
hsvOTrzmJc/a/YUCPaMLMHPA+zxqTLUGzflylg6yopRaJ5Mke+Yto742AhukaiLYYWxjC79ngWn7
Rzp5/mc/grQHXQpxMx7mOzuUaOsFV1rEqO4Gfc/iQHzRLjw1aiVpVdDu17UGAw4oSVH5L+0oqrg4
6HjVDzCgYbn4Ud88WvyC71O3IvQ00y7IxV4ZGYg9bhQ3RxMek1DQZque/gB2AUje9DERnQnGdq2Y
bdiOm4hXmlyEDfLicsge7rZsnwG77Z8EokWgcjpvkt/sZ6SPJykBRzYhaIXOHZRBf11OVLN+YAv0
d7/3gsXhj78f4LWnDOMgaj5/kyZZWojY2aEzvhYr4O0F8paDqtdlUnCyP+nK1xUk38gubhbpaR6F
dbUd0VBAyWnVsGgEfqi87Z56qhKv6s+yawEQOj1EsmmHMMWITmjp1+lVCmnCwwyjMD/wF+4NjnC1
1sxmscXxfALssQ4BSRYU5u2LeQxLXajeVl/NU12BIkB1yiKb5GTv1x19XA4HCYF3x1wL3aX+lWlu
hlLcTrhn5WzcUD18OmECW3E6w4GRoTeIeEoFXdgoVf569Wf5UrsaM8J016/Gp16lRcIaq9AkH6Cc
4ed9QtE0Uro9qdxZtpPWJNkwqAgZTl5SHr5j8Xs0eeoj1mgyGKC2aONn071b/Wharhl8Mb0GMKss
KZZU/LiXShIJMpY0Ou8kSwUBakR79sX++rXvc8o0fwARSWXKC4rlZCeeGMe0fkijUYVyeYc+k1AA
RXsIdNHtVSRaJGdAXYSskVfl2z01vAsrTGRJ8ipmu0wPSPbSkKGeqYUvT+t05NRHCTRhtkIM/R9M
RIoMpPQyvhfEXMDS9wN+zNH3F9YJG1zybR//OsUEyu1WJATKO+i/y5Yhh6MqCHFOM7/FL4Glk0Zq
rhcpGojOkCD3UpKMeSp0XMycTkMQyQWoRE3aVyjwND9qvcmy72lRQZnxf7AmkYCk1MjbiZ/IHZJL
/HsYu3srjI06VQSr4BV4XnQ9PhNDmmaGeibrVqWJFXPNKc2oMACas3u6iCcxgsOGoTUrcVjKGx9m
vtGlC1SNCh+akH2yejCNkZgEHN4hsH+Nu9Oe9Fr0oAHsVEroY2Z/sBlxIa8kbfK9SSvcoGzCVtBM
sV/WoVtm8ihKKnr+WnJYj7EtjXr8qdwOTrAR61O68R0WEK3yz0iUvld5NXuMqnlprAuutADbgYJh
F1XihU9RIr9h24hRQkoNn2Mjt3+PD2u9iz2WTz0BWXy2M3xgkVjZuNHuaRXoQhN5CAQRP+h+DOYM
S4+LBqzK5628l/RoU/L9nFjy1GITLPoSES3Ntz1US+EtiSUryvg4mlbT7i8QEKFAMAJX4nHnLhBF
f0L4W0RQz60zQhdurTm+hyfiRsahX2HH2R/dS/1Xw3vAstwwixQnJecO+5TH4b821hMoMhqanowK
RmnjdmoMSj1QCa8MScH4gSKzXQ7mvsV4RQMGDqabnoDwfrceBy3wYwNXTi2CEbfWtXhUJHferw61
hA0JcR7VUXgYHn/yBv8Ra1jyxft+sMGrvGMUBuQwXCPM6e47tJFSLang+EyOdPIJNhVz2D7ehHbs
25uVKvPOozwa9UMKPAL6M7OBZP5QHQ7AB7RhW063LcriExa0zioM7OzVNa6iGeGlOt88BflAO3Cw
lONT0ekZKfIqKwWtP0g31PatzTk57ws8cbmvZxOx4d4lEc1SaM0y6MPIWo0g48B3HdnY5oFk9CCH
h+KVIPj5PIARhdKKrnRAFM3bODL6wiYQs2NbaZtEA1OB/N2MGE3p93blH9uQoma48jF6N3MTeCNT
Ju3oIvpqcoNBc09oYasrkyXwsrEeMqTj/ZFDJ2Kn2dmXJBWDmkSXptDVeb/n2fYUZlR843nS0Mcq
W7ft78sfQq5SdzSq4YUF/a/zDW9BX6ssqfALtgiLXVtvVb8T+Yx60NvCREi+IKczLUZVZPz1Mchf
as/zHcvWB5aqAulsJYhpWzlsLdl7L75Hb4GUzUAwWsWGwFHYV1bPEr+AMsM4X345QWJgK/Ajf/zv
EZzSNAY5R5Grejp1NCaeabrJj3xRbLc74sd3rektgIjOXll27BYxUlxbn/SJb5dxhJkJbSPSZTiW
K2dbikbF/30jdPCH8Z570bXIBJNz7uRQ9Bbg11WvVBuPyu1dF7UBHxOJBRz3QJmbdv/tVkqlab8F
llNzxwxr18N5uAo4IWTnPdK17YpTKSMuUPZ/ugt4C3BfGBhSfWqakmfqAwjiFHCkynwyc+ZLAXGw
x8A5auokbDveIv4NNYmL0w15NkeXU3HdNa/qRyK9hsKOhfM33y2/A/5z+wHbDFVt9y7z3sBbK1Mw
tGHmbNkrSQlBI9zO1zi8QiKr5V48QMtI4c2Oj8HOCieRhARfRAyKCBkqYL9ItE0d7+hbYABEsVIk
/OwITpLb/GKbs9wRpXtbDqCF8ntPUIVJGYaLzVetq8WA+VGRqDm4PABLrizqdwYwnNzRf3SlqALY
ztwgNrvZXUKJjARO7Z7NEht8fblrHBKrZqs2pZUZlOku61tVZSyvxxvmMgeQ9Na98DCsQojISs00
MwikoqghaS5RUfUX290qGuUPZJHbTzcOqyBX+tJFeEYtOJsyph7bC9zr6ghj1uXWyq/xIbPpLOwo
jjIuiPWXEFYD2RBmP1z+ZO82CN6v/FLM0DZFLS+nD38UG5NYMo2zE2Iq8R/35xUVMVg0NCQK+ww5
CPMRy9D0yyjg6C2xXaIHvBRieXT42aHgXH6e7bhBlfN2XeljLgFKlsaeJ8pfOnTDc11ec7bPJVOM
FXLaoLfBuPvem1UTWlEN3Cx6+L52Ebb7WaT13qhV7VOWc3j/XgtmJ+pcin39HDF9PjnrZyihRFzr
aw6MH0MB80Yi9ntkFRzZYYlHs4xlZUGQOm9p6DB4s4GjpgqdmiDAEJIowRVKd9SYZJ+f3RpMQFXY
3tgG0GFxsLHO7IA+WkvvkhPcLoOpiFXuZWEYtopNFgQUEQj1HcM8lN6LKGogfwAigPQ1uzYcHCqT
hav58J6hRyZ1F2Ab9I207RwtrpgRTq4Gk1Dl/jfkZYUSC7ZnaGOO66grkJZ+WPohs6hoICk6FBHX
pPsBEu+egNqesg1xlqG8Q960zXzqIsp2Jm/DhYHjyOMS6Hs0dlg1s9LRv1yuzCPX8UuiEbTGOfx+
90xT6RMYsF8mSEedCOA6VOKSArP387BNSn5QuYlqBfPQvUgIIBnP8OhkpUmwAiV17gqlKYH7MizW
x77DdklY8ip0/hzznuSpGcUi9LhA59KitKqHNPVpb0qaoXLusIk95Ai6LISUYW2XjOLtU1iyjLsq
fi245+bXNVsM+MXj14oZlWYJsmODBLdKcSH9o2d+T1PEiNsHQMsL8+YGMRPC7XLgyNkMw5WpcAJu
gZaNVITeW0AtdFeODjbxf2TUH3s8XmCRk682lDhvaf4zT2DvA3c7I2Or5qjrTjEcSoP3pAbPsnes
8ritDAU81xkczouvUJxgC0BjoSXNFvDLDzHf56S+lBsJSiHFayAadbCtTvhxGOiGLq+UKCC6e+Eu
kaWCjHWJoSfrXEEGZSwQyVdqfsu/mHnrY5eW9xyN6sTMHUWUG7BKYfFgSaa3FsU41PZXXNvo0ATK
htBLi4uHpIybahuMfaE1hRdcaECDkKQp3WERjBuRTTjyIbnXLOnIfe6I0tngLf/YbMysROL5hZ9t
nZSpivXHco4OvVcETtLOA1PdMdMz+bg3mISgiXU1gnEUG0DV0R+nDwouH9ogvFuSBRZEXRDmf1DO
MJ4BWiovQle8iroFQY1xlNP8FrXxOW6IvT8irx2gZPqFxN2hedeoF3ImeY76AGvTOzCJ3wpW3OUF
gW7wLf1aI4k2B1TsyiSZO5fifIdZDTeBDuiXthEaIM39WRwF+YWv7bt9gMYam5HQPGOq0pjjyfFu
1Rjufi1IqLpA7SSDB+rsDPJ1FVvvM9fwn/AsMMU3F2xFhlqPj6OINbVA5rbCo7k5azJjstCfdPuu
wQlT23oe9SD3Jp4BPzcJUChhOU+os6uLr2V6Gunqcjcpd693gW7SZzXFI4oJYyveawWuBwwEAJuD
KH1GDZdE/fY64BST+ublCGplMhbTtoeYsWVIAo2uNtbfEX6qIQY1jl/ddlkzh+RyIFNwqOR4dr+d
0EwkAvFkbZX0IoudpDj/rJLZ1e+mwGguOE73gHGttK5gsGZUs3EJPZbmdNaVpZpTqnQOj2d2Wl1h
qK8PNfItAG8zbVW0Ei+Rf3uyIexgzr42cv2ismJyg7JifBdEbjs5/Y632a4ruzSum3jcMotSE43B
5iEF8n0Wdkmap+Gs8ouquJH4RoNy+bh1DuhgWSQ1AuR13GgJlVcwZgWzzYa+kdqpV/6bwwNkYrgA
wozA8Tv9SRPh9ujqq458/bNhn8hZzA02fYmYLojEVvG35egxbXOq+8w2n02FZ22YK/nFIspBRaZZ
CkzNnCM5fiv7cfV+oT6k+3maAV15Rztyf6nxXx7iEE6BwoTP7NhBOtII0M1sfPKz17uHAWevDG7D
ocogzk/qhz7PNN60Dc4VU2OKKKaG82+ir/uIzd9SS+dqFdyCHiY6xMexPx+W1oWFsCL9P1ESHsNq
4Xxt/4i7T6BYxRl1Ivk4ELJhG/q7yJrklSB8ZGqdDLq69mC9C8bsoIsX2RHTN0zOiNuKMIYCr/IQ
b3bHXSDYEeSboj7lDFagPYsG40bbOxa+gcjuakPfE5LwOX/nup9WFzDQbkXCxq1gVDYRgN+0mSsC
zFdB9r/PqEZADfpWmA42w/gkXvc1Hgq83KsE/pLItKoo2+zIewhq5rGXp7jD8ObSiCcN5zWGKcYJ
g5loH8D7OZ/s/udsP4VJf1fIHTCO2gosBxScYv5ntdAzHkBhBQI+YQuUEw47nohQs+qTGqN/7N+U
G/JPoDew1rcH9Kmdp5g7rsrIKcKkkk+lKVeBkj3btclHyvUgWYIKwPDBbYbjw3Jaix2BhLF1oBEZ
202aHhB2eggkymbprzn9wBPsU7MEi5WSV3G27A/Tw4i1johrp9NL0IY0uowauqU+t5Q5VSuh+nwz
FTrU8DJpnBwHlYmoQyzsg+z0rQf453qxHydSMKyiy41Er0o5LrWkjdDVIKRySaUpwC8rSf4nPve3
GRioha6UVSGB4KQKZ3ad6Qlc1Yf0ofBpEr2ryO8Fj7cRtze5WFESaot8rxjGcD+DwgWWxVpkhLZu
S2qF7oLkMpj/TpeH3TCJcrf2oV7jNdCZ1Ezf/kXNxwaC/4+4DZ6yLJt5emPhIKGP6X08HgleLD1U
qnIfmSmh3rNLcMfB4UbhYdBNP+LM7rfBwhJ0FMpBqoG+fNRmSAMsdNPISZ0AB2LpyAb05T2YZQvo
2wKQFtW6RIc/vTjxklJVzK1k8ztpmjQ80cQF4Okl3doasTo68N6u0CHwmkDKZI4e+qlKBYoMGhCt
SxHmiU+gSFS+bLZYXsEudZzQkgHe7Axb/24Bz97Nn41lVcx8Auurxh6S6fH5oJD9rpeCNf/IAKMA
F69AkR+TwedubqZfVHtx0cj0T1x52j6+5eKeScvCSCB5Dg83UaQrGoWJ+MqCbHCpTWdaJYNjH9Tr
Bh0M3LPRX7EsVPzwRy/fUWXsY8ucdlK2twq6Dg3AYYraI8si4UTqCvzhRTrem7zh8yQOxZKouacs
1iDEKLO6FD3+fkhAVUClTD4LbvhQv5fmBOnUKFmCsjnxzEJbPbj5ctQ/yt8uvGHy8C7htUY5CcMX
jjgwWCuVYn1r/InH/X7f4TW9LHpRIBwEwCXn7e22lF9Axw2mjD/pAY+CsvlPsh2l0jRvUwXYenXE
KEuE1j3q4rKUz+y8HQpNgVuUVFldmTqoR5IDhm27ZfwZyKnRlowEMrY4hlKvTC2RLzCsZZk8evdj
IgbdT27NAzgnm7HibF5KdGdCaBImlnskqh98ymyAySqeuKvAetVnmSVLA2iMYYGB4agiE0/0A9/M
5vOztHhymQINF4j62b4rBCJ56rDsrhOH4XjEgHoOn/Pygb/x13pttoAUTidkIV8DZAmJ2c1923iX
2PCYanbVOqJ91EKw7S+NoW2rgJg4282S+puIx7qvcNIRL5cgLnj1MMriQrF+yWCTveEp3NsUqlb+
19ekHZYdt1Bh6SrdnxH0PHaOM0oF/GXm9TfLfoDeAD8bkVqWg9Pz4FQlAE8NMyhTiJcE5HA3mPeq
yn/QVbUB2+NkuMOad8ziZTcLN3B14xD24ZKMNIJJG1ROw61TD1dDlx/677q6ltiqFFoW81JyZIei
8Hb7qAHGSR4W7DPaLItq7xeId/B9G0JAcyYBaIfaiCBDdJhTRnCAPOdpuVTuXa+nErsuQRhJ/Y5d
FYaUJD/M19ZUKecgTLxuD6kqaqF8ODTlXE+gatAqeFem2sq2mpAR6DqezkAmdjFGPpzFcJqzxggl
pcu3659vpXK2WlV4987ySPXJgQsttXEoFFypJqYd00Y3PYBFYzYDa1uOJ3JIMkotz6bXD/OZe6ux
SdGQvUXNt/odHeZMYnLoNHbBc+EVTFJKWATGVXLzAj16AYy1YV1EJUxt6Ah6Itrd4bgfCLf1unV1
EtB6bRg7sZ3fm5j5YqIC79gms8VHvum0oMjBRuMb55H08M59Bh8O9qSuFvdRHRuQyxsDUi1ZpksH
Je45m4zcsQP1W+y1/BizIoTpzFdWa8psT7zu4RCkLcGlIyQxRKtDccH4B8+2/cUmy5ZoJSBNY3O2
D+Zd9e+CuokgI3oFJY+vqv91fqz6YYhiKthM0tE3TQNqNTvw5QYgjiouIISvQFnQjn2r7m3KFK4U
OnWuoknygEDl20uNg2dPQrIxVsNB09xXcUzW/crEQXxWwT3KcP3jjDlmOK0vE/P0ihOQSYFi5XsT
zZuyXyhb7Xp/GCDdreqzALtmx8qZY5Rsb/pvAEfgynwEczT3LOawq40uQzYuc1nXC+ZH1VaYtGBI
5+DtnqMQarVzJKIsFKVLiXN6NKCU9Zwb6wmh2OuyeDJxEeZhVOSNeH2c4lbp+Qb//QmF+WHvVwVI
y6UMbIPTwRdrW3t/xQmUSX1d5Eydf27VFuuKt5Bmhq4ZOT75QpAWmZl73LqqZrSEUBhSmSULPOF0
qsngwZ6hogtPPGP2IQY+nftlKSdPF0rLj2mqa0Kd1XaTLQoOLhH+304RyZG69BKazxHlJiaVRRvt
dN7+ZccIpcCI6RafzL4rlbPQP4Zra9VF1oYUsqjm0/syDHefV8KC5zuc4UOxIYzLYW1n2UGRKow+
mPSOyEQ0LXzcS891qiWMx0NIvgH39KSoyIJaMmQPCTs0OvzaeTv4zfcr+TJ1cRpdM8etX27KD5sC
andSEWeoFPpJFiu2HqqcpGjyvDW+f17Va58ouX5dYuqH4Hh2EOqgdCHDw2zfKTTzDQhZVqwtlMRr
wz3RNkGeK3CfeRU68+ipgAuETQE8dfr6DUVcyoh2D8MGmq1ksPVhV3PN5tK2RPZfmvuZOM5Hu/ub
RelMeDZBieYxC39hvBseCRBXdEzKbYnomzuN/JuuEO/IuODndszVtZoo2+p4WgaWqFqJj/RcaISm
GoQHg4kV3+thYFMMdgDUXfZkAOUWtJ4uFiyDhFF411Jmnew/oHVWs340SWN58d/0i8LA6ChMjh6F
Ft9GmR+eJX4lgHCSA2yVoxH5A3H3vFVBqCgEr6oXiW5zAymABRSdSrJ4V1TveXnrN3ptX0TCDQR7
zqKIoNyUUA2fSOPHpehucAnCV3LMMW+1pyNyHDBxCWn1NVIanNcMqRQ8OE4ARJrlfeKwdJf9m0lK
P3eIep1ZRT8tFZEkLYI22c9C7H8YFWhiCAtUpweGQoBrrfjtYs0fzCik11KDgCTVsVu+TxeRk0gg
RaxotdfI/0hNEktb4/hjGKFldWSOAiksiBiVOE0DFjkRv1LbCA5w1dVdiUwy8yBtSz/itMl20bxb
jLaviPXyFYIVJvD7mLPf1L2T5yYkjNAJg/5Nn432RNy44rGjcK6HgTNeGg8OmAImzEflmDdUECyV
8fI0L9gK4CQnqvQ75AKqJW5pQBQQpHlGnoSxcf2v/JF7K7frYYCc9KHFSGNuZ9PeqUlakIHelc2U
r2tPost+2mAM76geFWUav80R4sc0g3xZXfnB3je11G0FOjftfMIZfbmNTEJ0janFjWOOcAcHLva2
MNHcrG4SYvvUIbD6+scLXgyxOblaoLJrtR0vAAZJVbcz/zU7/ISnk0Cs1/HEx/rDecYP7pUf8uio
rHwQ0hoTNA/9GUC2rw4TGpaiy+UrNIFuzNRcGKayfnvzuJiT9hUH92jprpDjg3NOkGOBaIxyTyCV
jDQROM+JvJdC3QLpEGGpll1nJf7joCoRV++jILu31OQRqBwj8qAwsLGe/6hoea7Dtcb9TGrLjhGe
t+GljdF2G4VOfioQNv5gkdNUBTxzs0Pzni1dYVG4qtZ91nQlPGiDK8JGfwQD4I4s1svF3Z9moCpe
tWMlkNIFLq59br5myDuZrj72qjd1N6/dydsTwh9b/F/rUkoaRLZAH3D0UHEH1CYZnP18j9UNIv2F
U2utPdemX9ha9P6XZDIaFsSLzTcgg+G1NIp8qOjmdrhX+QFRZBjRJxKuiNFbbeWvHR5PWHxvUjaC
6QP0mh6RxACcbRhYDDEQ4LHuSsoj479NC2TBuwokSRvkx1+NSgewgrkorfFjqJbFgsI8xOnM8UgY
PKyKBt7Je8IgcH6SA9CbqU49e9CmUHaaX4MvMQLj7UAPyg/ot/7fuL5r5DXJ/MxllPYPMRxPf12H
MJhyvuwUJYxLhkcKWM74pBFOIB9mnO4cozvowdrY85uxx3rqvFbehZh5n2F9eDral9rd3ykM6t+R
SJAe6gpjsGfx/KfnkLJwhLnN+t/1XWFGtXXyYB24+WtvqyuCUNZZYh1d/pcKQj2LPElvDTCW2fbq
ZR1nHZFnBq7rWprVOl32pKQQRBpkQGAb7HjMXNqSldgNEMrOeUgR9vyDh2M6d0PhJYV5Gttj/GZb
cnejm4OhOXlSJJDSyGL40WCppAOWlETA00UQn4cIUHGrQQcSseB/o3dEFZjxVq2h6BH/+kF3K1Cc
s2GO5hGqhjCjNQVpNrZfz28I//mFSdNT7nrCh237N5KBbs34L3i2LTPKWDRcQW2/iyn2rv2xlh0+
LPeqtpW8VNXAowZlIkL/lHxnqIoVy3f96NJyRSvGlHkKkVB0oKfKTevNJd3WhvCSCAyGRmwuxqM7
KQ/t1PDbdGHwcv/V4JK8gyrXnkIFIhLB3FJcuhdtrEAOCtKb7H0P5NIwaN+xmZq9Jrb06vb1fAf7
deC/V29adjEbPao/W0BJcouwEwcAB7o9shEBOfS1Di6Pjmb6l2htF6StH4rxTeyPJK56DIOMFEM5
OwgjTns8ymv5KCYe9lG1gYSHaxqEdmowgEl72RdmqQcyn67jV0jDMS09IgfZOwuejRAzap4CdgSb
unkpARxjTN39+B2pTO1OspaKrtvGt5CFPa3ez70RVwSHL8guA1oY8tRtgqDaA4x8vaNw1Pdb9aOx
c6nkM7iHMP/yA7LAeecYV7e8fskzqNGTZl5GY/6CPFRb8a8TGn+lZmICD5MySxPgh1o/iZgwv1jD
XWfeqEDIySiZ7neeE3PiA+HlceruZ0RuxAN1RyaS6DXCGR+jQtrgwb2auHuAk7T7tp+DBk+CX5KJ
WtsUIoAn2gpti2ED0vSw5MajacmV/Gj+l+q7h8r/mN0C5HKVo2xpK1u7GRVE57XnG7yYuo4WKgTU
J4pxZvkdKw5msheFF/97nZaPt6UuizBi41B1jAtaX+oz3B9YmYxj0YES4BFGSJFm+qUTaoiuuic+
Rw9/MC3QB+UUUIOwTa2X88fWkUZPlJ9A2+YQ8+hdg5Jc79Bp4uTCOsckbE9EyVFi+LRN573AQrA5
Sz1YrUI+yiXI1eEbFFjeTeG4Chk6mF/7rzlq8fcz7LK5ooBgj5FH2Y74hDBskno2tYWPnBC7lyww
4MWJT60CW0kQfbfXSltm6YL9RK5gMRXWvZ0DtVXDe6AP53tiZ3MoVQEEQ/lOERtlEj/6A17MQA8Q
dbtNUO7tU15HksX+ITQMdeaF71fMT+hGi/0kANNOO6NUZQvTD2oGscuVMpL4KULozXSiB1MUYntv
AuIlX5FjPjhpGa/V1Lr8MEUQQsLMEjd8UfMoA3IGa0myvyqVU89YhOJNPWT1Z3rve5Etw09cixnj
obl7eGafg+asb2U+1NpRFiIDTgGTwMlhMI/MNQNfif6t9uOGQ1jUa27rzk4D3+WYk6DTaUAKs4+/
Di5hNrNqDa26rtybZnX60biIx0t85R8UezTYHeTVsxAAfOj5wX6PJJtCJp8s0L42fWhvVmXLTPVE
E3T9fo9W9ZTrxjmdUrs9UCKvOfuvGPqctqhmZy0BlUsIgPa6A5Bu6eGApc8+vGI+aVGxgzTwZMcy
W7UAWYR3mtNwuLl7VVoKoe+SH9pMzRMyjy2JhG6M2Ht+GZu6kYweMKcuPflK+ltLBXZa1widnfAt
GXg+cfoEQZprtlmBjkCQg7hiL76LQIX/V8tQPkmEL5qCemOVDrRPazroePVNvi7b7o70wC5UxABf
MeXf2jPmGmJbmqBCiPm8oNsUoMh9wjI0wQO5hBMo+4N5fyGHPRy9RdOlwBQ+rtqnJtwd5AD1boiq
BqMEu5aZ31ED4vuLEzmL3lwFEQwz9BkURPCYGu0Ob6927FCQVPQ+QjzQsbhsXBULB0BkXgoOyoWI
RNwkV8JXa1XMDofR/YlkXMLys0uxx1UVupH73OC0x4CUoc0ryq2xzkYQ9fjeDvqevYH2Xiz3YsqV
ALCzR33BQ//kvBcquWBYZRBRuwCs0zy00eVNw7ycXArZz5k/ivip+ge21YBBk7X0yyASUmo0FdZO
9FSUU6jwMAji1yNnQGhUOmF52e/qUCYrAD5WACXfufSeRJgfRdorBNTXyoKuJzWN4z1l6GMF1lvK
yyExagfQOj37DGIlHv+3NQoOTvr9/VWp9aKqn9jIQXoDoq2B3o1L29HlXFTvnC0EYvTXQ7UBeJwY
wr5THBk0F2YY0XDMh3K/+GDZ/TTkLgSrj3oXymJreXCVfWG4rRS5jS9Fhsp4MFtwnXlC1/Ntfevf
8s1QhBZeHNP4eGnQK+HEHM8oCE+UFQK8/oQWDhNLop5mgUCnVg/8L919/XLG0gBGrdIai0hQAc3d
h0ICs8pWkdTIOK8NvCO2+neGH9b73YZjLvJWLNS9zO+bvCru8f7WSx8LWfyQIwk+1oESytmD+kK1
1OxgkYkVyAjrFJgb/xnqdlLscW17Ln+OhvCjiXSDz8MUL3uyAf6Tp8nXckdNY7jZVt2AuJjXnDu0
1erKRs85gpeNrR9GJKlbE57+du045NCNYtQimdZZR7b2XYHk6CQKizzUvTZ6djuslJ34301wkw0a
fgOLM5fB1GESQsbVsZJtyTm2sgAMJMDIAiqG7rZcw+sbnkA+LCInpjPaEhTxNxi8P+z4emY0K2OK
mV5QtGtNTnYUeevCFE14VWC5O4u/2K2OppbDfhvWoAkERuPL5NUu/lrDkn4BwyDSXV0mxBWBVdgl
7MQfWMjQn62bkG8gbuOSQnfO7PeSquHs6BPwvDztTLCbVUQR0cAPCLM8eqyxJ+78v7VB47zlJyzz
g78BHvQ33W49RDtZ3x/SnZ5BAA4fjpcdWYeYyNLqSnUz01Qq8UvSkqKIDhH+kEqJ8hiuyFPu9//m
cxr3YLz/mdLtx7uKrFEuN/kNycFWuXzgJ7EaYfOm0LgczT/v2wSs2cWiXWIwR+sSYke1RF0RUlPP
K8abYggSBNJgqrJtTnWAdeTnLeth2LhdrCTW9IPLTX297aoRg542z5j+YkZ5UE/FE+mJIvan7fev
SLHPkCfjZRqTvXPjAqcH34c6VsY9qS8xmElezNf7u/n8qewkVq9xrvdRfO6tNdOUx+vtdeQlQULw
48Wc3TL8g29zpX9J0NcuSvnJfthqLZoqAeaB9xBbOLDQZCI5g2eTgXRYfhchgdmxkWorAcHYAUsA
O7t0pe0spZtOqSloXBAwnS2rkg3oOxA0PgXRnUHAabv7fC30zeDC+LgUzX+CsanhKyYKO02/gJjN
85xTl0abSaLx+WOXWiUmInWrgta7D4B10GnIXXqEH1jINc6+hwn5Y83s6vDffcuK/0ZA7wy3WEl2
ByQVuXfkhHVw7sNyURiA4pCKh+x7hGkRpB5ONmxohd1BiDz1iLQYPqaF0HhHPAnUpYAnqLsXfBP0
ff8lAgLK1Mn7j5APP/VH0eN0OkMOK7jx3M9DXRjyD9CT3guhtrryCQc1oGa5IHNVtDCfe95zpLAo
ScX2HRKBwvzvl8QxQWupAMZJByYDNO7IQAhFBv4f5JB//zadHPuwZKPDx8W2pm96ne/fTmIm2KnA
OC/TRf46UQEFMAHjjy/qMPywdRsN87jmbpi6ILpkpYg9JHoRH7K7OlqYIzhV6Hh+fr5rW7ljXyD3
jX5cZiETfmVZX74dRAWfnUNl80OQAPaG3c4jSqt+n/Y1E60hc97ryNr/jIbAYmxJISzKRkhRQCCs
WQSD9RDwMrqr7FZcqs+tJ5qUjTfT6gBe8unnPbDq5poROSbTchHfW3NtilDkrEqjU0BPPiqipHK6
zLUSuIcwA5s3D4HcNizQblNH7g4Gmp61J2Uh3Q2a5re+yiNrQ9vujFaTayD1i+sCW0OI6MFXK7DM
jCEKa2felkWg2ZCTpgX4Fc4vnkTh+PdBDyiHnQmQR9ZFEn48QaBYP9o0UysKf6XN9RZ4C/yMW7Do
1LmD3YnMEISyXvHCs0qjHljGutrcuJMp+uX4uFM/LRTaM97zxz882q893ophQD75VSqQWyyl/SQs
DP4bmBdYzYIWEUaqs9iKlkg9ymO/++JmIJLmlqswMNAdXKmsRe1WgwlcsgahodUYLkRD1LY0TS3c
lPAAn4JOkX/l8u9515Qdp+rThFuMjTPPg4z1G67Zh47K3b7tgI2Aht9DFNcWqsPOUb5oAuK8pekK
IacMLMX/3HqnOdLQ15oEdBYqu0r/JMITsPDUzgfUJnCnoaT/g9h9kkUgng4c8XrYl/3UJ/PO3eok
CnRyQ4RfaWEyNgK5flxQxsQ05Sc1LmJaNfaxtHnWjyXAsDUX7a1OokVVCAWDuUs8+U8lrSN26XaP
k9aKtLs2j5n/qeiEciSWgw56OAYFt4d47dock82a2/0wNBquwf1oE5l5mvt3e4JjWLRcNq3CxBPF
4xRRpH5WRvD8VGBJYIul6f0LrXaueKAEl/n3I8CoKTNTG6IuZIowSOnINkzmwiFAX0BPM31qH5Xm
7IYHgtS5EPmXYP7AZM4ccXfAQv+ww4gm9FHFtSjT/RpYi2x5BuA0NGewH4BfVQVpkdoUo9VfoAVm
wSvetYkVAMM+XRvr2eMjFYOlV6J0rpd4zq+FUGa/jMnvL32Jzj37dzOzoPYaPHrk/5YXZ2ulSBdj
2xqCsN0b56SRn8mHub3A0bEDe0iVCK+Lf6ac7vEc6rr7ceCJpbn15JHQ2tprsWYFnzhvHzcaFQ1/
CFIYCgF966Xudt0L/QY0c0WoakUAVx0rVE1MdbXWUXx4Ab9G4Z2RPNo4OH4OWyde6LmHbcB0NcF/
/H9uU5o2DI5adUdHExcXu30Vk1pKqF2fSy6ToyU1lwwzFlTOkPFMTU71gGwwZm4YShh3tsQufo1t
Q6L9Nui5Es9aTOFTwbeIVM7q29OIqeWOOlGpCEHuqDUubeMd29I3hMHh4YhZOWNQEBna64Qmz2sO
mfp/lzteGZqLEl/WsQmGSKQ8JFJvxXhsqkODlsFfmA53hbQjAJUF3NdIp8g8eCgkqEJI2jSUZqxV
PyJPMkf3c/d2XnvAthwX2IIC/PSYe53nSqpWBHPUmQi2W3gHOhTMU1y+PmrgQxJDz7CMIMnRggmd
UdIWk7tzpujgLPY16lBO+yZEKM7To9fNhpVDMK9xEWkdKS/JazO3hkwPzkGWXr2sUHi3FWVVGyIv
0KDKS++ByMtRyn+KEzcasiirxgsFsUVK78PrKYQVdWMU19J6li8xPg6xLV0oIOZnU/SbOKfr+6+G
sy/WXdcM4wAWK2EO2ibxCF9QCW+/R0o5BemHijYEg4v+i7podzTAwjF3Oko/5rSn4f8+Jl1lbMwo
WTB5kldvZw1OieYKKoRxVhdA4geQH3SCW+vsIFl6V6FNHUfGPG3DZScYlUB5vw+38NqrYExGjBeP
0j1hp8Y59qSJaRcLkC4n4nI54uVHwKIpqLZQ5Av8va1ycwH79UDhay5y3Ao56BRQ4D6u31wfzEzv
Wc0k1YJoqP3WCM5Sl7Qa4l0W7SnWvi7Q74dNd8YnMPJc5FnMumc1yqIcsE0/sXN9V+/t/FVshaeV
JIwcfh4p2QLaMMiFFq/RzhWhM+k32CfYN3wuI85li4Bj7ooakVYbfICDf6iJDcAUjD10A7/Sfhz9
cF0g7egC4zvHuW8k8GhMaL2mVNfKFgKmItVgs6xGXlNbaEVgm/3hk+nLl93AD+uwDa5uIY6X25No
OlRhf4a1JRHroROMfBb/Zmvbcwgba4vWKL+00CXIhjOvsitDmeTJe73A9F2+7tFy2IIe9Idfjnz4
QOBh7Vmj6LEdH5vmO9q1awtuypxVrcpK5819CqNiam2AOPsKWnp7UN9X8xWd8lVNRNJaEmBP4vTt
8JQdjd9g/xSONpps6FMBDK1xkTms0fBbXgoI27+JmFF6GBtg0gh7YTUH3/DE4qZE9W36XNvKwJFh
XCTGetooiAcPoDblPHD4g5JzY777UupPZhAyCI+ltcDx3/e5Sf+Om/En9S/iftYmkUS/N+vPn0nZ
a4QminFQp/1rgvPsshguvtinGOvqunWyfOLYlrnlJERv2cEBJSCaXdvVSs7YoTzku2tfqFKddK+V
Wqx5c9t5wB07WGoHZ5W0mXP7NFJzajyJGrNiVCRfA1OFxtmmFyQpY4EuOH7msqJEgS+ZgXbERWjk
JJD/43lNn7+uSTe05QRHFAjjzLpGUwGZzaA7y7/kqZsZl0e9c8/CTa9tPS7TdokAF9nu+qZRdxix
xOkvw3CVPTruFtkpFj2Xjr5Kz3j8ov7HrobcXJRsx1A0uBYYnoW4QLT5tCFq4qqjTqrkbaolKbD8
2r+DQrf4fYcCXMTEGT65DU77V0Dgf37r52ZdOslcbK9+OESLt2uLMJ83yOO9OVI95j6btbrhXHlh
YKbZajV6iGiVQXAERhk+QQw0hn6uIE3xaydd6ORP57sobx+Lrhp5PM7e156pCZ/Sti1ED7wuCuly
pTJHR1sD4BzTa9HoFwyWIHTqxxQF5NEauf0MTyIQKkTAQzLdKBYHhHt8Cumos+PaUxZxJUHlQKcC
e1TZHXo8bmp0OstKH3/24cGGk5jOzMKuAzE1IiReBizoWfSxtMkqLMXnu0oaDGnqRdmB/tPtlFF4
0dACGxT8nyDKjiwnWZIsCSnLPC42mmspDOPZUK7nMKOiknIbblzxopvZ3TV3KiyKl/KT8+5uvkxa
Efa5s9+uxhI6XS+Qw2P8qXwzkrDtbJe2xKx4twb1YeFZ4b7riaGIL9XcFXTyi8C2hYh9jb6i7zSZ
3hb8moV9q1b78Kqqbay6Yf5yAfM+PAqF5WIF/0vos1H0W9OAdFy+1GCYYUvTxMrfdJa1UScM2Jcz
S6ykiHVX9ClxbhaZ0vvCFne+m5yVwF1tnRdL1OjRPiV6IK1iDfDMZOtQH4aHeF1bl7y05594jWUP
3c0uo0ttlRFV1tHviab6WnlHdLxbPEjI/Y27BRozDDJyp28fE6X0fk49R6ACk0Y005IzrSSCy81K
RbiV0rJkNUXi3KAQDVdnIfvaJ5s1jN3jHIzv/Ay9aZHDy7Yrd5eeUHndJDq710vWr4nB00Dg+w+A
WaoJq6aJd512PFcPuXcH2PUfw0E08Kut/yLOvvFI26//2ifWEctHFmOsdhHLiyaaMMPIAg6DXxqg
2U0UFzSkVJgKa04RHcGeUU+FL/Y4116l9c5oK4G1jxZY22drB/AyKKa76z8zCtIb08KyfRLkTf0O
vzmQx8IuR+Sil+3wD/j4vu+CEHURb6ixj9HblvkM+JXnO2nsbSg/oNswthwseQjNnwaShkzu+TtQ
CwVUuw0nYLkOpFzUmDP9eJ//IBHzVDiYnpXYCtjsEFW5j0uQVCAmUJOWK5SKrDIcE2vue1V/aQDU
CW/ok2u5fuOpsHfovTqeVeDzrlTHaQO75coGitPTk00xxel4WKWHhkX3eCrGPbS8t3XPjE/Zl7VL
fohsoOWK+cs5jiGaYN97EOIJZg6NB/SpfFp9cKNlbe4NXaa6ow8V/6OgqCY5F+59AfzFNzijvVw3
j87D5b78UxLVhS8Jt7onfZppS1mI46QG+vWjjIXQh5qbVqe7hkWDXkxewG0gT6XoNEyyjDaA20a0
lALyQY9oo78yohnq0InhTTH/U7p2DJk6w+SKy190HNkggq4MujNGUaF6sYDZ0hgM6i0F0vfKjvMR
giihEbFACbDCTV7QSYC66D2LM/TAH3OzD2YgXrJS/QWR/sGDXGZtpV8X/3jsn0ws1rRpUhzA3XJQ
WFO5TuIE66jEGjFr4yVbtaUeLG6Iifq7VmPsLEnAir4Gqps1L0yXFeEY1k2csbgm3y88xpCzTFkh
Dfj2s603GsebyRXiXZJVGg3bk7P4zvlbCt5ReeNfq4TCdfho3cjL8BkcWE8WQco6Pi6xtuXxy8IZ
ZWAKK1NSPYpy3jBYXj2EMSA5h8SXbe1SRiq1fXqkXpBbf+CN2QLNY52utPcRCSgZUomvr1iMHxgA
6qNoVdTfISipDLsuDm9+KYqe4Qr/zwiSsOfRzn8gZ4v0kWEr6pQVw3xPZFkpAZyIRchRUkFvrnfG
w/n4ePyObSUnWMfwlUemOEMBy05osDWb77PB2Hn7QveOX81riqiYUeUGeCv1VtzdWUn7ljrRzY0C
3bshlD72iIDm7kP4YAJ8McTak3KT4uejzc9ZE2I/tfX9M8BnEwyv8liXvOnjfe2+srRnuEKQsv+n
4GbNVaJgPFahMBdjSq/tJ5jtr6dwNe9soF6UOz+OoS65+Cbrv2COJLbXv8O+zpHGYGS7XO03IWuG
kb9+WCr71Ers6pDZ6i/oOmeWsCiS8cnVfg0+rHT5H//EScyHXpS0WdklGgqn51rtviRoe4oFeX3v
Y2VValiZNscXTQxRRoZo5jvtzdDEnErBD+rt76gGRoBGWqduxTKSj95T6TARQ4TC8lTPk06XSiwg
KnDstldmJbiZeWbXPhB2y/MtFYcjsVlQIKQzdUuxEZ/o6vSLFO/2Wo7d+UmmF2scdu1ENFK4C3zb
72GDDqI+FEmProegNNknBZ7xSnlW8TnLZ3w0YswYJGLSpvF9W1w89wKUdbwY3Yj5w/5MvvImvcPQ
NSKVR4sFfOb1Lg6mz5B3q34TYE2Z8odft8RYLh1apV0E0/bgelAPj4dJXwt6u7b3RnePSvQJr26f
cvR2c99k0vfGf6dyoiw2O7nScv+LnnfHfsgitvHIGf0GhfPUcgLwX9yCpCFxavHT7YokrgEeRXC9
2CXcBjyXWHdDpFDduoEqBpQ3LZ7Nz0ABvVf0RyyYXBrYyBKbOpFn0qC8MqVMXp/etVbSeGJ66mOg
QQCI/NDpSmzCkE1fIllpwkWzHqTgtCdtny7rrk/DsFSKwORZfbq+wkax0PRd00C2NnUpnYYCryC1
klzjw+VQSR//BARq8djg4nZaHjPuvlGDyVX2paEQ9puBUCVhcezd44duUmE1F2k9b49VuSQfK/Aa
g/3xIDpY649gquScC/ojUeczApmawEwdrnkyrEUsxtvPWD5POvM2Ah1Q9CziSrf3is5vu8UV6k4Z
/LC2k6P6eDBZw5Whk7TA6Jl4eEZ2cUTOvu1bX654F1JdN+gIC3CRvpw8N9qCiQiaLjfChBxL3CFi
rI/ZisSy/nUrnIzb/51x19RmIylCSjqxPZwfiYVhdbEyPTrnWHLpx0Q90ig6izyprNd9UaCq2YsU
QRna4x4srCUfGBBahEd00uZQNdKJSYDVLalfkh7lgo8rkkpvi2bCF+QL8XE3ZBZQ5DwIyOiC/hJH
cmYBMg2OxetOUBsnurfIp9P7jHtFeQMhXoy+49yYYuXiDJvjfRAK7RkowljzU6TBdWYqaGzRdgvI
FztqP1x01xIuA186epmcvdHiZfoHlLvLMGJH7rWtsDjdBu6+PR7DcPEtcVaA0g1CyPF/dlVmg1Q4
aJWztKdoijnJ9ad5Bc9P6EbaTBrfUCffV8NcowGgedRMNzvB8ycuVjRYiJRzfHQ8KP7omIWmGBBA
bNEHP16LRD+scbluWOH/hF+XrvBfWXubMIA9UYJ7uSbgE+/4U4qXKe2P6MWj/Fb8ah/nrw+9E5rI
SlfJPAmlfL04DOQVw7N6obIIhFelDcP7pOL2VCn3GSghxYeAW1jJ6LcyYjwi/fiDBcl4GJ4lohOw
/2BNwjv8h8vGqcGpSGkfkvXEgRRH4rHrq5wlp2fPkxFqux2DRbF7zaDakZl9Olb6iRpJsBQHHfme
de4WoJvH4FkWO622onI1QiCPUOzL5QZyi1PGNDKcQJpW2YtXex15Cde3+Lr1Ump1UzNWFPc0hoFH
cP0dlRkul548K2weVMIz4WW5LXSy8YoJALIvU9gdonGbNy9RH+xJypWMd/0KkXxkiEZRs2AaU+AB
px7RWF9ex4ddKkoYtLmF/hyFdRMV8WBg6ZMQu+8PP56QiMEkErutZq9cNoGm9nfTpFDl7/aVqGFW
yihax+Ya4zV65QUGkp5CxMBNQ93rzVGxVITfpmWGTm+6+bNmWC2lkaAx3FykPEapscExfCGqU7GB
atDe0HQIohmGErAMAZ41vhh2OqxW1OuI7Q0G51517eOYl58aB2mVP1y+w3xMgBRRUxYJQRp5B+2v
VbL8Te4XBwTHHvw6IV9UJY2yeCGEJb90HF/dNC/F525DdXOB4S5VgbS9yLElUy2R22N4anzdKPOk
cKzQBgGqIDn30H0EZy/q8Fi+wfvzg2mTWqf4TZy1BJVb9eYmUWdgAmb9aSdbha51dk1xPkYB20VR
Q21SfnK8uIJAcNGt0A9EhjyCIkRVboLNthYhbJ8KF8Fb2BnIg1LTHvlq75KzOBy7wIt73f8IRwhz
so0J5EEA40G+jCcFPTQyUteYhVZ5jPFuEl8nZFEv9QormX7WHJzSOV45M6nb/s/aJkUdcdiKsmeC
rTsoDwNq5+6QbI1/LZphRe+wQI+WvyX0SO4pwxUaQw1vjaroHGoxtO3ucIe9JFMrR63PS2hklhOM
tRSGCVCtF88ec85QuXnlb/A24MlGY2Z82FskE8DWJ9tRGcIdD3H6DtzT0ahfCroMcYA1r5glgaEv
ZfZHcCMuFmv+yFK6y6Ewmd638bP6dlqEH3Vl8YF2+K5B2QgIRdkA4gHrF0nTHDxu000xCFRHBn8Q
NEMi2TKYJlZr2QnHjPR3e+AIvHm13ehrUAVpbSHGUJEYZQJZWG4dhOdzWA7ODvYO3ImGgI5nhIro
Y72pq0YcmvWZFDR7fIX4I/edvVuIK7NF5h9VncwEZoGSkLAi5SCkHoFVhVwVHyMG+rt+/rFHXJYT
GSHovQIiUiY5wHhjcMFSNaCU2hYKrsPkdVBrVRlG9JeeF3dL3NhUgNQz9/GEukQsxiru3rWRlI3y
x1D7sq3/5n3b8kh4FDym/FyFGER6Q3JTT2CZvwufM1X5R/VyOKwLmyiuljOfmQGL8L9agLS3a5le
VU6dAxHnRnv29mrYY+JLN+pPSIlrrUzKlKrQWePRCMP4DyihqjJAAD3J/G1CuXGTrz3tMe3AkDjE
Uh7RKArKnycJqBj9GZEDOM/I2jNcqy7m7Bo7IKXSWyKltZ8S/MrPPAW0Jo1ex7TwpAq1MGg1wVzV
Eg5hiKABMis3qKyDCwkAQgNUKWaDoQdlic9WKJXYxzNbDUOnrC0DXeeH+B+ScWfn2Tm8jEAf67iI
Ill36xElBlFHqub3vP1kuUzOB3giRPocbzDXDEN4cOghz3qZNuCwGhQ8e44fZiDpdnUiy0hoOcMe
JWImozGbyhKwXdgoh77hsAjOD355zGSq0gNR75d8ZZqA/vGWi2wKURazTRswN/bQIhnD8rCXNq7t
hxHVt22lXINzgziN5it7gYZnTZC5qmU45QSqS3jq2anof7BlckabsotnkRzBLUr5K9S60Z/UHGvi
4uplywLUcbvPiYLUTYemzsjyKrn2EfbM6hrkRutuYnLO3rvvsRYw8RyQUxNX7H1uGzeVxwaIrMXH
VJVu5BDV+G1p/UTMh1Ha5kQ13nWooYyk8ei687/Cu9inpFTQ7S3rX65ThpNkhdKBJ0dVLsGXYnWK
8Qm7wTlAWrENas7legTyDDXz3AlCtFVEOWwoVFqSdPv1dxBxsMYlcwmFu7tK8HiYwhztYWFg0cK3
lkHz9rerHYw3lY51LjrYlGoaZWc5qHeVdUsDHl8u4cz9alYKzobQrESBRuHCuLjHU23z79JTqpRr
I1CmVFOtWl0UkLQll4uP9b0TEIA6pr2VNnkttPKDmNfXpD3ICMIcv6kZSsIum2W0GAlS0bAEiyfd
vrUmkPTSr11Xo5KbvS/P/4f7GD6kmJz0cWLvLTqxyytsqT+fHXyHDFxuJ5Cdd0DhM4Ruid7bdkGP
LWDmozw85ftHSspOcNjed2VkyaJ+Bc8Q/0wthtnjaCHKCZCr8ybAWX0Npp7e2S5VAwJbw7zSUq0E
lEeVegfdP0Af6+g5/Qjx8LmtgD3VRKSLfB+kuCNdKBTuPbyYjarc2J6smHhOgjidms+Ir42b/jBM
pBXzDC0ccKBG9Vq2TvI/Q0r8xepjnds2xf9nkYxVgNIqHt+c7oAUyspoFDJ+4tWkFJHPVCuvwMWq
3BvKwMqYD45VT1eJ2KOh3mDpqOTm317XTWWansYccH6HYXyw+7eCsPpOeNodbxFsib4X+TA7WDPO
ZSGSPe+gGxQw2QtHGln0zTcIN9b6mQvVJbMScyE1kpA5Kj+S8kJVi7kfypK62p1VhkXaIpskJrQc
KKASGQ6ZSyWvDYKG2orFl0y1dajH0coBToT+OcwoN0VcMbKYPID1T/cUf9AYla5VWKKISs5dy4BU
zOoj3Wb83PYYjHIV5w7NmBHPZbiHuyUCCjCQ+4jQbf/M9V52GdUc/Zw1gck3AzZUJ/NaZb1J2FAU
u5MAXcbdt45iiLEHYDQVa8tUBzm4ayTX37TzmRuQOyP7PobMn7X6zbC1VxeFcwyku0JDmI6d+6Pd
HPK7Pp/NakpN10DBgPhGdhp5cCjKTVHP0x5m79YlZ84sDszm30K0LZ7xlRYpNid1nxjRvABk4NV1
8CG2A7ri/joLiiHWB+XPv7bFKpN2eDHkcMj/xnxwFhepYD+Dr+JbjLnlOMEtcRP4NEX1MT8tyyFh
roaztvs+Pi5xd5O6ZIcFylZ02GamyPLBdWygjQDqRYgAftuuZs+AX+J8dWbHBqRorb42JGKp0LIY
tQnb2nv0S8kE/ka/gMzijQBIdwwyMpogRS0BOTBjD3K819fDYsiK8cnbGQz0DBa/MFm5Vo3WMJ97
4oWa0LqoXSQ/E1YAeBq9pjyuIRW0m9tDZKihgS7gWSsB4tn6+/tGnmg1r79JeKXKcBkww+8+OxXb
BuiyCBBuYrbGDckA7tRbFkYt0jqDuhFBD1ntyGI0iGRytzf7D47d1Ttgmbwq3D2/1AmE1ayZj8Hg
XnHTxIhkL+P/Ae8c97RW9IMvIZceXMWFYBLx8rqV70F67qIuflushUYcBKzvWHPJLK2CUSmoOsI5
cTRbEuaRurzyrk7+BZ+yyyKudrpNerMfuwtCWvQ2VhY3zmrXZJRZiaDj1RbDj69HK2X8tIRmq4JN
0bFOJuGg6+l1Apurcj9syjqzjjTNyfnaNFGjeduWUaLsU6lqfctZw3ddrxsQacd/fEVvARPJ7OuS
k1/G7sAWgcRiEr4uaKGmbh3ZZZuSouXjoV68PHea55G5N9sHxkHlKOW6Z7GSqoSEk8EsumxMcMzg
/0wZxLee2PE9zstPH02IbXk0Fp5uHFsiA8Lu/1sWOjmsnrYeGG6FCiqWrP1rvgkCAqSHbI8PWLdd
AdcqxD9lWbEChgjTZB5is3RT1gojfPNojbjKFgKLUXB0KlFGk45ndcGw1msZTUkh/a5k6hPtJuT3
EOnaWQRrh8ZsBh2Dbv1JJR1XioiPoRaRDMo2ZnxLyvXkv55DxcBRdqMXSUAmT9pS2MrBqsY/3R6B
4+36umS3emMyyC40fmtecJctrVAWuid/0JWA/DgNLmjBT2u5h2t8Jvg94+RocJJRrCZv8IUbnfbw
MkPoU+WrleBawfVRo0Pp0KJYwCa1bDF1XRoh87nflEHdCODTGelVjb+70bx5JpML6FNnerDejoGN
WpYre0ezmNuIUR/eXh8BiJ3zuDStC/Lt9t6FUy1qxGK6uRdP2LD60f2GeyRZbrnO3zlKRkNFaeYU
bys2Xi+QwDnExRyiZYwtCDQAoVrmEgGNwg0GsQWaXxhveYFZFOeIVmvRXk9CAS4ApqRkzWbQgXqS
dhj6jSawrhnpPzSMLpdpBR4ztkOE99t5UyJNJFJclVwF7bY2gpohoWPiSe9IGdnBQc/gghAiOAax
piUA6bslcub35UYJCwnMS1VFFDMOyCllBMXiVZ9wPPUqmnfwq+3VSNeqQkRGGiZ2lGlG7tUm2ae6
yTJ936O6w6gzS90gkkEXhHistnMuBNENcvVqWE57iWg7AriNHZtgjPj1f8k6uv/0G332IjX3Gmd3
pnt3hN6q7Mv6MzWlwJC3xJZ20nt0KBr2neCwAPdjc0ln5lvHDSDUMdXRnkk9bcUEjtxh98y60Qnq
1pjXvpspszN5qYBsQUmPE45b+H8bGqMmj9OTmcGvHGp4hTzDskO7dgjMYvDc/YqRRZfd9IOgh1ZN
dRg0H2wIE4I38V97ML6hdAdKAaNSQxP6vQcqxosu3ZrpJ9S/OHl7ZAkM+Dn+tq+BGGiUIB7s9jdw
ozD0gQh09z+nd1+ryko0meD6HIxTOPqW6BgwcePAzp1/N7nAM1l2+BU6UFQFSlwU3MqGCZpiqvbX
j/V0rCNWiD9DAzOrBv5Bozc5J8mGSjFtBf9x5qIhy8+SPzbgSEnWxsE0r/ROKuBflXwqH4h/BAhN
HU166nugvXV0mPtQcrWMANosoIa7vyy7w33NgcdehBzx0aI7ScgRXEgSlc8s2KYFRO+njxv4LxBD
amK6yOkCljWfCAgIRrBt0HXoi0nQ2faskTQeUZN55qeN56UMM/OiZd0LUTXheFiAk0zGtpWLvtlM
QcYjiRuECIDiBvxTA/qrXaj/ISQbrR1X3Nh3DDqyUA1mYl0uvFyC6VmeZiT1sfXA/Vg58n0Bb6yH
O5XQe0fI7x/WzNzFnfUhfEG2P2B4y4ftmEk/z9XUTWmdeVWTcMAg1Eba9G+6JagxOhIM66YABF60
0awM8nMS8vOT/OmW2zl6znGW+244ZlWZl8LEPqm8PIKqvswylvUfhTqmAX6Uz8h5gXOg1eGmUpHl
Y1UyAefUc1zx5j3oRKRGk71CttJ2NgExJJ3ZEejLGozsnT3kMdbVnXk1N7xxMYW9/eoGPhvUt12E
lpJ4vYpiVZDdZ3LIYFKNGY/xAL2cMqC7LlggXagOyZVmtKL5tcx/z6SSE9WZan8E1t85E7s1z6k3
+QCGY30wQw4gr61uLSuFmvtdFLDMuJZKFu/NH+GNawAdoR4wfmQkWqn0EsCA7r8HocK/01U9Lzs2
dhgIA5DmZfJhJJLGt0GcGkvrJAfvcN31Wsbef19Fi1ZoJRgRqmTyVOHkupZcerlLR6Gg6br0GrP3
iQjCGiJFRrCiSXG18Juzk/FM0Ln7JSeoMI61y5JlDzTMwEY1mkKOz3is8gESIm6KZdXvr0oCYO4B
CwEWVbM0a1RHHMC71Szw6jRHLcT5xCNk1jBdJboK/jBzEV88tD9UI2FqZ8xSEZJFXxSPD573bZ6N
NWdwgwIt9viVg8SpidptweioOBYU7mlhYtzJcS5+FcaQcoknIpDPJuYYE0g+jdmufk6MN/zPPAAo
llxrLzpX73fVz3Q/6m1ib5Zogp/EoyZ86d2yOSQhMoa3Djm4jJWA/1nM9gRp4Ybv8sq3HwfnzpJu
tHAj0SIc1m6cvz6dkJR/VmZNhVGNTjJ87jo+58alhq8SRXv43d8TM5sNibU41Ed6MXTGJ7F1hI8h
eNwiFm6p+i7vBOv03gY2gi4hTrW1VkhgsLXgUkFrsFvv1LO9HRTBN/IxhKbCMtLs3RLubM6SU9ER
nFTeQScKz3bIaIEb4OlISsKjRF4epJ7KpcJx8DhtIqMdOdiLY3J3eOhmBUi/pfVf7ehzCZqqrjF0
6POescqAV9p0O/4ys30B2SxHy6RqatXOPguOg0A6/uCvupuiFFfDlwGCdNSRM3JUvlH0C2uU+cSt
MWfBb2VuS9TVI2u5cAm+KgZMyfPYYs1bC2MTgz9fwOIxLEJtEF2VI6ooIBeLYdZXLccYjQuSI1nG
ZWt9nOCuOGXQ3DRnwAirdJRGEPUhjw5BkI9jUPUMv+6NPED2mo2FoV2hzVgoTgXaf09+fJ0haQRy
AJQn6gN7FfvX8dhKWFz5p/N4MjrmS6Bz28LriLkJOvfUKxtLraByA4yIOtP4d5FYjPcuaJ5CNCKg
BwQE9M+qeFvpJemtiRl1nlOubz6JcgczHNHPmC5bxdXiEy2EipSGugIPmeB7NYTEYNcnA1pFyAuU
FI+sArfEoxKkuRf2XWjj9l9xBLQL+uSz0JDUE7vxEkYM+TKIinJU345RzRSurOqnG17lgOIsb5o9
DjXhCw9dYhf6az2RQouxA+uNfh5uMfSkWwV82MHF0JlEZDun6v2KW2muCwWtPl6/YlFd0XoQcXN5
Lr0xD5f6xFrtegtSMVwyWQHquU2Os7xEJvsg8uqnlaM77BhA9dmiHuJ6+n8Rdu60TDMw+hMHrE0X
awLb/kBcHrmBNyrtIzc2ak4v4QHjKOr1R6h77npd2WiuUaR+hyIeRtBMPd7KHgP165I40wY0SYT+
ntBYnESHO+7+97UuVYNNbjTF95Gc6KEW5Qr5kPyRfu3YniewAqmkPnx5wdw/qu8mvSuv3gSgPawx
hNiM0J2X48/tbXwo5c5kosNQc0Fe8ZFhbrITTOSY3aikn3BeV5PKXdE012ViwHgYTkkxX3ihqpTd
1hg8jUb42oLWDKI9WUolnCaPmqkqnVdYKeWzAzt1acKsWhYzml0vtJQsNtOvD5KiZ5e9dQugkUEK
zT0Y5+2LONL5EjHFkDz7b2R/DMJK5Ynt46ZIF6ymQPa25JL7VsQho51PTJhMMKMGBPOX8+iLxncE
8oHGX328E4toX/qAZF16ooSjJZJZ6ERmqwEnQZm8DbgTi+6yASqXKi9hL1v2TK8T0vxm9grr8Ylv
daWR5FUiURXOWZpc3vdDLcLd25R5iDZu9huw7riWsNMIdDhRPRiRzjRHeussFz3A8PJBF/7k8YDz
tXkKpjMwPDzST8Me9tYWM4V7D1SLUfVj5nzV00VVzdHU0EKV/xeHXPA5DmNArc4b4kbnYSdPrCVG
bKUEWQZQwTAGgfU+3397HoATjk4rGUwPtuynZCHYmg1bWT8kQXTAHucZRS6gR+oWqLFTy4GaIPGl
BBvQ2kSGiI9UBS7nQDiHnIWG0i+iLqSlQc2qBevhpOtDcmCZTEBOcb4eDeWxdf2opONxcYGBI/n7
swSiqhyULVOQHpRJvGP6oX5ehWtKqU/5izw2hp4Eefs0DL6CecSF7E3goNKHSK8ld3O7lJwGElw5
0F03M3xwXOfoAegKnDYv9qLW7sHf7alTpZZ6ohS8xxThynzMiCe45SNQn3zKh9pkGaN5jgfTinAT
g7xR4totTeE7V7mqqmi4Rw0bY7WZEkNrUZht9657Vst3TsyjJX1Qi5Db3kVXEuhx+zm4i6UHt8Tm
8fWXlRpb8pRutsnTdHwz2QnUecTWg/kuo8tgM6C//0zyAVukb8j6sDCk7qBAdJtKoQrK4lNi51AI
9q9n67IDW4NOnR09fVeIgOvPqNBTDUcDPBVL7y5MhEE4zWAyFvlQzRODmELEfierWL2pOZ48DRMQ
iZJaumBM5uNKRN1H119hn8dFafS6bV/SccXsn/Vv/ycmOKeL4MhzylXZl27XBEqnYE2Wu+nh4Ey5
RnZtTmNJPh0nP+yx4WSg6b94ZwX0BpPWJklAqDg2LSFQVOMurOM/2craB5jbLVKodLQEWL1+DJMI
QbVCUjFrgUns+tBnucjOSL+ZyPG9HFdMYv7CZIk6LHIP5bwv+P+IEM1PHmdTGiFw1DfBFfOBKCMj
fsM/mWyOKb8ZcqbGtIIAApbWo+JqY+CvdnZNgHKmRgFvLTMzVT0hPclFktDv15b0FAoMFdiWjBy4
EQLW4/dqkIdcHMtp75EQsbgBwkviFPh0cqNoJP8ow1x14zvvMhUiTz6ZDPeIbhkRJPGRSS2woRhM
0zTnzXQZcLdXCjRwiA9k6onn16aLDYdcMgtzYDRnkDrSoaFde2HOMTn+glXuXXAbfQ6m+kCNXJ9u
tjxcTtakK8H7qeVMJkIcUBpplZss0BGlCgNd5vgUM/dgNAg+ClYvsZD1X5FbK+Bcp1NT0YZLiwdb
3CdJcAM8saUQZxyMwoB7wNXoFLpsqpH4M6LELQB8AhFBcfyOir5jOV98YncpY0ttQYPmFwwxYF/i
fVuQbe3YoSlMlyUJ+4Kyz5Ysv+rbu9SxynmpLFTgUu6eeLfa7aAELIP1dzj6N6+R4c6rpiDsjHqg
Gqa6Zn461QYuRpd4UHm/3raq2E9zDIvykB6uPKwc7CdSah8DN4sikoms7aLAZXOI9As+BXWTnznU
rnXfiFrgL/SWILhC91WqrbB54Sb0WRprjc0q7/nSpm3iZ35IIuehJvf+7zeAg49aHsCI9QlIORYK
eDni4/FXsDYBq0yWW8o85DRagzTkLIUue9quAK4EBZF4JBIWLl74XjuxNF/qzM6MWrb9G2vuJPuQ
N0lXRwM07X8RfNyzb0QFkRdYcUXyH6pzNmuvcuSsj+l/obzsW71FFeXDnhGfIOOLYUfujStPHh7T
LCK4fajQ8gMM8udZNPae/8GCcimzupqVZjT+fVxOJcLq4MYk9fnZ6cBQ8kCzdWRbd0owJyfCW2Il
xeB6d+g30SPUeNo+8V4H7bKDSsbl1mITO0nb327Elzo7miRHbxXKicz+rdimxK1uswvUQzZd+mRE
VDtLhdeULDV8rsZ28KonwXauYaEgmu7tJJ+yGfazbX/NsMR6P8rvt7YdZaV1cg85YgYQADmpu6So
k7sA1GlSNWmKwlj24B8VnyjgvUkAVCkOo2ZhvQi11K++tUrl7WD4ybQ9erhCRtFB1FCbV6McCPWS
PDFmoN6ux9HPsbV6SK8cvFFm+YQJ76ERzrPM4TfpTkKXF08YvBZEKWlzo6mZAsf6EVbAsflxsiXz
sHZQ3/1HQkAqno8ZvLm1UR98dEcUT7Q4vpRp4FFRch/n4QFyLbHrBcWUDDuFcALj6vKxM03ZSHhm
cSpwuXU22NLlWpP5FamNwAerC6qCWy5mFzJPQ3VqbGMW4UBT04X6NZ/ebNSnrZaqGfYXl2XwoXPT
MNItyugZsA4Yzk1VqFiPZRuwfGDkvrWsTL8SAmBETl7XAdQ6wyZMc/fY+gm985YuxEw//8YXWrng
EJrW4a2+W03bKfwAnRSxe+gNh8LPihBR1JxgX6uI7FxQRW9T//a4dpF0QkvchJmWQ/flTZfHjJo8
BjHKfpve//I9nrrlgirBZGG5ULgh/egB1NnAl5ibtokv3R/37zp83FVIej/4V1MMCWzymC6IGM4B
C6qGdNstu3peat7Sy3DyY6eKbPOglX/cftwuGwD9VvOZqsT1FgwQOX9xQowBzhnuNbk3VYYBzanx
ugNEEJS1tSx0+CDe+rSGTLwbpPJ3jsFjeO+wYM9tJbRU1GGoMVw3X9WnlhN9C7IxxYPg9/6dtw5l
zlbAyNLSklRt76T9xM+8H7kbpiRjgw8rJwDO/kO25onnEytAiAykljKmvlZzaFbsV6WU4zJKmelU
Y+t8acEEJIc6kBQSMcMa+RdVtIYoMs8VwsRJD46IoPC20cWjIHGulpWbs47Mr1kveWjSNlEmQBbF
QEVAkxQCWw4YaJOt9at61vd5zE6T+vmcQ273AzgJWY4yehk9P/utzoDBmNrEU6Cvt9CzUxLnHQm4
dCgWvLeSmT821iftk4xVYFd3XRuH4naeBWpOUh9qKnCarEZ+v5xjcGWjm8n1QdF49zSEsBijT29i
5aoppLo0wkj7+BA5YFfjDHA0SoPDi46ccuphP9shezpdmvQSrOcsG373Iszu79GQ4PypkSmp5mZh
R0jOsrvMzDPdq3eYyDHHj69NM0SH7+A1cWWGmBPyk/lt5rMfM55GVgiVvt6qSoEvFP5CQeI7UTvv
kxGG6trWHvYIdfx8+8+0ofXnKEyukYC4El/gngZcI2oMC3NqSoSB8pJGGRLfA3LE5UOTzYN60Vda
4gRmSRPD4Tql/AiBzLMIg596Az+7zy87l8KaKi3T16hr0lAWTRHeOUkLiUIhfDi4fvjNAnENIyTi
n35b62t4fDI3Inp80mYfLTkYbLqMc8mqiKC7y9JHDO1Si2gVFw2D/iqQYKq57QH50ZU9SzPp+z92
26SxKXM8egjQ5O3UyvedQLR68YDEaPZ4I7sZ1/R8hyAzVCqIPo2mZaYDCVckxCvKFZBWBnl4gA7b
5V8DjQxm0sJUq7kmSFATpZ+G4WYzXn4NrYAS3aUruMIkP+Oygi/n1wwd3KD4rHwH/rYDG79x4nB+
dmbubwBMx5On9FrQzy5yMuflxeBWDsh6S1XazvdUyPjoImFe4vFlvSsVETaV6eLE7gB6IN59V9J6
u0seIzcyGKNZN/+HDRS4Ef4pHFf6K2RCIkgFwXHbY46mMB1rzkGZN3XebFDul4u41j0MYcQ/2J58
G+HyBHaywoum1Be9BXJ7f8Osg9DLxiB0cOBrZExssFcPZZvVDPnLZn9D40JbKSUgH1TEBbpCRX26
aF6vaEzfSQ6g8rWj2OwWR2SyIf/X1AwFt2Sge48kYhw85eZjYqm7cWSQ/DXPXLd3AmyFpw02igrb
0UeT8spTdoLycKe5a2+Bp6E30uhTGaPG0Tcm9iCgSbzYq4LtPz3Z7yss3IhmMctf4rLfAAsmbD9g
QIh3PXaBuRUFaYSAdROcqKoaNRTuwH/zrwat4V2/QMDy3Gj78qnxGbPVTHfuRrnzvFYB2uGG+Z8A
wYB2+F7ajn4ZnR8+RNuuktd/dDcDZVOWLP9LRkWzFGWrjU9ffChQiS7BWPFGxGZc5JmXG1djuRJO
60HywPR51odXTOn79LDns0GA/qtUZDzNk0v6eWSP2qBQ5LaoqN83F1bwBGlnB168nCto1L3dLEmL
MPRj/7rF6Cumx9c0uzzAZOaR9mCBLOzNWIWYiomZq7Uxjte3eBFI1OBc/nJi3/UGZG1VFhVyUy/q
wpfpSstUTCfX2mwQdAnRuoSIMbHv/+VBxyoBFaYVOxGqOVYRHLbA+Yf8aujy72QulF+8DLX4dR4c
pNZolMvlx3d1sZ/3mnBovLj9tqJCimztk8gq0Vphy3DjlJjM3HE/RsuUE2Tz1Dq6lWcRFrF/EBGb
qVBf1M1ZG74tejMrGPde4YT8dxl0NwNvBHJjZzAUOfK6tcQAPl6OvVZLbPiMJnDrX24TACOZXPLW
WLJedRTKD1ljsCXZ0dxEvbasu1TDo2VoPbPNiQvg85q+mwbDauLGpNnz0JMbnR8jE5vS2jUG5sVe
fOOMt8SqhvlMR1qhMdZkpvgyBxPBUtyM5lC1wcLL5Nc1wI+RroDLqg7X5gIDNfdn1aU+H0uuFBhY
i43JcoJ68XMd4PdwQ9CgSTgws+VyR15sxxfhwaLkfX80YCFcZs6VgyvVNpDVNumeY6LVAwaSi0hi
QG1TYATED8EVExPMq4upFzeniDaJOPr7yvVyZHGmNa5rOaNfj7993krQoac4oWiSskzt8Cxt97mM
Y9e0hQ7PjgRjftmEIskk9/XpTNSpaaTTqKXRtVfm7fspd4nciTktRvqVBoO/tGrJ5tdesxOMQSir
Otyk02akulysNn5YXqY6cAZgUOKbEkAKC5JHBoZymu9JJaitkIo9wpz7YdXaxT3yNKrmyNoMBWSz
oVs6xZxhGrkGSRxJ+SrQt0UfwN/NN7aWb7T4CCZgNjnWLUjVsCR4r+COS5hV3+u5LhZaaCSnFzIX
fFL0wSfBY6ARIDD7vN3xEN56Cnjj91JOYrx8lDHsR/t6IFYsBwPK6vJXVqB/BHXRz1fPZmFNdQO+
/pLcVA4BJ32w25DC/AULbdPMk1S28BhDXfbUtycZsSta3PfxAAPHJcGZ6CwdJCT96Lx3XwrKuFD4
VvMBkFyBVFwHWxkyJiEEFZjDIqrqsSIMBEcEu4k/oZjcpFVB71DfECSMZ0vWcaVkalJJ4xX4QoxU
PEy8jm+2FwIuJZ4dipDLQGYuLO2Aj8q9QhRw/nA26hHmJEglEkQXK4x+4ykvCXqwo+5U8zko2a7t
c2mq3ej9Lgc97oAZbNPfmw68l/Z5tg0eS3qqdbMTEL41ZqElxRN8I+PTFkQemwJAX/WRFWdjRFxR
mJkwjCAwqSN4+kbeWfW0WORZUff4ZCso+qrkhZ04ABbC6iVeuDK5RKiDR5rFmECNk4qfuCY0BEwq
tqFc9kSQmVV7wTxSJ0YFYjfi1FIskCeqMO5jTsvdn4An40dYhSYIaFzjIQ7NQpOuXLN62d2fGg76
4ikrrnWG4uy+CKIt7cfgFobXKalITk6dKyjjdpGbJEAOwo2BERLIJ0W4NO60AI0rxa0w5YzoyMef
d/d8XabSGKvH0D+6HjtJ7eRL0gGV3Qa8jBSVngF1xbyKdiBjiysdBrh6LttvaSWECAyMfR0mbpHq
bHOVJtMbteoUnW6PPUsD+IljqThkYBO/0D6kHRDlfCGWdZNdjpMidQZ6XGSDYzGBqK8PnKJzN8Z9
OWYHEW4KyT2kOZFznI9+IkXDL+cICk6soepYJFEapQdRnzIBaKqTYGos9twfqdiCdT0Z17TLY7Vf
fUxyXAAbDIDkzTfSbV7cZ6KlDh+EGbPw7Izr+iCNsCQrOagvFCEf2E81Bzbxt15S9od8sJELcqx+
wrEbXS7QCr7YZeurmAD9QOsIgsMo+gmFW8UqXb7NveUydveC773gjYipccgFH3UgIvc91iF/ciV9
77F/+OwSD7uVuqyb/nCyJsztsX7XQeHADPQU9v7RpoRsACCofuotPHFxGmNUySg2XkhRKsNLGxOF
GaWmP5/vUnQd18TuHhYYtOkIi2uFZRqnpwvOcb+AKuB+5Yynq1mNnv3hBXB0m3S5Hp/nEGftQj4V
JTKHAWAuBqZteV8BBLc+HfgV6tlhd/dLJPoIIgHGCcInsuwzEt/xzXg3XtBBc0SZPAyd6J9FKUju
0YH3QJ4EaDePzRCm3WJ9O2TuQxMwqNmhganEVn5GRqo/WXuIVYm4uoukONDkmqsY92TgEKn/YWU8
wlNx7cFFL7JnM1gKqVeL631xza0KnJkJVZVIH4O9KtkEJymZ0ppncj/R1OVowfohx18ZLekAsMjg
SytQfgK1ZlIosabsijQyw+GkavHi78aesWDK1Ok8ZJEve13luLt13PcUT2Zjvx5i0FVXUSqL8XEZ
0pkynfLtbKiHKqRQ5QN0v+fId16sWQQhxNNuoYFFVK1rAyk8f3HqUyL+P09FG8bk/M+jzzMYJhGj
Oip59mCQMdl+oTdU3+SlGmyVZ2rC/fnPfAFKRkDEpFJ9WoYZd6k4dgM/gUNldHTsxMQF0u0h4L3k
rZk8lEKUYmPJkIviqG4Q1RcvSuhfJXUX/opHs4cwaN18oUrpJDGlu2oQbV8OD8Cz94Mx8twq9+g7
BHf9OvECjDzDxWHhqudsiSPpS8X2HH+oUY7k/qIOTiwi8StE9ix4Luiu3ufK+e0iHGtmEy02pjVG
eU1by8jKCFAvVousQg/FiMJgicV8CM2YaS+EQsJiEF8RColgQedawcgfucvrIFnOE09Td1q9lkxC
WMym9UqYnX9ouQP9WbS+5cprKsjwRj4fYAmborxhsVLi7g+ItLyFiEzf6O5IGjXmDS8jPPqKT7qB
PC6qxREEWTxVqzwq5HbCleNwercihCdUvsx9m2+6gp7ecvhdDTLSI0rcYq1SWyj71nFKu6YtnpOv
SW6t8ghj12Z1er/VtGMl0RXkXfYcTVIlzY1oOPna6QCcWoShvXKKWBt22ieeo+C+R2J4x4pB6OXM
BclJX91t7agilpzbWNB6SsZpq3EJ9sq58aSUzgTWeZiIhiaB0/xbauXmPKVZ9iTIE9xuBhLCLGuH
Y4///IMbCA5CHYg9ltqWKuATYTut5vmWltbXXXxcd3dCjcrECQAZ3/i1FLByg/2iwXK2M2uvzAPx
V17BjPBgNQu7BAkdERrT5tjb/ivTc0mpOjISh2nzjZ8pe+pOh5SjkTb6WbBsMSiSdF6VQtD3N1sA
xrgAyI6FzMXPUpCvbb3H37h0H6iLckSq1TGcOnNAzZe3+ug8xT8+qCJHW+MBhYGF2YBLLw8W5+zs
FuBqJTA8W6dPibr3wdtp981wdmNqLyla5o0JEFkydjWDorAvXig9e6jTR12zCGO477nDBI9m/ZKN
zvyr0tIN6zpW2CMrCsFLS+Xt4fheP/g3NQKzI5dZ9ifbNB/qAK9dJTM1QCj3Sbeg7hYikCPw6Ebj
VO0ZBaNkQVNkpfgNhftlVtnpTAW6bH8m43VdApVr+wOW+5fi/rQKgSfJW8GX5YKTbadeOZuWJzFH
enBbbsozACcN4ziigVNl49Gd7pxl1Yk+a3jQk4G0r7N6Aq4erm1kfg3ocmI41T0jf4K6gfExxU42
xgqalVcNqeC4Tsk+ud3oWDMw6fUjnC246yF1yqDSmMGLN2w4xEiJFwt8AvWXqOIGcte6T8X2wZDP
FjUJTcGJrLZagPd2/6fl2wkTrS98xUAzKqeCiDO3M2WNsYDHLwO4pJHquiWt/oIQ9w+I95G4iLP1
b75U1Mkz1AOb725Qmpnoj2lym/DPp4+IrtQPohixf+BZyRai4QefxligCkwZ/71xi+26LrA6s+UA
4RUgF9JlIxZBgsrPSiioDWwuXAFpK0pFoJyf30Go1+aNRHt8J3bZzYtFq27CI8Izuw+A71UHz1wF
7/M57Dedwp9E82xNm1KmQzVoAvbj95qtnOgJm3Vuf8h33YKuPfQH19oQFsdJUFhC4myB0KzifBG3
gznfJiq3e5G4r3TD+n467v3DQEQzByQcs5a3//YFSGY5ldBhK9W+kXYzG0u7utBZe+yKTdiHrrdq
+LkPJytFI5ICauHzXnVnohpr41LQ/tQz2fQocS0qt1olgNhBlLBIVsbQ6KtPodqa+SiKql3onW4z
4MzSHwx/ZzOsKayA/KpBLBmAk8RwbXztirL5hCifnq+bmYQEqFHasa5CUErNVcGb/6DCfkbBirh+
3lZBtmPXT8Zap5QCcm8Oyjx8k83za8tgmY0FYz0/tplrOsvrgLsPO38TO1mgv8WAlohhLr25dt0L
GPEss1vg0+etmZFThjhTE8BNwUiXBoeDXGzj2CM6wC1RUw++pDC0dMQacaTBYbU3VjE984Gvi1ts
1WnwIqW0Df3SZL+r1taquOOWZv2dIPi9I9GHLoJ6GjaE1trGDrVa4DllK92DuMJaQXrUWKvw1lN1
NErfcUPXQqqhbf6b9I7FC3hzpudJddB6sWWmDJgWcQFjOHgjAyEhcl537GTJtkr5RGM1sJk1lL4E
0LwRJ1VpKWkZDDCFc38xOuesizbXhHY+f9hdDqOicbMJpRPX6gUnS2VJ8Z37Gedy7SNiLGYPrS1u
7d0EijSvqjydC4RatpgDppP7O8a+DkO81Fce97tWwQXMcGjWEk1iG4lTERiacrdfrIXj2KxYHkgq
WHF4DZX5dh8ncm7aYI5/hD1Ftgxvh8maC3Pl995o34o6xebT/6g8IrRHstRWVmuz7c9SELdfhB2t
4A6JIIkTBAA6B+Lo3S0/A0bModaRG3SP54KM7fy9cHzuUfS5ToM7G13eIhuieArmV9Fm2V+F8Oyz
WzWCldSMG0lMQVVm8/IfeK03nZiz3CXXlnzZ/Q8LlNBWyF6epqDaIBiWnqbKH9p7nwRqkYRswp4W
9duxlTquMKDsyBihtPrzCAbk0HaE9kAtNKj3DeWOKClAhvXomDa6byELbjysG5+wdz4A21D+WIUH
N7jlCkzZ9oW62OTqWSKSE1KcFAxFlrZxPZz/XWTMdEfaH3k/XhWzeh9deG+QnBrGxU9Ahl8mgfPf
mEaazuyHqfj2aisYIS1lHdmIGAraUYshRLN/axHfOQtbBna3ZrQT7r0W4hDx+nGB/rQFdfn60BBJ
q8nF0cl/veRAWO9pTgfIWiV+xp4xo8+PmAVX9tAAVLuGbZmSNaRXG4YBaN3aqoI70Lv/5S/bIAeD
vh+8auxCju0+AR1+G6djxjigYz22dU1/cUV7mNSmQcdIBWf5+Lv6fakUFN4vx5QF2xxAZ8WRIzGR
bJDfTsYMTPORn0zf+LaHX5kJyp8lIGcdvnUHuTyMgU6Rf3/xY1KtcGMvc/vBDxClgKZfXC8Fp55o
HVNdRk4/rNxgo8mKXI3EECeJmGbo75xSBOA1ga5hTZw7saCWOMkrXJMpRm4pQU4+WoUj11VfTNaV
2RSxLWm+5OOmBl3TX7Wm8F3xZnaC1GFhozp9LUMSL5TSycRYXoXIVDjb8DYnxmuYNgxg3on4Y0fA
e7dPNO13eJk6DGfi+jTgYhF2P3hANkj1fxMl2bpk4WUKWrGfxFmh0kgCVfvFeAai4JGO4V7Vveuu
rDUaMwnWy+Rrxd6Pi6NrVFGH8huvOeiflpNfkfnHO2WxHusbjEjeiMd8gfD5/0RuYBboXiWx4zTc
aSJaDnTuQdjJN/j7IRnkaSP7gQvCAvW96PSNQ7E/PA/pd3MeNqSlox3TmPM8fhKYi5yk0zVjym6U
3AkW3ZeOrR9y/w+y76PlxpgBkkDZDteYX0sDhglqWzJAeNVOc0VFCpqljWy5Z3i3NV8zxjTd58tV
T5kr2CAWOH7Et+pDZYxEiiitfjb3mJWemovjbDveDjZnEQzZGELX6Exi7k8Ox4JScq8Bf1ZuVmyp
IlEDXfjUy6YmvcJVHIWb9ZUsnHz09MtZNJLf+NHFdOGZdRFo5vaDJFcNzDvbuHvGDP8FpbBpPrnL
SMBqI/VQPtByPI7ZOiDU2CehfIbxAn2wzM9SokGxpnzUF3LNql+cNncbMpLBucPQ5bv9IrXQKLIF
RSQYlw56OwKRhtdvqs/e9fOyYT5IVAMUOlhpqTQyyNGMiur6kbUR7/OwoiHeEHjqSwBt+Pnak76m
d2Z2csEfNZNfithgHB2QB0bd+a7u+pRTwk+s966xAlTTSX3c5lz//BX+w3gcUUf/XXRuZS9RG1eQ
M0BxlzJHkBQa46HFBLbG85xN6cT3hJeiwsi7yO5zsLvpWNCSe6oLi0FRkkj76OGVRu5MiQV6U5nS
URFDebqZHCQQ7JpOT5Cbt0uMZj95wReRyY+a/ClBNlSZIazk1bhqjAtEm8392+f7LZ5CbjRrwnSS
BKsLlWnm8J2tViWWimvnkwjyYVvIGpLhPYNt53gMLlfbg9jfr9qJeSdN556myNIfuA3qKAi1Y/Ol
k1aY0YN0824sUL+C1WXOMPdhqTqcahaFj9WwivhGVMf1JqpNaJ7PGJIZYOf08nAq58ENhHnFRHP6
w7/Sh/k8MxWqL2rF4HlSS6LYy01dOmt5HhuA5BUaKLMJdI/6hJxiHoIMeNo2yV7rkt0UG2xowK85
CKyFdr3FP4Q8Lm5WH0Qn0P+7Aeb8ga7TtLKa3NJ//PLe2X6K59M4pcEOnhGFWKHfSbHLzWFy99yK
AHOYVcJnLoHUUAZXyTLEdivsxCo2tZPaqwleC+OAC9WRJhv6Vu20gMWtRlUOhfs9Nv0QNhhYn07o
RfqDZhKZ+T7ecayxzQRuv0sk+7U0wh1rilbQwGjO0IYzS9dgsD9/gkd2QBBrJ76wY9e/zwGCLZiR
y/7d/IymPe0/NvAfZU7C6/n/gqe3MBejjHeUSjZyjTbrxK8di2SshpedRyLHr6MDg3QWijk6jmZc
Nrsq29iYGuDiunanl4QvA3JaZevKw8sBtYiIsV/o7xuAzZao9Gp0TzlhHC6DQryvRRJB1Nujjqw+
WZnsqSGtkT5R4fca3ZnZW9IN7AfXuXqRmEsDysAghWJkx++KikI2i8V0fR8GighZO5lz2ROOuAxE
gkjlK9Ad5DVc10hPNYSIjEh7dCbqcrUfUa5gOJzNehPLhhQFyqoP8xstuCbk5a3LUr7InoB1O2aT
2ddXFMidB3c0TPYkej/RHq4sApZ+24V8QMuAmdTEQjmG6X+MLHy5M56F846Un4kUOAX+d2cXGYQO
ivKd2dHS8Pdm/ia6krgN9kMywr/pJk+JhrqU1FIcROsoFOgP6vdVxJvfc1dRY14qy5WeGduwUZin
URNvrfb1TQ5SupyUd1/geNlXjxFLkIwnFX6Yryyc/9x8lSw8RdyQ20oFYqFUm64CNe2NV2P5xR39
uE6nCqX98LhZ1iottlxvoW7+XSZI9PhjLRErlImbrp08EUEeNPhHJGEmzjfWVnr6Yb7F0FIjRYb9
huzwvDTTRXA2UFK8a1wu7I35JuKnsxM6E3X512Ql1uA7e85HY913Eo1NPpT301lcaMB3bCTjP/Y0
mjLsnmbX4k35vriCWj6J3ThNrCmCbx9BDZNX3iaTmdQIAbLWxhbKYspvVXQQjEOrpV7VYquX0oCM
39GDaoaFeiqICMEvTg+rZRN++xIk2CFeJSEIWSI6u0NW7oMqLR5o36Qhi3QWZwArZo6iXRPOyxrd
6pwvcO91emy3hSE/20Ptbn9Xfmu71/D1wl9KQENjJC2Wwu1epawW/sJpAug1mSO7UFTsNytqq/e6
re7acqiH4QwVkDu65M1pmPKgGIQIQUctsje3q3pLdWeJsfNpcAJIV3TIfjZ1k5T9EgzT2yF0smKB
I7wbi1zw79efKYkgR55ejac6Ms9RWEQzT4Bpj2VfI/j6JFKhc7M+2DiM82P/qUTm4T/9/kIQxxSe
2tn/b71nGf/IGB9dyZ4jIpdtLb8VSfrJLRRyw7Gs+/b87SLQ3L8VfcjQD1ScZ9M0FoOk3fjGkfvT
663xKvI+vDqj7gElmZqfNHoec3fxByAbMnrYwx9UgCf24klhGKclmd46LCktbPdLQYv6k7hBoZR+
FuyPEjVBaA0d57mlfTax7t9BM7dZ2IYHWzVeSYE6vsgtQ9mIH7iX6TUL2s7V26PG8yQjjL8XuYdN
RJnZHBeCkDngGChwM3qQWgCVWw8HpaRexy6ff9lbuL1ouLrQw7YxpEEptgeHIXva27CXYSWIdoSg
oCZCrCohAgC9h955a9Zj7Hr+C719SXNwYMYK76FKfaO1LtrNiZyPKYO6T/hCkLUt3f0+AWBvJQVm
+4h6nNbrjCae4vuuGLqcrpYPlEkifvO4eZq2Rbq/1Nbd6x+Dd9l/3uyNxOJmY5UggNHG1ybdsxeV
cNr9TFvE12TKkDUnHggExJvtJsjMAN4ykqCZbqFoZ9RoQSJHMZ7CCcH3KdSWN3dm0sH/0s3KLxJ8
Bi76LqXS40O1yyOTaKFqoOzLqQZm/B20p0LRb50faS1RLi+C4ySJJTY6z6UIVcbCXluaOzh6Gy1s
z+iMWjgtuhOHCHtN0el0M8m+FuCxYajzM8cYZfkUQSq8whLYbxPE9+oLiFQU8UR3ONFsUhiQrmRy
rTDtWS/Fj0JVjdb9sgtpxGDzUM6W7020oGsDQT+V8IlrWsie67FL4+mPb//5W5wkG2BQ8kpQUZ6K
rfbNbuv5LYDEH92AFsAgQ3IJoE/FTtms3Ux2LiLvp4WSglnkC51P2SPJ9xWHfLuCIokPX0H/5Opy
VIGSuxj9LHIDIANET/jbbdiYEcenymblZnOByw9IR78LDRtj16g9eufFwfdwrhNtecze9pIHsfXh
VcOWSlOv87xEmrK7y7DAYPX8NRECbjux4y3plIdX6+krIxQa+bDsM1b9GKr8TZZO7bz3xe5WegPt
LfIaE95rtrqwV+ahOFy51CSlqFklMOvQtXd9eBaPN2jXxC6XuNaO0nzAf4Ss5faM9qHtvx7Qw6lT
3eQhHG63V6+j9hURxPXDbHkno0Pgcu7T0P00Oef2aLBRbp0SOXo1FBFG42Mxy+1YrsXPOupCfVty
RQ4kIhn4fmKKkh0Sh4BO0mBUSzATacFtzUxEzh1OANlSb9sLaOVZ2JD9gg7hsDWoA4dmMoAEOkGM
Kx0Ln2K3eh5AFqRAb7FtmpqiKTidsnHP0RauA0hxJ6UsZl2SUheKbWnxdicGB99KxIq05wxNpMeS
/V4Ba+e053AOF/W/7Qc0v/Vdiu2x6O0GlnnNilSvfjxTJR5YdNA7miUc5NWrxybuD+jT9IG78ScV
b4amIDpSZmIFdzY4WXWRkI4TobqWcdLheH7fx3L9l+2GHH9sYhi0xfD31e892N+Rvh+nH4AxNTbw
iouRwPu+ooAzNNq/MgCPM4+oKPQQGyEIGgpbgVmjLU6bgQFDcBo9wBu7QUxzXLWtCOLMLpF5KypB
seklOJfSk44cmgirH1hReZ39ESq5K9vZR4gTbU20YLxe5bICzXY5yi7ayT1BF/jUrWpurl94iqru
sP7vUuNvV0kUEc40QTdtW9S5smMvCjSouGFaK0c5/UuvFkF2c79XkNz1zVmfuBto7G81KAUpkDSj
LkPBXD1fR0ZnPDE6hXiDIh9bmUsFgAX7Z4YbBUYcYjSli0teKa+rbVJqtQR0IX9Hyg29iXA4F/Yu
nhF4jkOSlPtjf1RmrJTZzy5uUh9JkWQnxJWaddZaEV+AfKbA+nPiLlkfkaEVScyl7LCcbRNS1NRp
RIwDNjkrG+TZTU1tpeIEzp3P1N+q+WZ5PXnMTc2BGU+vE9/5E+kafSPUlcX4Sfm+Xli3CrHc5P0O
cJN1LgB39iqt42QMhP3sbIdWl2sEUpCZoaX8Bpexc0CREbLBzrfplkW5voR7TDG7nlKJyb4Q0pGS
KzIv35hkYtGZulZMzb1ixg2rEGIrndNjGxTwZPxffxwxn1Xp5QytFQV1kem3QMLhAN2oGxO5jZBr
uJmikTskSgzMjjLbAqFZIUlbLUGeDxEXCsbdji2VResa3fLNFiWziRQifMLnoyEcs8CWSs0Bicw3
d2g0gYjNYS57SUj0DbAYr1MVu6ttFy80LWLlQNXEj1g4eEKZ7bL5Ci4t1QxldeNYiZ57Cww0OwS/
++P6s2Vtw9HAEGvLzl9EfoK6153DcmW4N94j1rgyTVZVrKLVrTooK0aB8v6FYXotaMN3EDb86/k2
Bk5OYq7qKe62eoJsQUR3GaL7PHphS3Y6L0p3WOWPskHGG0IEjnelTBORWcNwk7YWR+zxw9Wpa+e5
aMfE8vwNFZV1nknZRG/1GxZ7dXzvq4xF1+9w+FGdLiJ57lFufA4vVa5BZ5ky/hfrTcdCV5eaoep1
4CRxiOTOTTehLMb8cwWHmTJr09KzqM0Lor9iEokM5TqN1JxqJlySzRH8nDOwwv7DgnL9fAeZcQwO
gKNj+2K8kT9FJ4hn2ERsdb3eYL3t1WLCJ+As84ZkpavJ4WE0/7BT+KZxgnOXbrr1SNul7Pr6rTDT
ox5xdFHz+haBxyHo+Cang62jltHXskvvY4uwX+1ulR9fJ8Z/ZymZHo2lBCUxojutci1oA/+LlFxW
DpTzMTAm3KTxtl/WQnprcDPxk9WKw6r1y4GxP4u2wLA95XHI3J4LvvZ6A96ubikuaxIo0NLdheS0
3RCNwgjBPOay1vDLdAx0dm3UoSmNP85VMbW9LNaS85xfxMcHgHXw3x451k6JjfUJzFX9VRU8yY3z
XrUIW8ESoVw2q6T8jz4LSPe3NEDDIU+o7eow77uCjQIc/qbwwIjiv5BqoOx595L7/n4CRneOxtER
MJU4Jtn8N0s6APaCGWm/Gup3CKeZxbW3wE43pqIL6xnzq7YTzkT2cvbjbbiRk9E24RrgADQNoI4Z
THRS2h3SeWumO3NFjzPxJlXcEZIcJTsDwXuhtavxRDmUPECUOV+DGneAlhVadMVrQcoKMrfs88/N
+vLYD5xZS7iVTBrfZ/rv2McD5GUXjdWztfBB3Uqq2P9C3PTGIOdD2W+Z/iyCsQ4+GlALsb0ye5+u
a0k3Y5/FJpstWov4EGbkdxxSHCRJC6/HIPqoTfcoiMQw8qk6S6pfinaEa+bd9ED6YDGj4/4/Fwgv
2wEQ5VSINqTrCVELya1iacTWrIZiHrUIBqIOuZsrBjbuKRCMj50hpMazoALYDDiofAyyH5uU786f
v4vR2TPWDX5CpBZizz7AZ2Qwe3TgVS1JUcI3HUa0g4K4xTXyPAUd+4wKcB5A54B13J6RjSMfbAM/
VXM8JXOvCMOx5lRZ4uJzgy7AHHlo5t3Gi92d33gpI/pndJeamlkC0XLxqyORwV3tb5p4DDgPhRbG
6WaCQbIxYYjnWkMu1UVO+tv1uCMvH1pi2spDFwCvgBmwhBD5B43i/z5kzxrD/7N8NdBwupJUvCcy
9CXdS4wBKjeIjS7nkEOi+dRU4fPPaAYl8YLLYIyB6Q3517FiZ+ZCh/oTKHswF1vUamFJFb+keKYY
vOjOKTVPXZkC1KfHb/obmhMLrROzQnXyvm/K4yMMj8KdPWRDbc0L5Lqc5GM1dOUORo2hSUEQbTPl
lHU7ZH2qubx2ivd6arJ1MhV8x1LOsbRJ4n11Gx7JF2Wvz5t8gmRCCGC0RY//sXGeaNVjhnDYG35c
8EQBL0Bd7UN44NrRcTjyqMg7w1Tr/BIUFaedWlki0poSHtojERZxWgnj/Lk9ZpxTurtMBzWmvZi2
gqlic1Ur9sQVxVf+uaifaMUd3CmxOWVT9m6bk/2DgenxcJZqHhnxXl1aee+4ARpzjt9JQ5rpjEA1
oFbjE2pIQwwUTKnk/VNuDqkSQC18Ux44q/8r8CyhLePEgxSc4oZuzyQGu+jyY9P6jgt+AVVoGXqY
C+bYNO/0uXj699JEh6oKzEIDd5bxiKTRS5HtcheO83vPxubPUIdY9Au4CbT2K64SXY9PEI9yurvu
ZxCU6UNUamFM90SXr3cvcwgr7/HshaExlqXyi2/F5wkF3Nn4vP2RVanwSoslDb1fx84fyl4tBT6a
3QUl1NZ5C4tv5rsVOBaZgNG3umfJgFdl10rIe5YxFzgsnfdMDYqaXF9qhobY3h5YjyuLbDYsoUFX
eipieXkbuAq3XE040OXQVT6hX4nXnSZcSiDfJkofC6pmVLaARCjQFBi/1tVK5ij7lZcPkBP0hjme
oix/7BJSIUZYd512yd+GgNT+LOTHclg55ybWC0hDkPtG3vIl9ZQ34YD0OJRSTc5S2Iq0elvl/2Oj
RlqycLFI0eQNpAlte2di1sG0f5CWHMtoFEifLNKfjxyIuJ52Uy0i9pzOIrIh9k7UQXJjMaqdSf1a
2sL6OnSuaf2PRaZTaJn7fax0hzRHknpEMIpDtDlZM1wND41o+nCbYXWW3F2jGplN7w5rOKAlx7Tp
cIQKR+qm+ORIe2hWCjv45r8vhVuB1BEXMf6+hfwxfY7QFhRXTrQJlzvzlvIgMaokFKOQ3H8ICO6Q
CHfmMDAMrqoWUAzji/WaaDk4/jr5VLmOV/dnGLVbBl1dZEy/eOpexNqvblNfYhFoCtsKgSk2B/RK
N/PX38CUYs8UnwEouk6bkorFk60PgoSrQsMhZ7FFG3UCMf1XYpvFAAtHuJbqIq/FeeSGQOwffXiv
6Rp9LPjE7hC18S+neVx2iDkilNeCwiJ0BPmGvmgcX41aY3vnCjowYWQdURi285inns0gOw6vA/gm
IlItwu7N2U20yiL6LQbXWEsAwzExa/ekv39+/jPxyXntBqG6q6g69eGI2XG497rSn9J31NVhJ5CZ
tjszVh7STY+mOZmqoOuft6l7OlU0Rdbp5bsTu3EkijWU/zq+WcGpDNR6l+NjGbzatxzH1j5V6Q84
zbGSlYtlWu8avYfSpNMehmhHbHtsQUaD33/DcyDqq3NOn9C1KYjoYPfR3wyqAqINdkoVDQLwqauX
j3UqP4xYe7f9hBaiK2XbfvP6eaQFlZRoVbgq1J46vQH93DS+M0oP7ZbV+XKyNFnf7DP+UMoou98q
j+rJeLPeQyh+Nc4oENJajGTAY8bVMo5gLzmFQLlGajL6dCcZBneVSVwdFf7cKTteJqZ9EYnzBq2W
czm3puJ1zriQPwYP33ceNdT2xJQh3SPvyhns366NrOrsFRRkpuEbt7AaHHwFdvSp8DUROIjul3rO
wecDCotPQ09jOse7af/h3QNNuscGWBODoepbEqRH1YQnNkQvGYcG9q8EGvoppVJjE3+NWhsbEBdb
Scd6ztOLSMSStfaegc3akWu4BEgKuoUzD10hC7RSGK+GnCXgxAoDDeR4Sscyb/qcn8HK22cd+dKz
8FkG5JSGqoSjQFJmkb8cQ48UgAHUabYZbhwHgtFeHChM49XMkmXHtFIIffVQu23ATLAx6MFzlSqS
Sg7O0WM8rVcLnk45aBlCjo1INuhydCiQdNAabraGSjd2oLSEiSTbPBkPMFUS4NCYOVgOqEu1gomS
rALMYm2GBEFq7BbyboR9vED8xeuhgBF+yqWxvFUFXZ29hdVPEu5bEC56U44VugPkZWL00Xu/oN+x
a1HXuel4Byg8X3y4ELIBiaZVFDBIAVktV7tjUVleOqTChO+Iu5COYx7F5k0ZODna9gQP3DT/nZtx
JPCbo9y31GM9pTcc5MQKo7xJlRJAmsn7iQgNYsQaZQNbnAuCygw1Kgkk0I8t3JOYZ9C0Oashi3Oy
JKPktTql+u9biMw4PExMmz7LIyPP+2K3SMps4c9Ws6OQvtA67vdUNtdBuZKl/Am/yEQ9qfazj42K
0B8zS3uYN4JCRPNBUXIU+vGzC46vICknFdpUbjzyd2IwUlmc+z+6eHxdPExzLVF6NXIUFHOMk4FJ
YXOsVZGnPm+RYpe7MVTh5ZcAkxi64bX3E3ywjHZyNG67tJe9lfeWKMZSmlL7Tbk8a8jDbds4SdAR
xknIc4KnI5ttnP/zSWnz1maRd2QmI+ZTSZBSL8j6U6c1K7uNEWWQ7qfZcSJ7jkMlKIkicTR7mWHE
+6jW3W3xWOJiUt6kb91pNAgyqKBGw559cXFhAODdLe45fApIpSA3/I4/ph3/utJ8i6W9/ZjaMNQ4
1jNK7OMPN3y23hXpBphlZZ+9xjoG3xUI6xMMPYoHXPWYaF++Da1AC47vNchu1HrYZk3gMiQxUFbO
dreczRENUPmWxPDCSBO5U2TQjlIXq7+cDHNOefA2dW9UIuQaa9nTVvuqcsOLANIyJV8wT0oMd9yh
eK//vVLxwCkzkWxnl5l8gBT3ztLH/LQEGGeuoPiu8J6a3W3tKLq5dg2tiVCCItvI8xo2t24Xr80a
ptIJ6M4PmR9vlUtRD1NhdYAavWA8muEY7ucwwctNQmuy3eClBQ4hadW2gpYq3+QhQAgmHSgvaPAk
+pMrWatqOLc7d3wLXew0SuRLBpoNuaiyw3DxxRJN2QptHPPYJ7WVGvqE46W0pRFmjx3FwQXkb7KW
nlDrJSkjMBlkoonHhMzh4mS4nBQaUvI2La85cOhw629hKI6a3GlhuB+ehY43I1/jQ00M8/ethFSi
NITDSr3XYTQZzLzqKE3/E1e96y0HvVwNwEwSHZ6K/fMEpphDX6PEfYMBilzwtDVmW2A3udTb10Gv
b7/eIxMYYtX9YfeYJ33z6ygRvRHo/aflRtP9f2ChECh9fwsGLpC6OjCBhy2N1W6bl5G7A+Zszwil
aDAgWQek1oMpPDpIgBgvLQXYw+rJOkQq5bFugOXKixovoIR2YEba26vGhhVVsMYLqVOsBIp0xSBZ
h2XO4RQged3eDltYXsHNEYeMEQJtk5Gm3sznrPR1/T0ozE4qgkBr93TuOseJPGIK3VhK9+7gsslT
QKIAKGofDoSIc02KNAqemZ0HepoBweEhw+QkrMkZiyIVn5zg0E/36EhA14AQyL+jFrW0K4iwiLCO
HMG7cPNgsdZbg5F6nFuVfq/fNNP6XFL4N+DLX0Og5GMKrfOdCywF8DaKlDgbq9HJMy9Pfh7QuZJv
WV/ckktZ8Vz+o6kw13m/GXUmEOjna1IB5Rh3Oo6gI0VniTXMzgOYMe+RxFMs+p65AktG0vADG7Nd
8CLcOK24ajALt4/13DEqSB0am7XCSQ/j3t64izVJqSalQzf70JomkLLo7naFrz6Y34eoMr3L9dXN
Pzo49LHYR1ArrHVPFHv1qxbXWxSo+HMbpUnxsRiAh80OytyykAPuXeGFDHngpWAZQCQiScZU9sF5
rPE+5hZGl6MdSxE6QQw0LXtiCNm0Ee4y0ccwnVQ/tKNEJKFrCP6DfXQDRxAWbFvSMxYPHbozAHob
rSJb7A2JuuluPllfEIR00dhIroMkZ6p3LXHV7PYkNI/kfyj62Kn4JyTWJALGvLtmcTC//hVhT/AO
lJkAKAtBtvUNsIoM4/YuO5vLDwN4jWvrJdNNinKKvvajW5/T3UE6cuXquvneeXpu/GvCuFr+58Bi
He/YJMbg1G4k8eQ50Ue47ROIaqeu00mLsqXqi5AicCL0O0QB27872qEgJt4MoKKM4gmpJVLvuU/j
Z+Rsyl8DPeQ/BOOD4NlcaozJllkcvLRZlEygBV8RxUWK20i34lAxxLTaNFJ0eOnqNbAZ472yqqFu
uK9n4hvJm73KODVAIwPXN/AgklKc0fTN98jfyo8EAASe2jomx8P31Cj892SyKETgBd8pWSaVr4Rn
rVTRHMgFMkwW9m0Wjv5S66KuvtwL14PjrF0ILi5xjhwgYh074nTd6yle0DkxIwdMyM5zuIH6ZvIj
YLkcJ+TFchFEUq19x8SRc6k5MwNC4EgUfENIrLV97nbqbHsWt+n3hyfbcLPca0ManSeeZoU/aOJ+
dHE7a+quKgUreKvQpSKki5e8mZeSWbd2hcwZwyV+32BUo3gzeiVoJ5UFqceEgpSOGzZmvO9IJetD
DEL/od4mIFtvZBSOO0tJ7GEzIpbhI4d7AtwTiAjVgCzeEIV8xvN/22Zi/fA2NZuiBuGzIzJiJJLu
6UAs+3h0C/3Au9B1pprzs6J6qNl7C+2Sx5+jv7GuluDb2a4yTEKLX02rZ/Q4l0zoH1Vzllup3jpH
cqaHSo226ZsQmM+VK+afZaucHfHa8Gwk8P50Gn8m0H8ZS2UaU4B7xuqW7R2JJNV9B2gpcA0yCe1B
E+7JctbcN074TJIt9CFCg2NCIuGxx9O9/IZ+1PvxilI/vN3B026sYdv5P0neJBA0dtaY3RKItkwD
WfDD9axZbfRWtlFbCNXW48OebjuQIHynAAiLLe0qiIIoIS4bCtOtbw6eo+XGzLZr8NXRU+2amhMY
dyfrSx35MOQUVqkNIC+a3f4Q/Ao0nd7Vx78BssQNg6/Nh3ChEyiTGFeITNYaOX/QjZHaaXdtmXz/
uCJAMuTY1zs/a+MAojCcksHlkzEE4S2ZEGhx6BDkLi0FKFKD/kBe1PXqYEBskHXo2fSr6U6mw8Nx
hT6/7wBE2LstEK22jFWATqPOf7ih9l+0rjC3n5eNPh1kuOyMEMv6U4bOtf2hdGI9Gfe6jcThqtHI
RoxKSdB0+du7zLdDaynxJGjnTVSDdTDg5adiDkErDnK4l0SA0Eyn7dSprq3O/aPNVH/S6k0VnXjC
UpAMu6xOQNUZVjvTbGHQbUhZ5Mz7Alv/T7i5+ZrVgt5Jd7KhXrNJP8aJDhQn4iiYDB/NZIfB0eAF
bN3F2Rohh9kKrdVjlsp5Vpge6H6gFbl5nhQqc1OAq1RsnVHo8hT4JSbVJwr+xREWpAoslWuUNjGm
mFKoZtlGdYVK0NzwxHLH3KEDjp4JCO+HMGquSyZf6HOykzN3NMAn6u0ZbOC4BB6c3NMT5BRAdiJq
ZY+JXciXXGa72K2sv0TDCRFaRvEfpRTfFip5WCV6IjZPgGWJYVLTeJL+hcIthyJ2LmnTCWeIyx8l
OOI2oL4ZmuljtZB1TeGbc1Ik1aLZ6DAhCUKYPq8vNe2C6MHjPgn1qvl7KNZtGA1F+76i3EaYxMXy
QVLcorXrYhdJnt3ak1Aip40PBqbBEilogAfO2IUFlbXfAUh+qmm+0DlVPiZaGOKs0Wldp7ntiF/V
loEcyhzFBZbRH4FBTp3i3UmuPdl+Kxkm7O88/30M2EnUNWkvyAfaiTU30RBNU3U6XK9DNmOXZGHh
jP8uI2iG7Mf2g7kFvv9EQYgPDZK1Szd2U1eIF9q5Q3ZHqzhokMMZixBfvcVNALO+V1B3fc/8/59h
0x83TP/uEqIUmODhTvR9nc3bB0hWwS5rO7uxgJS7vcgTp3G73l0l+BBAtWnRmPSORPJJHoJ0CukS
HJ/6RCPruaPKwwPUxQxGHoapoB6m5mqAy1XVKkgqgENqgobP/2jXsqkT8BcrZWGi9jQFJbrnOCsu
QuM9dtiTFnYn7GveqJw0E6WIswlq6k2N3TQODJkyCcFf21k5JUgQIL+PYspHFljanjzILykAoUwj
WbYdeH+nC5yUlEV94OSADHM3FDdyrtw00xWT7pLhd6N6p7PGy0aYQyoKy3+3EqOYRlezPxNYRpnO
PfsI5Ksu6/0aS92R3qFhzSzyz8qQZSmvTcRT1Rm7mzjMbY707gQ0oarZa4SqcD1v7J834Q4y2PwF
nB6nU53HsNHFdgXm09qQbN7FAKk7r3J83sBkMzpCEgK9kE929ZfpEojrG9upsLpRq0DKzMJuHXuo
miT+1CI0K6Xxm/ohHJ+yJmy+JrjlkrLpe8kQjvTBfT8E121GUqTSVwbNC9t1hWrlpRROfRaLKed9
an0c4y2J1Sd9uv/ERMaUpqprHjfYpetHAekEsFYM/uLEU972MgmaB4XZClojf0Ule36k1Tf41byV
IFP+3KVc+hF45tlgM6EdJSpM1iLPzddRVT9cZ59YAmLiA74QLn5+AWmGbLcosO8Q5V9enJXglAxW
6TudNPgg9zUU72L5FfYYCvI+E72KxUw0Tkr1sOQmu3WeXJ8qHyLf2sqqSvhpGGfDtAXDqjQstZdK
mYCTYuqKWKTCOwsBODv6yE2XEppHiSwriCtSv8mHxgdc+lSiNbMMpv/sXUSfhgXSIhwuFe2ABPxG
CFUgNhHxCYjkpYIuC9F73ShnssgDX4BTLxMuzuXrt09/EsjPgDfwm7Q15fc34HVgxTIM1sIZq5Wv
GhxEE1oBVTFQOeef7Y8z/wikyNWLqlcK8njeG4uaE7Ue5E7X+WiuTv3TkmFanMzPJOxarKxvtIQO
y3cjlZ2wOE2Bj37UvFpZDstDflv+lcmhDfB86LACV3OuNg1VU4tc9vxDrjYkaxK/c9p7MZ1RtCtz
KY7fpFbLpNMXfCdpjl1raHmK1CGKAizhBjOpXhTVyeNpmIDtkMML8+9vXNjoncpxmfnN9NscRPr0
WOtr8VYGlSIEU9+xE7RUt/4gWNiQNsWAteiTgX+xYvz/icqp1g+a5HyCvFvCV08cjxEpcv35iE3G
FrgegGM6H2GMbUDinJZkZkhcF/Ibo0/1Ta3uqjD+9ygk4p+ki/+1ZrLtxT/XR0NbSvxy5fPlIOUe
TmZXDWxx9rVCq5+MB6NEosbM5SXiy9v3jlr1WKvaeWW3iMq+64Y+RkKCrrSzmR9qEXo11j0wgwGs
+hnQotfc9hpI4r3MH5anuP8EFZj29wWQ1wkyEd2amw2D6n7nebQnxXAyqb+TbmSAFftp7iKKvXna
vzPQLiSUWOdgyvY0SCgm+K4+UQDm2HzBPzSM5+5iOYuqTFPKQ0akQHzB74+iTbEaZfAITQcFpDj6
uIMC2YWMfh8tt7e51RExIe/qR5lXa0makjot2jicbsDj2z625QyZVf4+GPBHvNkG5YEL+B/9SO/q
b1tgBLhONBDCa+jIsFp/Jd1hL25v6pNSiWkp89n3pC43K0w5CB5GxnFYjLZFG9E5M20E0zrb8H5b
qK30/VBbjLmdCPr/4jcTrf+StjirhkL3itm199wYxOo0V5rCmCrlU1yikV+c9DHt5I4cBsG7k6Hn
fsr6EFHxf3hnPEK5vQwCl95e0Nr419jQcTAnkwdb6Ev4isVEBhhbvPi4/HaD7u2C80hLLSc9nUpF
5q2U6TnDH0YLt33s9hjXUjN9N6gJE7Fqk33Vfw6gwgMMsLWWUeVHboC+WywbSdbZTRTJEf8xKu4S
Uo47h8SxjDnEssvE4l5DUF7B5PD4flsn5rMnZEA61XBt9Jxede2FzBoRgr3z9kjZSS2ypvRWGCTm
JgSxWkMBE+RhYeXRKVAsOHsIbpUATLNXtSBolF4y9JcIQQESVHfDpsmGlOu4tPC3eTy9V1XRzmVz
DCOI2hDw2N7GYiCxkzgZuP84wA0gqKyKP9Ayi5ejEVHJGp9XehsUWwHSpuea8oIShode/ibOc4+J
eFaP6eR6hOmTLh/7kTqbG8KzOXQsZbdB4RejZLmk5MLa05qBzD5Wqk1KxX6EBr1Rn4ZSizkFAVfd
yf0JZNAD+3XF5IB7nqvQfytbOlRyqrTU/l4hH3XzX9GmEHAVFMTkpmW0B+tZSXU1AOmHY8yFGlg5
G5q9vPPjdPpwiC0TbF4jCblPH3DFFq1dMZu6Jshbun4pT2Zlmv+ykY/2qEiOZ9T0oULO2ocU7/qZ
dfjl/80rOpCUHNouDAAbidwmJww6pSeavbVTTrcA6dMGXN8uzsx+fsy/s6JtvhC+NhVmoYtAdJLx
jod7pGx71rOES7aa2aPE4taATyJFxlHzT7qqj7YE6+Ct9m2r12Boi5axO/sjYoWjCaua8pb4Rr2w
Z/lsM88jBzG0ZBvNsmAIWb2MCdw4UwTdRGdD/VELIzV64XXxPofWmM3KTq78vLNyf4QwId2Y3QMS
zvz4pN0ZbX/KvHufbFoJvuIVYlLS/w0v8Kbi3pmqGwkxhJaEp2ruqaPh3TDEFxvm1zv/38zxiUha
ge9ZvG3ihKum4a6GmCFt4jY5/B5NTa1uvLInZlJB8XyaCzigTAAJCNl648kY/30uwhIZJq79Mlq0
4SiGLo2/97PS93ut0L3HByWV0Rlz/TdFw3acdLnWJHhZroDhPkfRKMMRsetQGLW3cmgnsk/w6kxQ
87ViU+rkDOsUIM2lKr6UrRkUJkOTjqdNW5rb+utuqx5nx77Gqlh7eBtvSYTTm5n/ce9k+XXSJgY1
mQAAXPhiCvCusGOvAtlZJ7+tMNGQKo94Y9yXxvQcPoywc8fwajZezGldzRd3FNpWxaatJexBcNl2
UDzAfiNOGVB8eFnJPwJNmxQmeJjWzTvuTBUBQXUrEMqVO4yrbjcDWJWiZcQkoosPGmqyXkx6dM77
4RZVMEuW3HKPw3NCMQLZR6Ei4b4jMsrxlRnO3439btPTqMUJzN88vZdEf5XZMrMWU2svm2nt8O4K
M/0NDaN29KAEegHRZsZUoLPckcPr9l8aV2YVQawCv+jRVRi/0tuUDx8BnTzfpOADd/DrD5Agcup3
yrt+7PE0ryAqcwwU1D1OgJyQ8O43VFl2F0tVD1hGadl6Tri/kFf4awRDlbpY8qj9f483Mj9iU1Jm
xzrQZ1ciWdKEVqxDtLh8vKXj5kmxqQHv3KSDC81kuXg3uSlFgyY6hffKjsSCpjDkpVdvhBmvTsJe
nZ/oBl/hWYTNPNdj2QZZmgCimTAWpWkMN52ZpOi0ykkry6RfZId0TZp0lXLLIuqWqjRclShZtKgy
QRuqHP+Bwe5qe6XWrkeBTTw9r43OXsGWe5l1MycYGL/Np+mhH+uYApl1JjnfTrDM0gsbpFBj7DpL
T1sscMXPfNwl0RLmcH9E85K1wWGqLmDhDYbn5uJmHI/6RHyNQtz/qVQmHzvrKH0fbHW4wtphY1jP
Bol1RqwKDzpTNUs8LKaMAIMLlUlVHyFpozlj2LaQOYB5ZXplZ6VxOYjxg1T6BaSRk0WojeH42NOI
ZfgJIMkzEidNxYin091uaSHRu4rUeVlXPXrAcjj/xv8wV6/KSE9TjWdu7UU+E8Ro5zjpKNHgAscl
DYg/NykcZhTbgG9BW4bBUAjU4+LPB3Unb/PKVML2H03ZxQZIDzkHVEPF3DthENxMk5n/5dePGdcI
ScTTdyxvvbCsYMiKF77m6exDceRxgZfPGcZhgWJDy4jSKAzITaX4XUe/Hm8h1TifKmrDgyysgT5o
TqmRlAfd6ByL4Ckeljh5DP3zyaGDAn/CguwM7XU48gugfZF4vZpBn3Flpmgd5Ph97MnfNC7h04ew
TENGjUzxWqTT7eB255I33SNJLbz8S99FeRxsMw1euICyUbJHBjETpCWiUQefUWqlxvaKiRwHqgQK
Dwc+zm5c81GACpITNgvSWCVYu+R4+T5Ls5/rCAW+ts2RxYcBKU7IO/qbmPbTbYe3H4rxkzPkawZE
LhRS6s9rMQXNn7x2116+Ua/yE06fmatJFKlL5gXHBtFsB+Y82OoVtgyj/o9hUyOcUSFtjg4fFRwv
wLkUxzpVu//Qg5Zg/ppdQJGJPTwMq/qPVenpq114hkniZyvYtQdI+2dmj8RVkeKnBLyTRvrrrJMP
fp4KUaGvFoAJTM7CN9AIhrFq4qht4EBvzX9hi0K0miO9wc4a/tXa9i5WVvX7XRtWnUqn1uSb9rNk
ZcJ+/1+JwmTxvtessDUVKLCQWQTMfSFRYGMpgduKrpBKsZRmWneiLi3IuCPlhCBIGjIxylkJo8Q6
on8HmcYxH8qQxkwBrY/tDwWn3fuU3SbDUPcQFB4hF0Z8qY292n+JO7z0xtjsBeYxOg3P7grCmC9W
xW3LLRTnl5FHnfe7q4/osc5kuHKj1dQBAmszuLW+8qA43sn1IpYpj94MORmO2/phhlL/DVJjqXhA
Wkvsl2uDI82Yk2WtRHeLpBmTAI+64B38f4Ap4Fl3xms1I/+H5INZ4qvYUmpiqbiNJEvRHdb+GhQQ
HVglOGxqhgSmJmSa5/YwS2HpIFDG06gXHg4EG9kwtWKuvFZjF6KL88TYUrWtzgFSj3L1C+E3Rrwh
GFjwKP6L/oRVxkBP38J2gWY3zBckIvRUbUahJ4woouVDq8Fa4Nvj092t08arSiB6UR61gcvZnhsQ
NqkxRmv7UlkAUPsgLXQ3nvW2viRRzp1keET9Awwb8BHiWRWUQAUXh36Ka7F8xS62+pKRIFhzhZU0
Fk9bVK/Sf3F8O6nmu0avKD9E8IJYspSsoUwXcIaygGmVNsldAUNm0Dr3Rg0z4/gKRoLJTcoAaAC7
cXJh4gfwf0tQZXLF0ipybGh4tePH5HCJ2FbS/Fv1BH+x2b746mkRyuWpG2rQkcl0jB1con5n378H
A7Hf1O1TJt6ac5kMAo6yixHRSPb4ZpSAqtjd6gBDXtQJU0osKMpe99K6mMzVUh6okA2BEpgdw6Qi
alCmjf27OlG+rfqU3sfQIrM6XsVnW524SdD2CV2YIPlS5ZJkB9RQoNH6fkKQbhyK0MH64jy38prN
TWX9hwV5XrE90Vs5rm4DJPzglHV3sfva7EBWKX3rHJjYNyo0R/jjaTf5tFEDN738DNCPtz7gnpqT
zlyVVqzOIiRy6/Tc917aBMRAg1ShoHKpC95iA6fBJCzv5UByneYGdQJYRXVXoA1EtnmzYLwrTksG
N4dJqZqjpcdiMbkMOBOd8qbDjjtUoPEOmnMdQ+lNNnABAfHofyERxCWW9tmUcKfZe288mbRDsvie
tiAVj9JUPk7DNwBWE1VwonHI/NRq7EUKhB0AOwjF6Q0e+5to5/0J0jLAUSPYq3oxbEbVbBhbljHd
QMQoeoH+hoJQub/HXuiTt8SscOdhBEt4ZoiSn3Ykv6zxIBnnDynyWWdzVrWKwVf7rycqIcDroDh3
qMTc32mA5B8jK7M1sEj7uxWCBRJd5wCIeGlWvrnE5t3f8OziHmXNomrgwE3+2RxrvSEsPbY//RPU
NYf1DbUHOpdWWtsuAkQMDB1PP2eXhQv8vkjyUXDpGSWVVYctSSsEjqeKv8iQ/KC8D+kd3zfYPqMU
pq0FXaND8xkb9BfYfkCW6e66CKB4bolUYlR0lE+9xsfQgWNFVD9HAsHKBnAX1bG8Kb4h/U/zozva
TK4xD4JSvYXPzDXUpAePTpb5CwAEqYCBLOw7qQ1+AxA9I1VftInWjwa88ZtmgYjixoGFG7xIYVru
OqJcl1En0a+8LzSI/OyxCw/KRdKH9Bp9p5MQbssy1zw4O8w+a4J8owU2qJiH/KgpypPmsXydlIkc
VuEUgcyGcGtUDknVeMNHJ5VU80Tkblvi/aEBKOxeeXZKumjWeiqM7RlKo7cAYIX7DpPGEnZ6FgeS
ATxP+/RWwvtWm6O/b7JqLCQIq0XgZT+KCYPXMxxu6el1fPQo3x0ZJYZFPOAFznq8HQq1KPFdvWlb
WYfBOzVrXxO5Qk0QAu86+OvK2aa6FX3tU5bN/xc8icasVFVTzZEUyMc0+5l8XqtEC+f7cPQcZDg4
ioECKer838jqT0AaqQ4Yze06XHlhFsnn6RMDnXgfTwmVFlQU0lbzX+9zUc7VS7H9EphlC/oKnApw
tl47XLwaPFg/Itp4sJM/J5XrQ5MIEk9UoeMiEwWTq41FmEEVM1yEkN3k6PScIcjtViFwUT3G9LdY
Z4x1LvsFqCVeWVfSuZ9ekULQvnoy1ZOoD4r8BCrDqXcl9mGhjv6bVz/76oB58lU9FTVnQSoJ7zy6
9ubeQ8M8zWP3x8EM8FZ/GE7XzOWI1BJl/rNHY+C640u0/xvrvtkF0lg2fyz7U65yroY+Pp4rGW4z
8x3qRQn7vgmZSikHMHlR44bTdo2dO4gx4TEk9VZugDB7EwwP9A9APSFx5o6P8j+m+q2IbpDHQ4UR
Zy9nW9jfVZ/iFqyz1V6g61BZ1E7nfjIXLJz19iEMMs6WpEW6qZjr8SdqYU9oGonbjtyiYhGGzwW3
yTyUng7qJzwSgmm8DmrpzcJJfQA9PwpF1se0hzYKLeuewpS+UJ39ztA2GiTuZXthsBcIBHen+CZJ
qTrx/yXcE0pqyIFumQQkp5J4mijI9EFeJ7XXAxsfsbd36Ay1q44Eb0JT4hGKWA74ACi4EZyVH4nx
jLS0SHYSXUUolt9/fWvhKSMeFfh7/u9fQfXuS9bHrZxn7YuXjkNEVJ3tCruQhDiWaFwj/lCzAXnj
KFmfLnDTjyj0tTNeRzlbZsY0/Mq1neojZ0kGdEIzby54AsFVAYa2GZmNK2PI51FRfKEhBgtRvueF
5aeN34tDAnEJXG87rOR8JT2g+UDxsU8SpwPcu+rYIi2H3X/2AHcOnqwYCuefSdTNCrO+aGJLBKJP
SBPOhOgD59WH869NRBACwcyf966iw4k8K8lr0G2P+hmnVhwUnRfp/PcZxqLm/ee0yFYHH9eM+nXt
n8Jm08jWwp+mfTlMX1gUoBjV5gOmEur7mC0ZEFpzbgWG/WG4g2SsDXnWvWS8rM6AHxbOpva+VH/A
9gL/s6xZ5ZFm86KRFEDZZV5hB+/k/6Sgl2SJxMqm3wKUrVhJUrrlHQdr0MJdMxfJWV3Qj9PEv9aL
6BoEm683aBzBKkhkFUHxlx4mEUyExSNqArDkpRRsnBs4YKxXmtGHurs2EgLjZWLk4lcvXfvmA/KH
MNdg+qfuUzaZEc3/H36M8EkOoFhiF0SIFEe3GIQMyAVyEbudugypoMdCZ+AxNWr9INfxhWMN9dev
4XIM1x8crkVKHqNVmFMkpohmvvMTHcKveR8gLdB2UZxXHxGPBj7d/RAwBDMMsGUR9HatJe/ixJZC
zrH3sQL2/HxvqJ21UVdiYplmJnI0NF5HHdgqTZ9YRlHASp9C/u0PQba5qjjb3ham9TeiI/D/8bIy
appdqyiKwVm4IcOJQHYqkEF/Zj1LiX+HrubwkNBRN4DErW688cZAV9YgMZ/CnjZxVLwfmRTjf3vD
Bhx48B6XTEwzFla1xePUiactvZkuxN4KMkZ5+f3SmLWtJE7+Xg6ABWG0eUNgMIp1HRBH1cSqfPDD
FALdyumIIAiwxwYXLaDFiYdZmRByfdqDUinPCrWIGp5LStN5zM3PMHDfj1A1ceSzaMmhIKUA8nyW
cCyd2ZmziR9EXEd0iBd5eGYuhELDRTgzwDl/4Ip75nCOISA9auZxwV+kh1dtW7SBUUowvVBdV6Wf
BiWXJmx47mcm1/m74xcXzItjCrtGWzG6hAclXgemljBulvSvku9Ff/A6r2BjTlobcCR9/jmu40qd
xJKTwRXTbzFGnS+siWEHINosvCCDLmLEBj7LnYuQpiDzBMcibACaCJAOkfvuPyv1uoWrCUPP4uY5
LNTlo3k9XlcAb2BkdD2bN48l9unDY41lWz1cBzl1VQN+ixeFJQwUWiXhv1DvJnkNNWmybmuh/NEE
JCmQfENpTHArMdLI39J5gIikIWckFDZn4XkQ4+U53aXr0syF8QvTV7iz8joV3bvUdGgeESNYcviF
07BABklV4mBTXIhnUllpED2427GB6GL4juhUv5mWG0Z1UvR8WFyiCX78QCLXpdevcGyjeimnKbQm
KAbVbui/eTcUjnmZ8KBVs3OIEedu0W7lhmnABOoSt978TtiQV7qLBS5y1Il0sqGnQpIOE0bsqoj/
ghWnOdPrSK3weXuGp9iYb8j2z9BSKZEpjCxAtbQg6p2BySi5g/DaZAJDgeWfYL+VRC0l5oDhfcWD
8DoIxzJ5fgyxboukZMIVCLX8pp6/LvzGwoxvkXabK8BVa6W+WcD4PYSISZk70TBU2a7lVTBrTrHU
tIBYrl7lD8XSXSSplrNbQNFU7tOEGDRRfd2WlHeQxnCrPAsjrU7jfWWKDLhXxZm6RWcg4m3F/C7k
M/dITO+Wo0a8rxyYDjAeg0CcN/rH5Qdt4deXhjzr7nIVfofbwTOrvj/d1QZ3RhM3KdYOm9KHPBs2
fzhVnr6P6Oo3165CZYel6VyknjJe3Q2PG5pRrKhjJ7jUE+dHXyKR+AfD1u7ISdceCbW1rmJhdown
TJGUt8jt+C1TRiSyqBaMh/U99NrwiWV1E0V0BKvbEPHtkk/kk4t4vbmaZJe6HOfIlbEkkTBVXEzE
Spo59DG3iAMCXyKz2wxsi/rMC5BlZ9Z1bVvrBrQW6RNrUdfrbTmqrEIY84x6QGAPvPEbeY4tfeXX
VqIuX+jR94xey4cu+taZGf2p3W1zuLoB8qapTu+MzW74Y7ypRahdDlIbS4uPgT+6fveHSCqn2vZv
s+kLW3efGyft1ieNJ9eFFSp6QFBEaOjCdZpgzQ1MjNh6E2zl/pudbN+4Oy8d8BwaXMtakddZ0/5i
Kj0diKhZgSQKIjQO/2Iq3kj7vpWkPvt7lqBDywd/RDZUi8TunS1pKBfxpxNPMQDJrYaqCU9aSiUb
MNQot0YSGbgos6M3b1f4sWpoM9TwoSTTx6mxFln2PvhZM9Vm3u7Ht12leDbRPEzi4h8Uun1hr/eu
sL2rLMmsht/0xVQ3Gtn33Z01tGUEZf/V53aLlI+mo8zaoET6kbRi3+al+Ri9HApudihPa6EtuC38
Ra4y7EEdJQ5r5tQquq/8Od9h88+Gq6zQOlkcD5xgPKFzYtsuxkzCf5Sp9etPpxD80qJMu0nvUdT8
lRHuDQbf8coIa09x7EilEkrMIuV9N731u1k9riZui18zsB2L3ncSPSe36bCFcR+2Yt5XqB0gNUSC
dMbfhlC8PptzunWA3r3nn4U0A9o3pBG8mjqNOV69ek9CcuLi1zERDj0aA4zj5TAHfeq7JjYVAuCK
2JOCae0UY8UrNqpCQTJKTQxuf04TzAn8KlTtQufnKl/7XPbw0M8wwBDvV3wghYf0tkaRRnS7vvLd
hUju5P1YEuwlB5r3ajT9eK5Qn0xE/dFvS1DBl9gO/FATuIcT05nOXVvLnrbDimMYuKLGBqHqlNtm
UjI2jIBqT2rBya6gIPxMur4Kr3Mwp5lkNYkRNf+Z5NHueWOwyTtDDFmjmWWIQHO5up1DnvM+QCxT
4neHKFt73/VQpYQEJkh8n/VSED50Yt+FdiC6FWLZrVBzEHp7W4q9n8/cgp0B8+7/T6Cw9Yh8I253
Rro1gKi4kqjyf95ZDgHBedg4lQBFf0ElnIqRU0JzVojZQu+zj5Zcy6xxw7Cy4fN/YvDtM6KqaS4W
c5IUOwC78Ngbz/Bfh2pEA7HuRJO7yDT6mr0xde02SOxI6UEOUh8wJJbDRgXf+kaiJcw94fk63Kou
0f5uuC3NXQJDCLbBd/CDFUr+TDm8fh8VdODgUWtG9Ks8VZuptimYeU3OLeVIE0jTPIyhdRl98ypZ
lRdePD1R/UfbqKLS2Z1YVubkjF+uaYPkqspR8GZWPWaPhEUZWToo+D9kknKToBDkO5bCh7Rikkm9
gFWRCJvAx8hjQpHojZoEaWwqumHUJCCigZa+29COCJ2AeX3lzihQB5kWEqxR6jJAf0lGlk1pmA07
RaD9WO+xAmPOk16034Ti8hZKjKRAHwuW4pqBChPtqVwD4hqxT9kUINzaVv1SdDvMZRUCghMAXXMW
GiD4z0cbUEMtLjqEcpYjcAreWfb/lUpwke90PFHFM/2VnD1wHB553XQbmrLIHliODrQyzSpAFRtm
LbJtwTFJ7RUd1f+dGgckBxZ37kHD+ItAyIBac7Y7Sn5d+sHuoCCLinjjFbG0bpfDU2xPdU5mp3Yh
7R1z4/DT+iHd3P5eDSljexaK9xEAAfIoFcZ5YAElh2vuPBj6gWkUfOnFD71I9hohgXhFZYeRKlXN
kB0tn5YytfVKrJlBSTtXFSKKGpAjiYz6NqSYrKOm7/twLXa7G+fiAwDEtUwkXFdShh05WHBbURZ4
nVqiTebm/EenJ8wNd01nmhV07SSQ11BvdDQS8e7BsE3+vWu2EdItkT9GIGZnMkZPN5SNY1dY4hW7
2WDQL1+MEHHQ6UKM6VL0+rs9wqNzXi+SnZ3Xa/bzzCcMN2kAgfOKmMEqorCmjRz1uceJ/grPKGiu
bHHxYQu7rYofC/9q5t8wkNAGAShiugCzgIF1KSb31TczjSsD2dy89dKcpDHo1d66uW8pTzWWU3qC
E+/bKqAYyAXU8I8yX1cx0dshQzMe9WL7mto16n7fIJBW2WeQeYQKc0GRdq+DWNbTGWB0DvHjP2+N
szHcvDI/D18/ieVivM4a1MS+YSUvEoUfSczSgIxt70q0nAMHHna6L89CWeZiixAliMNTn/2kiRVF
Nh07KaP4x8WwnZKV+bJ3JlYJqO77WNyYyiaYJn7Q3rtoiWk7nC3uAXe18WGv8Z9gbrQsNcwOIapV
mkTG8PFfiOaBUMutd46eq5+HqJ8Nbx7Jv5TD1a64X/pXvy95KDj6Cp5Q6rR5jULIPY8phhwwYgdr
lq9URkuwcrwYsoiN5iHwSQ/R4KcpglgI5dOu8ORnFO0gGvQ7jyGk7fnRmvJIwBTBBBU14hgV3mWC
99hSqZ4ZEPbBsYCRCjFzCUgjC6ubLaOAV7iEzY50j6mx3Uc/6OwbTI6GLxKVTN0sQ15iPBDvfV8y
MZ2O1tPTJw1gUcDaVpl5mvRW2Qmst88hdo7Ywb2/ZKGK/inr++vmq6XYwcsUlKpiXn+CmFIg1djO
ZYbTwq+6JpCpMONUIzA76VAphtLno8lvNLRYNYhcMKdsMOyE6bmfUblmS/zZtmbUcf5i9nu1b973
TN3Yio+El6amYHwgNJ9N9Ok7YiT8mD8LiQgBXPkDMP8jIAbnCMr9yNwbygPJY9FDjiW6usaJEyAh
TsUvFOyMH/oMH3GGiWXNPkITqjbgFI+2DCOD7CmadugfYvMH+QvRr6Eas4EuZk0ekMgK55JZ6Rk0
jdivglR9XtgKMx50ouhD2sqwp76QwdCc2XOfGTjLpAbT5dY77NDPbCduZyphcqufwJOdvVznfxok
zb49KXf5T7MKyk5z5Mhw9Sh+2nVhnHo/HzjB9oBNyO7lVqE/KahoOpRRtZwKKocgPwIwZSPQM9n4
+88hyWx286ETYo4kSFKmQQgUt0z7pIkrVJtv6gmivLvFUKyNBV8HiaHwHG9acQYdBDD1AMCAevGC
GCeUiYz0Lzey4t5M9AGiGam73dF6uDwWl7CaE8uTCWfR1QhhY30g5am4zjTdHFdaxRCyNmZTun3o
cH/9GxJghUDHyjiCah27s5ou8WAI2Rex0QDSh1MIiwivdExPSSVwZUperG/4OJU/9N5PMkYW+nAG
0GLP4001mxlN6z61+xwFtOhb9VfmO6geuw9+5SAP1rLix5c3mtsNnvkkFcHqxWlrSnppMH77K/tB
ZgGBZUghC+R6EMJ3siQKPkGIMoWW753Hhko51yBbQSd3pZDQm6C1jjXsv1Iw9C4/ZtlRBRN8g8Wt
3CaF2RJ4wK49NPJrn+QCSF12DuALeZt6v41xuTai7PZryIlLGjMzMEUVKpqGuHvFTbo1JLpdB1al
RcseTmKwJZLOB1nyTSrGg95u02eA95TfJZHffDhry4yKiMzY5IkVeh393QLKi3aNLWP5MW+dceIt
I+bUA6LJbusdRzOsfwnlNZ1KF8euL/XKm3cJ1FfduYaDJCzKfLuGVUnDAIb0zAyDSth7BlIK6CUP
WVpnwkoz0woYUHniE9t1mLpDL9smmt/cr9J9GX/0YKDpvkcmbaNfrm/DN5hGMKN57S0qs9kiJQQ/
niYcXQB4jU6aVAaC9W/SmDdcyN3CrzNKf2X9N5BF7tPigwpMU4aicsWYZ1rD03+CwBkrT8P3KFuv
BngrjUPY5kfj8NXd/4xVz4+jS/qJIvxWma6t0IUORiigQWy27tDIKwwsGubnpC/d26D4j8B4jy6b
nRYCuEY+w8+YDE/qYTVDF+Xv29gQhvaJAAOs+YttNHI0CFm5mlrrOSXVY0Bh80QXdd6NA+htHW8F
jG7SYn/j9x+oRJSvjVH1JSE2dei2YXoGGCJaOWqy17PEBx9zq4ZyhPOIyejLAp00ZIyJoJIIkssg
AP0x39I+oDz5yDio/ZqBTp34seh7N8iHo11fhsHucVaLQiM+KnCFx50pR+Ub95rTpWkKLEuAIp3F
YodR8FFqEYHZDUk0MQSvqLltlc3KidKqbhOukZhtLvAbD5GqMrrvS9ScTTx6pX2O2rCaAedh8h/S
a0lE4OxXRXDmpoEJVUoNkj0Qi4i92gz5bEAkKSu6Jj82cXPJsAHCFg1BX4x4s5Fw5vbBzpv3oD4J
QuSyEAzz9PaKjpBmdXP9n2v5XPBfMe5gAMBYIbnc3oMIffPWiwJtXlhJRnbpbgaNKwbDGLBiRyOt
M+tOfoVx4MVf6as2lgYd39wVEV5mmBq6r/gRg/NA2fqpY9S/8sy1Xi/+9EDbHNB6Z61m1ZrQHJy7
Lq+JM5cUIpAqmY33j8mBHwU9hpxvNnrXyA6ko4BLCeoH43pMcJnJnIBpeZRH1YwKfpW0EdP3856o
OuhWrvQeUlONgEQnSUAFf9v+MRNtd6R2TN8HQA2/aiR45RXtnai6yQhinZKCPB9fEMwVdKXLABlI
ZSlfGEfxmjA9HXRaQh8ecBB4N1CiJiGKrAis00X6Xrsp6r110I1qMcw6hWydWBtZPJZNiDF5c1iF
JRxDwKGIWOfSRctiVkGz9YbQOJJjSGj1/QmE/9wyyyDkdALv4fqlzssE0b+14Wm62rJ3Ar7okzOp
W/oiqMxiRAILw5FTG6QLFutG27Ux/hbRBsJjjKgCE5HmDb3Ke01dUh8lSpVtVMeazll4VHlx1iKs
n4Wx9ganvheJT4v2f7PRhg+kwjiu7remZ4Nkbdmac+jxvfRRDMYcBJmDap7t5UPDtprS67mlOIVP
z3Pnnm8m3RMffsbPkHSCdIvQd5D5k90+UUai1tKd33UOuDRwpWJN1bEonrJKJzwYzWoIBZDudTdb
L4vwyVQ7YGkoepCm9u8TCW89zP3RquW1Kp9wFCXIqqyTa4rAWqJv1acBDO/Am/Xg+7SZCH3XXzDR
wxWjnDaitOLF5VsTCYJFrLjeDYPvB2AyFYIVoMHRenkJNDT0Tb5OGd9JNg0dxuTL/iDlAnTL74TP
D79f5SKmTTvuuBY2GyHkzmgRH2atVjJXP5UATK3q1oO6YP91zjsSQBVSGFdlkxVyBqWN7q5yGscM
Q3RWtETTvW726ozs8hhskp2ZW7XOJvUf/j3BNaoGUPqTPG0weHb8RlqREAbu7v4441bBY63IHmHB
zjzszUmCPpdRTYX1mM+28iygeVXmoq/d160f7hdk4sK/tjUb33zS4l0zixxIVBd13sUW/rsVZRH5
EoG2haptrE5LD0T+221mpxoy9IVb9sK7XB9sj1bnX9xAobiqyEzK5nmpDoqUTe0Df2LVt6VeCReM
teD7/WmoZo+H/3HEQBD/L7s7lqY8IhOQLRXI+LaJRiWqJ/L9Iwj9cPSUUZm9o+T52UMDl3vX5MJi
NZBR+mQQ6adeLPJpJXZ19nJN96OvVL5qmtwZMxnc6Uek8ppn+Xwu2VGP9c0tDs1y93PQ/Up6URzO
2xPclhawwMiHCKXR+Fspk9phDJ/zAnOg5LfMM3OC2SgmZHvqBCBFHsthijgF7S2W+/fB2WnpJKKJ
zvprT2lpeyA3YgD4Rsan+fkB6tzH6fP2qGTF2J8++1LxvrrI2XPzYpjPtl0umyRDz7hcSg5NRVCq
B0DTtabNwHTo3bAU8d1zEEb9904w4GO7G1AX7CNy1gu2oMaxA/Q+g6jaP2r93uBUa8RS2ggyyggb
9HNW3ep+4N/AKHOSNgM/0rjZMzqsypAlrmoYyrZIGH0e+jlqDDW0RyhFMoqSUgCg1vGd8OTpdhnl
CpgZnoirXlby78oYS1saYdxpUVDi+oyxdsbUQKQK8y/8QDQMTzZ6bjCghDwE7AZKSNRBP6mD4h9U
ysxYAdgzrTF6XYFzhpNwsG/3uRl+X/scPYeDptaNbBRt9DGusrTjkTU+fd3WHyGbX3wLJaZdopzI
4UFFMBhY/p5hK4+lVWTrX+0YWUSYTj9tXyft023QnJBxdmiq+4DIEk1w0WVvKI/N6AAOuka2jZeo
hHz8cD8KZSfK4ZjVyZJoROgK/HyWphur6/RJT/u96QwWNT3kUsic68rqxY48t0jRwgkTP4TywxyN
IMTU+H01rI1PjhHoHR+riBy/1z8hpkhWThW40kZm+KOocliULpMQvWb9d+vGN3IAdqXqDMOyVutp
uljRjbTj5ekPNCJrd3aJPRcgF694upD0bKi6SD/6X/NIvC6m85yibojciOHGs9OKOJFR9/4SlCep
HDuZLlFWYmu2jdylmRqn+Hv/P/VznphBupzY78oj4CdS06Swam68a1Q/pL7Rvr7HliAHcZO9C8Pg
OOjjyPh6PWWC33TRwNm9UYtquc5PZnwuqrOSulDo7CcYgmm4yD9Zf0abTcyahUU2FE9a4Qddi4jE
4ztlnNsQCK2pxCd5zg1I0TmJnBbEYCnWx5Te0Uh2gvswK7X7HA4DAZOoU2fFjfpddW3FSY+JldRh
4UXMTnsu8J6QtYjp0iU92XyUAlBCTkVQGyo8ZbSk1Z9JT9u4aQdxD2vR3Xuvumrn3EmNjEVyZo7h
7nl/sLV6lXsBaiPwb3fj1/zY0n+BhAfe6I8fq2MjLRjBOjuFv0Hw9yIKV8TCC6EagLRJuqGZRQBp
DQxhnO3QsBSZybfop/T5ylC221N971OI3skyELUczt1tvzLHSyd/xrDrfaTMNAxPa+XvdKE9qJhr
1FwzTkXY/kvu3MadRf5YBYXah95Crf3qNjvpRO4VuNH/42mAzZekLmURr3pTGiGGLYfoN1NeveHW
mRQ48yUHf4+PjhM0OQsidBc8XsfQGeSA4k/9K5zh+N/O2/zksilCZQ49Y/PvUzAt4WwSPW9h7EYK
vwM0fDXzuickLukCh/eI/EqfmEvavukzOgzQDteCSiIFHfAp+ew2mzKUa0zMv9B1Wk9RZWtKKsDz
ixKfmc3uxYdR8uKEg3DUPVP/L6fkTYip3rgafKK4XYkpQQEJGBqhwhwwiMmTh58LxAQ+iU+z2VN8
Py07j+5OVKD95jovSvX3WqrGtSvdLGsfZ3G99eEstGAngppJodFa9fczoWqMBIYnibvmsdmWqI6n
OYP3ZVSpXLqi1rNius5QrYwttLJkhAi4XUQ3ybLxituHSAb/CwxZ8hbOT8WxxwGK4A5hqWGoL9DQ
6BdhNuxVaNpaXf25qzfQ7EjjpZc/uzPTE3+rdgzqoNiaLoiyO+9zdXOqOs/kX0wcJckXUGi9Uc+P
ekY6fC/x5pcXKPFeAAEulimgH97vFt+Cls5yu5UGb7IwhbI9mMYctjyoJ4nGDycuBX7tS23QgfqF
SzUSD3fvknwNdnTT6KpJy1KdZJiNN8Wv4ypEE2x9xjVecJnH1/nFyMGy15GBg8aFcPP8FXj1Hi3r
zI3yD7B2yKMc0yZ/OMEQIZDMXZ8bdou+1yOZ594zJ9lwT6nDb5R4egty2PlQtI3lraR9PfokBfbZ
kq0zwGU3fQyLdiXkEMCBbMOl9ZW/FL0qXY+M2nOBL87zsmrVGGMwN06RDI6D0VZpj+8MqVmPx4XN
yo9IYZ+aa7+ZUdfWELqz4+io5ddoi+1+1OBSAv0ayptyXXwbVsfFL+8APsvIfIOtUILMyQqcdJ9Z
AWz7Shhf8Vr20wdPqzv24/PRcYU73CJEMKe3eHzIYRnBZz68hvUTpypEm+YnMATMhneFRbeLOs71
lECoaeyPVCzwzO5qFT9AMfl0GLmFiv4M2eWHffnphC5z2xSgtP6btvyQOw5bu8ZRCAvD5IHrzoq0
s0npCcbpwo7b3hTFmW60H51MxvzQFagM4XVx/Mvieue7qMiNI2z72bVNaOFszk0ts5OTflVrNLVx
PktrLSkX1ZSwe/LgwNPvQSy2ivyqmG7YBqUDvwvIFnEmHAyMsErobLx8K5waYXL/HMunTwwcwEaS
IqiFYa3jntwgLPmTLZ9wQtcx6gG6G4UvUK6w3YYTeaWOgUUsIokko+5402Gb/lVCptGrhqVx4RUs
ML9tgVmwwEfiYTnflBgAB6yKuSBdLc1NiBXZsJjdwClZ3ipdxZyOmviLFdvZp5Abni+9HRsH27vl
4Eu673wsO5CtQLZEAq0m+tlyqtxfp/m9xUQ2F0bV+RuhxNL7FxqvOR5T4vGVnIQKrx+1u7BqCXx3
nwyUSE0sBKchv9AAFdQp52qstqXuibyk2yqt9ZmmOfEZjdPb5qvkIjsA7FMD+A5m2pWH3/daQgTr
B62U3TZavmh93ckq1b4Xe8HPZwjxyOQYyXQP6iCAyDkmMvjoe/+1AqmzNy3XamBPGkb4ex7e6J2m
juSkEKpL0lPFnK1LFTNoXMzaDfV90wuRF6MPRlOOXDVmWcHbLG2cX+5ay+5pLGjv/fNdMVYMbY78
5WEidoDH1hX80hrqcGf4Ty3Z4ZOhGbhZ5qNgJxh10EC41UvB2g9yKSKfkylrWTe23sjrA2A2nFuu
8QfZxhsuP1OVjOS77u+NROhfZVvZrwruWQVML00lyHMiLNpAMhDTnuiRllOKjstdCDA/MQbfACr0
GQQuQeHb88VfRViSAFOi8sNeYzdNTDAJlv9HcKhhA0NG9OHiOBDPNw/8UP1QUcNx60pMyMyht6ns
LqwD++USRQ/1TFVQxEm8kSktQzRu4jNceK+TcKKlgtGGF9HFhWGxj5XxtWNyNKfhiIEtq9zU0XPL
pr5FLG9NXd7gKB9GHMZVT/3/35DuH7reYm3C+Hd+VtIzNfG5qh6zC2M1YruRLeacBez1mBfgJHWd
8VmotN0UKlO3ssBNSzMv0kE4z3vb5bWoNvYIdYoqBO+5eNwom0ZpXMGUppa2p0/HFNcomLGfKCFN
94bFkyGMfMtejFt3zRMVzxN06W73LTtDKkdjQ9uP962+rAhwkd5ijg8XI/UCChI7ul09hoz5yca8
DmptChQOTwe+M7QXZIlITQBQMLm3KYf+AdLFMCkXnoOQ0+QK1yDAZxBKLlF+TlS8p+nwNGjPOUbk
p8pZbxID2JAsk+4AXlvtoU22rvmudpWIOXzzABI+E2r+TjRJemNaRbZIgfcNDF52f7vQ82+9jHKM
w0mzFmgxfR4m4QwVQAocmuq2W8I28mbZc/cQdnxW567gR4QfqSJ55T/e2voHmST7JKK+GJdyOxzK
S1OsTRA2HrkHcKc1yuRukdsfEZWLINyYtBKIVb9LA+IiJDYxbmcYe+VPW3VOg87EwUXVcybFx75O
BsR3r/TViju8IhybUl5hKajU0dP8BMQVbaU4sWcXFXGzbXqBkWHgwK//O8FytUBTYuajL/wQ2pDy
EUfOSYDRut1UyZmbzmpyNCmq/FTbyUrF1UP99ts+EWQ3Bu8OG90ub9VcJQuiCWT6uzBIj533CH4m
45I+f9D3qhsyXbKVMZo0kVH2tXmbocXlW97fjVZ2G+dnzEw1cS2qe00Z5ko19+X0KqHI1ZiAy5dH
uzI0YMwNdgRLJilZNZsdTJ2DPX3qykMXIgAV3W6wql45qprfjB9Ykvy6e6g1xGT/G74vSJ7qzzCf
VmeQnSmnecDH3OKMj4X8b6iG1AeDvVjivOapMlX8grldD/6cX4/uJ2qyAYo/xH7nOOl9J99SVhT9
32exI5Yllnu1FsdENyIbRwUS4iaUEVaYc2iZspQ/hN7oLLFar6Pewe64qADEMdfRt9IumCT+DGSn
uunEZcSxXCZ8iXcO29LBGrrX3RJGdbzW+iIXapFZ2cLS99GmG1MrlWYRtCmC5l596ZruLrLbw9kE
+WO/2WAPPMmso4TjmiasAR4BFDUYpGMRD0jZye4aJdbPKECRsEAgtRgsLhzMs19fdjX3lY3S/FYJ
tifKgUZwV5UV6e517QoqbVV/GUe+wC0a0q39smFPbRa8JFoBsL5PQqfU/gf38D1kuZ2Bt7kdFYum
wcPHqJHIBzmDmjD5kC/mnTdJcR6nXGs4uVnItwfwUz6BctRIGSIY6nNx0j9W7QCKBZbL/srQXQAK
hu1Kd2qaYmtU7JfbufGSR+iDOVQvr/gd6m3f2i5jBHrGfiHZHXtlee3cGLALZHF2GYYP+varcbw/
rbJWNjxIjYCMkxt1ceZhd6sGU2p2TI58WmTS0PA3ka1spCv16Yra6jGPIF2TOVk7/Dynm9hDkwZh
4EebNc7IiZ1euUz7gjJkQMwT+w7Sd+lXowXCEXtPBlHbgjjrLizUj31iCKpoACpzEgVwqGt2KpU1
Xub32kYYjs2uw4TPTWKfnMb3sgpw7MfCl6vDXkAjsysM6osQutmy/7+ogE7zaXW+IPJSC3G6eOah
g0IZomHOo6ZQJyRNYQw2ywCmf54kUc/RNYBx7Hf3fk4JF4zFohr7iKKF1GztTi3Qr5BJ8+mf7P/M
moec0yO8AXml1h+zVVRrRIMEifTwD2AAlTG66gu1sFWlFbH320fZOFeArGV9wXQwc+p1wQ9OyolQ
GLs1c/sf+HcbSQH/3JoJ8UIcsc1kuZuqYpeFi2i6AAXTKJIAUXHzwpxcTf4mSxH/SNDb4QoUyHlP
FXOng97yT7jbZs+oelTaQM2abYQU/Z+YQO3F5lVglF4Qdenon0+f/gwc5lncXhHertB2806sbpNg
tvEWNkkY3945oOnTQJbm3MtkpYdWjQyxHVX/BNkSBmPUisLRCX+IIj4TYY/6QwPCymvBteCfVAMH
/3xSgfLvNUIMUyH0gJZqodq/XBKg7MEzYoYDLhwFBFzlV96+4M634VtMSfQ7ncTfvFC8GO/YGKrX
csEb6Zye69r57Tlg8OYLg+9Sf4cQ3JfIdCEGY0hNSUi8/m2OQ3zNUg5cVoAXJDXQlNUzVICipumG
4FLHGHBZ4XM6OH5o6s31fVtIaxPF9wT2yl+iY6V6h1rgvsVhDYPSReTS5Ey2MH9Tf4ecbjH3RMZB
KkE1xG4laRNPMR4KJ1dSRlt8Cj5tTQ7MwKjBzZGBl78itDVXoFWUSG50V0/8PnQU4OQUxbH2LSj6
YBK6lXFJUxejXHhqxLriLyCC+FpH3F99HJXYZZGSAaYliUDMyQWVqzYkJsPMRUgZFDNmoOk/M23X
h3hNXYDutDWgkiMpUuDuS4x99Wvizj4qE7KYKs6s9MwRpI9t/+h9khpZHGoNraVD0zMc3x6bR5+N
4itAbcLXUCekLmqfD/FrR0TjcV8QGFh9hluLAjJECw6+J06dD6iFIImR4w2xhyHzWEHDKmUbPVqY
9HcqmawmWJJJwz4XbdfW78zf9kusJh5hxiK0+pksdEOBXeOEKoA42AlSxnSrogBlEPJg4jjHL1PQ
CwneS8KtROpRDN+xsCysF64edHEvuKzq0JVHBacHFT5Dgv8mE9ZdsVUB0SY46X0+fc6ojqXyym+S
0oVzC81vxzjA+V6Fo93SRP+a4FwLpJIgvXuVMugXaHjNjJSmpSeB5TH6bZL8o7P/ExxvACkPsSW5
JklQJNVfsZCZodYA6nz/GTbp+muh/X6GgrjDLBDkbZxmSoytOe78xOzjBZk1t4F8SmgK7hBIFVYV
axdx/oeumqBOXQQaFFlVUrABDeqwyvx2kBDbKAOYHQ3p6sTJhMMp2uMDzK/2fWxmwAfGKlvGf/C7
W/LQrh+kmY7vTvJT3BPmOL9muz199vQRMy6AXlmn0Zf9QVQ9s1LbmCb+OCEtrz7z02sUbCMMNq3O
exDjAtRZstRelpF3EWCx+wPe5JedXyP3vsBjMKr+T673MQVPx3dkUvCSdJCK5/vA4UfqrvZibVk2
nA0owuK3YrVzvM3jsws14q5Si9VIslH5mBYG131uzRMxM5vJskiDQhYDalDMtdxDGXewFo7PrFaB
BGG89uFQx4Lyzb8H4UU804gOsbJoYmmt9Yf8Jqp9fHU4fsdhV/q4UdQkCjtK7wTINS06iUGw3SJL
xc/gctkmAl0neBIAmcDp5tNwInw53mTbDopRsOW0kpQ/Z6hCdYdrI2D0Co8TYFyY6GJiVaqZ7zuV
zGOEUNLRsIyP71lNtud1p6Ic267kaHTVUbWC5B638XcI6tyW1/I2nVel4FJ3bcdVQEEV8YHvkbjm
FDqzDeGGIeYlc17SGIuYyJh/X2mF0Ay5I3IDt3OEr6m3YRMUu5kJz8mTix0PvHIgzq1NdUEXFOJf
gRrMcJ4KOYR8r+SMlxTsbodvKyv7FwZD/qeuf+lDYF4dCQ3w656Cb27MSpWFWdNk5zEuKxxg7c2i
K1MRrDFooC0P3Z43GtzB8GuYZWk0b9dXJsg6BWnIa7XRQiRSeUHnCSvWmF4xCMW71NdLPZlsgu4B
4l5qZAmHSkK1tbl6MF2KQqh0yPPa9mexcPbnDJeuSVpNcoDHV0p4/Phpo3gYybAC7p3KVhs8kyRQ
n/NFydH4Ehrf+HlsLPuk30paj4J4AMKewe5qlGHQMk6FEUw5HugsuBFMDYWXw6Wxtt0ID5liIIcG
SXgQAtlDlhrVHhSm1zCKreiyNBdvZIfBcA4hNst+COEbxv9DgRydDe0a5g4hKpGaqBei8mtoGtr9
VYTFvRMM8xwz182nyh44DUmfJZY10K0F24ftkPdne2ZTHhky8JOgP7k6EFEEvFRxhiKdUxk3mRY/
oPH4Uf1cNGREZ56x5HCkK8HHjXpoNcBboieJQT3XnYi3laht+c5I8Vs3dJWSyQPhLOyqcH6D7rOi
6Uh6A11nkFbstrdXnVhpYnz1yaRsXRd5i7Wud1el0ZjXNMWAd7fIuJx6+AnADxzzIw2N12W3C30c
pJ1JXf0KeJALQ5D/k3pY7AmhCL0hPiD7fUiuRS2qScfLat9/N02N68NA7teefJehU44FRjTsoKsm
Z58VDtwhCvPLMW6kzPo6U6DLrNTkVSmHTG9FJj8P/JP4WcrBAicfKJ742I92jbGT68rsOkaFX1Kx
oMMYjxo7vG2k8hNk+sZ4Ju60tYGVvJHmNR89CmwT6B/OHS0nlUb0rBSq5fgx5QSQouQkAam3cdOg
t+x85Olm7HFNzIoQnkgBy+ortNqRwDAPzb4e4JYtIKiFVLHrDLa4+RejOj73+GAevWBP9NJXTCII
gEne2CA8Xi3QFsorzwKkS9+VISPtEgBlttzXJleKu4Jw7gaUldX5XnBOEac5mlwtpP4e/8qnPvS2
C+D2q3/0MNLynxNSaVi9utdyzmq4VVJHVoMV5FpSUBBFzLRqYbkphwV/F083qJiwBr+OHGJrLrJ8
dYxPcGxq5seLZTJdWLtRtXn8z4p61hKcFr7PGCGnOz8jz7R7tk7gutDA3uXYNwEq9oC7mOi9DGIC
W0aSENzJWgZigCjAPAwdx3OyuAq4tspf0QcZJYEU7lTIEn/uEIfUgW1BsmxIwBXPUVMu5HMaaB0l
rLapJO4JOzOxYSlKN7LT+1dtT1B6sRMWvRGrKmpF49T7WApwFUx86dyjpW2IVzbU5+RYbVmSp6Ga
MbVk/Hf9tcM18atpbzPiwrsBLg++kUXqGG1TXgZ2lSBubb9XxdtmZndorY2cwkJaDOJVSngyee+J
ROYIuV+hQrst+QZRqPfZRdp3E9/9a16zxwET87hVNaPCebQ/oA6zeSBeMybtt/wEAHB9liKRirpX
vdrD6PChV6wDf5Bj43Jkyve92uNOJxK8Ypb4pcfgANiAT169pDjoeS2acaL4BMfKuyY/K1LW/7wy
lanc5mFgqvPILumQbAvHvM2tuAWMCYmU9UNrbzHAsxRDQTY73v9PEHkBKecsSRoRxrC5RaV7mYyE
Y9PBFHuTRjClpO1JQjyUedR1hutHJYmWPrshgps8uFPhiCNHUAd5YDaPkWUDCUSvUEpoYa+6+Uz9
P5Mb4N9KAj00gRmPDNe/htBY0iXQqHGxm6XvddARCeohDzAZjxgQuO0V1Rr5JN09/9Ki1IO7nCjz
m+Xm0aUUME7E+7SXHckAVeycnlLJnSwe7tfkaQNXhYjba+TqYCpjJimdBa2JuYYPzcpotNg6wVso
EDpdk1n+tdmc2BF5SkvGC5wrVd5FoH1s6NgtX/CzoUpVliyC1mwgAeyyLUVbs6LSjqC96wngYtn0
I/GAmN4uAe+oIlMNCISiyYCdsB3nwdmQt5TX6+RKJnySZewqBIb0sfmWnF/0hRsUNEk12OY7A0S/
Lc6k1O4OmR5QgkwS/NpZzfl8uX3cL2IlGfSke3Hobsb57We4QyZAqRGxxUPjyw8noocYJxbCKYXP
bITwwYeTzaE8+cCqKOTduPtWWAqhTT9rvgkautkhn5JtJznVH/q6DEpabItYFhcl10gEQqKun3eR
XibMjWivoKrHaATtofD/snvCwkpTMoar2IgIiDzIQKGEwaRFlQjUT9mYs9JKB4yThtKTmCsu1fCv
5eIHJLCgztzM64gxoMY1epLAghNV5M+fd0oULsPGXkr6h9yS/8CkygeDLEdEbGVmkJz3yG6MdLog
+Xe2i9dLm5Hs2a/HB5rP9WPH7a/s5BSi8Hxdb8sCRPE3Idnmhj+lCQmtKPddXtmM5ib4zAFSExi5
3IPYl6wsM8VaepDOEc17yhd2jMPZ8wcPcRI4cxB24wFbBqwMvYD1Kdko38sACIIT3GShpLVYotGJ
8BGuLbWaFCjYJXrp/GrzzUSHpP4jieYaf/ie9qKicAbBjYLd2/aoi9bL0h/lrLS2SsMGWKeuYQFF
HrgpjIsTIJ/Da6KvaOQnFqFzBiOs0cv92klX0+Qu85ZQeTLee/EQa1cAbRJxr9ALvgK7wtfo3xqb
ZcafxKtI6eGg9bzwEP7MFlbqoxYOzqUEEVsjHO9b9RrsPhizXXf4cHbuehe0Ch4FgeY02mflA31J
DzfMy/9zLqn3x+gF162qS1V/yk+sdqEdiAjNe6B3ExiiYycsJEck2oWwQ5k04GKMFiWMta2PCmZ4
+ThGjK3g7yCfL499FUTC7NLDQEvP9Wm3TXzZo44cQQ0WtcZQhYx/w+qtkNsnTZ5gaK5JgFBKavpO
DyAmG/EiFF40+7s0L+uFcJlaMrd8QAGo4PAaB9RM85WY2cfNtBW34ETcsTPyF6puhsewJICSCjmx
Xwu5dfjYkh3hWo5eFF6cx2yrbggiYSbOU6MFvHGF7SwhfLuwdqxmcsY/2MUQ2J5hCAbpuP8wjr9j
zUaE/P2l+srV812P5T2tzhWgnXP33mu0onhOOID92fZsfUFh4O2rJe8LF7jfPdT2lTeWFMLEySbz
AsGOghA/Hp95683th1sPlkSvkiB397E609pKSnYu9YsJ5xveVtpP8Cu44o2g0mgZHWrpF84sedTf
xbeRnRziJsuS8KezUddBGHNSFyjYWdEz2VsTa19uV36CJg29bJNKZ6/A54LAvOtuTp4udZ1aAHzm
LwtP1coc5HwqIYEaYssR2rk9qVcpIpzYeqL7Vr98+N6SH5wg4nW+D9OqDcK3Bz6gnYOVWZR3aI/u
s8YNBlAEuCmFVLw7MaX6RorT7GFBBe8h486n6BIvlBeFxEltRTYutEhZ0bFj56DvBsaFlhtjiK3Q
e1a75flRk3mGVwO2j6H4qboAc85xG2VMzpw+AO3k41QR6+kYy8fE9xHCmfHWcs1HPAUclLFtG5u3
2JceCFfKcKZbZCkiQSa5fruOT8//yGppQ+90238OdumllOUwj8uy7yxfh9vfj0o1ODDRGUw2BScv
qgRuzno23e4cQhbKcosYOZQxWYbt8I27lZMdFYUiKQ1EEtVzVH0QzWUW3TqnqOfXZ9WSMrgI1pdT
R5h7XHIaB9jc7iu8E42BmfphHQK0FnZ5WZxtYlB8KdNqfo9qMbpwan1wsnHdnRDEKs7if+2Ho4oc
J9V4HOO44kaHhaBcc4Hu96Ri00vZk0+pLxzgumHd+jY9Fgdfv063XBACDT5ajfHVc0U6r1LDq2os
oAVB5K/AvjjPUt79xeNgb1UIDI7SS2loOS1SYtj3PsgUjZNHV8ESjSz+whmvA8oXKHDkbAXVaSKr
ACNVtMwOQejbicg1XDqJbwg19vFk5R/C/e8gpTMbRWBqhqPhQwlLLQfh4GqPY7RgSi4Os6zMe+LL
PbHIcCnMDf1cqsOYyJghnULB2N+ph2wokHolBP8ogdPSf/oxuZV3ZKZm0ZVAparakg1+CO11b16+
5jKMUmdl1zL6P4+jlr2xa6ZdXou5gOYuTKGjuN25Gp3k1E3K38GaT+UADOdIsSzSGmR+ddl+3pKB
6jvBJeo2rEewOrsqdabydTtEb5LGCkeCol6M4LJnp0dJTRUhAXNGD7Cx3oBtMP0PzqT5DwzH+CRL
BSi8uFWd0IZyxjMqhWq3XRxYgiO0Lvx2XCVVMl9RIJToeHlu7+aHT3HM6DpTOcJVO0Xms4or0Fl+
GcRFDEQDzQzP3lQKRE3ox/2CFW/nzPWLo3HBX+FZtETGL/1BycGfbgfLEpa70pACcsfJhEjWhhRP
Sz3WuiZNqOFlg/8LSUNR50wTOTJxw56mpFmxGTjEeZNjuqJzPOvweDJDlRWLwGcyr+k6d5o5ljik
TNcvu5uehbtfHQ6Bu/fxDI16BIItQmT1TEwEbatrqyxo1+J/i0Sj6sjOEb4QW9z3/mihA1vljuKx
PlQAQGXjfopW9JEWwrZTTfkeXT5dRWVbXA5+fYN3Kd1ArerBVZUNTnmnx+ADVXd1ZlfeJ4umIffE
zs8Uir0kT1I3NatkH8mUmiAdknULmkS7nIoptKsVCVxR3mM+7sID09cnzYGmrmu3DZAH1wuxSrll
UPbdMCsVxzKLan+claXBIpIbuamH1uTesDdrOZkkhTWGaLBRZwlJE8/lem7AWg74nOggQrOLGgW/
iqmNmkkM6u/ScfQ+V3CYZR9mRRnSJ8qbbWtFoE8/4GF6LViImtYyByTOF297qqo+C2OGUgSUMkm0
Su+QrkdVCjMeHhVz9WcKlx93pVb65c2COKR2VkBzNz7ZdwsJ/pXsHGkdiUBstNZ9vz04GEDcsQLm
U7DmzbAl22g3rPf7kQ1vWtdP4f+qeZL62cF8mlXe8NrOVjRWLTh3H6Lant+Aq/w4aowOl54nJqI2
Fcfzdn9S4VWJ0Jm0KXL5Adg1iMS2fyOAJZc4K/cpluiJyy/sBnHUrXNFW6Cunz+sA7U5l5aVxH00
6V69KZJQZAXkFzU+k4qeZSCVYuCaE9hSiSHHNQ6ku93d1zYVjS5rMLv3gnwmpkc51FUa9dp2VKCf
c8THIhokhtbceQCQTC4QDnCCWmQhJu6CmnO4Usgttp9hpXMjLrf/ni3XOybKkrNDseLBprWlUzPl
RJDP5Oc/F16rSSuGexrsN87uNUD+q2AcTxZpOL1tvDNYn1jpKn8zuTpQNTf4xKmocYsCZhd8ygNQ
99fbVT+YH+mlS0i1/zxJn96FB3S4c2JQRWWOKDvAkV2HNndbAp5TMdTaVYWdU6veSZSgVm61QJqX
3FsLna/EdPydwy+aUDrqTbIcJqVDRw7rKLmdGDBxzNZfgFL3500ypOiBOa8NQszRlOr1+qlpT9co
umE6RJoAmm3DCRlddY9V/8p6njGQZqhtiu68pKWgcAaZ6xFwQ+Z5S39FQqINtCGhgEHXaEQpbRwz
49T9DYCMhRL2uoV6U2TSe6YiluAE0DWupDW5HeQBWzSd9go5y263TmA3duilBsiRh99ALXo1StvZ
kFzLwirdT9dfbwf5VGfuezK/ytRFb5zw84nBzUYKi+1aQhl1J+PvQ8AUAJ02bwOgxglhimNSG+4d
dvTDpz+niuSYxZePbL/ZaEZBluoBrPnV/2zRpYC786+k6lFnEopT2F3qHeGXXAZWEOwWxc3eD3Hs
tD+GlxYZI2gy35BkQJbWL+hRcW8zK5ygcOqChC7fqIZT8F3iA7v+XX1VE0FVjlUkiyYtrIfAT4At
qs+PjzQABDVvMknCuqKR+PdGsJL2hDs/4qlXdSZN8qMdfFFrc0EvdW04tAG9WMhCBGjWRQo49DHK
Mmn2qD/5TAH777gmTnOzYsWYZRQZgPbqgLnbUtaQpI5pt2BnVh9xyqOV/f7vP+hwHC12TR+wxFdA
P8ED7dKL8nCTn4K24pgbeFd+7E4oVC05quCPIhJ3APAixOvzp4bX6T0lKqV9aBsQR3nS5yDnRFKq
D3TKCZLwwvUVSW7haQ+DxLC75AfyUSeSsN39upunigV/QOWtzZz/LR2V4QiGtLIVxn87X6MuTAtm
QFzOUtIMR+IXdTKm6WalCX97XeuyYC/ViZTl7z/WPkpH6Wqzz/cjc3qlzyCWoiUFKDAb4yI412Vr
qmN/Rzk/7j4PbdE/nl0/TgzSRQMI916xmNqB48db/kjt2XdHzo/lNNb/l0jg4GvZXIvmohQ9j0c9
jOoK6oumuuvwCVsQsTQIyOMzGC3T7VuUnGW2IC216Rxz+QOiUqpoJI3ka43sXJINgUsy5PBqI6KV
+uDhE/CwX7Pm0uNL7Xy5ozIQqrvH/1dj5KWmdgUPtdJyD9sRPfayb0OLa7SmJe4XqpeuFkKw+MHY
7syqk/HZeWf57NeDLst7f8PGHUxlEFEn0JhxYoDie3fZV5Zv2T2Yiiwe2KqPxm69FBmimi34xxH+
sBjDAiewRWCJtHn9ZHkb/hYQFS0rzyarxWh1rJSCfYx+BdygP8xUQn4M6fp8mfiRBClyXVNiwuFY
wZ7XgARyxZyheYdbCBuYCfbP1Sp59mJtOpakWsbc9hy1XQjvlDZdyZtHDVEf7K7wQnsnloexc62Q
FVAnp55QG20hWBLSM29jq9HM50L7krJchmV+14jEsPmlFYgdrOKbx07OPh9gNLPpqnfw3Lwm8Mqq
9bVT25U88PetJgA+Tt83Uyjc/pPu8/FzhovUBIQ6zvEpv5dTUDjz7j9ib05mt7O8UdtJtp0KRbVo
vA+iykuwcQEgcbPPYPKTEcwzvq0NgwI4hJ23xxRcfuQ1MNfUupSuBZ5uaZWi3Gjz/Ceck8ZEFrZc
gTjTOCu7UQrHiS0B0h/D0XNvUHAXIslOHcOz/A9sK62Sw2pFOUK+shspXQgwvCw3fg/KFn1HnDZV
r8zCr2uHNrA7woUkS8RQ5W6DUPiF5gnK73faIFgYQDVZua6l3MJtmO4EcHImHW/mbGCofOWojEhb
spJSjSxH2fUOA2W3Ks8m0fqpSBybexhcfCUmh29g6FPAmU4+Pe0u6dREicU1mXHBcM5ssU0cO+ZV
sLbgEv2QZ8Z7mrtH7HqQ+7REn1qT2rZTdY5+03RSM06cbXW0ue7vpZT67tMtt4EHEDJiEC7A99C1
/hYzC8iGyBGETrGRdcgZGFZJiZ0BRCRxW4r+HZ8NnXX4JqQG5G0bRy/mMjhd/S5gnc+G11eSQOrI
97y/ipIaHOfXRWI0cV1SN2xrPf2HtaJ3nljE0hMqy6mJ5h/Xzwc7mnuudJwjE80+3vW9Pua6moap
okPA+GrWBD7zwJssmfFHoUZd3I9ZfgMmZHxRY92m00hCVTx3pRN23BKnZzQfkdIcbWubDDJ6OXRb
/U+uGq56wq4/KDbQubg7K91Znj2BzLTGJsFnsUxOiQ9X/aYd19Bfk1lu9JCHSiq+2vcgCf9ACPq7
GDpSpbZELbFFlO5mFE1O0FFDdNWW0sfdnMdHmYA5y7t6iPGXh2dJNcWSKB7/+0cetsqvByS1QBKz
hR3Dg+vhcv5ExVjc0sUB4JMsXXNBG5pUqKEu9weJknVjL0LMSIJc1A0iE9UhJoviLtFx8iBHSP8z
j3vBgUooYKDSNTwIHDFvejuV/fAkDcU8MFQ5psQ6fTy9vUUk/qCLejYs/MFc2Rw7le7YlZVFxRug
PXlJCzq4wfScwcRS/9ST5w7jj1Q78Uk/1j61yZ8OikXbKe1PcQmrXC70qzsy7HYbGT/MF792nQd0
qAFZnmeHah99inqpK4SxRsuQU3rTPy2gbbNLv4kqVuDY36TIBKfii8LDV+Quqak/0lnYmHWF5inN
UO3faBB3+uzQ8kyKNyZQ1VbA6/badqlloIS5dgBU90BQ5+vmODIwSXIRQOJ5Y6PG9mlzq73gTbL/
kB0z5vTTYKWXuFomuVaTb6CldY4bKcv1+g/HtEEqDEQ5nXYq+YyhjG2YPl4hBnleC28wq2M648Xp
kIIGROA+artdTgx1NqqJ/NSw7/h5WbF2JRKSELDhThPq5mpl0C2wmYKSotDhSqDSuDdVoDezIBQx
5EzE/23cLgb2xDQ7+pk1bmJazjSeaXimEX+b/WYjKeF4yrI8dFY3M8G551xQOQ7IpPBTKcKwVbUO
bElJHTd2OfCRLnXXrtIAy5mOyBVtY4yJRwiYdRxNm9dp+Jjq/rgZaxYLeSDwu7R5w0JAPTHuXaIq
wBbzIJzpe5Vxl+Uo8q/EDHit8PPB8cYH/aVXK/GdvRSK0ZEeq/On7E+OOH6YgwitAYmr+LPITp8e
O9qlgInOxWBnoMn0nARFuCheWvoJNv8NWL836Ah0Iq8scm4l5EWiV+Xdsdht40i2ZO+rpP4tlmqH
BkmajlcUOWPvrHaLCY5NzipUzYtRtaVfrt2TDx2ong2DIIe0RAtL7RstM1/VfgAcG4lRVCGMYinD
vM7kqAax7iqc9tlCo80huBGCBGVZg5cCP89C/i2c3XvBv0NPDMstDzvB4mtP5NSx/n8XrQNxYWXb
8WTW3DOYjffjwtWyXLc0OzpuRhmzbNqMJGV64El32gO4Lld8hpq3UB/LY8lk+lFQEYG9ze6NIl5o
AHch7gYL7P02AM5929A2zD9NtztOQP5rnQJw1JsvWmUbGSOdKbreiA20VIdGbR4mDfNSlPsbOy7P
FOzz/25xD8RKHNaTpZZzVxiZmTvRU2wUxTVEeH0aS95HbPCEMnlQU/GH1uUxiHKRrYmT4pY4upH1
D3HBSHzJ8zKYjnSgakhcRr7cA6mRips3HZPIKDqs+9odF7dbjn2OfdqB4IGDlgJfnmZgWXluk5pE
+cAIehDsIvHw0Ik4u8m5qJFUnz4k7+e7HiOCk8fkSDJZw9Gp1VojE/nHRgbD4wLYZkTD15jRRESZ
BsTm+N3zEJwjI9M+2zCIjisdXOUPtxReB9U94sXQU3dElBnYphw1ucHmxRgfbrlZ1spLN2k+bFmU
vuHO7qOU55ybTOt6n6t034z8ChkD/Tdea9zpZtv/fI4H3P+1EJteLSmWajO2tgWZwEhEONukZqKz
8o9nVy4/ynL/CRhLTJqLmBztFKahkNddBOX16AULU/GbKcE9UH94T1hVDgwxZlwd9n10Ydb147su
osts6heoZII7Ulzs35ALLAWcuS77y8Ackcej1fS2MESL0IN5snurMkSDYdHL7YKVkj3ms9LH4mz9
cTTL+X9WtQS3jF9suqHKgz3dbuaW7Bim9YPNw3RzYrq/E0JQeVJRgUtF4XsItcNnpO/oEFiR+RBU
TE4TwYTg6y8XQ33dR5p+gdxVCk3H+McwhK3H0Lgoqv4FpgAdcEX1erPd/BuBLUp1kK9Rr03w+qj3
z27haY0zI6mmmxRIrSM9SLjrytKWJQKLnmfEOO95CXK248He9vkItimr4sJhkTFrsnS7fQ4iIKQs
PZ+psk7gaG5sD5IlA5Yxwh9rU3gJ5ys4tT6OG5r4rps3safAOwcXh5KvGlEnkTchPrn2VvMjciMv
YdWS383oqbzecC32kEeijG2qvqIcwwQopxfdxXCCqkqpVGDmeimZTUhoAUKtiigoZ9D9tXRl06sX
bijJK5kDofJDr9ta+cK6EWvqFEc0pYYj+/HGsNT+Vc6T/tGk/FE75qqhMTng32isnpVO0tZsspYn
4EFAOr7yoYWQ+pZcl0kmVVAPmt49LEKwVoG4OQOD7ZG5wOLORtWZp+BXrwFJS5ZBSaMBsPi2a/Gs
SXMwps8xdYb86fB22kTZvk/83ru55/H/ysHRuhuadOFz+wbcKiN/OgyT3ymVm8QQFIDb4/G5xEsM
So21dvkty/aPJ4/lVpFmTP4TedNIU7Hcfccfeosp+ABKJ7fenZVtZpjRVbIrjXiEepauBKpEiUbR
5HsDn02tOSTLmSKwc8x1zaYIb0XBNmigBqSfaIcPxuv0dOkw0D0qE8DkHx0BMmJZLQwWp1mlG6nA
x5dJO8xR9HxIdJ5asl8xi8bsDayvIX5qfH6Oowpzw4GkFBXKzYM0KO6I0PRLi5p+FLpt0YX0oRp+
Wow/VZvgF8DuBFA86PtlYA5xUz7VP+tpMpMHGATaxUye2ZRfJIaTat5A7T3ipypQ3o16DyArG7fu
bU8gy2PW9aHCcZhzcpWJf6PlWBkDor2Wb72RsG1pav74nTeYLzs7A0lEO10vI94Bkj/Tv5i7YwAd
i/FYYtgAFmebFBtPojfg+4OFuec7VhTDkb/QH6c0jiSKNErEShsk+DUcbDzY2K/pWZII9kjxIWj/
D5oLz7iTi93qaTdj25E0pnfPolBk7lsmkzEK3YoHXTpC5yDSb+6X7PyaWyL+Piy/g/zX8y4TxuG/
0G52OP4qy7ALH1FQAHOVN2mamaQI8EE2sUcF6V6fJ/9gT3Y9zVYFgww2h5/WRnDt5nKlPdXjeuJh
+FIWyLuAiacNg5oTzeSqOYPB7IU3tEyfOERtKKlC1xVblV3ffBbX1bTphnaumQ523gr6409KySp+
RWnS/jMePAso15PuinflEjJDhmmvURNH/X5IhxTBprkfiZU+b7odqhULzQdpVt1hg9xSxOhY6Jj2
/vPqcKkzfpj5wn/AqlxlgAkKM7/Ai0CrgcyRqVAiDiV7QB9R9hp9WzIKPQp4xHK3EGuMiOIG/+gk
8VBz8Wfg/8cXvcHDoduDzPA5B1SwvVVmIR0K+qQDv/WikSMeXnXoorEhVcEg7f4lvkBUByvdipj+
WQW49TFRi+E1kI6NszR/37Pe5Ut3H/dCK/1ugmfNOPD8860sRA484vSDNHLGGR07GbDKpBD4CFJI
Ioe/uBMDnt9Gdo063Qkj0SXy6kE3OiGNLFxQhBXeXsc4M5FX0HZkkTDYgODCaXBsi3krEVBKFmK2
a092mOt5A4eUxsvfHc3StHvRI+ZJ7uE0Y/undmPGoMSUgTamQXQRMbKW+x5CyrvBzTLrWH2X6Psz
piZ6UbJ2aXhezoY4Rbp2OglQYi8T44VS2cVyjL3AQUO18JywjeEyvZPj8/Huz2LVwUrafcI2Znff
YvYacOc14euZuzL1FtkZdC/L7pcazZ2FaOQIi5ueqow9p+lvg36PG+G0y7ACAhfuTmzitEcHL2Q+
r9S1KwFo0VXxB54Z2hGMxQVLSQtQsamMyxr9sNwA5NOeS5LDzQjkem0Vpa5aNJCwC7hNEoFu1XcY
FcjErhin0na+5PpMzXE57O/xBtEKcFW3VL5vBSE1/WvMXkYb2IpAcdiw+CMXsavMoJvyHbaBnOwZ
H59ly5V1cad+21HViv4NNfZuT94Tw9WoVwPPz3C/vbgR3lcrtNS07S8fvh1t9tLsYecrZ7fG/9Wj
/DVDqm/75U7OWGHOM4ftXVgW0BI6hrs7vMdYUZXK/ZYaoYCEqPmHAy/FpqU4a1rn6TX8IIqZ8WZ3
GlHuqf5hYlkKN+9La3Lr0wA75BHBw3Pd5/TKgly+Ntdndv5VEk1K2JJf4BpIr4E6L/1BBdYMI3B8
Mjar12FxSJzklBTYXUsdc3IJ/THp1uuRU0RYXInmkiXW6lrJteZaY9tSnQnyzsFDShdbz5RkVwuk
mkzzd0LtSpCsO1AzFnbkXplx7trnGwqv9pisINOsz5K2hNA/TQsglPRLsIICHLezpnipgKP9K8QW
aQWWAboEt3Mnpd6tm4qEqG7iN0YTkzVGOEVF0VF/X+todMGi4u2PNMtxNel2dHbiAZVIvLu+t7jH
AgYjvVWHPRf5kaDNofzn7/R5BitH2Te3nyrD6sjy2UA5sPc6r72uVhZSCnGHMGh4MxTIUaUbkF7+
VX1rk5+b+oozxbscQBy7cunlq08Kz6vo2mam+7tVEdjA4nzIOWZExADPlwN1E+oW9nJ7zFD/IetR
5wtTmrkyXhsspHnGOqHd4XnDu23xh48hPci+na9nyL9pKqnAJjq7V9E2FWZ+Qibo3w8o7v6Y0FGn
++hYWnL3GdByXY4UKjGJkx7gy4mXH7rAmIK8UBjVTiwGpSNrKosq9VYtwzHrb2ifCW5VEgGQLIgL
lHZEL7tqsYMEViFUGhNeTgum2u1ZMO7EjK2vWj5X/PcK2IpmQyuK/vXBQYtkickFsy5hg5YvrlHe
hXfYysO1KVdC4IAppBArg9q8XutMWRBruKR17sItd0pCCxrjzfIMQo8bR9P1JttL2ksyYz8kdyw1
n/D8y42JKjL5ujKcE6nD7B34X/7RFj1gJEoe+8o+pTj1yL8O69bQpgABH4SH81x6M4kFtl51Jb0P
FR/kGkKl51AZzaRtaDq0mStwo4IGTBotcITFc8n153TkxdQ2zElR6m+M3nVdA0F85KogGeG2UxIn
pSLcDAVspuuq7osHjtBLaCvIGldWdScJDYNwCE9qgeDN+L8vImMD226UBnPENzXmxhG7GZLZfzY1
iiTJkPBiZhjftNXWKWmPmUdh209YLB6LoaYmZakLwAFIYG4/gqZMAvVdgEA4g+Byx23VqoGBamBo
UhhLMjdyP1AyJQF0AqjsYPeIyjPCq8giMLpbMX3FZUuEVkna1DHAMVYQO0fAuLRNMQzpfaeCv+/z
7j45KRriqwJKm8lR6quGSxI/7I6MCOeGV1PpI+w3ujw5sz6/rsJkm+yjNwEwV9Ed3P/Xcyd72R4h
z6wf7RR/iJDRiUrT2PgRTWh7/0m9N5Dgq7y4EkqckqxZOXf3NJOo/2UWS9e+6vErsacDPETClcQ7
N12BHsek/VVweawQJawa3HpSYOdYznU0MLSWgb6Dvj6IfDjoGGhRUZGZvozGL+TtmZcr6NwTGhi2
9aVa92luPl6fmPsTvD6QWYWRRBMBAqktY5bE3CX55/b8CEtGDFBS/AYBBN5grCynxpCWnbYFRvGx
H/HSi1xtjAHUldzvdp11jmpu8izgh8guDEkxrWPF6El3OMSj6KOC/8dfuPtaSlGZILFlWgvcu0Sn
N8OH9f+Oeu6yxDJuSHxuB5enyS0B/9JU3tMWcM30YHYj8pBbucZYvkbgcPLB3GK3BK4NU0FazeKq
j6cdq+UHNOhUYh8E7Xp6ntUHL/7oBXmf2m/PlSqNnf7SyXcBcU3l/uA5eTakrRJnzstSQyFJb37D
h3RvqFjoVpcTH6nQAFI0ANA6MBr/VsP/f24r3k3ZLleE82i866vLmO/3x/DTTZHc5bDL/J3R5StV
LkCRRZL+6RlM5lK0ivfq7YfOKz1DIzjGJN2CDccmt/06mnH+NzPbkHyd62cyqBftvtbEhCUCrcql
H1bdvs1/kxzT4YisMkC5LRfN/kwHEmmxKOpwfRua4kbGUWLMEVrke2KYX4IdsvC+l8z17s30Z0oq
rAs7rRAIfdA+WUNZcLOPSGXi4ZfLYPj3WpvZ95efuDjoQfuSy476NJbBgOBMbxRbO/SSFaDV/rKp
b+3A5IAW9oAazv5dH3XXQSHjMAXRRRpS/kBfXphCSu7jrexoQk9LsiKRydTcduGhXINN3UZV14WN
L2EW83RXXKR23NrcR90vSSt6d3PxG3cptKfSm/8gbBIQD6P4Uwd+A2cWsR3ne/8TV3zOKnXj/SSJ
M0IVTGHXiPMjl5ZQLk8ee+lL9uNKbg6fZknJ4mIg5ehlCOseafFwb0qJSrKnjxlg2Zq3q6GnwhTu
/XNOZS9ydfNHf/R9l0CbaR9wh2RTBXgHKjMQquuk89tTMLLVB2rj3Mjxsu+TS6fMgy+HR1hgLEsk
nTxwfN3se+Zk8vi6rJAcvLrYwRNli6bahbz8O1/sSyC8XsVQe/qUMQ+yjN1H+qFRitAN8S1zG2rB
BntxU5gp3MpgJUurHGkXrr/KZc1RC0Ow6qsehPbMVMcVl+jUXCVIIFzWV3zacA0Ot0TZnMDTVmeO
/MVEa7krgFUyg8L6kha8ooLgVN1SwUYfNhT4Jbhp2J+QlxzXH3zVF7y6+t48BJhppLZKw60im02q
KqLLuheDCAJTX4dLUdYtFwv1IqoALwslk3Qw9/w3IKgf/ME3VUgY+rF5hFZkp8kfADA5c0g95JEN
EojOjChRJJcrTom5J2kZJSvNiRTFJTYnuCsdKN2y597Hp72FIw7J9x2eMIGxbMykcfVJsBtBXs/G
eDnWTsNLJAJbqDr60iOy6ZtOc3XfQKrgeRWuKz1At3i7/Fo9JIiA0yzBXw81wVmFMNJeKPvpPEFx
CSVye9Q4RQBh0cMMJFHtOi3RkRq1PXBjNEj8WC0CVpJwy3FNFVaKprli8++hZQNwbE54FGcmRS0u
eZQKFuyHCfQAU+9asngNn4UIRB/zqmU/HPLMEkXGkOTxUAOOjJfHoOFq9yfFS7q9g08nJ9pJILPb
sTEOkUkwJsdHKBGm4nUFVNpRiqfUsfnZSnNto5biudbtsAsuK/JYdgfO/D2rqBSsDDsUPZzSaxSB
VAn7X55Br4i58sbDBYY03KkaRtDCr+DUpt6hXCyJLQHFczjvoM2L/EvAtuRTbbebcKOSb+cxvV3N
xiweHoRAp5Xcgr6u19vUelaCYueDV7EBIv4F9AjCJQciPm38CWJUs/qhMuzIICPVFi3rTJmDztBv
Fjc6sxn4W6dQ/jfZeJ0UN3DR2U7RSV037nceFsg9fAy4/xYOR60lUK1AVqbOx3I6rmCW3cwMTC8u
4803UWvd5ZA+obxbDyJTPAWmDnH1HzHID2B/tEHpng+akWad9Y32J5Td68XURfdrUvREjQRQWxF9
Bw0nyBKkEDcZ1CHHdB2XkewGrgBZ4panFxFq3bcYW4jf5w9zV9oGAZwFnKUcvIR56HQ6f8XlswJj
ZDJNPfgfxEV4v73DVb03tTUqqXqbn0dHagJqi6iliC1RYO43C9myQVrC8uBYfwd2F8E31fINTdx+
CdtN6S88Jr1unlHnDYpjXeLF/Vmez0IjA+2iOBXrN8d48rrbeOSMI/SXzPQY0IWVJLdSWbj1s1R8
R2b0s/AXcx/DqYSfwTipP9GNhyJfDmEIlSPJZu+FtP/BCsxuQ4aNryA4TYxW4h7BP9usL5ed+7MM
2McrTtTDZFeZ0lvurym6k3xP3o/E/DyMGtCKZ6DXS5NVDHvEqbzB4PT05g8wFQ+ooY1D5EiqFHWB
S4jQhnvH0x6XaeecwRpfbU4Dabo4BxKB+dWaaGU1KhHgCwoNFaCAOJ71gM/ROFVmE2LjMfdj6/+O
UpY4q6EzwiFvg4I1wv1Np8y5OSnOdju4kkBo32s4e1+F9lDXUBXt09oz2naIreE9gZqZyvZCUSC+
o+xpdw2btabvim/HdqaQP8v8gxBiHWzTd+GIGHkJ4Tu2NOyYCw7Da1ZIfL+5zaMZi9y4iPsEaifK
qTQiv640PL1wnaEwxusJCJgKhH3pn1PQ7RqxRPHmp8kFapoqK56b5pt3M8OwMhFSAVL8uco+6wz9
30eyLhn5G1+zPWHqc09idbRJhnhoJXGl4fVY48ZvGCL6KaSa/gpoOl39Mj7ezr9xChF02+S7+rvV
CpC4M6dMOXx/BiojaM560eJ7snC27OrIXZrFE6AyyEeJ6lfMvDc2NuVfSQG32j+vlBPjs4jed92E
wR3LSxA3uRHT9OJHm2wJnmMQ/ueV6e+sdPjVt+QLyPhi9fPlK8HGm7r9vdChV6fYXRFWcTwxftmZ
bOoQAenxLevtS0Lg9qDS4g0fDXQ8+DYR6oBirSEblNoXtI64D0YW6aSM04RDG6MLTAnkj2fBA8Z6
0wUJQNFC2J+AzzNOjZnfBcEYMNhxNurGhPObpVixsQTTRBuzUerKju6PT+lYTbKzFS8xeLlxdO/v
EgR0Xs6jP8HqnRU5xef6R/ETUj3YBdyaOJgBIzYDd5R+4xwlYUniEOcWfm3bWgc8d6q3jQ0xgz66
ZMu1YKb0Au6CTcit/8FhQg5A2K6+daiiPa2cTkJhnjF+98H1xS4nh/gPQ2BKzWyjOOZPlBZHFH5L
LaJ/rRmtMH6lQsjXQ8yc9xzHEkV+a2IdIS8EHXBgz5jH7K9arIWDo6uYODfTAyZZNQTvDwmvYZxS
Rn97pQQaUE1UWYbsaIUEMSo1zDFbz8oGZoV8l852aN0SAM0PclrOrI97nrZ669ijafFcCSq6loff
DeWk14qIHn3wq1FPQQSlMaAuMvj8koK/98tlpAwzj0F/fOolT9VKzWfIVrXScbXLZ/7qUwDcm62J
dCbY6H9k7AWBWoTrATfeSCwhIbYO2UE+V98ZQGgUq1ueSFSdudIOnxGu4oqSRVkhMhLScSjkxVCY
EfKw/VyW74S0NL2MlqEI1up8WNAkrNUfC4Gm9zd2gPsudp+9no1E9B7zbjXxoBDFl121qUwtGGkF
N8//HlSvaFRDzeAIeweZGatNRvs0cPpBIBLuD3GAax267vS3jL7ILpY1iUJOTZ1DyzL0yfaU6b51
JjZKHldrUvtPMoyqAn3tgwHFjQ7jt2bPso3SlDX+1StXM5AdiHuqw1UR10bLDSdpBYjXN37+GfqP
g27OU4PI8btSLqytAckJD4kkBZwsWvJEEmwODrgl2FD0RhBNftcycT28ELTGm3xBhpoCL4Q+oaef
ifnhiPpCqZIUhe4xi27J+Bjf4hhPQhcIOD7x8ur6yuSO9nOC+CRUjvPeEBE0+sGAIkmmAel/6sMF
scpzJ0iOkIVziMvChT1eqzCGC2O4LrIxbD7D8vX/gCQIGK4sXfJaH2YZ4qGLroCFL2H917Eu+HBw
nxCaJZALAWsWhgJV8w+kbxpPAFFnA5uXf6K70Hhixqs8NsqqhYYITrWwYnsLAFWr//LNkdMiw4H/
dyat8AeI+PL84VaqXq//leBGFLndueOS80NdcHlHCouBWGtgCUjlQ8cYdhzO6NMjExZX/D8XtwVw
Ns4uhV2+Lw14p2nCjzExuLuw+Bv805vQHQIb/6qNcsx5LefePGloKepd55Km5YhZOxni1jFW4Fzu
OWPIHWNINdW+/A++x6sVjHXOarY6oQPAVG7r6J9JRXcf8IxdnRn0DS+8ea3x6W4b9ROrQEZXpY+i
RcCJxn5KM65bNYDOsTlMVUOgkaCF7PeH13+RN2bVz94dgC1r0QBxYn322TUlUS4R0n60W9fr4iCj
vNGW4jupb+HjZ7C2NRM8/fYIL4GBXIkd4EoEWnSBQTbLRG6OajIL5w+ySdPqJjAGQx02Qt5CL7GE
M7QdV8eEWLwR0stgoMsUhpo/2EmW8u1l4/HLgsvC+JTTcM8ruhXtYMf7MhtqE7JMw4/MVBrHBZLP
OslXqHMwvVgTAEM+QC2VY9c3BevwYSWfICxzJVmxSBW2Y1dOKmxTqA9sXuUK3Vt6WES0/yVehGje
5ZO6aCeLHK2KFdguy2FQYHcZAByp8GsFc08s19xDVTBC+kkRNzVGsZiSr0fxMO5ZBbPoWRmzafK+
ylGGXJfNi6rDFIqF2Vm7CC3ZfGNHE3cmCsaAyfHwNhvMhYb1Hz0ozcXrwFKOFGYfc7EE59rwwaPs
I/FPZGqFCNlzjPTjTAhvwtPmOSYO64DoPU+TJQ4OIygmtr2qDXriKC46HQ8oLebiv7hSrkqeucjP
fHLAq6YZnjSovNS8EUMLBje3R5Oncu8xuiZ5wRqRhlVsJKSr5GMnOJBgQbrPhLRELcZVbZ3XZHqj
nLanMQ1p4+kEVVqEOj6Js0oF4Himukrc5tKPKLiVQakvdnMKupMjCfWysuJN959gYMl/IYxXQ/3s
RW8P2wrdo2UnDxJ20s5L83cskfS7KJ3jCQsElVTobsSASCK+poho4CXLjYBN2xaZ/YkJqw3SbFgX
0AibViDkpnb5LNE5QDCrcuNNxqHvfURKZXeY0GmEI+NWhivBW2IRu/bY+dLRAtYA7/UP4Nxyc/D5
DC5DrEp4LhD0jpm+lSxI1msCaXZGGsN+wVbkXsoTqKRzQT9PuKDqZjnx3yutV/0RH9cLg/2LeLKE
GVsnjYFeEZVSoRJwt8Juxqz2Ga7VGBnE/yYaBcWeNpy4j6xrvTGC/lyrG4mTQPnKCD2lAy9D/Jc9
4u5n+bxww17IO2GmURqjUXGa+dOfDMPTicE+TzVZbRoULp4MdUJtgnwqMT2e/3NU6DfydLrImp4b
4/ygiAPfX0RJGnVSEoIauQX1wEOUnpKHfTZPd9L7vs7R3pPehpznPSWIldNJav8cP7BbnmwC3lMe
8nTxtIu0Muc8X9b/PXArCSYg3/Y9VeMVpbZObbJWycodI8OfzrzLC7gvMcOFBTczRwTIIPzoEJje
c5zjuPe0VyYW8KgGKsUiplmZlw/u+uywnqhWm33sRCYF+RdbwcxZldNZzcIjBw0UBCixquVuaRrP
kMGYs0CUgIuK378x2laQISOvBUS0Va1GafSBQndrFgmHUw4zED7x5wQ09uaETfUzv7OUgrTHYok1
fBWWGAt/WnZbgVP76TYRJdOSJCjO++CRDj2fHu3UpWpmy4a65aFyp8L/MsAiVM10ZJBsudxjUbVQ
7S/wxmmctnBaGEsviSlo1FxQxVgj8HZzxoyUm3hVcGsdfK2WGM/8fS7sVc4TZ/pHVvEp+73CWDsf
+UC5uGfD5KVARsULjUHuhwa/VLMC9fccVAwehYnWBwVHnSM/cqeQIH4acUP7TIxlbM736e84s4Js
k8nr4VaX8hjZwu84jlqb7eihEKC653Vhxcnldjo5Gag95uvO1B6t1Hqq9iEVucct60e+bBrm2cwg
piWD6u0uh1ufB238l5hlS92hq+OM3q/dUDY7pl+lE1ZZ5q5bqD6G2sOAv6n5Jc99FiYvS50/G7re
3idkN9PwsRNUrxtcara34qxovRwtAqKlJW42HXdDwUeUm6BP/cKf0QLdVp18F+yHHX8zr21eWvw2
PGoz/mB2lvkZbOlhR34F+ePh4b25D8JDzrjkYb3wEYTs+n+kF2uauxD9UyJ7/9ebv0r+C2GGf1Pu
K8IzT2nhX+jgwgLOpAh07LTB7aY5iyGMn3Zm8/fRFaQV+UykKXu18ONHabz71/wuVxInyFgCgyJ7
z8fMEnIiuicVtfZ828M8lgMoFCOjI1af6EJouqmXsW9RaG+W2rQEpw5amC0ROLCjX9phUQCGkDO+
6sPbL/i5dzE5tWo6Qoinc4qBW5NHOsH1G4pQUtTRBZKD6b2YLVE90ncEgwnqBfcDePVJBVzkzg9O
WEfnMmhoEZdAWECTy9IQ7BCEAHFJDh6XDmnxpCJvYRh35DG5Yr4X807Fk8PcM08Yz0BNsfLKlxue
onAbCSBbdvwo2uTo6eq1IaC8DI57DS2ZPfbM1+PoPucdEp2Llq1TBY09kF+jCcIJyWGsAGedCs1U
4BKno5+srzMjm9Tclh3Rnw/Jg4LhQv77Limz5B66xyyhaHwzQl3+mGGuPSkafnwrgheZpatUHBE5
J3B7tXM68253K6Mvwm2yBfMQOkhcrH40aDLCdivdzEITVPIPN/wexwSOfmwMV8qI+8v8BMpTW/dF
JNR240n/5OpKwcevq/2vhLTur49rPgwBCrZAialYI8f1R401w0T7j43AlOW0r0ldOLfqkxmelVq6
cV4blqDRFSZAHKsQ8k0POQw10lxf7gP3QCzKIl7CRofkRY9+8N/R96OGgNpj+biIZoeF5kwvIS98
SfR6mZ8NwHrGQhPD0yfyqvkyXAsnIH54d25NwsUcXEFF24iZshBpjFd6vgw4gILGvcbt9M9+/Ccb
YoC25EA8sqGYmH5oBKe+XPk6IXts+cyEN0ZlFT6tGzt+4mFKc0x88MfD8qmVRAUTDlmKWRjdbO1H
tze2/q2Cu9LIbxsoUDsCMWLXKM5MHeVhB3gR62ENyRW1ywaxYgCVeOf8BoVhEU82eEEAY5MEJ0Kl
BIKom7zdSFnaIDt6rUacBL8kzTnLO8P/4aDBM9TM4qoiiUBJajcp9LGxn93gvzrKJDTpN1GqHIcq
/orudqfqJq5XzPGzSj/W0vUiBunwOvCBGq293yAvfnD3fDwTTyVNmuzayKX33odhQk07Gf0/KuM8
aLQMQrl9+NdSRvnqykNNERdbjjH64xq12uulBRnQO7w03iPGbWgn7uxm0Fts6CbR9bugu9ZQyk14
BdXfjpaUD6QsALpsGjZlirWyGMPn4wQ51qJ5T5mOH6Ygcjzqz9ZuELuRT7mbccIsdQkrvaNh7CJg
AerGOn0ffVizuqcD+HE55WkR6Rl6Pfie/mDksKEsjT4XPniwPC/YrY26c1VfuIh6zH1bXd9guQJ4
U2Yk/tCQati4DSNysaMc1Mw5oENAsc8eyhWnNnLOuuzI6FcYFECOTR1AFuZai2O8d1ZzYxD0G8d+
EaVaBTzE2rofx++Qx3Gc1Ph0EqhOESUXgefBPg0VJdK6XNg46Gy48xbSwShCvFhrTglqF4dLyPCe
GU/KOot/p/9YTAD+zJWQeUWzAaq2G0SOmYaRzukfWk3WkEBNDfb8jtz5mHIM7QDHZpFL1SeIhY5H
m5cHiVA8REpYfiAo/STgsk3nXOf5oR/8wF7e/FH+UoI0DNY0mY84pgEfE9xrAJWNegASuuOxZTPS
Nc18IZYrYWc1RMn4bRYw47bThhUFIH1pQ+GDWlJKw+7sB4v4PUp6t59zqnN74G0ibJ23dP/GzmSX
Dh1CEJk0j44PW47imn/XY1RuBmjAMjfHPXMD/uu8Mytl9SfcTTV6QGG9YOJruLwkwNWowwI8sSzK
BccU8nRSr+Heye4OT7/xO7TD3EWILRI47tHieUhH6+wkCkiyDb90QxE5eGSmi8Vso9s2+oIW//yQ
GfzvwR0bPaKftYef6h02+XcDMj6XArdF4tjXW7Iseg+JlkoQ/WN87QiW+HkqEkUZHT6E2orGtQ9i
Cjkpr+7EpfHC9psTJY+seSlVHe1sxvUCSiUYxy06D2G/NcYUiM050JqCKG1OAfTD1FQgQAEA6qNM
T/cEgmpd8dN4auF5lT/QR/ew4YOtQRi3PXRl5iskU25mrfubeKd4k8t2ntrJ5Y4YR+0LJOAzc6qT
gPVAd+ImBarac+9PS+EKbdNQF++wpImWrZORZFj78Y3UGNxawpkvSOkojRlzqMvKC9KKie5/Bi5f
AVvjAnPCpiUnlsetsy1zWehySvsxcnlMFBPRywJImbJ6uhdzdhBVOLD3N6Zgt5XFOHtEONxMw4Rw
hM7uDQNrVQnB0i/cvwB++U4bAgKeCwZ1PRR4F0vhg2+dv6bIf+y4doUG5XE3DQYx5YowTBz4UnRe
91nNYusLTBsSoeLUEQQAA8uO+fl0+xCBlvZZWQEPe450NKpfLvJ16tasys2BP2JRa1P+yUu7IJO7
klkiPgCfgAx5+ovseu7lANzfBlfdNZxezCgoHzCf/OtGqw++AUqUL3C9/Ghlmo4cQ/+HdU6sqgYh
C3BQfhNlKjzqvZvd3vHL2rMhTS3Y4TjSLC44HdxRtQkAgiqfttqC1Ubx3g2hb8cOVd3mCWEKOa5q
YPURKmrJvvxso38JIftQsrl1+0xdti+Pwcozo5fsiTAmC+HK5poHOem1GFqvghc0vatNpze23vKE
lGQ9A60zbwh51uAiCVEdngES9bmk4iR3mtlz+ucpp2TXAG9zYy4nIjlc/i+t6nufgVAGO/QdBj9F
Mgsf/0Dhoxi0NWiGIO+BLP0jKthp80schHvT6xSgHRWkaAWwdmP0Hc14R50NkzzgWtGFhZCC/V1M
jY4xotQIGyoOw49RKU+dd9/fE5IeU99Ak9IruD3lFNJ71/vCel/RhcbZyKIZuIFioTvYtbqVytrw
KrFNJaUt1skPC82nohi0+KpoB10eBBA5D7VNqaP9UXUPuJFF48nk0W92c74Nz5Dc9mADre+jNk5F
yP6SAEEKduYmeWSGOdh435cs73NY5tPZnoq03qKDPsQyQmCYpdVjpX2Wz6cIo3yckE28FMJ/n59r
YMOiOwiRLLp0OTpcAM3cmHOQ1JtrLixGd4ZfHeGzF2V5dUW4GeHimhSRfK48saO4MdFBFVOfmUfS
Bm52Q6M6vVBVI1E27oE+xsmwrdjpQFwMbfWLoMguThk7qrkBBesSI2sSLyZfzTsL+8o/2xAiVnav
4B8IQ3SAS65uN7G/I0O3E9iRwFt1iSdvVIQktJdV1g8Rr64LVwhVHymBX6zGUMcFfbz2mcwdiM6n
Eq3PuJUBaKcndOlMcm16joADMVS8+Mk3/wvRWFo9oCNde7TnmY75s9kDdRMw1taGIfTYEARxozw6
vJVyEXW5iGrlJ9NXIf6oHN43dLlOmmXoqI+VPkSP//viDjWO1i8Wpm33GuKx4VgblQ0r815iZ4sp
/c5FAm3Ra3V/yJmpR+i+U8Q2WB7JMFuhVWIV8emT13y/lRh72pT14hoVlG0/POI2IVL2WatGfSIr
x+b6LKzF2UgJEzqdyn0TJeYt9m5dv+tHOZG+taenmz62EZ8qfR/SIJFiPqPU2BixctHwuf9bKtEm
CsJxBhPQjskD3La8NO7Q6HpX5cToiGfDn3ZUx1e6GFA8iHvcYRcTx52V3c4hH9st1qZni+Lgdqo+
zOojurQ8PZcxp4I+45awYXd95skThZqSW9cxRMjIQOoBiDcUYPQnTxW+jqVC8Z4Qil217ov/nhwH
muTEd+t9B1Rjl3x3cr3yhVZHWJina7BW+ixi0p26n7jVX6Eq0U7L2YSJe4BeseYwfJ9R/D1k+9JU
D9HEt0xID2bc2gLooxfuqVcpzJ2ACbOuwWz+D6o+guDs47P2LyzWLtneYkamEMBXuBs/pQ33Gxwh
UGCSyo59dpfJP2QkHVHw44ty8R2t0tPYPSI3l8NcUKCrfJYduKW0+M973127Na+XV0Dt8NsEli5R
XWR7royYYVuPB4S/RwGID6dlnKWgFjCw+DYM7HzsJlwh0mA1vaSq0Dwn9CUvD33AYpWTS3Sgnohi
rtzeQpnyIWmUEIrVLco0GZwkrAvGIxc0e97Sg7wemkKBIGxiptokn923r0g24nX2NmwwAn3bbTiK
vYrX2LXRS9mvtZiGO5qnUBW0SLEaoZPHp2tcxG9oxu489d3EiB0t3/lOHm39GChdYJQUSpOGeS1d
g7xzm2zk8SqRz7HAB3XeQ+La6eZdgsfHbN+H0fH82U8PhoDW51bwo7yAGslRS/zDoWiSb58LPqHA
+fVky5Z/vanrNd4bbBifN2Cg9WBmENHfz4sOVC8MiRnL2/1TSLpwxyKo2iiyPUDPJPle/TCm/RLh
U0NRhSOClAA4E5A7LwQmQv+mMV5ixPgJwlXyvVHLOeMSYrJV2q+dC7skjctTr8GYzj5+yCmUA0Le
zLzcL2jy2JLjEFDhuofxFTdJz1rG1vxaRLercNlpKNoP3n3BVuIx/6foq5TVUU+Wwzy040f5nPed
5FVBLfHF1HBnhfmxIZ/7aLVfeRuRl5QOGTvASPlHa2LEMv8EIDxleE4mpl5rQ8AtuoPvqk4apG9x
2rwzHGzNpv+niSfo2T1PgwStoUyYNJHDRbLCu7VPB5fumADGrsbNKWHzKZ1VqtrOkc9OhxmxQ/Dm
JUGyDTAHPLxKl7wow1awTIOTDdcNs//kbKL7/+xgqCC+8OLOhSzMjRVq3i7G7Y32r2yTHHpQ98RT
9M4+YnMXTN46hA1CO4JkspqrH0UcZwdo3jzfAvKtOjmpEcsDTP9dIdufGSbwlDBfozlu87Q5LuMV
xoG1aqcSNqJVBJnKJS8bq+uwDs/UXeOdY9CvXuaa4kIGWV0JrKztMNaAGZiLu5cTfdZFTVzZIWJg
AC4ZwOPvQIqdynzZI3mJ1/+ZzYQTo4SauqYpd9hFRVyB/v4d/W9aLENxNcdg80cKMgwru/9ZRt23
OSkmSi7eONkpxWrtnu+m3v1HvD3GQGOY5Ps8Kk2fSg8Lpk2DLfd7ugt6n2s4Z8KzGnYYnxwDtDr9
IFottg8CuwO3QFxf2DrhnMOYVCuNtrmxdeN3Ql49BQDuNZbZMT3d4Ku7DCYjmZlW6tCAvqQ4DzCU
r2Ye4KbgU1laOfOOOciDou0xHegFhgw0miRjERgF/6NaTvZy6rKHQ6D8PZrqqR/KvdigDgHyb8t8
v1nVsTm5c4qzm3blEhLxXlIpa5CxEF/27h7RB5qmkIPSj4qoDVUBZxSrJm3Dv/31iB3iuwLHjsxL
UcHk8Mek05IQIpe6ij6p9hbwK978m9Rdqa4qZmRlPUHORTSnkv9utKyUVrx1+q4Yuz7dG0K19Dcj
HefcH8fPnfBtJci5QnodA6TWPfN/jFCdsWWGPQDvAPgY74kSvfXvB3z4F2tdGEkL7j2HF0ZHyLDD
VrsyDl0zbX/zOqbeEuZ6zGUeP4CWMSNyw/uef03VVKAbPmkOIeG+5T5VIQV9SIjqkDN0W6/1WXw3
KUD8vYQlQTdzp9WOd51U8T6yLkcKVipVaeZG3fJ+MNddtbhRMWz6AYtE5e39SedQccjCqQ52ugkO
TLGn74VLMl2wPwVLBwPSuwHLNcnEGwlszZ0Avd8iJIupmUiW3jarRxgyt09vwObOVUoonTOk/HdY
72uz2YDvRxmfn0GT+YWIMJh3E6JWCTRkgCZl5meP8Zt+v7KEsZ7papG2XZMO+4SNy/JCpmVXuOhd
q5vxriFr0sUkyWsDqZf85hB+3B59Adza+GhGW6j5j1TZpnDkdLHLydWqMDjStJGPF2pYsMqLow1g
KkGMeHRqirE0knYs73fpGMiHUjldWHqRY4EDSLEoW4JXCN5AIAd6g5pwUbW1zLe8dRiAYhWb1pMT
2n6QzG2wj6xfNzRTHuBVqnLTpQ+GfwaDDn6C4WB8gRQk+EcaLGdu2PyOTetv53msjO2hvE+SnUqH
P8F4RmY64ozER9Pa1hmjXkhzSCmJaLd/9rkVUreBrR1jUY/84gvr0GPndQo4isyGkledVaVFOeY9
PfGW/WZrBLt7ogex5TfC3vQ9CN30APU8RjpNxnc9lnJjT9qtl8e3Oh7bKLzP9Kb7JmP4DFtdBbq4
9mqOY7gj0hvAbQanVXsAPJcPIodX8WswpPC/O7a5qTbvvrIT1IIkP7taqLdM8qnTA0BowIuvhtJN
rut3s+5IjayPvIrwaSgLIqeRYn5wBqK6JtjV/KN5jNGFB8MX1lxpBgVJieNc419TObgDTSiSrNGr
zkhtjpJzhO7kwIP6SVKxNa+vJX5Ta6WwfpjE0RH1efVWJaAiuH/8u/vINfkdTTatoQqdrfxu2wLx
OVRoL9zUsWa/kGq6a9lR8dhUwaKOzFB8X5gQzLlsjOALVAZJ9ABPVh1jd7oR7Lfm9vwraSpeplst
ltCcItjyRc7WssEg+hszfUSA6mhx5o0j40v2FcDWSccHC7K6zzSn75w4dVcsndcnm/RHqJjI/6eB
UW+LLMdlP3Q43b/IVQRHFS6Ojq/mR19Au3vFqA59+niVm09OqhyAgVPYuNaYT/NPumXsaPRrX/wi
iwwgGK4aQ6/wK0tEyYk5giRMsC4ao8GiRj12ZKQMkwdXo6HwW+eo5dhfLWNi1Wj4/C9XwUiNxruQ
VIlDPKIsLKZglSiQNfpProvURv3YWixnE28TOentIDKkqjekR+CdXxaaP93YqkZj/th/Yt4PbNv5
pib20aQ5plS755s3MDLj2N3jqwE6Nkaa50hLkFESIJhaMGXsSK8EBWG3zQ3EsHgRqqR60I2Fbjww
zIwG+G2HAZRlQjZ0COrFSnBr0mJ5MFGBeg//bnwH1PynbAdirX1NgibJuoCcW722ZLNYpFIdZ0+k
j73RXorQ0gpc9UA7v/bDl3OlIMFatrdKN0n7RuAOe0ZR/BjMwHabQ5AX8/UXTGhAM67sEL57HL2Q
w8d1/zx0h8UaZwxTw1o2AHzTERMle+elJJy94FOw7koygPGtpVLl/2up+yV3sp/IM9LAvwMkNCkt
q7Dd8CclHOcHwJC23zJrtC1C8MOtbhwGD55uPv5w9yJyjVF3z2kZ0xFofvlbWrSWEPv3qgJdwYhT
J5bVrGmZB8WX49ybtFQM9TDZUaT5qyZPCZwdA1E8Xae3KcN7wbvKIeZ2QMFMpfI1/RkI30ud4GcI
uG3ComFPA0jUEJinUDTxwPzEJ0Bvrrd/FSFpe46b9TUN41dw6F26R3u9q8DR39doe3N9PI1gEY8A
MWLaCMPCzs7eQNeITt5DmvQVCKC9UtAU0fynUG/uPqXc+BeYJBadNgIS5O82Z4LfV7/gZ/lLQCFn
ixW8KlnmJrkwa1EZ5lGqOp1aUdVtDnJ1QDkXZN3toOMq1YUVWa3uNlMi7MPCTh0TKY8t1MT/u+4S
QN147wEkeX4Y5gsebOccFiP1CYS+P8siJJUnjwZgBA3ORkqoS8gDHLT7NLMzdp9GhQDGnyKO/BRD
DYits0FNLIjxZ3snoiCH+yVgdFVWioA96Fdl9bXHRSej2erAe51QXkmmIczov1Df5akdrKOHlqkD
fmVKlHm0Hya2yICtMwfoSDmdUaxhsR+kD63l8OWFE1Q41Z+DgP84X2dswJXrIakbwH+2wMBi252a
Nn2CbR2bK/fRWrM/L48HsakMqE07O2uyG2BvsDl3uewOHny0/pw9CUolbFtVwkceEq5Jc4FE+b+P
7qgf92wppk7SGn4Es02WYhGAV3gWuuPVz7ToI1ZEnUdZeYa1Qxn1MkVzydFsbuJc8C5PTwEhUHC8
MkIbTZR34JXduqnUOJJELzZGnG1vFcDZyfDgI5NkBCfz1F1Me7tu6jE4mOAjeswuT61HtA8U7yIr
suZruOFraJuqWU3i0jW4iHtrPbfP6RYM2L7aeWoMHceMVD9iXrZBkElgZPC/XLT/nMHdfe05V8L7
Ppg8ui7dtyE0/XcUlZ4MlzBRhDq4C2sAeRyHWMbW7N7BvcDoz4WnHPf8fRhrtdGPBLMy4cuqMOHk
UaiCe80x/HsUTzySpO6IS2tQ2IY6IOFA+6lxm0qEeM40uNT6VajLLb0Us/mllms3gOfXsFy95pi4
agvhmLQgk1HSMzUVJSXkZZE9Bpt1wnpSljMETHF4QMErldWsHlbCO5dyDhvFRSJIjwhm3aU1yqSi
fuYsDcP5SV9btn4eoUJzJRwftBYA7xj7MJQ5GLvs78QCwQwpoXHoiWaK8ptfJdM6uR6NBeF3Vogs
lWHMieZPsK8Th+k2+47VZexjzLVERBzjdzn7umyM+aD0IfA4PJikKjo3ud9/0LisXxZ9C4oz/Q8s
wa/Xs0izqnGXSBQ2EQjvhsFEcPqZeD87Xd23jHNudlnFiF7HlhZOzWVuPhSdsOoqSAltgq/2SOu6
LKbg0N1hMV0AvwRI0v1GJNTxJAvk+lPyl2ZFd/fmDVrdHfOqaJFqZQbA2utn43+3Zshd2iITeJt1
aauQgBiEYPTKGjhEPZFd5iE7Ys693F8VL3UPJ/MZSXJa+IyjA3PgcBvadMZc1kfK/hjsck9zgKhq
Xug6PQH6SP+OJn+eBdK7QoV6dVQPEC/lPaZqsb6qrwa7nV/aD+j1kBwiBYmWzzR+e+w3BB4BIAU/
cO00f1LYfcPpWktIiRquiQ9pKsw/hYG74C/JkoBPJDQJtp3T59xmo4LBzWhOb+J18Dr6RxTq+Uj4
+yzlcIfE9aTFVcr+jGjgahyMOH7Q9t6kKlu3wMHDDIzKob6XxgYmNleAqquoxllpCrFdjm2AJYMb
xoZhj1kTWBnrDjadXUKoEQXWelNP4CbdXlMBXP5aGwnM4ZLD8A2uD4UQOh7GCyeUPJy0w9F9nQUy
73z54ELs8InZ2ZGjmPemU/XM7PEJ4HKyCGKrrF6bEdfwNRMrlu3vuXjvXpS3P7NO3R9yhzHq39J7
KMEG9V3j7c3nUkNFVJdxqQqyETGXu9drp3ItWo3OsvE6pPCvXjuHEMrP29iw8Yo4KyHhLJL94lp9
9n3PnFeEm6sm/zT6j5sTZIws6jNFz9Oaefb30+We5erzUPcceDUY/1H9bMiyxx/FVCOYn9HCS3w+
aRZ0vzu69IdJZyKkGarTpwq8bh/jQhbct45Ffk0utWDFwMZ0wATW4j2XoZbjM8CGvFNWvsTJsypY
5xg0cwR0Qh7nJ+un7WutlN8G0213IbsuNswdvh3OcPBVBwPJtqBK7gaTzCMbJvBhIDl/XtJ3IF54
UsOt268E5xdLIcioui/3tNz5WYpm0JbpNVt910UySLbA2sClqX+ifDQHjdgE0NaAjYpqfOMhpVQb
Yz0IqlbB1pdBdYFYRNLa04TXM2PdYmsRV0oy2+DWKwc33ASkDGRtV0x+VgsHr6AQZ9xfqc/3W8Y4
0/6lGMmIHCHweZqk4NwpQzglQfIRalj4Tv6N1fu4DsME0YQnSxWnfQbjv+y/k8Ko7PRA1TxXmTIE
6sSV5g9iVOfPArj00wAv3RIVnrZxsiOjHlED+89y1dRp0AZuB7mk1ZNnCWngVaV/O556V8gTKZQ2
62bwl0mHoAEXMAAqOdhEbu14HWyFzkBp0foKHFS3sjZZYJ54d7UyynkDa+PzcVGckOo/3mtfGP2A
vOeIW/a6b2e+UVcLVXJ7IDNhUUo51ljTTzyChamJab8s3DiZtaPH1ELEH2JYSwbjGghijPuCN+Uo
6XioJPK6g1GhTHvl0b7RdXSKDdS0dBqAa0cE6zUvhouhYx4fGjIgrCNLsvSLo9Ox+MQuBwX4KSBx
VytwYQWle7aObwrNA1ibRqr47tc8fhp964EMPtcWjyRvJbVrRGtMw0qfXAcZEmrVpxMc6qqICysg
P095f/c5USHsLwdXE/K7V7CTQrjKu6XUNfuqZAcG9FbApC0UqoGhTDw6FpMkuiS2fTJDYkVO6gU8
0uQbdKXadRVyMMQIPfBYB39nPWLg4uiOoIe4biP/0mLl7xlfl2+lVIcDEh8kZCyGTrz8IH1tOUTs
OLmMrzz07tliuCX9MbdzkIVBlb2GuxlycIqKBD0daYOsSA9ys0eK3SgRXRbYc76mh53NwZLROGH3
SChdXpWbjOy8oz2FV/SGAn/LwC/T+7APGTfSXJqYonb8JXNP2PD2msc+i60NBZ1IZj9cr+wPQdhY
A+w8vPfuv72V4vnLZ8hyuUj7hDnzk9SGR2PfAuf74Pf+Y4QNm28MT4YQglsn/SZwaIMMLwF8wdqe
z2vm/YYst9Y0r3ECe4sVnFR/JiDkWMYP3HJLr+ehfA3xHJpL8TKLRXzvvNNbn1zJlXvx8mcA+j+s
5QCIUD4Hx3tU24TevfNgE0U0Z1sPnzvEQ3zL6u3KFK3Ao5AhzYtltDgK8b3X5ZZ8bq198i5+b/Wh
vlhJgoRB80tk89V6Ut6mZ7bFx17psJcdY8jdiDyw8QPEFtc3hyg1YS8oVWO3xZOX2K6pQwSewpIr
IjG28knJ0/z0JlP/grt1Pp0x02P+MNt39H34VOyBEdWqmBH0TltCLvU4/TAxEwZLVTqWCcF4aunM
K9uzel75zu5oFHQv3jIHWAAQ3VIHZYS+EVLLNBaE+eYqVEuvaJPMY9hJWIjyhNAk7LAoxtMU3wUL
Nw1x+pNmTk6sq9FqEEOeMxW9hzbWMDb5tUlpXl1RgICQTxHW2IFaFKBDDkhTB6f0kSFYJDYdMnfi
OVYGFv1WQda9WbfrF+pMabj8h1Z00WQJw+2FcIgLU2RiCX2BqvimZFCjOkVnwdwDXxQ5UmcxvbkW
QWynrCvt9tZoL/AKyy2MrZrzswfgrBanAAUfRXDwcvrnuzQg7UZok3fPaagCAXM0ucUTpAxomLWO
31oomM1MRRonBBZY6uNl+2ZGU6Gfnf7b3vNrQc8t4A4wxDQ6rqftar6Pd43Vgr3StsW643QUlpGx
r98Fy5A24kqw6fcuKf9Nu4ZAcbuCjPj3eBwNtN195l/LhaMwVqrsjdK4HHfej68hTLCv+oW6TMCG
AoHcOScj9XwGz9GEUEFPv+yFtq3zFiTRxVk56hA4dX+1L+m29AbqaTal5hA9yq2tMSpZDHWfEWGe
pKedT6lcmluywPyt5Ij7JzXqK77L7zyS5gzEGnC9u1Yi48QpHlWCfXq5nsD9n0HStFX45mpIBPPK
g3RWxRYQI/QMg/KAVV96gmXD0CQaJeFuSYtwNIB7XB0XRbJ6vAycyMrTN2BT5X26StHkolby6sA0
muUOGKijB8QgnUh9cq5irEUI38hADYQsr1/ab6wfFi0+Ck+n6jtPuiONfgfGuTWmqPO2BTRpoSBv
4EY4hZv55oanQ9eCRCDozUIU3iGa+kKzfx7oJqvrEv6/JH7G0h2O+IqZHefj9mSJclgg5RVFjU91
aZ1xSbnVE7xPJA2Al91CyTCyexMkyrdquhAkqJnQd5fRcqDk+VbezJqQIQV5NxH2ip0gvGYbTLeJ
smALM/c79RcCzuPGRqOOoh9Aq2YGpbF04hi76r2D8eV6sLXAa91qKIC4JasGm5ON9CA4r9ZcZvRT
GyQaJDhqU1ifgbIt0czO3XIrkXVdAxgVL2hqhxNv+ohJYn4nLKotGmUOQj/tkKdLH4YgNhCA/39w
9KEiowqjSIbHdMwcx4gx5GUAfKzo5CdvlVteMxQ+C/tEnjHo5K5CcGzXjCNEgk9AxruwxlE5uf+6
oZvabFjZ1rJmDc6qCyxWTMHa8rDRCtMU/s6nCh6ScV+0xgig6rMcH6vsFSuIlCLEV7W2/wyo8omC
I/dVjbMZEvREABWQbzOmg6HR2bWtANR9+niJ2uSv5KTNuDn1/zINwIU0hzbHMAZlXAxamf7GT5xO
m7B4khE4gxf3Bv/3tycW8W6IXrOwPonMAd75lJVgSdE0m3n2UEaApFY/yuow2VcfdEp15R6T6uZM
CJska1Zk7M6cXgVjJNFzohHWRUroJYibM9w70iw0rl5rfcUhHijrYx/Yzb/rTPM3gr0cuC6yJ944
VttQa7+qvowq0yrO5QdoarWimjLEQyL/wZ+gdfXbn7W5SCzfXI97Fif4elAZYAaKPS/qsRu9NoWs
S8AmFI1sPjcX4C0Z9j1bFqDiFrh1kMYXOj20ez1i21fUHlyN7IsVxwjT1Lr/075V+7hETYTwcTpN
tl4P+2FJ4dbYcxnZWfWb+UXRTDb1aLPRuFYMvEpcLM7ZZuBGFbeUM7xSl1Z50DFw1KnpWKYWJ+tH
Qz4n8cP+enSX2gtG5gdDQicuxCNa42CMaKx53ZQmO+xJC7Tk4Vne3ZRMCV+hAGykrxBfiPEPHMeW
aAYa/xZtmOzpHaHaCfnEShM5qQ1tNVv7rGinXP5FqomhZI5mvpGVjE9vbo/PNvDUKQcRtaEnMqzu
Nrn/ZbkRjOSI5Ga6jd48hGq7EzWh9/YaRA8aClpM3esLtBKUAEgDIRzfnNzpVfi1Qvli4vAH/7zI
9OHFn67pJ8HEnTR2/xhraE5rMH629BQ+b2hQ1vNYjU4jwucYi0CnDSyTzc9E3j2BVCqWxa31kgeL
hjufXMLCea7GWooPPd3moEMHdBncK89OkYuunJd3/44XDoaikQ2nHYMJ6LyXbOfMEaltajeE25pk
dYJombQImBC46GTA/edxDvHz1FWOsp4KPGvx+vJl9lpbNNMLR25UvOzLgetq9Ssy8hga8WZA3Fzx
gtb1I+mIqAsvo5G6jlAiZhO3af5oKJCqfsH1g8meeAUvCJQcyUtTTRDhp+MiuRwm4zisnxrSTHXm
jPX/9fGu4r/R8uD4hkYyDqIUBv271cM8co/sSeZXZLGrmLiqQ/K6Y6JWrSOOwM/KSgywUSp+Zmuu
3MERNupmD82BuccZP376oggDd1Tan5J3pTTjcaU8+r6UCxnQTvyqFxVIVsd40ryrcdlswSfIo/Ws
KSSQN26FmlpRyH+a3+L8RZet5cB4gDNhyUNQ7yYsgq4hdVjX8g4ECxknBxdoIUfSxXhd4+puBsGB
3SURSMKRReoc7Atr3fUJqq1M0KGlEvEI1IbpbVuesuyaqG08uqukW0D8ckjPyeNwYchUTkoJU9zP
YSgJYqCwyewYTdUMDboQdrxXlUqRh0Vn1q3RdizM4tywGhTwkdwTGf5awCuCI5qGByOdKV3KnsVr
LxMbviO9uUyUelDF1CDvXbkHyqdzKeCtKfgGynChJA7zSCgb1g6edcyxtFGBYs68X8chiPiP5vjX
RABBCIXS1emjV1ENdeGy6sn69isYc7vKo9LdbG6hqUpbwRSqncjrC/FDVmd7G9KdlaD+oq5a8gsC
j60M84V4xPGoGoeinDWVz5E8Go16dbMju+dbHB7gxzQDs6QMBN8ju55tr8kMgaCfsAffJsZC+WJn
hTaYmQsKL2ZveO/6afhw2sQb+1HQ6/7AmfmK//oIjWxgsnf01feeMtKTp7MdEclVgq0+lweBlpbm
cIxRRyMYvYv3QcXDr5Jj3XBqvsZCfYlLToRRoViUTT2/y+Vvt2FhJe0uh0Ekgetvobn7xH9bJrMD
nsqbMAd5aIPQVEoZZLAc0yVZ+RMCwMG6sgtXF/WPnfBM1s+9QU5A3tMv3uGgaTDUutQgQO3NJwPy
ZnvVpDEIf4hWMZVwAyE6dBvHvuyhwObyGV9u0sw81XhW38FV5/7CFdGiiQML/aEAQ90YaRAxI2mn
REU14w7EMyeZyPrY8iP9Jp6sOkUEz4Q8+fZUmT6T0z3aiCzKLmAA3gcHCZ+8yS40HZ2yWTHsOA1m
+F2lepqY1jUKWRkSh2fh/T4uW9KC1685gihKZtI1X09dwnuCU8cAdcbQrHIlORyAqxpiLQ2qBsdy
l3D/GyMFbis+66BDfXDB5l9bGdDSdtNHCG8OsCXW3Vx4ceGcaLUXvgKmAUBw0dLmDvFAidN669AH
PEGQsdz0UmbkmE6vus5IrGvVMDnPT59UQVdFfebIOYTtK/IIkK3bUzkxLkqiO84gXKXFx7l56GGl
lhE3pKMaIozxjCYeu4+VxXdCdzYHXheRi5k92ZvtsWUBquR9YJ71UMSeLzULEsikHIdt5GRIqRB/
6KQt/OdInM2U7unwMlV2a/wOJPj/YGNwOVk2MVzDr4pa6AqTxejQXf2+0ji3ff3yOIR2ZqGoa4U3
fo1l7Bwv4RJS6HDOY+HqTRg1J2zUS9wM4YQ5CuPIiB+zzhZynr16dSADeLKJfBVjVMeHhB1L8RBj
Kf0YC6tA7PQpsscX/dELl0lGSKYpgX02rL9l7gTeWH/i5Jwl3EKbppZLctaV1M5IeAc1CxWbE0Bo
xiI/g6lV8haVxUKj50XekJtgCFLn450uONlC+rYT8lEVUtLtyaMcdAahuie2lTXGdMZWXMKZ5fWt
Bd2S0DjTfpjyZ2AAcXkHAD1cUQA6LmclAtXcxmNR65SCfbgccNH92gPQn+pdppTuhu9TSj5O6haJ
Cb5OmwQ23coUa4ssRFGHBcBVVzsb8vHHfssGC5umNk6GHafEcWM0JwwPp8k9fs0ZeQhiRWfHdKg+
dew0hYxqY1KCRxX+EaSw3xoj3FvlpMQT+FgAlHilmh595FNGJrGT4wpc500nryp/H/fksEAzQOUG
yV7lUfjbNZarWJw1sbZHUj93lgjwKvgUV2Pq4uZihnmZmrfdTeE52249CWZZVXolZVLozPwmNr6w
lgS4GNSTmT4ItSqsV+yNeO15CsUv3AhHh2RsOn8HKjWa/3YQJ0fAB37RiX7zkD3UVrYX19DugmRA
1h1bVEGk1EGUl0eu4tA+BAoOPGoiJFakblFEjPLgaJSIArVf7EIvfOGfErO5Me9DynBz16MJUJnR
xO5xIZ0mS/KqJ6cuhxPipsMUlDnzMBok921b7FQieqZcu4mJAgVKyHKf5yXoQpXUO/+Hpae+u/U/
az5zToizhQnc1PwuOrywTOIW1JjPbKgs1+pBmpQOuXPPhAVVH0tDuWP18pjnihjSDNXZKPicZAJw
hbGtjnEmHoW6tRt3vQXZfdcMape2VBDgQp6Q8DFsV0RFNXhMutpyeMKSMrRuFE1jKHRzvI/UE1ka
ByMBhuj+1Nibzq4HtNhShadoeYiZlfQMDuHV6XozM3swFqzqxHi9oeKg2UHtpnP8R35e/1zeml4i
oF5jJ2CzE+vqPLS9dFuaWbdIWSUaskfq/Xf+MGLqsMM9ghGe6V4JfRMvz0dWfo8aehSyvv9kOnLA
yGyvM0u35Ihvn5gQ9E1vuJTspb11KdakqX1UKTbCmSwydODYD7dvK8iO0nWy6kF0FF4FzXbIV/xx
v2rV/ctm1CLmHhJvo8Kj0qdf4ywo/v+JwbMbD1EbvN7nIEdMknSN4/nQ1iZ4hVq+hhFBjNyRzcjZ
tUWINU71/7hX1tKbJstheX47oguNKiQ9I4Jn9OODcpG6/rJ1zt2m3Ln9MclbtGQzp3JJLUoXmUhw
GRQ+y4xp4/muuuKQSHFTtSvO8UivaRBlrmMbYQ1WAYh/tvElwOcrBdd9Bzn85Laf/wItxmYWF7n5
1Q04CbXJ9tiHSXgOT/ooq5tk1DK+5C3+JpGQ9bRp50qoYY7Kftt7feqMsQbkmEshMjrDIFmJ21Br
e8/LzJIFBnnhOClWz/CyCMdUS5aSsVg1H7lKRT0I9lC04KaLfH3v3+ana56XW9viqAC3GDGIH2OA
70XXD0SKiqzyEJEqNieSL6pFI6J3joe5c/FSyptlRUJVtr8vPQ8G6p7SHKcMzvbAKn7+V6FCLSSP
exumX8bPtzz/KJnDFQ+a+9aM90fIWEgYHLeLzjfwgWSbe1zBG+VPpEyCw2P082AtAybdmkrN4rpz
yp1y4wu7rTVi7g5Mzdc6LwEBRnojqF7ysph3YXcighnchsFojDF6cde2iG1/DRmBTYNOa7jjvP4c
wiX9f6WPiJ8LA6r+eyOL78sOz71P6QInU+qFie4808YC3kNK9etjWDm3oDlE3kaLspawho4daWSK
Z4PsTXakchcSCn8mh5gg+0BZ4nPnsw8Cho4yB23giLBFnG33p5F7bXMTKJJaYN6L50kDI5HsUVc6
xOdZyw4HAB+BEFO7Fm2WX/CXY7qZ4aZz927Wj3YBKsI2HOSH/Vcs8CCmyUKKwmCoHi5iP3ZNiyBQ
IINEmxz06A/rcgTz6denHDb0+BfOZKI+9cjC6M/e3f+Bt2+7DXYGvLRojvcJwdc1nOiSUCYayv60
pBliBN1qtIC0cfXmlmF3DCJHnd/2U4YTBY3zaye75C29Mbr2bPuapub5YbXzBDtuyLAKO6E4N2T8
Vn4Xoc3UrYqP32zEs9N0hR3QtjbqrLeuBqSWyI6dwy3CR5KMJ1v+2ZcrdLiy+6MnMu2w8ywcAIfW
+1UbwHyATd/ZvQus+rs8Q5fFfe9qSPD+0BYphNfYyc1Uu3OD5qjpjIa6n7SZ9qn4H1SLC3AMH9rS
hIhX68U/y6yO/GMBUTDmuNu9XTYjNtVQLuCZbZB5gjOsh5qcmRtuyoiqrVYl+Rmev0jrCuqfVdBy
QsP6oA6Lat9pCAxQqNd2PvCcOGhT2n+oI4A2KxkOmdXNW+NrgfQ0xA855cRgEXf+wVNPEEh4c8Bu
XIpR2jAkUz9cuGCwmnVUO7Pa9PgtlnTuzdfVHGVsXdssjX/6MpBSSc04j2Xr9Ws76fAOrDb7vhxB
StijVHDO9v4h/4lwiD4iy4gwOG0IgOvKRtxs1qAQC6LcYpQbh8eY3nLXDWPIJZOCU6tHw7bXiAP5
T6XIYAviprG8gaeIip0BtagSpsh56Z+YMbP9QpTyqZEILC1E9JEI0nxh3UJrIPVA4hnkS5g85tX8
DJqgGsAjRobLiszs6lTQhpDzx+ttw7lLx8zJMHKpanJJN0mZafH+PGHS34eXuw1HV72/Da4VUsm5
BOZCtH07IXadlO1HjA0GE2hi3bJFoeCymOMKDcm+Cr449EpRsgO8npGHgshvQqfHoJmcI6/z/DsG
E2/LHlPK1/fGRvThiHgsiJnMrnaAXjVBFmINgpA/0SChiinX0BKXB+WnI2kruBmvqFt1gqwfJWAQ
6kjG2OUi5IfAU2MHt6pDD16cyCXsIQULtZIv65MyJQQk3wAfdpZGWeGMTR2PM4xf5J6cR/jGQpov
WcZlX5BkppRp2twHhbz+fqHDkwJ9DlN8G4mRupFeTAVGdjioqWXnagjeDZ7XsZ1/lBAwYMeVsD51
EB3HfhnpGwqgQ3rQlK66RFE0Ivk0bK4JswWM12zEjTXUVCE1ZRhI+5HOKFfv6Qm0bb7qg6mK6fsm
lqVXjRB9cWtLWQQBrgxPIeRAmBKHVEXSbwhHTLWyi0ap10hDYGC+nP1fA8eTe5m7yHbnFQZD+s2R
sP35HqIVOXaICHP10dic7dt7I4QQ5WwA4L1QvoGnuZEUr4ElmZ/9kY+0XUX4mkbZkcg98KclE2B0
LREcjebv3l+R+Qc7zJEN8HgPX+s+3kOI3KAc8Qsi0k7EOSa8gX8WEj5yH1E0wVvAUpkwW4fZnoDI
BGZdbPYJm5dLCrXpz/yjbI87N1slUopepRzRqtA0ieMlr9JxPhZ68QjLSG6qWuLnW9PqH08vjF7g
Gm8YvOxJsLSIy+K1DdwOjaVIa16STcz5JPpLwqc1pgFp+nAN9KQsV/vD/c1uq8JSvADnxiwd98Rc
HWQY7kprcocZMkXu41w36mUJ4Ux7+8OfC+YQyWbHEvew7XAbUWvpqfw7lXmL0WvKZrUDvYrOOf3o
cbG/yXJiJcEb71LYXH+9W47mRgplchqAYUTljx1vBSlo0qXs+4PjKkbSRC/Iu2tBY6ZGbLYscckb
IssM5uBnVasCbxOF7bvPZvBqgsVtsuALc8XoA+CtNrplZUWsgyJ1dvsTwkl3trnbGy/zjoUj3j9C
FgQECIvf3Zp0vpW7q5BrnB2vDcz2TSeRl5Pv8D0tf04NJ3OrI/H/9T7WRjGmBWyeyO9+TemUAA+r
3C1SsZmkD8UGfv2PEpuo2jHWYnK+gaVof90WsaCisogfwVDbQlMSOkhP+n94cqg3v8Ns5q5a0kIu
sEozJjX35QYQslOylHFCBkHAX88bbgHC6kqMelFIW/hERmm7PK19kr1mLvA7I1vcDwOyZxUoh8/K
sXkeGOdweVYbrpoy3dV24Q0C/c/9pNE39/NB7Ry1HmzvuCiHFwcQAAnSZc2tCUmfaJ/NS3uE9xsY
dunhr625PyEL+oUq85WlfhcKetC6Q7I4iNa9cXHEvSlSp8WDQYTpnrGxjpgIkQ3US0u0+JLyPIEk
aGmSvJxcCpS3AXZ9tJGWj9d4/XkYAiaCfRIQrqiJdJrXovrIJaXmRd6TOhQK14Fchy4+Swu47qDj
PJ0GQUSej7i1boExwuwZsv3HJhkSvdW5DkDD5nLCghQEj8vGC3Y166CPoMMD3p98Z+Li/KdB+hNx
FJfgnxhx1mxVZLvCK3UZEH1IlWsOxelM8r//zirZJC7gKjUJmymMg+MteOA6DAH+Jj0ZcI+aik0p
Bwpdyy8SflcPZ060r3UTcpS/DIHFS58YJgNqI3B8JZn+6BP2U6AiRroWZVtuW9wsC8YNSQE/fAHI
Gn1HejJs200rsTxTo0v9T3EDASpQtvCKHgXutLFaiOf7bf33ttUkCZVNHBR7UYZeDDE8nHcYbnGN
eawl2lveChjjWrpPdZrGV09lcxKpdeOdPVfhf1YezsOSYiEnx4XrqElzS8JirhycAIor1/IsAVcn
zyhQjYbNnbGan0k8uJ6R5h5koT8qrXgboXhPBcOnkv988E2Mm+SlWlQFYY6Wf/4E1H39MFPSFLB8
04V9BTS38MOkN1zEeuZ1IsDs3RqRfEu25k9AeIuYJVWsCuSr9HvvnFvmWj7+9wcNYHiOlhpuw/sz
X7L3A9bpsKyYTLyXhKmxLJX3EHezJwTVMaQArcQhMKSULCYXQTZDtJ7mT5vupgwdzJb6raKFl19M
bhizapPY3aRE6QGTvDwoGQQiFZzl1V/EYx8v4YS0x9jUhNzYcS9kfTvO1TNLoFYM0w5CzTa/j/QH
9N0EQdhYPdnXZRmeLzUdCUe5DKMX5ic1dlznHTIo6QfJmH0tq62s1fO6bIm19+qJcjaFgJOarqx3
ICCMpQ4znkkK02Mxxp0XUUxYEebxtCSrZHo1uzkpLQ4NxDLYTYE0nD9+9gda2gv+DoA+kptpSZYt
oO49HJjJG/f6hxraDX8nfPA5aQGs0CZoRMoBGR4kaxLxiNGJ1mmVKyLFS65eHFQixh4pgnS3ojE4
BIblbuBKVbsP46HrBn4PpGQPhMrNItHBkkzSKQ/XEQzaw4xiCOIGeSWLva6H4WATtEIFqHCBYgF6
JHlAT1T7S6As6MlxRFJ4xxqq+zEJCk+3N+be1TyHBzMtZTVpA3aBeqjWKpwR1S4G67/z7Ot56Y1j
8p8QnWcQDyzmhFMU2kayncCuWDJVxyw4sFCVJy+5997yA1gXxhB2JKuHcVYNkh8byvHIakIB4Ghh
OrmADmkVfkNyLG2LWfCmoLdop3yArnDo3Q4+vgA5P0u6WiLqewHLCprrMGhSPVbyow89AzoTJx6d
D0dmhgfmCZMm6oYeSBTarNquy6m16nJOgDfSUPNPnoAks1QTu/hwoPMKsj28+h1/mtzXX3yzEE17
PsNqSFyxuIcd3LOhKLinKv8Omr68kxN6mMyPnODZn9DzLeYjwj28wvRq09PCvOnc9nOL8xPALUfs
hogXLP9iUuDZmWwu3mfgwtnfv48s8nqlwfGRuFb+RFDL4xrrw0MRzN9KTwapePYa8mJNauu6ZnLG
nS2Wia25X20Jw8XYqOEFMCbjZIzTA9O7MrAgF7iC/6Lhd4BGbXvdut7xZHdJf1Id3lcTOObwJon3
tl0rFr7IvoykRqmaPDH5GaLWE4QwuOppTY7HdRlSWZ/QtoIFkNnrktqs8MBtcO2jW60wJ1z4joWC
VsN76W2cMvMcXKUw7LvQZCh9cuQAm+iKelDeP8nqMC7KBuC6NmMTqWRV7dL59wiQoGshsE9qHEUg
FGPKHkQCVX9vDERx8iQh7eu2vzfReeQMv6J7BD5H8OqtGEZCTNRfbUqMB+LLyyJoHUfLY6Pt+qtj
CgKT+pE10UdQ23L+ko2qDrSrnw5EvRpw/BFVxN/WolUB/YVDqzMHpAZBUBKtifMalaNKF7lUKW4+
ze2rF4IgRiYKZDhtP29HWlwivc0tBvykxF1GOIeO4luIAAnCIb3C6g4YmUFW4GuDf9m5xyaNadJJ
4cEO8NVNLrmyfDw/wMYqYRjJA/Wi+Lle1zR1Y9pFVUzDk3oUWrBv5ZMR/R4un2yNSprJXymxdptD
ryZcjTf5W4HRQDcmbB8iiLRnemxVGFktnsMg5LytyKlVwlW1oPrvtvOe/JGQ6CujwPpr8OlkSlMJ
MiIbzm+AtThma2vjBi3Zn5mJu+ANAaQbmJ0lGxDiU98MQ6/xPYNHrSonmnhnuNFrwn8HdXTobFtw
mHjod9zu4/IRyB28sXEHubKizSpHzBt60MEywBjh1mVzk2m1QF/Hq5isyY8rCj44Xwkz8PcrUVkd
Szr17OUBx+2pHDFUVcOaG4qnHNJyJ/MgIfckLmNfmhhOkF3QfpqZ9QNAcUHSv8ambLmMdqeQZqKT
FOCTPUzRoNTTjSfZurjPUUWeKEJUJvZdDpw6pwUfGQD0Oqbq31zANOY7O2/WjI7JpWZ+FaqGFLqO
mQPsF9ZtcFeNYtlwJcSk3QryBiB0SWNrIAnTMq9G8OF+ONq1vOQXK0Fv3HX9/B1wzkG2Vy88YLNP
Ra2Sh9k+wW4/xwm7WJooGlOQqvpqSFwTbGwdI4jx50/WCzEUjCddLMGSxcSV4dtlLkSfCnPTNPMG
p0MPNVOexry3hHEmEx7cqd+Q3AkBrWejzJYRCRyu8nAiTLWuSjPQNGYt4nHj8n7fU6wOUQFWRN42
s6V4IRrHm8Lpz0KWLENwy+0CJMu6+ha3QBjgxYgOElljQlTyqlZF4xvL3fvO5XUki4UyRyAfKd3D
rTQzkSxIoJ2UZ/2G8zlKOKprV+mSy73eVt5K22+4e6LCdIAIPnkXRIOdSfVaMXF4prd92MTWQMPO
gCKW5+PcBPC/29CxG8YHpr1kjzbsRec7s7+Cjd3/ORvuBGC+ZSJ1ujkHXNfEyYM3II7tgflCKMYP
buiDxcsFwJRsTJGo42K6lvJ3AAogTin6MnkFdRY0crxH81RxkLBo4xlBw1h1K8BCnrYfa2m7LDVw
t6uuFj7SMT6L0adyHEWfUBQ4ar7wwETfpWlMe9YWKn+FSMWMEtUomQ+nvFl3bLpM0MpUBE2jtKA/
aW2/8LxoGgfadQs4O9jpp6OUa2F07qzhX98nDVm7hMibLt8q+h2VaWRkN6OhFSTuck0pLErmUyJ2
RWfg5U7c/9ax5yMBxm6Y9ia+sf7oChfsoagzBaCHOZJO7ByBDDTOpgWDACc5IyJZn43VlhIdFZ/K
GDUpkyqvW5GbMcyMR/oT+ll8gjW7yxnxH9ZzSBSxLK5FPKPIpqGO+ssFhSZZ1V9+Q/9QZqeurGD7
hSY0JEs3/pVOFyz3eGyTCSZPCHHKYpc5a2DGIsG5IhkUolXCIXg9birZOeezA6aJgiqmTqWD/5u1
+rmUEA8Hv9BR/Za2aiqPjRISJX+yhUF8drb6b6vHRPTExCpFbuZg9iT0r3aFAnZ5XYJdaMJQ5pre
7zfBkQ0O0rggAeULI4ubSApwBdJS8CP8tCU0O8t2tgFBH7KzKV/56QHVNhORtfogFNjxGj2X+T/M
ZrN7u2QgPvch6c4Cs1kDEwFu3jc70/Yq0kigWd7PbLcoWBmM8at6VQaCxWR1TmSwCYUeCfbmrxbo
Mr1UOaFMkNPAvZnb3gdeDk0DJa6f4kVsOuKSKRNa/y9bdZZytNSHn0sJUo7A6oLA/KosCWBlgaAd
QsWJ2g1MN1p4UG1Fx2PBPNDWrCpr95uktsJYeCFCWEUV+poocUAFlI8swMGmNWHEi9AwmYSpKAki
ThAZDSTnQgX3ZnsM1NMXm6C1NDvN9AvDmQbvGFvuz/AITPpB+7XTJ7HtbmXAfx8CagJ+TN5c8Yrm
I34ucAAQshYUnVIlaPtPn74Ic7al6/cov2nftu4CELnHAqzlHaHhmRvGEDabjKSaHm3U+GFVKk/p
Hw0MOgSeFqTr57ljZUjlOl21blfsxT9eLGOJ4NfljPCI1vtbdwPVQcMHQQGXfLBZiFA38c+9CkIY
07uyKETVbjxukBsnttI0AvoWmDpyJmWwlB+1sZZ62TmTyEjklt+FPgOGSftMQQjXwL8G2JCBarIH
0cIWSQ1V5YvM7q/mcs8deFu25jJ5IQEV1GFK2kEYUMxFKPV3MmzSSVQCRFfqSxmCz5ru/B7CUaj8
6jfx++54brqLM8jM+D/Dq83DF8wK0ullAiYyiqQ4GJjKc+BArKFrTlPZb0uwd+fLleWnGl37qFNf
wTCygfYByneQYG/rHkKSydUPa+fAGBsq/OyHdsRr01dVlbIwrCkL3EC1ZDY9ULQJJh1CXk8Xq4TO
Ko8HGJ/kyLgshDOa07jFU4co03wIdSNom8Onch+k9QEwypXRbqyK/T7IgUXyq3FqNXkSK4M1UBbV
/G/qKZCK+ygyrjT6TGeek6oW3+Cv4rMmuynHG5JudqBAE5WUOCk1ceK63RLzfrJu0O9/lFK50+ei
OgR2gIVii6RpSK1YYMJ1Py0bB/1jYeTh4UnbuT/5AHnazpjWAbR188LkinlRX119+Sjc75Copqtd
g8uKj3LO1hxP03FVTu9n0IPWwvyXWevXls7UmfjsVhC0ZrbLoyE6KvNbJFkSzVdmgGpOFb86zSMy
UjF7DyVSnKQ8gjTBcLE1CPJ/jDCZCj1J8DgpH28joSlOpGEUbJ/RLFP5PJGnoEBpA7rtvtrNUyvh
ADVv4mRwEFuN15EHE3uLZVYGV5MhtZwF/pKCQKXnRlABWNJ6tK92LX+50R7j9YdJLB+hG+WaPRQ6
rLk1eOV4oBV0a+mPrMg+it1zKiHSLWw7y+jrC7c2uyiwAqoE6mJDmqyG0GYOZKFhfiOrL2BIObo/
btqU6qgoDb9UNc2sfHwCNf2+SJIcQB8q417t4fMie9wtoWJHID/XSWdGYWZfxgc6xA7O8x/P+RN3
7afi7aHCop3u++FK20/xO6X2p99VOxz4ijOO+J8U4qV8EXV85+2gZwCMyaQPCOFIkvAbzX/ZcG5X
aO18TI0ly9oGyD8vAbwuM3XU2M/r/V3NQg82zKtElbpQD+a5JYpL+MXu71LFd61DkMJiHhY+cuFe
NQydj6zSQa7t4UURjY0IarV1/2TPdYxOxISi8PuoO2D9xJUrNZu/v3nI2hjChsQq5Pu79QId4ydI
jaQY0DWyNFW5yG5VVjhFcy8hXYV0Fd3cbk70MJRbg/vCkR/yj3PEB3OWpCFqi3qpiJVxrd53MBWn
P0rSU+Ft7SHqlbel4NzjAh4IeqzATVmm0y/q+S8EF+stfqtoDmsC5l4PEYkY8R44W0/KUaBoFyDb
5VPPWmk7YCZa05zhAzfcF84h18Vt1ry2bXn9tKWwnR9yo6in3XHzl+zHT9WzbD3TRXuVaCuBubCp
5nbIEi6lsNUufkqGwN0aSF0XsR8QDod9LwLxj366b1hREnQfyUIbpHJS+PRVgJFluw3ymJpcjf3w
hhqUEqfTgizCjUBVWO9TOtbMrCyQI9WPxj/CVCsR48frN1AwUT9x3fONMcEk94fSPMY4PRi99YNB
yq/e33F2yimE1WXcmNYboqUMtMO3NXXVpsQX4rFA/Nd4VwLlyoe6djY4fl8QoFpqPZP63coRNRGy
bVKJCPaC8P9UYgwIoEvjxFiHsrBu9N42tzCdx4l7spqbf8rAIRuoRn885oyxbh8cBWFx/UsnLnAB
ErmV8gwwg9ih9loFJ1mpETdEk+IGzcr/S6mPbFIBi0CmgFC4aQuISmmlqM0CK4pyfRZMSwz57SRr
qtYKKBR1z+MDy6Oi80iIxmj4sVgJPXOBD0nKqBs0Io8Tcl8UWzdluC+F0PU0I1q38OUCsw75Lqqa
L537711CUTMwcplqIOGBF+9lOX7HDsybkTjSgeAqbZvTl2KAFllTd0gz8li5qMdisHE87Jx5QznO
ycs7HJ6zTYdIFc35h1DOlNxwnSY+9aRS4KzAIIVHNz8Ka/yj4CiWgPQ60KUOOyMTeUImDtE/pTig
+N9cP/KpWfOzxSJ8xD4qLnPTCAVMuoKPghp3mMMs4uIFbX890waeuY/qLcgS/3In771tEfkncBdY
9e2oqgQOQ9r95yO/ex5Vvvj8UqA5c4G0IwpkjqNh43MNmjZip8Y4WnU7WvcSwkiKC083wy8shqCo
evr2E+cP7RHz/F/RQiycIsgK8CE5W1mEfkYrpVZ1q5EJxhuSY5uyXjl3L0R60a/kFRfl0noQftQq
d6mErwtPbaYkq/FrGXucr4hC1uARiyX0I2VJkkpvj0HfMVSVVAmFyG5RuS3D3W8/tlkOq9y8b8yY
xXKrQV68tM7Kjb0dXhGOqbRVeYAAJ2EmlGgyl3flS3AtmpiIqpJS0snqiEv1OCe+LOTq6FI/f+fn
83reAJuOFOEYm9SYsMQ4+qWNdpPyWDUhWWvwHupnPWR3c3BVH6EsozEPYSe0li9Z/U6GVcqlg5NO
TZn7br55Sy23HqDxPSqxfebNmcei3ts3AFmxkFQ+pbveeBdbnZCT+iIa4WPDvebBAwdhiF1If78b
6z/T0RszTU7TVvqI9hXfzUBpI8WK9qLpQEqiso06pXJwURM0ldAFhTlpwIscuUm0K84RA4jv7OT2
uB/DekU7duq8EcosPriY7Qmqb9ZAfPcjV4ZjDuVYJ5CfImRxMReW0K/mue6XHRK9oduTCopX2bdq
woBCq/RnWhJYStnLus+IAEHgTM7EGx2Igr3h6Z8uFhINdFrIx8oeR+3hMQqRwRuqlIs9Zew9V1Au
YGLHzHImCuWTyGBrvVa3+03T+oU4xsFqeM9pfBEoU5uE0PNp7Y00wSt8qz+weGhphS5iKpymh4+N
smhPcjwzL3sbH5i9mAb9RxYoX2K5NHwgPSb1LVgEpCWR2q2X0cs9JM40VBOBMc3grLZSd11xPyTR
n/y4jm09zRY1U+GH/SLSQ6xwLrSh3/d/Xqwt7m1ZfqiePSSafknKRQrumf3nfQPXsoZCnZyB5CHp
I/pd9ABzRBdTgU8zCD5Q2Cmp9Hu4WmUONVWC3qGFGJLj8axQWf2Oo4I4L4hkzJ5rFPCMNOoVyAPp
FWabGr45iStB3u/31vUoM1tF29WWUScnutn/OJYa51qynp6/b3jWCeVjw78l6OXnt/3LYdVrMrVf
XjUrFuUg9/f8fLpPhXOsNk/PcCQRBxogvmT3qvCqhSaSvPO0aa+xrfiUNrFC5hxe2kpxnoc9QA9e
yCmgPle8u+DQXQePHLEVoMdMMyzRwjXWAIdFhd/J464QgkOSJ55z1xRLofXjyEYP/A53Z8FicA8t
4mxi3P6CaRoO/gk9I3Ir7Fz6rhscePy+C7WjBB2hCUKx/Q6nxqI6V5dfc9PRgFSma+tJ+btDhQ+k
y+8+ZBOf4kzSG38wBuQ9Yjcy1Uyz2j1Qpd6LUr4VTfkGHBnKMvwI/pYvAcNtj6CM44fUVVWLbnkO
ebgPYu7NUQiHR/J2TQOjDpZ3nZDhC5j/c1R6zZOo6lT+vUASNiQOUKbrgHgS892tWGS22H7RJFhi
I4I7fEkd4Jlq39TE+882p9tPUKIH9UFiCh0t8HZH5jrRa2Q7KWibApKvcBvaX/io98Ya1+CGAMw6
+fryt+4WL4JBvjhzfNJXTeAyTh4Rp/xFX/t4bRTir5L0lVFtWau3qdb3s5vdLG+jQXqwBE/g0wTt
gLB8ERrKGR0zvcJNdgPwhnjbpziWO9bTP7kD6oOe/nXTCGx8tvS56YVEkGOf0gSH/f0xowWAffeW
GSbGg89yJFgHgYCKbgvV9lFMW81f5XUJPmxF1FpQy5cmiEhQgWHhw1WH8NeTRR4I0Q2M0lVBbVDJ
8POvpSAX66ah2fcacJOXGRgxDDlbPdi0Tzw3Byu9PiPZWl0zx2vNFQPMZPIVX9u88tVdQnKgTwp3
e/VRbmGmMRaSyYiV8AQrgUG/8cCB73h9XnIse0vPm8AMTLsGSvFELe4qskUGqcllFW1UGUKws33b
g5fxdlLuhQiHaTs8Oj55l+lamFbFQdF7HpZwbMCQ7j14SLfJ/c/TNh6yBzN/c0CfB13BJ/AfVdH5
Tr9C6Io+xqCysSBXFJQKxvSKXXOW7JD64nDJg/V5d+Vjg101MD7RBGEscH4sT7Stg0zbwhfS6Gw2
XlQHJBrFwWY8YoLmIyHtmIkgLPYgvHsxotdx7obEe2nP4b9Vjnw4VTseV/CzjgyQN9SQnxpGhOmr
kDBEtAWGHrKkHVWBltDRQZEQX5LhTSifVNQ+CCuJeknOceCdJ+mXqvunU4zQ+YQO2bOcPGq2W1DF
z2ZbG1+D3yHm1JP0x27PltEpJfTl/TqX+hNVH9vcaho4CcG/odF5bC75pJof6byfBdQEoHScqcdM
phhgLh8+EfpWkGIQlkuHv7vBZjUb+2jj+paS71pCRCDVqiOXHC3JOjnD16/eQT7DKIWh4s3dLF8H
Mia+j+zt6tCsdWIsYllhetD9bWEzidrnkfM7/VTb/ZjTJRcWiGJIkHtfxiuc4UJhhLZjXq/QCXaI
kJ19CHIGCHZkch8SaTQpmKkefnraiEDsMbrV2FzTIJ41EM1IAmjgcJ44tDPetUDHet99XCYCqxa3
UkWUjYxvDGWzCANN4xaWH90l7nGZm3Kw832+zXKoztCBWPSfBy74lM4/rCWSViSTvEqCWz56UjHR
IMeCrMOEwLG0d04gSszCp+sLK5HPXHFNzt4bSnt7xuDti5yQyKOXkrJlq8QocEX/dw8AvYtpkb6x
VtGuQXQlMRwO5iDhc8wBJpshzKbzwptPh85BCyH3b4kmWCAZJ9I2lUVOt+/in5kvRWdD4s30hjLO
j7lN/11Kl9ZgRAtsfrWUmcCuO1eBZKrSlQilvH9zTwrzJ8rM4l9L7hLP3dwWrETtkuUrUBKzFYq+
sJfmS8La8OshayBYSxxM14yD0QUA1+j59nUUf6uhDpGFqglo7gjnOXD0nAuS47sYup8E8UWm2Wtr
PcCyz90sRYNzQwykdfrSlLshWZyRkTmTA8XTmnWOyiBf77L2QVSK/vGpx+H6klBoeSln0iV9JnUM
8+kqvlzZTQucIwEMZlCZ0x84DVk/xzoL2V0UrLS6n/vRiJ2De/r+id5uU+L1eNRrrdD4QsooW7RF
gtbUOsl4pvZgQQLSuw95MJ4ofpNQF+oTSMb7BVDUdxWPQbO4ZQeAFUxRGzGtlbkFOwDinNUt1m9K
Wz5z+n0jPOd9MC08Tuo5S546jBRnzju5zTMu59ikavPlgH1HcThVqYcp6ilQ7ZjpgXJhyFpF6QBm
Cikt4Vx8LV1Eo/r8UbDkjRhblN5wTFtlNjiQtvorxyYXdkcOGzbPCWAN7dlKRUg2PQaeHxnaAMZx
LzCht2QO9DBReev4cUaeOdWveDS4SdN9Pd/ga/tEXBI6Bm8BUUN96mGs3/Tiepzq2JYomvxzNBwI
stJC++VJj+POtZydiUH5uqlH7IrsZDAi2J1LVcUTHPjZc5a0h1fqaaUMzxgqmigFlrbtIWyOMOji
Kx+4tVz6NGE5K42Fn9RErN4Lr73fMCdZHCVhGDDW29i/zcSJ6SzeqAoFCqCTswgve+wQ+NNpQ0Ip
/XFKkhGhpCrrgHsjxgHtRHRaIRa0pcSWBfTL0Fy9JaR3V1xir8RjTEo6hCZ3056U5a6JK1T60gBG
aqxbQAEF1I2bl8gIRFm4ysYplIaPGuHSXMIGB7mVO9J/GVKXGxn9gzbdFLca/K5gHZvWvbonvumZ
+aQBfOhZRPIeMQSHg1Z7xCaEY0R0POi+tQdHp3DxSaKMFDMQUp6cBdU0FiqEZ5QKKbnRgKjxCery
PhvScVIew9evXSJqGBwEcpdyMDgP+WWd7qXNa6yVRn8/7xLi8vxpg1PYnI/Jn/0qr7vz1ozCbZp4
fs2oyPstgXOVdf6d2MYIW4lYxxPtaB9sTQd9UTWxKY5JxhfvwGnt100EYgsx22n9JsjR9qpmGS06
jGJvMEbEj52hmrtp2edNnAESlKv2HuaaFCWr6/EnaNq4iq0sS77sNKG8vW2eq+RALFFQD4xfy6DJ
ym1ITGP3Gl7ouIjFn+zLm+Exv1lLwgkpaPK6NeNr4kbuZExTygXrPt5AqgSHgpz1AGLiQdrzcUD6
1HUBCeT140U8kY9+0ymkq3SrfimancAG5PoEenhB5wxwWHKI+4OHv3ImtY/IGOK8zJXgPxoeFz+8
rFKmtVFlXJnQPSrCHDaZ5MM1GvE7RMBIvKu7v7BdWWlG+jX9MbqYaoYWU83Vgj6PGEVf8ArQaYHE
+Gr83W8u3mNBx66W2nCBviFMXRAxFcIP8U+gH6YjCmZPQT+5VAHUrPslRRKHJGD/jZkFTLzz4nQC
r93nCn3rVOw+6GnjYddrXikNr3eM7QWO6tr76wAFyY+cpXhdtUFQALVYUMYrw8So+lsp9BFsqgjQ
9Syvm6JcKCPw64ol8u2S2FVIhDrz/vlEIpBJ5yhfom5V8+h+Ezz7EVXP0rUsQjUi6NoGiEajQDEO
Db3GhAUbb6lqXq7VQ3qycWugDRHHWfwsuVUbvGSKR5tRfxOD0ydyehM1FV9Wa5nMT5aUUDLNZv5C
t8Lw2+ZSgBwFL7O4650eSYFt46yvFk1+7gw+cOhGonIMwgZ4eVUxdBsGEZltaoX3ndMBsORYdLxw
2rNUTKt8K+zW0jTFkQDmaahoN32YDVYbVM7KGidgVLjxoyJvNevmOuc+b+i3dR3eKc3CHNgJemEK
NCDXZxQoRhBfND6toXKREHBUHCS3AvhVD6uHV0hQX+mtQ7hsTTRAdyqObAxT/K3Ff7uLOJ4jxmdM
ah4mLfSnlwAb6cqQ3GLGP1AhFw0JHmRf7eRC6kAGKE8Z5YPo5cPLZPgi8RUmkJKZJG4xwFPnl5/2
AHJMlTajuJ3tA+8per9oTfvcaQ5NSjE21XyU1WNIVetLGd4d14YyqSZ0rp1ICgb6Dburzb574Sqy
ftGPUn5d5R1Ih0ZycjTqdUusVqtFELQv6JnQl64MxlUJF4UO9ZePamRcAN1hThXbYyukMp4Y9Prl
w+X7uLXpZdS7xBCu0AsoRZFquUyvcBEW21/iFabD4ciopoS6LEkrBhmG3KQWIZCu7AgpvYVGQnXA
zEbTV047Mx4apRDn5oL+1IEM5irvefSnN3r+cYxNy49ey7L8JeBixO4CFxHN3KCvjskxjbrHuFKv
7uB4hNIdQXUqCn54hEYbQwW+u2i3PsqQvgzYKfUdmpoK05K/LEWz/omlq6WsfctQGAvUWogdPcUd
NiGcxAUG4ego6+71U+vDoMOFZNIOYCPWgfPIYn+PGbPoXRPhrDi4LuEyYG2hjNN/pG+5KE/Z+1IC
XRRPnueyPhnD+okbsOccDoDMDzAVyyCoVcTPylYZ4ARZM9wvaq33y8RL9OjB0rd8Bea1Ep6iCIq3
94sSkutdjhTrX6fHBX0AOuK8YH/4geG+1xAhBKt4wPKDQGK6nUNrnVUS3V3KRnihzblu8KIiA43F
NS5EFefw5ZUVVw5rAYLh5MSfyb2Txr/MZUc+AJ2JRCUCbDDw/WQ5Zzk34qSo1KxPtW1RiIiWWwOk
a5hmVJFxOBSBLnoJOiGzZ8XDAbmr7BXZiJHqVEb7TY5gDIRm4jTNiu6dlK0feN9dv3DAMUMxcvRU
aIY9mPS8MtTxSD+b6phPYCtkWgewPTSlY6Qcar2GXmZY3y2/dJvmL9tSnWYpC+gBjD0rfCCT6k27
A46DmuWFqRWnvChrg4DUY94ZeGMX3xvrfjfZQnG5qU2mEvIKfQdwJM7fSm6ihrNdelzBAc3Lhzkq
Us5+4reX9yzTMecGKcJBAxzdrpVL+DNUMsQ6G2pfESMsL3WPqARZ41SlkwQelKu1mHiYupzoKGVK
zAs1tv13y2qDJXspyZDLdaF7AbzktvusuQGEwuw9/BDLGJEY9t2H2QHvOpftWdXwzWkkC3nVPvAW
kwAkfTCaItGh8fpR3tU2mSImeX6nJMn/8j4UTnRQdBYjb0c6YPhqeVx6i+eCY7Giqhp+XJWOpUYv
fVntXeVlSkwHe0rSBI1ZR70VWKAeJsAuwUzWR0NDdzfBC50CEQSnEdniPGwNFHq8vMZtWi0AEWr0
h40FuyXYe8PLbOsW7E3mgubFzsZXT67ir4U4bH6tDTi6JrCgSaY3YK+Cmr0jVSm0CpZbYWo9tLXj
tT9G0U86g+oEj2fbDDgo+6dN8PoNMo3z+RfZHHu3rkc7pakb6+n5NuaqPO3lpAfXbVSRwECD8YKV
3ESBSzSDU9Qfbtu3j1kJVgMSaDGHkpKcv6GsYBHR21C02uB/MW2uoOv8YMSPCyfbxpr4rERC77ke
VxtgYE3Pvu+kyqZEPxO9DZO4dNFtTTLCyqvusMKApTiA2RmD1fOb8N/aPrTIvc7i1hiRsNMB+pAN
SsmVFdzjNSCoklTbD3WGcGwn5zuKqFpPhAoH/lhPmpiVlLVHhCIVXx/O8Sh2oTi4utGmpzlcxx4P
bm2Y1m9DNcgNkftOljj37dhPv2Pqk5TgYQvZ/1mzHSaiiqT8YdfXXIo9D2Eb4g+9TXudhDEQDLI3
GmtZULdELoF40x9j8T4cTCSWFewlt1ZzA1ignWVjchFvik6VsrMX2baqaPhZOb69rVzK2+vxqz8m
TQmiCB9BB/7wOxuCET+EgdcGWP/En+2ALnNVI18qYW7dFawbVx/rTBnS5pbwViQEsOCzEMUW6T5O
ZawuEwOqi4tF5ulEwj6tSfCtbl1ulvtUt69rBRYD9lhE4OBSVh8ULLSJO4ktvz7evfEoUeX3B0m/
GI1uZk1pVn2W/S3AmMQTSaLHqEmGPld2Uu+OWoNU9iBbjskppIdg0HBzgthP0INXZ6EonsT6OAIr
p5plZ+GQOl0Ttutitzh4oEuVDU+Hesn+F+EeyLIWAYWx5SxJL6Dz7yyWKVxDLDKQGuZ38O4rUBSk
sbDYior2WWkMX1PoC68v6u0XOxJNWp+OnMKzhWwxDz/KkGqHjwZX9/juPcGYT0hJ8Hh+7dZgW54k
bY7hLG/cxQ0/us/3xmrLgWJEp1iZ3RVnyVQOsGN3Oy0/K7GdmL41RXeSK67Q4xTlO6y8bGGRT0xu
3+uhKCKEz5v1S0gTJVmecw2fiqPeOoLeDpO1uJtB2e8DojuyD1NuqpoYowclUwHGpEboeNDfhqL3
wbs0EzFC7V5qumu58ZK0gWn1zmkTV9ftxr+0uopYOl+5LacigvxKFC2D55KTVCLskoR/0kPulBED
WMrvlIpM7Qw3+P7e57GcnMUBPJay0se9bDiPwpZsLYb7UQLs7gmIgxreRr7n4iLKOR7cVVIK5tAX
LeKJw7FI04i6Kg9hS072uc4zwj6dlMbfnAf0GGc25rLCuIVI6ZDnscLkGoOv8rWJqoazHIShJZxW
845Jz6wNit+5qRjS2J4wZKS+plcUC0ydPwO8dYTK9LCV4YZhDJ1Nfzav2DnnPJGkWH3wPj4R26uD
nRzb1bEagZ79c7cM3AGBnxpcAllWPI8lK5SheX7qaNX6oNd1APYP4dtswhT5emLmGapep0eS8ep0
gwrMo0flbsXOYD9sGt4wiPHmuw4HfFVWYnQyR0QcQdRorbhQ8NDB9NsHvIpzvd1lLhn499dmOPg8
sxkuUML6/i3oaQEaQu90kfmMmZM0/L0PV4I7bMftCbOVkDC8yMiakiPOwgOOPFqrS/JxOPDWZ1xw
HOR7Od4kVD2cSJlSLyLjPKVH/HH1TAZD6ZpVMvvHIE87kIY+tBz8MXLVLKEGiGY2kglIcANP1QIf
M8yt/h+GEswIlgMQkk0kEHZS2iClSTP4LUmX7kzr4Or2952iXrN6JsuST8fJDBdOKUpMGucPxFxk
OgOJWtRKxh5UVyZYFWSnFwnDvIFPLkrYlyIp1ACpGYgi2yRlveF3+Jp2n4Px6qmUNZocYOEmw9aV
Tbzgl5GuVAr8V5+U8or5lCyXsGwbDxSBS649o5JYkdIyBQagvqyrt2mvnMtSoYYBpdvF6lR1kYJJ
GTXZhP2zZYtS4hCYRvI6lpprsXfx/fS94zkrEExqdBu55wXsOZh6fYROda341Eeq+tNazCJah37q
RP61NcEmJ/YPZUUE09Qz6ph46VSTA6zkmgoih/UoMzYcjFbkB1Pild+YA839vBVsxuRkeVpR4kJv
Yv0a9rvgKpYY1cjaRfACzitNEz+RORyy2WHY67U1jV3HF8y2p7HC+HrcutDMZvWghXMMeaWrxWk9
1LcTklefU/4p6kSG0Wl1BzMT1+2BGpNvp+0dh7KSJ2Ibxa2Uaktyevz8rwSAdD2FpZbO6pRnfWns
rWdXyLrUsk2WjOP961uZAtuMJoPDUM3D7dnG68KNiURipwoSi04j5PVTAL1syo3n+SQwl5ZmU1ZR
DYmw9C6N+MSG6b1rjWq4bdk3FLfoY7JmtisGLpfKIO9tya/QfGHBiFnD1ZJ8eSSZDOSAk9azm4XF
ONnQqsNFoH4+hosct9ePBqIpTkFZdNZVNzFR6LcH2ZXQuxML3rNsUkOBtL7JXwZpVfrqJXDfpBY0
4t0H+QF2Qa6bCRSh+j8CWmf2IxyWw7gHp/zLCW/QzZ3iY87srRD54lxlc4t3H2TJ20FOncqYLQGL
WZthxij5HnuHcgXO1c0LkHpDl6D3bfcNkXfUM9T8j8st/huwHVJjl9WeqpJ2rw4JHxL6vDmg4r8i
v4xg2BS7a7ttJsPDUWaaXJi5ydVwoyf5jLwsMvCgZRrVnbJA1XBNph4nIuepz+QnaM+ot8itzEv1
2EzfdBGnVX/pe49FRMpyAbhzSH/8td7SB+exWbjRzo0u0w7is5WyIkwzXxKBlNpCW/Al+aFp0zU5
odIjBw+cIKtf5fqxcfLnUAWnDz4sjtHfRWGOA3R6uA7UVf2ZRz3O8ZY5GloOkMbXOBofHku1O7ZK
0btkjfOtI5A3BUeuYqCZv9tBKMsMFCLabikAYELd+NDfuYtDkyYdBSfzQJGscU/1WSJoSn1lgxs/
9lkEDrnKNR1U6WD1j6U6+30bhqp3Mi/0HWvPD9GS/BPLQAmJGN2vjXjxqpz/gbkCm+jtgP8C6E7N
LUVsqdtaLvPMJUeZjhYemDgkMM2375NZyRt+HjXmavI55l8oCYLZ7qtMxmGyK7FdhsxeuDX0sYM8
yZ+qk4JYWCAp/nYFhtz2a+zaTli6WhlS0ArwOYoAl9nziZDvsyW21jo9z+rOPuB9tyzTlD/MlFN9
fshNGSln1LCL7KKbfEjnxelMV69FMH2u28IxrA73pPXnO7A4f2jCc13MUS2qduFrQzZDhsYLkevP
rT+sY7izGKUY8maHsJ9WLAA4Q8n3X71ZbuwzrKt8lDW3JuaHgMbbIfMJFit6G98l3h2Z6GvfrSKo
hySCDelfmnXj3HvGUtFReVCFDll9YiCYg/ve9LEqfQ+R0gwJwrjm24PL3KPsVNHhHTJfzMCjoPl7
qzjy4pSHV3Ry0SVVnTggc1HScQEe85ukfX70Lm60N89XcPtaWhwUyuqdNpS2mn2HXROYU947IW/J
lVs8Q0eqGCGCqfGoe0BMpyVVehss/h+kmh1bOqiraDy2caB7Jc7dX3YmvQpBZjCE4nxCcViICdxr
R6ymuiV1wA5PyE7j1FtfFYEncKdpTd3y4CdgM+mWRnv/foVcBlAXnQQFRXebW/HIqBGcps9KOP6M
AWSGwLtXBneVogvDm1cEq4VLq9miPamksoHWd45O/nYE284uz88EvKxU5eCtmTpFSfWOAOEGrmZJ
ekFPHeq7UHciLhrrSJTsCVyCAS9EwWUvl5uUlbXw69RYyuno3jx+ZLf46GNcLdF2ykqEK3BEOA5n
vKqSzuePiYyZLMGv9w1Diz2zzHPMjS4HIrzYLLDHYYkaNHE+xCD38JFDBSZE+EhybxNz5LDBXrBm
/fVXuNkxV2KXuxvtIsb2nkmKmORZvV0fkYuXCEDHdbbOo4SWqnh2173zdku6ZeDYkan89qcaLxaT
NiOtH6Oivr5DU6PnftZ0jZqRp5qlFHplOIbnrbcqUE2I2nMIhnPfnaANILNIi8LmZLUfxzabffpL
oUestLH8KvTd0fNylNVdID5q6xo2cQ4gnqtlwdEeAOkIv4KMCyE0tpNkufqP2Zi8loZt1p7mV4XU
tFj8cBXdo8BwQwmhMH+zpgTwcDl5LI+sCCjGf8efNoQJBEVKUm8v8UyOYa+RB9HA8RgfIq5vK/Ih
2dxc4qzBRbjZSbEdKKQQXhWnZZ5ImWnbc4xM+/I6oL5E3Jt5oiDclmFnpZSQvIlbPXuJdslK2r7X
9JKaEFXZMwg1+0hFG8yuVF0O7xtFRSzRBZPHR/oBBa61NeKmodZRvHGOLwdqnggp/bZPyb4Jh00l
cTGNfACsb7E9zAI9N/Jfh5RhgWvx+D/mLr27s6sA5EH9oukUpuczHdw7T2YuEXuPcpK16+tb6bJv
TRKQXdfzYIlf6UZCxMJFE/Tsbt6LA6o7V0qDLKJ3mSD4zemoRTqCRGLBrZe8HoHkhqQxIYOpBflJ
JlEbWFArIvIKy3CGw5DbBE+IaH8RKr/YyTJC+mseHfX7JNz8CclCin/aR7uQ0ptNrmsaGuVqhBlv
N5ckkyFSvCcbAxGFY228C2xpBlfoFBLWLHfELMuLLUBY055aW+nz9Yxx4X+/3UMW/BIyytmoIn1x
Ghfqf+ECXWOMOjL89IQMz/YVfYvmMq/F9ugF7/Pgg4IqSJG47r/Z3B6J5L4ZaCLMnHwwmAr7hK7F
aq0mWPECb7B0bNbt2qQeJvsbwA+PnHVGXaeYbCdFD7lSrOhZa9qYWNfnoiRD48cIN9P2GkbQuTXz
VQfQ7ZvRW1cOJIOVYv1g4NqDcPRpm+v7Ulbhb9kkrkDSfhFSaZ1lLE749y7Mu+Fqux8MLJ19z7lq
kuZuH99BHhEKRWrmEjFIynO6klFQoozx6ck6aKSGdmfYHaIb6lQXf5YFFgJ6O0FfZujCV7hZdxeI
wcPS+GG+Xchrv2klO2o/nzLvR/mrqHZUN8/Bm9f1zv22YBNT4ENEAPCPfz31s7MbBPxDEdwe3dMC
UcpISG21wyiI7lxHXxIp0BcERr9fshotml1zkuL57HwTEpdG9daYSoFNxaRj6GEqxVUqLSP/lFtp
tMuP8rpoB1MNQlADOcXici715PqRs5uXSL6DVPQbWCBfkTZkWOzeIu0XVxVxpRLEYlbPhqbw+4xv
MvhMDWWAHvdwMKRqZW1hR61E1pc6gxXsb9+15CG4eML2fPaSHa8jw4958iw8NHfcAZNF00qDxxb3
f3tafNQ0lY30E8qmCzw4e8XtbqyuVYg0Z3lID1uQUPJkrv0vCFf94qEhuSspA5EGkeM29VCrfNfe
O0P3g261VDM3I6g+feTAR0E76q3dMi4i5ndMZDoYC2lDYoi29ARKfGGA93VO2km6R2J01ajShc+0
cAEwmThWPevUdYQn15LbF7HEFUivjCt032DNUktE39xKvk/f5KQ3WuV/o64/U8N1H1AgcJfjju7r
tw/uORtwt68AY2tsUTI7oUISudaYp3jmO37D+1WfdNq/OjyZEm/VFNiFrTRbrjqeOZGsBGN17GLc
43ZYLayLZFNgq8oPuZwCo5wabsJSnAyjzVabSMzUBud0yJNXcXrKFfxx1ig0Pkkk0+a6rFBzWv65
DB2jTBdsEBnAQp6GoVXquIE2eeL2vp7LROeEw5gja6oqk+6vLI8OC4mc56ET0Qw1348lJsZtxT5X
jF7h8TQPU0NWluJ0Y2pZvze94QhawoABLwPqmDgZQ2YsTRY+c4B1eOKlj+44w27Qv2WySz1hvo75
3yyD/QSbfFlc1ChToLNGaE0fDHIJyZjGdOHbozs6rPnrldwAxpHN1x6juNA9rseNJjG2MxVqoAzo
WqVV6+PoStzNEpZHmKvqkFVW13ytGruXovtXLCQ5tO3JnAp86f1tF4UThJWX3ieb6/KsacWUP1mJ
hBTv4wSM2SK7fHhVWCL9Wmmcai3zHD5XcIve88ccSWr4PSq8AOrrE8xz7mAUerDZdO+9ExQnbO2W
+AJJ0iIHCwqxLLX3MzmEefgDzuE2XoYDxu7liXnFQDFa7bf7NMfJLc64XH/jE3h4eaBqsag3k+yu
P+kCy5NHVMeST2VUzmoml+z1VvHF7Sy1F7HYeg0Z9K0jYUAZzIM7rYdv+15NnRIJylY35FVF0kZN
k3/mhrFfNpSmfmr1RR5Icw0PTQyeQpDh9dset0ud8VpRoZoqDBAjkc1nWDV5fT5tRCSgxNx14CfQ
w9XDsewMkazr7h3pGqsGboV3tI579vbLBawNMcb2rPjortWaL9mDz8EgPPU2sXJaZV8imXvSwElL
KXUIiA5kCWawQbkHPLQQtd0LxSD4HTAqX/jqQoj8WrI4Q5tjs6/7h88EHE2zh83Nk2dbSIvNLIrQ
LCmqvnpd/g0eAjep+aV3XRhNjvJQeWzZqgZZaQ6EqZizfTyFHHlP6/A2qJHhycery8efmWUIaSOS
/yXpPe4VbB4Kbkr6i8hdox+W+q5nMK3n8hTo0CR+mGYBFVs0znBIfqqhobXunKmxtPrvhGJ3R9xF
vave7dWSJeahmvVmIEU4ije8sWVy0ZSHg/QUlcEKCdX/esJYPVDM+VbGQJILEofpgVHXR/YXDC2S
4/jakRzVofhxrj1zHQ3usrRkaDEjzfC19cxStCiMgOrp8+bZLZOXNDL9ZjP3F7oJAvWkxT92tyFn
i9qRb11gIVUBzlqhiiAs28Mefz3sYPPMElHyjetevLeH9gbhYJOHdB8RvRPeRPiHmKwJu1/1D5GP
RFIQcBBDl8DK8CU2FU/KKOZfPpIwZ2k9IkptPs9rRLv/hACOEp3+upstS7p2DBbUOerYba9O/vWZ
JCUBarBCcRGO5iqJ4bvrroJyCq5NxCfQJuaMPki0y03DbZFe+U631bFAM++hAH0f4jFS4u3DZuW1
wuGUlSIVJNooNHvKpyPTUkTRa9fKWD1yge6pGt5/jwVqtT+AHOl+olPsLnOB2OxLN06N1jnexxmA
xU0ZGGDqEM5xGnkbnKAM5/GEkIyzppNAsK9uyyUv9wN8JIDBELgSeUEn5JlNY859AenlurJNBLbM
Q5KO9g4KUMn89OkXwYLRtpaiCTfh0YXO4wzRQ4Q5G8BCEUBhKGC6EQqL1zLay7WiYbmBkGBVo6Ex
9lya4/RJayitOz/huBNGbQsMnRSo49G6wJRKKW0ij6JP845cyzNU26r8f+FTkPYn1OpytcbHTyCI
r0sHRu3oas2wd3iyBRimHMCJM5sipgHZbdg8ioFARP5xOSITtbGMQeGrhYj6gzv7sj4GyDSvhuST
tItCIw4i/Q2RZzqXHraOpxgWTWHiW8ymqtq3DrW2ZxFCo+80jtMXI9DF+fQYZECr0IhEBBll8ihZ
S9NkXEPERA2AZCLv1fqbCS3b3M804Dx/5jBtYMY0OnCw5j9iwp5YA54KNuJ4HUn85gD+FX039J5m
Fbcr8of/KB22sbeWqeGfUh1YCEXIT9OO8B7BqBaxlap7oI/6PuIpT/j6p/8/S9zDvb4j6ZeN5psa
IYXNuJI65dT4GkWYok/y9w1cZ+xtgtiB6AAu6E3m+W2Db7hdCdTlePZB4NiEr4xR2Mi6bsBRkj7S
6fnZPa3hTdeKeoeNrhCBmsmuB6pIlE2wH2ykdlcAFTkJGuPkYUqOKgURzfLypd1PF+KbV3Q5GhiZ
zLEkivG7QGUOHOsY/kE2JMsSBjeAYaMpmc4fhXZsUhSbWDvnEh3yb5g9Xl5OV92zv/u1vEwmNNz9
Ujdn/Jk3lpDM1iUElrldpXDd2N+wv+3fFWRv7CQwHInO8potEPfvZXhflh5OOdfSsL1Sl1ffQYUu
r2W4nGllXqiLZ/ZbjxykcdKwa+aM9ydoO4Jk0G8PsljdiFtXwGj+c+nSkGuc2ErlAMixtDhv68kD
AOb4WNEqr6l7d6PjAEWUy2/Ne3rEN3agoRIE7cKf7oCclHBptdodYpaBmmDuXTOl21fxg8oUXsPw
4sdUkoLBiKNv7AK+7bx4xjPhJc9YYERGAbuhRO+j1nebqE/VMQWcSvM8weIpKs6XMj1Tp6L/vv0W
98oIWsbgvokC44FlTLXAEex1blb3jigR7LKABl4lXwd/fFUUOKJ+31smB759j/sjenX/4BRVlTJy
kQ+CvNSCgi4nmIqhsDcS6NqtXvWCf3L+MV+UEgFNTgrMh+41/aTU0o3Qt3JMgdW/3IqOhO8TifnN
QGMiYyTplyo/EXp32lX6J4517Oox1ytybsATXvBkTJp185d2lQz2yx31PlZQYcmvhkpcXHDd9xO3
9OlGX99FF/dfnF0nqzwaa8Tj8Sh+591ZkiJIrXMrTUzw8YN74OIFBNhWXYAuot3xP2L7rKuLF6uN
dxZF/KqyCrpfHSBohXIJN8qrI0YvFKeAeQgFtLdZ2AgLWCMAFrrDt7dwEqXaMo/4e7CBTYYWGe9Q
52c5YyITF0Fq8vqquRgT+RArdPj99OBlL3V7qUPNXECk7XqC6pB/GA5t/T6aGcxWgUOn0SHlJNGO
YM2UuGHyuFRJowaafr1CXuEVLyjV7bhwObgv95NvgmbjDUWvY17psmX6nfazmKT+R1G6ANDehnwr
r1MCX63G6ARWd9dnpvWEuSsrZ2n7YRyUIDOfPLlVgFkBxpQzdmZt98kwIMRc0ts4u+pNlCpEfCSU
oVhVzxVm5ZUB5vcK5wIk5WRwVR8Z/va64gSWZeoaCSfhi2h6VT8HuDyaniiXosyS2czrwDZw3mhT
OtDgKV5VaByXZMiq3RethoundyiWDhKIvOMEuig3L8CzCehZLUH0pf7rW8OFFzfMmlayO3b3i7nW
HOL9sEhZVE72aWk/DfkzYVSHUqb8eM0BUZZz/e21+LjWMtzd83Ep7MgwWPcUu58o0s0WGc01r0F6
JJsaUWGTnyOydmEX8mTFTDoGc1KkuB5FFVXlp7Xw8m8g3mv4kSbAGVZ6WrDs/GlP5JZ0hxwLc9EV
efI5U5h74C/3TmkinBSJ5EIVpa6P3Snar240nvPMbXZvQ7sDvhXzVNRriCHMeKyGrPgFErFTvuSq
/ueAA6nhx2YAj2iLHhk2jV13U6FV428SHEA8O3K6kz1ubFx7kZN7/849QIJvonPW6vF4c1bpBgYZ
qi6IE6DefE5nYcCDrNml/2iBRwncjZvdO8h1DR+/5IrzyjSfX/MErd673nbQkcqLhk8sdf6ufpGy
70+qNhFO/9WQAmI/lidir0oe3sQLJflnjix7R6KUhy4Yq+B3yclWa64kKdM6yJYLunYwyS/od7g7
uPTa63+cMDoI0W7V+NY1ZjqvRFEH4/fbph443NPPZsmeipbBdnIbFlTv5htEeo7j4qeTo3fQ5Hxy
rAn6KBWS/vk2r4hPuQ1HyTcHS6CqzbYCVkBkeosbOpq24ewjx821G7fi56xICKYZ/w0B+ifx1NEM
yYSpyY+Awjisf6q0yEdEm71TdssWHDsA4qXCZ3zUFPMZjvW+D3ACcG6qieXI6IrBUcdm4JPMq8sG
xgE9hpnNk1rXyVLMKmiPxCbhTP4zQ47fjPWBSGAZfG2k+yZLVJF3RbllD9y9DDvvQwjRgAFjYGyV
zGHtbDooxCcCaKQJnc/8uon1VU3oSp1IowTll0KTPJQLdCKNURECbL4a/0/XJSt2dlLEUqzyhHBv
oLF0J7uwLFdff9D4JY/MXOs53I9rqjT51S3WWhmz7pzTcsjyGh34WpWGrsiWg2ozKB4BubZ7hR+y
CA/yZkOlt9BR56Zr0EwfjTBe1GTW50rVMwPAOya3Yn/DpuwLHi9/4zpF0QEcqcZWeZzdKqQrBInL
+mN3Bttd79wNw0l3Uch+RceM9FKtb3GKIg+FRj7ODjBVV/FaHg1pq5MC40nJAi8kXtYcvSZEhm56
WJLgd8MovSUeddSgYT+0JBo11Vl0tWs4Pkv4lMiqSywzvkeWhXY1rUGZbbA8ONYJ47vubWqBtOhU
TTnB+Y8tbnL5ZOa3FExiaupGde0j7At6UVe2LvSx5RoZlE3PavtwCGc0lagFYUbmMr64X0beWM06
g5Khsd7ztRTPHupdeaV9CLWwcU+sgEXjFQ6ECUfcbCm0D8HkuTg3DUsR14/sIxG82ZUbyKF4BG05
5wmUzpSyCWXqXjULz5DNW8rCOu9xbWWHPlBBaY+p6CGtupt2KtmFC+IWN23yQg1+RFcVk514aDRS
z0Qf/itkNL2YOPwyecC9kqSiIMdBEKex+4G+0fJm4Z0RCmrcgRtGapxocFpO8N5CCYmPzbemk9Zp
1Icrgjlb8hYoceeUy7qN1dj4ZsOANC3QLGrxjOJ/iymwmPy44Xu2q0eB79hs6/iF0thBY0w4YLCe
PdHldGPHNa6cHsa44tv2qXL9s/RWG6UMtqPvvxuez9IWkvGCuM4+0UOxnFSrgNA0Nk3J4kyBJBO7
q4JOtX/WIdnmiU/DGkv6WOqenLQaI7LpLjbH8ulpYL4S0bpdQ/vM7SlnQtW+q96gMfYwV5eFThq3
jR0HCuGZDegt0B12Pm28SUVhhVPayZjuoRH+f6y1ZLE0ldjZazNe0rL8DIehZAKexXodnfHU3wEL
N/tHm7eZb7hIiZpqGeFELH5vA1xSRgTaRe+PNn10YP/F+p6lcjtWdLtteJ0eb5G0v/TnIxwiX+V0
atef7SRCbq69Nblbwnw4TT2fdNe5ljMkVlhCTlu2Xu9CWsHGo7wFibyCKVlIVnYAOidkO9yk3//q
3CXqOsAiARVstKefyDjAarAMghC3F0JGy8BCQLSSnUL23fI4lJ5nd7ElE7yIQKOzw9IE7/10PA4B
XTE9taLMivTxVufxVOYKlWNYBsx/o8y+zXh/+qBs2TRi0yFBYadeLbE+1+qe8wOP9maHMfF+7ozf
mjCzmOUlRKsVGIZ27SIrhufVwfsxPaWlA2tnncfo1Swv1Hnl3zNLHUdzQq54/e5JiqmPhNeqZRoR
ttNWGbZSJB+9f2QsNrFUMsFoEMj2G6k4fX8j2lg/IK/1QL+R+b50qrRcZyhzxHVxPDgJP4QMGHFF
vMlrbhwZCbIM8EM9mz0z1rVIe+O2Ww9auJewLd7Vpx3YgnH1pjDeu4QM6PUBBDPCZetjOuGXIqZE
c5V8ijgDgZL/VSB8Ht4TKbXF8VtISPfbS9u4XcebrGEwdBj6eIpyXJkLIDEVXqu4TfXaVKdBBXOG
v2aXvG4XVbtfC+RsjYbjY3V/12n8R1hq0fM8w4yRpQNiQOdNwkg4w1HDq57u+Gc8hqR0BwOwudtQ
XaweG4r2SV7+mWQG8JM6sd3TE/SNI2NIeC0fpAvnxxdxBKcO9KCxJtK6N2O+Fz0fL7GYNHW8pyys
7m2t6bYjGmdnrzcmcmBZSsdn1Q9YKCpZB3m8znBIQIAqcjTXthvQ/as2TVze+4BLzBL4EpozLUh6
TScVzkooMxA7cdf7G3dARAH+okv7YtohhdloWAdep3Bh6fNH7AdicbHi4IaYa65SroepAXurMwH6
1eE6kvANWFlcq3w8VfsgCzAHtc1TFSYXd9/8L1u/AjQjIOc8xK5f+EUTB07F8bA6M2yxDZXTOM/f
qXzCjZCpLT58YS46rMo8FnAyXpKUO9MclzJo7JAmKphtsMXpaCCRbY0NVJCReG1+ceL5XnkmmTHf
t0PYUgQ+wvZyHu5TRsPaofd2DhekviRLYaqY9CnoYw6lixI7VHVildbt2ubmd45EAB/HqF02bqi5
lfGsJwXC8z88ovXateoIELqdQFgTvfZtuUEtVC2VW4R1NpTd7ll8PDsigraxjA8r+8+PKnPSdfx9
VAFas2zBvBafdoy4qtbNX+XxgPsl0AUv5IUU31nUTh8X69aiE4ehK7ULSGA2QMzb+e7eFbvIo/eJ
zfAhwVnvosMJ73/CoWLlFYRYbyGGlGL7yC7xTTyKkQ+6gSX+1FlRJMbGBGWoiSsy88PGM8OS0beL
MSOCZvZvohQqbKSXKxggOyaE0tdtRbh78f2bnAnIYPDMIcPWtiaOg3pgkdW1whljTNRI972qb1q4
doUF4Iqv/FdqOoBmfXT+C+6eky7YJxpxKcY0W1nIjDWsqIWNkjbXMIMNi+LEuIPdA95YcxjQo8YZ
hURH1BnmAQ8dMBI3zllu+4NEQ0++1g/8DP0s3lJGaCRmpdwWNkWSk6X/dzD1Vk51QPFSPIHQGfZO
Bi5v99ckXj50XduGTFy0KL6HM8a01dL9sT6f0TjKFtVS6aV3++BI7tpd/KIChMHG7EHsKNLt8kCb
gKJngwx/Dfya4UmTVL7co3MM0tXnvSLiaASX10UCetgG+gUSmRNnnkflWAqS2EQpPQGmUd0ukcXw
qLj6FQ5tl5IR9nbrKQLne6M5ASim82rdm/HhliiN6+EjgggGwflvjqxeqUdqqFMDXoNuRmUxQ7rw
pSRTKhuXRblp2wpn+Deo0C7YLy6HHiD884PM/4wKTYCBe+A18tugOAbwred7FjAAMDDxbXsFKCcg
h9vjp5lr3aIGhsOIq/RO4Dhwc/3y67Kk3MFa/I2Jl/f8D0k+EXfO8DUOsxXJr4DUmfiAQHCcCLtk
ONsE8dp4gqNAB7HMRozkvliaw966jk33hG7MaTi0+xOzuQcqzm7/g8whTbbHC86VlTUVaV1BjxM0
1g1H0hMrXCC5u9yL/nM6MI/EJSZbxzsjf965JYjV1ryYeQc9XA0mTAswkQr/O+B8iJuwF1Mja3YA
eSazbbDyBsJNflsaknaaj2K/Bgh8cPXA68w5RSmztRCfdTZkTo/fOQJsY4jMsLz29Le/KJ8uetsB
mSmfM2zMmFfoTIZHPPFEMZ1PyPSZT7yP+XYoFRvabR0bg128WqeFvx0jLDl+f33L0BXLiRzlOOqo
kXrosHhEcAm5qY6xTDocvfP4enkTEOFjtuJySgOQtzZgUae/RZZwGz622D3+oIjSWDWnS4C2FuDf
gZn1b5VCfWxrkfz3S5ff5CQqOlgjGHz0IB3Odn01PBQe/9wHrpx1BGr5HcFhO1Z6tzqkvfp1Bqtb
AiJ6fA+6HajFS+qkjZ5jNDxZKPd3EnOY7SFZs0oONhmKBw8nnI/MxQ6DtHLlzXWGDDs5ym0n1vhQ
HlZf9q5PV6jvDWR52G6PZaXdNOOlaMBsmsV681HXU2NdpBakmCVjcoOs2U4Lw5334nbQTI5q5/wf
sEZkCNsojElCV+P8PBrIqMUuoTAii5V4ErvLx/ECLde1R5o85sAKUGoy2X2UC4EJAdGmz72kvOaR
iSgcJzJPOYLFNudT/SJ7ZPIG8E/oVyDW4nNkMRbgC+7Ai//xWblLcLBNFbBmDfFqjYyEeTA2wuZD
zNIeScdkSUFCCxW1+NoFky8soIu1fEuE23XPUj1ON4OG2M+Rw83YuVdFyNhFTEInk00rmWfDsob6
uQ7wVs+fY2F8iQqxQSnmN30yo2yv1fEiDsUYthnDBh60+TmMacvccuji1qHBeOtWOT/HRYLR119h
4L4zX7tZFzVqDug8xhD8Nc9NASGDx7elrnQXJNHpSaeGCSpQwYdbwePn6Q4/pgCkL3aMt/YEr/W6
xVe2pO31EWCXDNhpxmKd77I3m/hXqLZlwUkiesGFjAFilOVrsOnUR46v3pr2IbeWXbPYrIAmf6wz
XtokmKu6rPfdFWZROae6s8ebaR0uiA8d1kouKsiK8ozTfd979H4mwSStsY/oz1p6CNYr+5R0Eg9H
Z+4lV2VAHAalkQSHgn6oEuzs+0az6J7T27iwAVabp8vy7d4o6s5ocKYSA+hG0GPYm3mrfXT8qQbm
Gm/uSDR5nTAA8QLabJiQLjdgKbd2+DL+3tOKFmGEM5Y3tF3g8sMBq8xM9HXACUK2lF6uKM0EopoV
iPRTFbedkXHV+s8aaQwSo4tYlHuoIyg2BqIfVFikFfljE0DLqpLMliobhIEJQczB2iVWsx2B6xX8
XhpSikFFGBp0kyEh3Ks8YyqVnk7G4CYGiTfHi4n6DbMuJ+c4nJGswo/sYGj56n8kJzRTJ9qS0z1w
bSEiNR3d9nIqbAdm7FlkDPrVKSS1slxQM6DKxrMansn4+YhEl6BJOIjLb0OOiSaUo9IUpDsgAlob
rDaU3D601DrfotTh5YMTw2HvtAqIt/6BuWDmJJEkV+wSbwPi56x8mm+WL/FugYb7KEw0C28vkrGr
BWyasrpUn+lEtki7FVXyN5URcjeoAlr0CHFQrV/7zL+9lTAvfQ0Ep1Yd2ny0h3Gj0Cy9LIYC8fSp
VAhdur4WBnNybv/isJH6Tw1Ej0VzSaxcRoRPEnOCZikMzN7iSgNGYBMb/ZA3SKwzXrGhKb+talJH
u9vu39GBM6kMFVnhaIqRM5RKjsKcgrt6ETGWMhEN3M37VBTgXVVrEZX1f1lOpVubmSKwAFc1hvFw
OOU1tZ1R4mj7oWgYdkF8vfYvXhkdqP6IoMm88snk+cRBNn9xxdpAN/Pb/SZ0qgK3iYG68bGmL2ZF
PRsEZS5+8QOKiAgXCRgb86r2FvrvQm8vfMxNdqZlmgGvxAiltIXVDEnoBcjd2d8QDYJEtNgZdfJA
tCa13fN+TkPVYY56j+44299sDP6j8RuzGs7CVif23wTBANl9sR+RCtGJIP6ouD0rXCQNuFL+fQdq
4J2nCs5fTR3xjDiULnvtzxR6HYkKeTSa9NJL1hIZxsai8MjlZzWGOsvCxCJbvP171lj+5DsJyY0p
PObhbevZNtlV8MdyZilfEb88kxaczLnqS0wYEEROK899HkCmek/Z9djC7R7DzRDUZKST5/v6BPvE
kesb/ppIDhF4R1DTuatioGTN4OSGPuGqM7f6WD27oZSv0sxNthMyiDrwKAuXzCNnj4/sm493oq1U
umI5cJfMT835IdZXnlpFAkH58QnkHrzgL6iR1h1p43IPvDoBTpfTjl65yxxYwD8J0/Krv5hCrBIq
uzIGCA3FrTFpLszzOYDIyh9nfLRm8klhL2pJC2PuxsjHCM5O+X3+aK4KNk+8uC0W8pxhEsN00ooe
Q7egDMNjYipTTXmVtF+ujG2DHoXWxPZu/aM6C8v2mB4DnT8LeCF+LZr2qVPnZbJdfZ3wWbm5BmrC
HqO32eMywMH716YnJlRhSTMz4Zg3J2pPrHhMliK+Rr2MSEzDVm2XgxJGKjRffv04DsVw2WPEOiGK
6/n27cXXuKGv6v589m9Kz7VZQN8Fz1kIMPd47c5UU/w9QZ1xImv8eJRhveLv6pp5+mFpzdGnTMyZ
sDjQhDTyOjxDkruu0RWb3B8P14GikhJhejRsqpSU0WCEU1qQf4H2Ab5S2M2bVquIb4QqJXJo9hj1
Sk2TyNNCQs1GbAkT2TTTDOZ31K6vYRISB7AhLzNPEvvkpyGLd5Lclw6v16qmjh97yJljtl3/hM69
UHQJmRgklQZhtFo/wKSKiv6DzFSSB9Oy+SFC9/L8Wg2ebM8xzK8vAiUJsEXNl1UURJpP1veF+3KG
6zmk4wqmXWSh6ZiDDDFWdXXkv1H1KgXBkQAOIPqq/Z4kZTtT/GmFpbtS9RKVq+Y01M8evLl2iFV5
e0tRxJn0C0ALvf06ouZiOdKeosQcIkaydhtARUbFJ6cBPIZEvT10Dea/QQ2k080QKWyZstpYlB4e
8XGZaZ1tsi2zfbdy3lF1I8HKdo2i5WsVyMuP6b4qMEVuVW2HTzKHJZlqMfYF8NNBJmHywYCLOvm3
GcQ2UJi85D1eb9gIrd72BOtGe7qy8mC5F5DOFJrB0+JT5LUeCNa3w5LbAoVTTzAh2QCWgELx/e2+
BCF7wYKlnvlQwQ3tBnTFIYrMoJClXrkItM7mtjE9T0lDTPqkAvn8wnzUmcQgw3RM/OiegBdLXX+X
cShhXyBvet3N2FUNzZETRW5VXncNOldlnRQyOBuRWX83TpxqIh6Np6Wp15YJh/YGh/btfEU3KTQ3
mxE1JtrK5dpJqVnHlVSn4YiBQMrObtjDmDffUamJsjefIark65p8p9njOgMaGY7A4gZcXRnxODPG
XlhfoMIHaO+DnxO7o5ian69YFraz8HK79K/g7vMeQbJ+w7AGstE1JpquHmE/PcEBxZ6XJHhggF92
nUKRgPe4I/gq7CvER94bTwad29gAUEcos5FXADWehZ0MIBjuBEzEgQ9hmtgW1DMYyH9HcIgdT3m1
aXdMKxkBs42QFz0Wr/PqOV9Od/44oIq80nTUpI7qVGy6+sG2VI2GeylWsNmnZgaD2uhb3EuZJGpi
wHJgh3Go7tuMEN6cjYEp2ejdWcpQrUR75ZTGTzR6SfjDnY5DYxm/0bvllRRfVqAHL2zal3qmjp8i
s9K2XuwQoi+NxbE602grcz8wNvrZ8QVPXraHMkhnQVKQApE3GWpOuOjCgC4HfcKjG9rbw8kgFEDb
c6/dzYK5q48jqKWkeOVB4FJI53uyQPfQMaTQiwZ5dUnIoJk7vrOwA5GKy2+LrkT6rv0jM1L3/bOb
LQOI6hSoAM+fL68P8TCE/rtitQSha8BsB9KdmVhslRU6pHZ7QaIgBVIKQyZBCOC/aH/P5JJo/lUZ
iXtSMH4TafVPnmWqorYZqhf5g4Z0pgYfy0fElYbJXrBS1h9dElVzlvgk6Ym8F0NgYJv342NXIRd8
NRJkhs8UcYDW2v7j1K51NfyECHk34oN0YO2pYSuCWG0HZRK7uAY0Sjx6HZnfj1PfjQlCNOaQC2/L
zR3BqMNfttsPVSMg7nIOsAZKMMG/MEcxre4fD/1IKHfeICF9GGz+mXSYOGIhorOMDbqz8jGbLSMb
NpAb3//8g74Wc03mH2PE2rWm61vA/JNTwshrQX6ZsNeTN1hLYcBSgPXkrZ50g8kLUXQi/SsVoW2K
yEtLdtWyFjQXnq2H/ko32trXGqcQCRxdxzhes3/1sx/4S3cc7Qd6HmLUVqlqW37G00Yy9M/Jtqgb
auzCjkhkJwbOXWm/YCbYYEcNGdNcZoBGD70x9wI1PHzQQMzZt+wQxSlpbwShX5T4qqevGRTdhQHf
PnSjQWRsyr4/BJVSejZph6gi10aBultp1MxkVWFGBcn54QO79Ru/t5v3g9uSZY3i0pVpoYvxr0AI
9eN+oVEP8sx+ee7WqHOlRI/WPtxTjoGHyb+u5wM0dSu7+lbUq7vKhSZdqmEcC2dhPaw9IWKT5fEq
aNksSLEXIYsC+Dm2y1ZXQ7lo7ZG77h7DPpEsXjr1S2uVF/WTIGjBUhH8QUI/oFbg0hXWF9tYWbzx
bM88Q/f4aaiuDmBEewHZO+tcxxMngdy8iwp5fTfm6XS6ZVVBJEamXEVxZn3ApFwsGkYtvWWiZ/aG
IaAfB5Tmhl+NS15nyq5D14lcYWFJPiMqjIBNxztCAwnkl7It7GLybZdXfMpipsEsASAXuo4WiT7A
/EwUaLQV11KWTr3lwC+nOJrwIfMWR6GGmZlh/p11zWEOFN8es6k3dUKaldmFHG7lO3yq3CGaot+W
Y79SnxeIXR9fF/NLTd9qn4gd5swKuKqwX3GJXo5m+tnGBnraV6g8xlmYAJ7llkgkGwnQTcxJD5BD
mtsl9Ln7GEfgaR2Xh2OhD/cWFB4toKRSmpnN0EXz04pqWmDP0q9iTDH94tnr0tr+w+9TSX/JXx+P
ie86a3BnyhRmXp6POdqMqhB9uoeEGlK69jGi+1d27XkjAdKPDWYCdfMqIx3lR57SVw3u7J+G6JDA
3Na2Y1ohM4FMyLROGRZH0TBDpTF2CKLKBOvHPt2pL8SSrLoN255ORwxkt8FRtraO7n9/wHXEasOB
PnauCKYUtf4eyoME4BPEhV2yl9axo6b7MZulDSOKmoKlBrkUDSW/4p2hJGCyc9sWhiLUFGygK+Bu
0aIjiVr+lzUNm7Cr/VMpQo+ToI+Kw3ljDjo9Ig91oTotzJ0sndra2iZpEPjvzAixQ2h17Z5REUwM
LJ79PFLQN8ncsPbZoppiiDNwa+V4xZknwlrQP+Wsjc66Ec23ETxWjWXmGWKvgT4tzzkwKp/x7GQu
78hYRmW9pNBDfIxAL5UmNc8jWlHgXTiVo+FEpDjeaU0Qgpvzdog58QPT/rzl8sOEFaz4qwfo2uDB
ybTe8oLphWEjWuKNrRryIYTgHCrPqyf7wR57RXiIwVWjM+UvbRGJVJnJi4a4zMdr33nsE8FgPWfR
8PDYKjShAuWyfRZCvwmkjqMzx0bEac+dGKI+1gcW2VvWkllfSMT5l+WxRtDrGrf6zJcYhndZ1eJx
hq4Xf1k6shU+6+cnkMFOODyQzulJ7LSomrDdwgWgfzr8zhS2vDMWqgTBUpGEsFuYfL9tRIpMUJQL
NbhNfSttO2DoWb9ZWKb77a3dqooH8Fl5Io0gcEAQY+hjlap4k2A9X+qc1nbHTk35yjIOTwBabhEW
rDwhF7kr0CtGNhZMyuFCgG3aS8fR3UI9S1ohK+rGJm0UG7MUbHieRevsHLZKrde+lbgS89i1Eh59
7O6ZokFx2Qdui1zT7rrxuphFfnFX83A7GV0duCNciS8z4ELHcyTzePW3FlIAipTc8HSTFi7dbP7/
fHdlhlHGjglQyU9hfrmqoYuzdusNjMpIw3TajYNzhhR3bgiiPfqS7t/dTgBzgjzGJyHhYw5jalOo
T/MAeR/0xcmam5jod+xlc56wajaRzio6/Zb16tL+ijBLSW2Os67fyN88MRooE/OWG5pL3De0GsB2
dE+rzWV/2BQZw4g6osNQBX6OF9vlI9N2k/cP373mKzLxvJKWXKoJ01iXitJnRyvC41/65e2MN9Kj
Uqrp+khz4mGEDWOlglCRJmETP3wjxjzkHvTtvilZm4sAY7a1lgOC3obobjyxfd/6Xm9w7Fe2w6LH
gYcQOXBLa9TKMQuPhH3trg7uRtvyh3SRyj/XRxIVmS22JOgKSlYU1ekfR0X1M+WgL4LOEi7UlOcP
0/y2xnaKVnjjyxuffu2CF0ekZGYGVrC2UMojqHJ4uc+B8FO+boH/AuWqhfQVpFS4HRb9VNIYFiNl
Wop1+Vk5LqiUHtaBes6VAdRD4VxzUyxius2tmcEczGgzxf+UOX3b8+xEpUnBOJRlhwkGd5iXvYUk
W1qQ6uDI/dt1C6CdvBwfBPMbR71k7rJ+jkUY0TZ6YS5FQSs8HNy/zgotPPAy0fnhgswec7WcRLpx
qohHzqwetQztWoLBgHHX1G5v4KzY6U+CHPZ9fF6e7zcPbJxr/ydYtgco6sb7I2KLVXwpsPjHSJS4
mylA2fnWAyTqGYxOmmYM3Pe0IEt/5M+U7V8RsMJWLRh7R3qBF6i1fIKvl+qwzQhlu1xu08N0Omt2
fJo1lLnKB0K6CNbCdq1T6OShQbH+rmLzoVLxOOeZyAgw/X8cfwm3NAPQGuX0YG07u0s36tOa+rmK
F9D9/5thY4pDwhJc/bstjVWeYsHWqDM5g3of7Wm2pCAzVY1ek6X04WvGdKBC8Czjq+qyEB6b1IVb
aw9HFA1loCghxywW+LdDTXigQL31OO3cVkw0qiJRFLhLTD8Yw0AXtCIw8F+aOpHsTHlFOvC1xWfQ
dai+j4ylDga0RhZDJlO94bFnqgTWuPh0ZaGkpZxqxLBAQ4RIvbCLiZFyRp2ZORTjiKoDtPVMpoxo
Lj9dLlgQVkYpSpouBIC5ADF2jeTlsuTf+XoLgijfL+ENbgRz3MlX2t/ZVDYBLZWPJRpdweuWhloZ
2M5iXm7ulxSKA1Uxajgw08QJl3D6iYY4zZncVxMtaALbHJkgaQ1dZQM1muls5f4n564zOTurp0+F
/UF8jNvt5hpVSZpS0syqRe2NcPDzm6pUxSl0hS4ZMxHTrQT1DFo7yqMTa3LLQlhcYS8I9k2/jLcO
gAXQoZS3dPGtlkp+rCc3ONAswPL2ZT9Ikf+dTIDkuXvZ/RWxKpV6mqbp09qGBNmchCRqML9pQ29q
znhBdzjjvrLE0lZF6FUHzZHRcQ/S0vP4h0C9+HD57FYbRSKvqRsIqLk7nXpOFJtEX1nFUkhdw/xD
1r/HedJOQmgKbFlXr8V/fMBpN8LzjDwtXDCuaBhPPQ5F4gboFa/b5dMVf9rAFE8i6w8XX8pj9k5N
2lOjMy51096hrly66Qw8x6h//RPfFckOhwvlv9mWRf/LellEr9djGk3pN5ShM5rXaaZe3mAGQp+8
mhH81DTnblDNuYazAVuyAQuMs2WHzLCEe80doNRR2E/JG6MIhwE0Ed0YO9NFR5PIrlW++iC6mGux
jQYyPaB93zYibWi9hNfTe3vO8WjfIlmJvdAOdYlaILFT9/bRWawtKN4nnImLqpz9cd4oPtTG1tJ+
ACAIAT7epuyxMSYrU8U/W4JvdVz+xVO07R104y+wD3ci3xTiIw8sZR1xrIQHpiR2Eicdhx5Z1xmW
mh/lpSpOqvKJuRHtJh3AnwrJdSyGXaJE8fdlZYW1VgOWPHMEQ/MmAEuA6JryZjYTM2qlxNwNiVdd
MY6RSpyEYY3RLa/GTLTgr1mMGZIKx2wM7+ykPosgqD7Bxeca/I+0r51F4JoZLyD3dXSYhixBvoAv
7W63QCQtmMYfL6yqnTGWhtGNCTSbS1f579/Jv7fcPxQlHaEDekV0hStqkzf9+DEHGJ7OzrZkV8BA
g9DiPFJXQjoHcQh6wv1UhHWLvBvbsunGPIaqwazzeTJQ9PdQA5Kea0AqrZLGGsemzvXcVAgFG2wD
TpFNh250R5D0MPjUKXzsuaIWGth9Ti3JlAWo8G6BdHDJBjgBnm/gRCOacLoER+IkuoHidTeNXAMl
w1gm5OXcL5D3OjprXNCtvKZFDXYfWHCPl8ipJDPfDZSHnzRdf+bXhD5SSUJMkn6tbGyIvMqXS7au
mIoI/nRcBBkzs9STcCStIVwwtC0kooJShzO+y8fyuWCj3pjnSP5k+OIZxa/TlVmhmkaIe7PvqYFk
lhe9yT+B5brxqrjVu+IA1XCK8zbao/pK07alhC/Tgmo0dQKj1lzDEgNvhzjc2ams/z4otPwOXeoL
A/z8wi+sV5NtOA9hej1hM3bY5CDLbipnf3USoVTofzRwv7JzePK9nk4qJm7ts8mMN0USNnGuLfyo
NPTqMs4ZLdewoK3Co+v8+n8v3wZ9UE8LKLiw7rcYaXZ9GsaWm3mHvYdgYJoz1gPRcM0U3SKbrC0K
fp/TwpxfoSoG53YLXVMwi5uWV2jhLbdWq1cleoPxnsdQp7o9NJE41ZjjrggnK836ExT9ZT4DPzlM
wcYmjUQndRZywYF947uH+WxyQpRhdts7fEiq/30YVRWMDPmYYwjQp5aF7nQ/qDQKeArQ84ucxiIf
R0WpxqewL6ENjJPqMQv0Qg2c5vDfAdIebpD3LgdAA1Jx/TSt7bf1681eV8FtLMpoBajUk/ChDPsD
8ooUQzSS+6qgNP4qhgtQePgkFO6dgz3aXiAv5JAqmz4LG8M0HtFx+HmEsHJTZe9dL7qNVKp5I4UF
BfkOvHZE0bs9h476qWj7Q4pFfosj/uwfRNsxh5GaTsFb3LJNkzKT4SnYvtrdsoJUpoN6gIG6QtvC
laXw7Q/LViDIUjShnQSViHqSU1mc1+0D1w2BhU7jtOjEAz2EMzSRCIhciju4dWUkJ/s/w9Ou3KQW
1K904TQiHvJhpMlc2ycQ8j0Dsezayz/Q+v50mMRsMzT1Sl1j4aO+EluP77hNBk0kXlmfHo69j4rC
vz+3UMRf4mACUrLOum6xOqPnYHGsxbO4w8Aa47scz5upy/rzmaDcGXm9J11rgQrYcb8Q0Ybd6DON
hgszf7vP6m11hm8kIwmrDl9s78n286ib1SoJk3fvvTH62AkI8+USH5MiWRlCs4B+FljiG3O5faF4
FpPB3+LjAZZXxUAh+bjJGxcenSiIGrb5G8Ov6ACV9MVZia3r/nHVOy67wWjZLPdHs4XUZZNxEjQi
7nj+1YQ6c9kD4UpJFMKle9YLTmRCXpqS7EgXIPd7brC/r7yEyAP6aicv01ZbbEvaxsNqG9z8mi90
HHDAFF8V5wq46pqX3q7E7h2BsgHAZS6Egi0GwKjvZSZF9gcZ9ZNtKOm0JGb7LwAbhVKDkPfbFmU0
SZ2Lt6zPw/irtS8vnMgWWilzeuquXob7jRJGqrkFbczQW9N7+tZMESMawMjRKdjWvnbMl6hnIzr/
p4UZShbgq8widD0LBtLEvQ5lchFWRn3ikU3fiFeH7xAsOS0JPYUizMj9W3TESTi6Rr1D/dqtr9Vq
t7MD7D1LidI2Yb4UtnZxF7TOXmY8cyquB+L3aEGBZ5ZdI/h49MqJ9fE0vZvQclky/6EDHiBn61Fi
uEJBKFcX8xc2ncwEi7+gB9OhDFUFzjWomEuFb0PlHPS4fwaD7AenjUBWa56Z/2GTYsN3UtZhUtnm
PG8kJPcvqlzfFkrGw5NZ5k3y/yCelOthUtnNlgCKA9E3cIxVZue84xlBK3a64wYcBA5VuxzSexOs
hZKbhXoWMsYtylcYGk/Mfp/bSXJIruwiwLb25hx6pxYZ4ZNm2eFKLX0EpvG0VrRN24cooyR17pKZ
FAQOLfyAWlf+0JjEDD68uYbR3b9iwVk26yhraZh6StDfASr6ahRYZvPRvnHZKxEWGKcTqckr8W6D
wWXHRxR+ld5WlyFKsSJcdEl6HxWGLDpBpLSKNzuduiIGOC5Kn2BMj2m3hJnhjtlKtss3FG7KFCr+
qK5JGtqxetS5mQ/1dEr72Q4OsWZA/iWq1tI5hQMtJNlCjXm+2NHTpCBUr2ti84qMjgby513ojHvN
Zw/KyAwF4hAjPiijljNiEVo1pq+39UN2UyTClnlW9vutfu3jJCv81FcziejVa060epYkgvFPZGhH
LXDe0faoE/fnELMZmNB6ScbbSHXEDeDvzvVdCO3Q0Lzv/7dx5imn7fgEdrburNwpwSJvzHBVVfo1
6DaPNLQx+bNb2gZ29iv9feeRuvTfNekp9GuNT2/59xRc0d16CQbQSpq62yPrU1wU394d+injqQml
8Nso8ptWZd9VW1dx5fp9Z7skmgyJhXBkuC2ChpmQRJO1kD6VMjxPGFE2w1xS1u59k3BCHJOw5tEp
hoKBiDYKG1jqzwxdVodJXrK1Yiw9Ghbtfk8XwWL96tOGcAioRp9diXk6MBJFNb15nhsvp4Ocsm6K
TPj7PDT75tReetwZF+o7DYhWl+U3FRzoQfpxMwg6cwM9rzQMVkFhDxMcCt8AhQoAOpzmtyXHAlgU
dtZmsaXI3G854VfrK1ijZHnLSJyrKHbyZl1KPTaVSEefm8EMZYooDkRDmLDNCSdF3axB9NuF81aa
1MdfqQRH1MlYyG+kqq8dtcfJEPuB37W/10L5uRngnwxgeXqulgehTpWrKP+mibSOlGZuxNOW57jG
fYBMW8HzQPPwZZvXw/bL3c54+rZD054OFGzymvYQLr6NhhWqVvnFgng1LiE2/+FcQGnPz+R+MIaU
UYir841hWZjfBqtFMUgmf3QuQdq+UQ59SXAFxnO9hhN8ZwkhmBkDhYgH3rd9NobP60nO3qd1jgF5
KtYyylpyJJGwdhGREOLiv4cTy9gJC267Ki3gPFZO4Rqu1VSE6o9AAWZxgHdfUV2opxnVu+0NQPd/
T0CiYy2ABNz1A0IqOGqKoN7+5zWvXLSBiNuhtpIwZIJ281FVFLVcpIwRkHTQK/Kico2sGUOvRgOT
ZjbLRB5+fUEAx6np/rm6rry44INjetn+8Xa4Pxhw2pnTYvVyk6jgjdDQSUvVvO92Y0eY/8Md5uPv
y+fDRUwUUIQUYZj/CmRXK6mUTa/jrDw2yrEyMTGelJkc1xRv6PcSJ1kTIyt33rUAO0m+Bq4ai367
1eAkm5v9ddmEEkSbk+WAVNjK5zziyWHychzFebW3ZNY9obsfokoz41oMqLWkBzIftV7PAIEydjZy
sLPHHHjYEoJX95L2lt16NfPga6pMITD8rJuepzLed30gR75SmKrWFh4epXLWaHEC2IOKr3eOj+H2
Q9PCE4KIdDF0l7CA8sFJCDbYWpXDAEMZbt5EsDRfFSxRCE2JgvdO8JW+GavJZFx9or+y8TLtjUUO
2PTEJwZte8ITV/PXQ1ondUnj68EaRkG+KnFpI3NHCeOKGGquKpY5CtgTggfLCz1OUkN5/eaVU0U3
yymNgOiv1PFVuTjnnOpWleNJcgKw6FBymuet1JEso4Bcz8NDITG8OA0zYJdEJyHMXGxw+yOh/Ovm
nPD6uGFGQ1T3sT4GXq4fuasa0a3uDXmD5sAH/qzLpGJ3NGYFMp35OS43emi10+UeJ6jTho4IdrHb
h+/goFHzXv9xAqFDzuvOy2Z+A+aBRVJKax1zZdO9zdM/kNJQEDsWFvmaYHRh8H/dzNKd9deDJYWP
RoVSsmgc8iod6braPGcXbBMwG4mWk5623WAUzXoArydWp+BTQjuxaBWMuQTZ8Mg8O/zILoh4cvng
VKu77STyHw55CZx+3GH0uEz4OzwcSzvr+cCWyeHYKRlb71kKl71MF3wHS4DVzdOvRsWqwKPezUEX
g0BN48JtOawCMP1DkAMh4jCjzh5YJtNkJfxOrzRhiOXXRXchLwvepJ9b58dUL6IpnOMZavxQxYGz
rTEbr3kT3XkqaBu3efU9E+Km0jLICFQA+qXmm7Pmuf8/yHdtojhO6xZ9xsxWBSYRh03GF7X0OG9U
83fbLwtnlrX9O0u47kwZBn0lFvm5TLPNO8d9aVmas1iSmtKxHO7uJeSHjFI/JnH0P8OG2JYFb1aZ
5A28xxCC3p+Dr7MPb3fdZ1OqWpvwy4ci6I295ieFesZxF35OeP0pHsEmfpnnekFaNo76qC6tL6ej
Qi7qbGS/eKXxvlNlIOqxkCiPrg18NFN2pF4iM6NiO323KQH3V6LjYxK1oRI/fgGehYorDzLBA6S4
ztAzLn/C2kBAkC1aq0FlSceSZGP40tFNqGLqYswNkePcY096c2Or5x6ZrbdrXrIwo6h02x/5iqqd
6q+aEEAJqamtw2IzHM5wpb3rH/W8iPiq+KrWAG70/EK9c4tX81ejfOTUBOd8/R2r7uamy8E72CBn
xsqtcbDYx9OeON/0VnrQyVFeNxuo/HdUkkAFBYOvaymzUjHkKieUR50ztgh/4+pEp1caFPxVPtew
KGIsNMfQQvLocVGrjVwP42sWMcsbikjtvDXw46m8KYtSgPvoTs8BDbCx9dEvs2ncUmsrMUjx0edE
txoprY7RGfTDbbD2naOl8yejq8dWPj2Ymx+lwPYdJP1HMFR5QAAi8OKzjkS31wu8MHcSNSlRt0Jf
U/6+C4pmhw58RHCXiwGccdri7QqKwiMRYAijYhJ46KVo85BKUjTnM6FlrE/2efYHFc6BQMCRRxie
Y6CI8yT/gvsnh/ON4iTZVv/mRMsJnTgUgSUs/CmBhuB/kIBWtuHbVMEiqab6ZvI1veHUUgcLPyZ4
0siyVhPzSkYEQosiJkVy4hG9i4Gu+n7lJG0OzLvudlmtErWcBQFgLMLNYEEWxque7Dab+k5dFFoP
0WCdR1dwTML/k88oJ9juRAIrlRum7kjMQOXHY1WuKKXGkbmJN9QuZIE2YZHrBopZpU7DZNr5EMhW
uqRcHFMEgDPm8VyHhvzZyYH7uZhLSQbfP4lwjuJh6evxhGPNFsnzt+ofG3cbSXfYVooqzZdpudrR
CMHeuRtLmAc+rNxtcbHZtPiPCkBABltWWZOZ1b8N8n9wUKLFSU+LYRdvj6QbNTexgyFuzGN7BBpv
WPn3A1B1y7XYgJSjwqocOHzlLqhV/63RrgyKzoFsGmG/jVN/W1M/91zUggwrO7WE/sZUKTUGhuKU
fDWVmyEtATSt+SBby7rJM03WN/uZO7FD/t5xr36DI5EmzuVREszQRH5YaNX4h4rW2eiVI6IIasql
uN9CD4cIhosskUHmRr8hi4ZVfwFSoq1kAcnxS2o/G6qjXOLKbEB8aKVVbb8OpkWYQ4qkyIEHqErF
TjmjwZJlvPPMJRVDmvQpiwfRoo929mRepvx8k/Id+FkR28AcOvqrrCn6PrVFxpwWUx6xaZDI+Saj
UvmjBvpymiRZetw35RgDsftABcs/Gbf8+MRfCA5qfHyFfxm8NIA2wdd0vsk8LOAFsQe1pgC1xZ0/
wGll/FI1U0V9+vPeCq07f+zvjvYOtMaotlQN4GDYEw4q0Tbhq4I047oH+5fg50y8lcnHbKJZqWPr
E/CcLZmc9UoFvLBaTbLYax6N5JJYSgzmVzCj9aJMEjqy1wwCVrNotk8FQOBH7MV9XoQop3AXaPPm
G816Tv7Qk+bNCnVLzrm55ygE5IrwF0XdbgNvHqpoANOk7ecRvacwXfmbCofaZw23rLGnJK3T4sTo
VKIWvaIiXFc9xXG+JSoZIxe5C5qCxXFHa2C80UG3T68agqS0z+Z3kcynHBjVaDJKh+LQwDDfV8UH
l8ZpPDr7C6nVhLQFnaKmRUGTy0U+50zexj0/8oYdpnTzLKnlh3k6ZFreEbYPR+FlsZYXxqxQTwGr
5tMkf2R6hHwCigQbnSgxpllv8WCCXn2iExGRG/kr7eJVl7eb7fonKbCqi8tTS4+aRwlDOzK/d8cm
uSMP7mjEImZ/FJZaWVMiRU284wDXq8mfAFagH5k0/G0UTiAvCsRiMLybEqTssX8AnVpBhaNJ59AH
OVuCxyrsLPSA4SbLcKnO1xSarVIPjfN1TLQhtisCBc71LcHATK4IXKW0fPvyDn2ljm6AR2c3+Ytx
MqMUft35WqAK4i2Az5Rc31Da2QADkoPObnUz+xu0FDFVvgIZTx7+C23ifAEHBkP4rcfzpW7RiKA7
9o7CYp5BXxZjPyHEAwXw6YJW+CkDI+Y8/T0p54AHCohGmn3TAKtMr2EEs2VG2Rst1wSkn3p07Fd2
HmSIAFr7p+DHovKkyfQMLgngN80b8yJWky3uiCCdI2AQxd6Uy7DT7Y5QkpbLwCLEbD0O/8l5vrRP
LbUYU/T7Zs0t5IvJwmIPobrwPTDcndT818nQO5Cg2QNNaUGFJk/McmbWNJB3alGNfe00XS59HxPk
oEd28oZE+rGleHlPw3lrroFYKFW0f49nsTlTmCtaG2BB1lpab2rPf4sqzgmggsh7J7/cbmTYv39u
t+gPHevjrfYMnTfpf31K67tZsSmAvfVhM/3EVxK+MgOvVduI0KQvz0HGL2elD4510EvaAlWfp3cq
simTYq7j0A3PDGxOggpeBU44rttar8nd7rAijN9eUKG6bZ6FMet4R3le/gWAEmlFG1jOFTqxdvG1
EtNLUlL8y7uzCrRHfr13DzeYubevl7cPWj60TBoBQ9AJHp3hsx5dRhu0qj+75JHB9hXtdisT6UUr
jSospVTlW0svEGSPXBsqOTARgh0/LiebYAi08cmuh07CaQg/YvuOW0TpXhYQNjNicNrTUCi4KXoF
CWDO0xsBQL7XUNMU08i1OgjyYUBaI7Ml6QhfGmi5+aPgVPL7blYzGlJBZGaUIL3IxNvrXaAbvZMm
kz+0YICoRE/PKF4oAYcfhY1BMkjypkKd5v3B9yY2f+/20D7JC1w9F0FE3cMSYxjLHLw2qjOZRezm
ebZO0Wn5ouMJwzHKOYMvqKb+83EVqyFFq3JpLSXJrlkJWCXXNv/0PmZj9gAs+uysMEOuDcpCxj0B
nRw05z9J48G+lObrmeWdA0gwp3f5zAZQI+iV8yBKLXk8O9cptU5VuDKhHHtWI6vtmGldCAsjx4LX
daxzkBXeNZzJ/MVHPzQqkflrAlrPqW3JpTx4QdfB2thECM9s8Seki7Jfx8igB3zOSOw2Yo9LNnEH
JCLJtk56xD2yRKI2f86PCz1Paxe+M5EBa/0r1paiQSM6OW7qJSC4VZtFYypOq8wbKJAvuuCn6Ppp
efvgngV0sSwW7lP4It/wE+2zEDnTXeSdbNbt5PPjOegRBHrn0oh/WWn3w4wSt5fDq2qOuTtoMJtq
MjFCbOU92NXBSZb5XzqCkNnk4J+vBVqpR2LgwqgoWtKsXFyLprLRE3DTUOCzwCKvmjnxCaXfvkrS
ILxV4POlkESRWsiZ72uypWgAp+KQ2wmQkLyRTgu4alP2PkbnE89flFCs2XKSzqIl5stfk2+EMMob
SI90yslfShzcaOY0mTDx/dC+GoGDJ5l12lpInSDT844wy3dhopK44uDT6zFp4lzQHnVxhOdeqjBn
vXuhFz8zzlAmBg6WnhBsfVea/99W8Tmal4wSph77slbeyPByhH7DPNOI5ajEFIArusPowjnEFkT4
gGTAaZ0DrWrCF/EgY4gcEBUo7c7E2xiHC63zsdGE27hodumungRS410M8zTI9y0nHqkTvIJABfx6
nf+E42WkEJyFKo005wVE5tmgNQYvX/1iHqqm8FL3UAW8Wjb0mExGQ5/MF+ZiXQzp71+UWev1wAw3
kqFdMoThCT+Uqm7ExdV7dTLHZg1hm1OibGT7vN7uWdEB6V4LU8qv/rDku0w+KlmgZfAVVRY/9796
9zGzQmGdrLfGeUCHqc0HbeQNByblkWr0+V4v8k5mrwEu4pqO7u1Jy5816Vk8dXM/cdkvs5NmYvVB
q8koMAUhcKGS1+rZ/EphAk8R062Ww6U5QGD7HVU7FzDMfeOGb5/ttDjDTftq2Y9UCBzHxJ7VYPNs
tx1O5H51qDW5ze/pMcbczLv4YLRUNkBt32qS0HjwQcV7kzsFa219DhraDi88pnODH8oAU5O2V7Ed
eNJXk7d36LGwFxj0TTnZiZ3k4EGSOfaCDkYawHIlan/CeUcTAr6oSZ14ej+auVqJild7INO/Vn/K
Q1S+Mkph7gKh88taoC4jt7XHjPzxSNFid6IIaJuAFHXiXuraxtf7BhGVdnYpyp4Oze6GRTUcnQBR
Y7ka0RzdWQb6lVnzgQGurMcAGS3gkOfKnvEswuAxpCBzOEUmWv7KQQDRWVw0JbNJ00t2r0ys8lOp
++5X+swVS/wBb8E1t8MuO3zh8/ii5mQe9SAFNv6KdTeeE/hpvTAsTB0w+AVjFwLgXiWF3DDcK10l
Xgnn43u5yUPqXUAhC9t/8+T5Q1i2pTALuquaRn5eb51Ry8M/76t0YZtTmAnkKQb0deSBmh69+vW3
Yf9yoonto3IxU3r0j4L1O/X59mMONxVW8wtwEIPNVruvEg2kzGarLsmsLEkTWgdXjAiN29yLOvSm
mYMLZGO1zpV8ZDWLu3WpVAAvv9MnpjJ5kkAmroVagfa1x/j+Bfockt7u7b3sGrG3kPphhN595XAR
hBv2jzFSe4O01RwmJdIQ6CoxHAv3ciblmPK7F//yo9nIu1/CfHcEZ45tEJZf2toSRv12EwXWTPmf
LuqRyW73swBdkhnKm1Y5NvshuWhXa/e6NnxhnGGuFlMZujThdiI1M4DLtyAsi1p3T2R6KbnE9O9i
VvOYt+Li2Ufr08Dz6gcRTFS7cU07VTIJr5aYtd/d2ocPPcz1ZL3NeSroelYOO1xGn+rvv0NqL01S
sGg8kKby8vjdsWbEcmxo+PFb57ahcS6uCci/aSH//QTUHoB+CbDTvmKLYre7g933z0o+xGxeXWCC
c1mz5gfvtKB/o3CWs/JXIU1WAhlgt7HEpIBbIiTxb2djGfOmaMocNP0FIFj92I3sZtb1ZbU0iMjZ
rWEDgSKbgGQpLtBSon0/kTOFEPWUMypYGWQIgyyduCOgB08ClsVTEU/tb+4K/BmlCmt1LO4tGKt8
R/ELgREzWFO3SBIwDWbxllnvoI3gFVevSl2H8w+06znFnT//Vv1/0Gv15WAr4D+Dh3BSN/CNKwtS
ZJlv7SWlArRXI2klHMpsw75AJfrD8E/PRSJHOWa+ds6uOSLFOyW9ur6ZkDPlU/m3MdBrR8tQFu+h
tsmI1eOtt30aPT4R7C+qpXssEPIgqu44cdMCom2onrKakTQ118r+PMNFL76x/ewKYWRMnLdFMjAs
fxGHbqDgY54EwjkK7V/0/kd1jsOvdkoeX296nYIM4oM2dGiuNMkoT2T4p6hJJS+aZ+n3MD88Byr/
KbgAD8M1wTPmghiBamGfWErdbQK+Ipvz2tIqZjg47fXQchjC3J49Shro2lhmyr8qRUyZ1B3742bN
HbtYvbuk3NDJin1IkRfhWoKUF82t03Limmtk3g0HPutMva23AYe3usBuEFYODtSC7rlee1Mz2gPT
Getj3OsVCAlSJxSFA/VKD/yKnIXJo1Ws3D+eH8dDcJ2WWhCaxq/EoPoOHAFgg2djxaVdJVE3+NNh
gDWfE004U752tI4nkhSPZyguiNptVYQ7qr8OPBCCzoaXHFMswlR3V8e4T4oyf/sseHjfaHajdaX9
ZdaGWXgAfwDfLkhM507Sq/Yed1eVAQVFjl3EzClBVI5W+3QtZ3W6MzIv8LGDWUlHASiWOWFsKwOC
aqf0JtB0uqW9IEms97Poa2+H7yxFwwZmJzuMt63L9tllkGezARt5aARlHKXWTqJ1BOY+4sCQ4xdn
unpnsbcXn6UKeFIW8B4/5LeCY2TsEbjgHc6kmc9PelGPFsGntuJcLPeRqmYIErFVrRacRaYQHKCu
mCBdDU6mzKiLr9AAOPf1zfX8PUfdJgBHfnFTJe9nr4rvaC+X3y/gRPAAzvLMnQrq3iyCtIV6xHoH
V5dDzJoNqsf9ShpJrh9nhF+3vR1K3KgORBgQTNGaYFEcmE3Yor5nIODqCGMDlvBfvTdGI9fvxcJN
16yHWxwaGP3UVTFtDGExmFaPX8S2VaJzuXlQ3YvAZxogPkchiake8SX3qVnZTMZPhqpBqV6d/it3
6BUpYHteXxSOAmWX0m1Mn/6qzhEkzuyM3xqNNzmA4O8gb8kzyeedmb7E2Fw7sBa49HghmeEUKZp5
0rA9w3jOjESBHWFjSImZVIQdFrC8uwaOHQgI2Zat4xWGy2C0yy9KanlJ0wn9WfCo1AsGZyeh8qCO
VU8i6h+oBEljOORlidJ6pyN5FjQNQFXH+9BLpap5Y4Dcbtf4gZNnpzc4+YYi4dz4jSkIPTVYEXGz
9Lgqf3HbIZO6+74fZqYcb1+gnaXR5kdshMsDvZ7ADV2MTFVdlVX+2OVVd3bdmK4EJ7ivE5Z9jI9U
FIK8JFCglyWOcU/1tWkRmb6w80i+zE05a5pziwXtveBFgjVw+1WzLHa3EKhUNJzmHMBF0Jnzty6b
wY14E+9GFgLxxVAdqIkKo+pHlhERJBKA9+Ay8ALxL3itjkxI/R3pu//dwv6jEAfilI6fYne+UQFM
kjcTIqwIeTmcMhXMQ1o5s2hcgZPwAiBIyu6q9p9m6NY2/cdzMvI3IxYfEpeBoL7RXlbYiNsYBMLq
KrZsqQQL96EY8k98wqEWbJzZnZL+7bAA2ZM0B/Fx/uJVH5F28CtjxMBh+ac2+Okiw55RHV1T5Tu+
IHZzuoUYXXCvqSJbUY9cdZtpmFgm62eFfyWQ1zvP6xgTmwZ99BkXhfvwsafv8sgu1EUljGrHTDVT
egfnxocF0jyrExvruB3Rgba/Teekq5h581zkRPmaE+pxrFz/z/t1Ikv0tVCf0oCyKAB/QsQ1NNgL
zKpdMSyCAMel68xaLltd7fsGbLemEN+eroZ/8XWQ6Wx7+kDTKrmSR+cu/q4DGj6BQmNBvvdengbo
28Orz9mv/Yr4GCRdX6R361Cz7/m+24dp0K4RddM3KN7mAeL8PGVQnw7dZ5TSByS3kyaui//XTmNG
8gJOx7drzqiyacNTKgZ4ceAnfL90pOlRzE1bb4/tU5hpr6qVjV7gNW0Ez+L7wng+ogQu6fREy02/
DJtdYBfcbMuJNxnn9OJWWT1EaGaRNwEIltXAbrrgzMudLJTvngkzLfAnRUcb14as4wHdVhWk8NWc
pN3jEDg3wV3MUD7wZ3oGLAH5hLPIdZk8ld+ErkQyNjeDH96Ioal5ZvK14gucR6KLJl2OXSP0nHXP
jJmTgIm56FJmpa/Set682uNotMh4GfDIN5UwwkU5GS/HZU/5fSv2A0tyVfAFHAHoWmJxNMLy67uX
LTZpJa6Oq4j3jHRmiit4qpOzaKDW9OKL4pt6vR8UNd07WzIHEVMib99vhrong56mPTTNokU+kxOS
BrsxnH5tQxKqUlfxyALEdp3ElzT/HbPpLVvlo3r2Uqp3SRedEPa7uOEFSsmuWSfQP9JNhqqQYhX9
ILAosq7lcpfUtoptighU91nVnqhXOobvCF0Z/SZNqSYWQ3pgAF67rTEE3zHIV0yyj0gjDEtCwW11
0wwDWwgjUKRYLBLHwDEtnBRiNFnJEKZGUP/hgCmYrJlEvbpyjlThwe7Z1ig+axruX+EYY/P/g0pm
dw0UTLX3YP8j0QE0p/6nPxhRrplGIOKINUDi3tPomg4ULzq212tFt7nyvGQs/GGJzn1115bHkGvW
m2ZP8TdK2kg7EZQWjGnGKuMZRkxaME/DPeI4E8adpcidnYbYnw1z2cHRb/ZG/ATJ+UmQJ5bsrqZC
5f65Eyjd0XsZhdRWmzafYBDK8GhmoUiZIQeEnWSa2LYgOaRN3ssBbXY7hhsxIlfkrO5k9Tv2wEY/
etz/McYtVR93OkEHrnUiMi4BZSJgLTR0oeyaOMZsJ+Qsw6VQzfKJx4NLl0+FG6XbRLKvevlt1/tX
vKkcLrYQoSxAGFip9wU2fgFd0ODDB8K+Y/4o0Ew5WMKr0q+ZNDZ8ZX29E0F9C7Npd1uMBLo4Va5K
uXUanKusWZyZcmKO28I8T1dTddGuCbqtafnB+fFdBhPk2OkQrl/JyQyXuN2vdSflkPcTwz+KFZnm
K74KpjAWsjXYlMBuIVsGyPxm7zWdJIrBXCDl0jWjjcWtroJOxekYrLy+aWEGW82crlYWFuZwUoLt
WYjPNwjutfAHY1CxEiJw/knygGfbFYAb46ADbkl/0i+lmR/K3ZEOa7i/Ud8c5moK5A785Pk2EnP1
AOEkQdX4ZDigpQZ3Gq2uZM5KM0oNE4IMIFAc1eqDV5A3MWADJXHGanrlqpfjhtFkzlSgdTKmniLK
NCubQnuHdY01JQsFFmaPgn/TbImC4x2hPPAE+RO/0kpXkybROlekVR+XSYMPi/sohTZLuZEmS8I4
LMyqtL3GcdARbUiCV8dy4N0ZF6pfQktqvEtvw59AdId2PyLVohoW75iAcD/b8YyrJEH+yrqoeBkz
Lp2cKoOO1ddOPn5bAOUdwna2th1K9KbqDMHhobW2+UScIw6rTo2p9ZEgYAeaLiRJ5DTxp1uAuM7G
TcjQYNoIEKfoJvYWzGr0wJ0vbo9x3415NtGsxs65AkuNnvlp/732c6khb2XnPKElAtW6XjtOokoF
E6AmZMmt5dmxgY+HYgQPnlOr1g4QMJ2wum7I2wPc1Xm3bhS+1G+V1ZNRY6WnuUNzjkQYNBpbVHfk
3z//YqMEbmQ/4XE6FltI0uhUyhZdsNHfb1t8dIyhIzqEhaHj3FINWscjUmRYWcpqD+xJq+8K5iTO
H8/LAMx+m9bv1cv6/fPg+G+NYaLsy69RkwfAHdVFzIlvFyi6VNJK/sFlqW0vHj/TvmdG9Wrtj3O1
WkekYuVgUeUcIu4FWYQlGn5Di6jov427CLt8/9pJNjkhH/W6som4NkfJ5K+n9isOhd0x6nOiAVnm
xOJ2lGttkzX/P1UPipUw/tsBsv9x6YnZMus9pf/qfd+OaJQu7/OKebINmQGo3e3HWxN44uKKLeRK
UPtEZXwubda+qJdFO9xs+fPNFxKvhdr8CprcdXaA3m1eriTpiDxaoW/huYLnIvdYcLXL/4PgRh2p
o4Oscv0MDIxerk3Uh2AMNLZCr1OHBM88QbeTZdomp+3Dp40BY6/a3Imt30LqPSWtGhU3TXXUVSMR
rL63RanBKDxcteIFOMu9T2k079C23PYARcYLIg8U9rWmyp3G5rWA/tzDZ1m2/+yIiQGeqVYq+nz9
yT7oeMvAGTda1LyAdYFWvAQyPxMUDhttsYumARRkxtlRsEmNwZ5Rta8VygmpncIzOk/CTcuP8PIC
OhGy7yJPZpEEcWrKy37ApWoYJ3tjtuJdFS5jTcsD5GFUqO4CQ2LvGlfRFsqmiCDDJFkmJ+CABDuG
9XZKo4NmocshFQ97XYzoOjAri5d2D+nAr5QbTXopJCtATf8KN1PgU2hl3gSUhl3FZPBUvwJqqfb9
5A8wwhtqdnZdL08EVuQ0t5EXOvT4Gy/Ok4L+DatoHLUWGkJ49Zl4/55UXs4ZCWGOBimu7/jq/jV+
a3dIoQP25yLkZOFZBHo1z0/CxEzQ9/yOf3hwpQ9ieF6bg+SyJlO3w4jehi4Iw/sJlh1mOTGe2Lzo
WYhTMYGg6DTZlBugk/ED4BPw5+ioH2/vv9JAIt1iwDwthLcqr6Mal1iLXtfos0GX0ZSTu9IAxVc7
D/4/b9xp6M0T67Ut13hu7XSNDKor4M+/MbiJHfvPEJuV5B99qiO03vpR9y6EF6SP8nl/Ccqqd4KK
n6xYdvx8TWwFSYKv5RvxnTGH7JNfBgMyU+RlSb5YyQGxikdZhDpqsiFjhBP3kgobeP8/0Wvuw0rM
f5JdwPGkFUveKDOvd01iGrJtXRG1FXIAaOwL0TS/9b48aR5z978so0lO5ft8Yg/CVt/mBMbZcajk
PCfEz67n6D4+zJQHj6k2HUJguNgl8BTW+7WBRHY+9C70vc1ba+Q/wGdMzpJvcF4m8LCtVuG+l40a
V9Y/oGlwnTZv0v545/ZjMtF+0Y1T6H79uRnI+cj6iLC3Ek5111qJ1hVS1pO81riFROFFnJEIvPXc
6I9DF6IP+bTm28bkSKWvodFPw2SsJKb81xx0/V0nZLbbBX8YEmczLPlwixXO/yX+0fPaRIvq9Sdr
aL0dCssn5VaqcRTAYIIsVLEgQSj91W8UoFlv2XYnSFqSHMdLdxvP6xGm6gQGvO73gn4kcmgDLYdC
mVV+cOa7dVQEK8udcX452wNlOmCFVF5Wkri8wJ7wuPoRpl8lRxi/Ar3oZRPs3/pcW4Seqe8GndCf
gsbdJBKYuiAdLRi5Q4UDnSZjlvt1axR5z/S9Ds64ECb9hzujMivUW4FSlN1lvPaccxl6x74qUpLW
4kMmx65g/mJlgvc7vkCWfzmmYr5pY83qpI7ce9yfty/1/Zd52N/8bYZDd1LLZTTNvM1zVU4p+89j
vFqbTGj/8Ledjngz/NiOzMH4xWn1MMNj+4qyj1CeKZceF7JP07K3udECJl98p35jnZl/qbIJbmqT
5HeSbck4HR3wmxudGHuIPxdAEkTnVraA7WAD0Z8XSmbGhCbHQVk1sy9MRtmsnOKCUgSgoTm9H5vA
S46rAy0/tpeUxsAfjREzkGT0Bd/WUKdxSYm8VXhNK13+8qdUrOsq6n4F1grDq3IewraWBmJ+I2LL
NO0hf/mf09gFhVSvK9iEhssQq4xXapJqUPhoyXd90D8aA+IIt+ZlTAY410v/lLkG1Cr+ik7UGpLM
+CX+Hn6fZSMYWbSznTntBbuWnpTfXVAeLBCYINp3+tEp0rWtHJ+h+MQCSpYqjQXw3YmH+ENlK+HR
ZB1lJ91pC7Fy2fx1V9WOBh1gQeBN+XYVXU20CpgjcOL7qyaTXVCITWMYHLXd1n1ewohLuDU3B+hi
4FDasX2jOrDdCHI7Y99zmg0JObXV4jXbR7KwSskO/vXmQYOJFHToYhwp/sCEIyjvMiI8bMz2O1Ha
I+DulgU2r6hybRe3U2KFvNfan8gNCiWNOO5vrg+fH/u6kFrXvzZRk+gD9EVy1Gq0OlGEPzr2A0zM
ro09JatipAVpaaP6izQvtKy9dIKzOPXL5jMmNjV43wLqgH+5BcalMksQlzLgNHrgoUBAURrXs2TZ
Q7dN8sG4m0B2hjBr/lpMcy0t+8ZfukgkvdUK6GMQfOrkmlTklEweKDWkYNICOQVwH/jL1PLt9+04
3ETfECSZlAyrXNGZElTdhTy4DKw54w2+kaqNUtgUfB2Fb7SzsQblPuCTs+lKpVf7ED+W7EFKg2Hm
3vPykwu5eoweANzukBj3tRHPRTQCVJm/pzIPq9z/h99iSabcBxbqK7GkhbVNt8Rs6kKxyibMbKmK
p0BLdRpHRFLPqcnI3UDR/p16gYLDpX2GNjcub6q+xPWGsSY05w/Hnr8On0i+Fm1TZ/wPY6sMMjSr
J9Kov3etQRX4RuTQ2ywgYNpl3Gh84nTTBIrYSSIs2fUlO1p4Ypy5xIN2vOrNZ3tlXEoc3TcWf/HP
k5ZaMRJY4GOBNF6dJ4j5HoaSpMq4sQdvTvEEI7WVqQGwqvvpdN9zTvV73EIgeMOL+c5SuY8MG0X8
rYdDRIM9vxx3GYASSb3Ys2JVDyLYiv5Q2DcPbBqnZD/E1wMNZw1rPnoEAPTNPaKtFa5FL18Zw+7s
EXO6bgskvocP7P6Bj+m1473SnpeLF6bf5kVukX7mxgdhsa/Kf8eMT7HC9X1EFyEfJoy/iYmRaBeO
tFG1zrDBP8AnNJwxlwkVNnCUhyK0nyAvPnmh/yIw6G1ndWxbsudirrTu8npArVQrtZiItnE4PM6B
r5+eVIfXOXt2q+9LsZkrv7p4mWPq2eH/uWayh5kSnwcLj2b5m1NN/XBiYjGgKBnvuOhsOk341bEe
kGXf+6ZQZ2/BcHQpvWxtKpFwHO0kD3zIqfrUVqfduXwhqT+kXgckcqsiBPB8SjIaSVC5LXrF0wDY
XcVXT1urXkkv+d7UBDUQjHzx0ebkH5CeZef8QZ1BLFybnP5b954vd6zzppMtSFD/l1ewXeXL1wzS
B+CFnBdUeFR4OYZ4OSt6UrWEqzW4/I8/9pPzXgq1P/Z21XK/ndL0hCR0u4Fy/TmppTlOIJJO3jqr
WytdvgdBd1zN/Bz99JKMl+Kq6c2KYGpGkXjM3Ln+5gG7VctRaLpfFUC4fWLxXUYMNDZzDMoPDzEs
ycKskOwCMI+sy3ISObAtjJts+3tIN59amlsUIYVBc2dR9+xWaYu0PLJrT4DcYUP3iu/iaPlUCGRO
oYsHRQy6w+OzNoJfFltTUsDSgW8PiFObtggjYcujmkKVgFcg6Ep7TivhhuUmGkORcmYwF8UJGP+h
swALhTOlFye2LSIDK3BthS4kWfS/BdFj79+TEOidszSERofQZYrltNHyraXY//DRGwXqIwBcTQ9m
BFSRurojvR/qL+3Ofn3A8xQYkqHkYh6PxhqvL7afdDNs3Ky3cnD16JSQZU6druh/niyvd3HagNGx
FaBW8wR/EHVejXm1VSR/sFA5pzdWJ1eOHixHRt4RXO5c7d9+5BiH4yHGm3+RiVnUZ0mJuq0qa4T6
j/QBznA142iCZp2x5NJYFFGo9B5/SNPlvTlxiCXsUwlVbvsSyqI/HqNsFDkwjmcprt01WI+ww0vy
VKi97xBtOUt+ctFOf0EMqBFxOFOgd5JkUb4gpnkgwALBjJyKLBBvALZ/jmMe23iZxVnmiSrJh1Pj
Vazwb8PItuujzE5AzaBbfhGgdRAeTJyYjPgd2WBcjq/QtuM/KIBP++n3taf5n6INorgWVu9OOgVt
3b3Rp/3uHT4auKf6UY7OylgVJe6cuvvUvWVN98HV1bok3dSyt4eDL/EhgfQVh7YNWiHC4sXmZdF5
nBfc/g49emLG0yIryrHSdHZHSVuQZbKM9/xvUc3FxWn4cNVxpFV0kC0pLBQqwl1s+rBJcnAFy3/d
gcv8RuVxbMJ0r2v/oLkg0pEAH/V5ehm018ftum+hjjGMVShaN/OJecmuCPQ5XexYmtHx3gOq1RY1
IyhVPClGSmGjeqwitVVtReSZR7eCCDE2uIQQQmmJqoQGEFxOntI5JwU9/yk5IGzvhvHvGhCNV4G1
s2wwkHeYmJGxyK+JMJN9wWH1CGBZrBJZryMfr/5wmdnPgMl4/x00YXT5OhZu7iCMsQaHNtp2VsJi
d+yg/Pj60TuK/m1K7bmnjqFL7OcEXWkFjK7xCN7ytmbiNfovksGvJP6Uvn+1OuzJ+Jb8Of5BHhPc
PoEoSHOzZa1vbaWzpn9HgWdmOINq4Alzqg0gwcrvmVGKXetK4tJZdnrInckWktHaJOeFHvz0Pxza
Re0pKdlw2Wfw8sEl7pFGzvwB68YmVkBOGtWZkhvu7UaKL1Zw51/bkTuuNjshTK6qE1WDACW+bHdF
LF4BOaNaXFRiz6qQ7gvnVaiigSfx9ZnAQJFOFboG8xebOg1SRiMssUV2yaukFaKE640S8+3c+bax
bz6wFdSbnLc8ywrw7CH39Jcamw/E9It1WSc3Pk5Aa5ImmOpg92FhUif7pQzkryM6y3OXYrCvWpVq
xwNhnwJpBpawsSK+wS2xGKWrWDJFKHRd4lgb89xkbQt3G64WVqIyk1WfsJ0BYxY082tqaOBtKmDq
VQtSDQmQIjIGEhSk/HO4tcVP1bq1HWssgFN/E33dLFWx8cezvK6JMUtD0G9Qv524QW1Pb+H+fzOH
8AsMtQ84CBj36rF0aaJ0eurFIzYr/pLvJXgvGjLc1pe1RXIg5Bx05+sFmtKp/WuYIZLcWlnKL+Pq
u9OzltJuzQoxgb4Wm00wJR8AVVG1MzI4RSFJouE6i3MIlQUy904Ck7lYIyYFn9jlS5nLyQLLeS7X
+dg7A0yq8Xjv1kosLKgAwtQyOoNEm7ZYEa0X7y3aM6HfyuUKnbF0ClQLJpNAA+ari1FPvIGCE0KD
TkRY5CtB1u4cOWfOTOPkNdeihXHs8s9RKARP36XOOqI8+GDdKfLNyy9TbU0FupiFfHz3baOZGfw2
Am5L69BPWBJz0qAcr24H4Lq8e1Hu5cbFLDK9OGzT5i91ENmO/fvwJUjbqJpAtZW/UK9MEuzjjQFz
gbpw7HJtJzIag2KqtlI0iBa0vrIxbJiZVEoMg6UiRPTchb30/MmG2TPYTtAthRaI3Ds6WS50NK/j
88V1bqK/agie046D9EPbwjiMeS6KIonfeZDMJxxtRe884ptl2rPEYWSUHh6T/mx6Rc1CDRtOuYtl
x1eD52NKu03mkKVCS7W6SRENczuVIplKngal6VQjOTDYu+yjhuPAvPzqfejPjVNAOU8z7+zWhxDn
PF2ahtr3aEIcUYijvPE3LpN07z5evWHS6frhcwYRu8M/2Plts8RCJRJ+yStPYcwic4pWiSd1MjKl
uyQo49id/wCzUMLqaPv6KDm6mHoLm2Dv5vDlrcMzgaHW60leNXJkBZRCxPbtoimGexD+vRvEKTa6
LxJcd6l5FqvgbYZk5q8NmKpD0WmGE2s6qFQepLFxA9nNp5D1Khy8F+/cwRHJu/7xwcRfmDth4r1e
w74yAfjEimN4EnV0qFqUG79nZIvGCcKdCEP996w/ju27YFK5YM8rNFQWfkEmRPCOs/GqOPRM6Rm9
8ZcASGeYKz8NpwaINAkxYDfQ9xqOENzLCoQq7xyAC79ZoA358k8fhGad9dDzcobWtHasoartuScL
c6GTXDj0x3GWxm736qZkvKHHp9U737RDRmYJ7+ajzsr/+CurFo0ebSvmxbcxsJUEwpNxxaMV36/n
1BecbdnKsvG1QK1RVhNI6fRJAJEoTFbFcxMFmHjaCUuYZJ6Rj6Awi7twHVyCGPSaVOoFrlLQo8t9
lNleVl6C73xAOj3/EZaxzyb9iXRAhyqiYTc0wMStCawDBjNe+ncFK9lc76roCHotz7ABQTS+1mXN
CW2fXePq1NZMfgqKsOLSfQSvBioTvuGwGYGbXxai9oWAoEt7N1N3Y/EFbzLFr6V6pKUK8rJZQf7T
WeqtdSuO2rAqzXr9lo/sSI49C0RzFW9vqKrNmRfdFNorK8MKP7PZd9UEFyI7al6xYl0ffvmeEo6E
vAvOVz9x7auWq280J+LsD12+35byjyDvdUQT0zBV4MayQsFN/BUWJ2CvGEipRvIjdjVNr2785EBK
MK+RwDMcLavv+5ugCdmz9y7fn4ruNjzpQ/09aTgS/vK2g57Q5e3+sx/dRivD1JG/RuXcMHA0RQ5P
6feJC++sTqcVgdoZlResXOV4BVqr5yKKgpKc17L7q1dttD8LLpkBgXp1XS7DSATEwJ37C31L3MIP
jmHubxCt/JRyAR/kK/w3sUqsriY/eZFEgV+zWugdeOyJ8jRGXZh5oefg2ktkjIJj2s1YZnqYqZ4p
3h+TFQgiKSijw2PMp/tFm+6UrjsCKNwbzQI0IJBaMR/d4pfV4E1Oi3BdlxDS6DWlnQcCKvNummuc
ER/8fxZd/CaIbD+Dk5aSYphmcHgsRwy1gECxlB6gYTzhx0o/gdOxi5HtwK3aBcmgtl5Krp5Xl4qN
UyT6yhZ7qjTNzW7E5AuZi2Ibz2Nh+eAmGd0ylWHfIUmZgexwVvT6qhr8suYg44tIMCTcuO500UKA
wVXwyYSWsTLR/ct38Z3jAfGqD7Y8aBAfQrf8NsdJwed6p3iK3KzgqdFrDcb5F2aj9fLosI7YD8bX
VvHQRVfoKEcpnWeap7adhqYM8I8YVhBCesGkYNp6DeKrfjdwC83Fq47fC3//u7WBpvfGycUqbano
Y+TFN/5ELVTZS8poYeF7Io8r/GWbk4soHGatYv+cTsrfw3Pl+3JomxEbe7lt1VFsEuem8Mmmkb50
jZfNBXyOB6lH6L4UvLY6wboKDEMROW+eAbeNpVKemTjwvDk0EwZwcpnklhe7D3SNMnoI2K+LQoGy
uHagoPCc8yQN+Oxb/lxzvf0bAx4QkdQXNvxofBs3R/11Bmleg5x+xs9vMrTIOEXK70PvJmRFMBKT
Rr3jVZegI2dYQjOjbfwK8KEvWGzqSDiNw/45eIOX2HXA3mZ18FN0KHH9bhV/kAuoUDKAAHjmBL09
m7/aQtpfpD6zzAjJXj4jbN4sHEprr/+uOlqWtNBzwWcz1iLXv+I4TcIYY4Vh+rTH8seTSi01OH3U
XWy+XMjMBKCNYixnYNV5yd/Rs8BqAFhPl1201W++PrrXM6mfiWc5b+S8RzsG6I7NqgZEz12aJGyS
VBOV/5t0N6ci3fs7o/3LweA5efGKoGp4GcTJIZZT8oWrwWEnXm7hJ8SzLow5Me+tzwNyKDcSazwi
JDP2+HDoCoEeGJHWEZ6Eyuep3pMiaf0EN92uUSvP2kxYzAyIdnYRp1XRoAsM5sUhMYtJhV4V+bFo
0Qz2aq+rIamX1jS4G5qPEekzN3npI4MutOHgboMHStCiK1q2KVEd0ZYu7Mw1pCtaXr9AmEHkuNpT
scJy6y65/s2cUu6siFCcb8MlGsz+GVfc0o8YH4/MT9e5delSEY+s8ZluTNKhYBpBEZ9ZdvKOc92g
6/wqzIb7szF7j/GVFil+ZRqBHtRO2fa1E6pHy5xlnCgf5MIZNK8HdN5sa5ApSwbwKiP90vQLgMMy
vZWzMqPunE/LLAtAuzv2/Rdzveq9KeCLYVXqEm/ymUl8/E6kt+XwYrUvheJTaoBp3MqeNaRSsVX9
TIlBk8KthxSYZbPxHRvGms5ZSGaaHSpJc1ugsLbC29UOhrCMioH42RLCmq/LGN4m3Z1qNiCRJq0v
6+dp06ybkayptwE7kzPJ8b0K3Rpm0LosyzaDt6Icip6dluQ/xuCYgm4VnGORAdcXszxiwoEozUeG
euF4V0dTFzyRxWwSR5izVgVfIZpe+wdISziwONZWayGjFRcP++tkD3qYlG8Ln5lN74TYJBIMBxEl
Gwuh46OV0o2+IDsJve8aBo4h6fdm7VhNlIy15KGDe2r6FYAfmoqRgCJbqELqwfMO5oyrk5cblvTa
HuLGGnr5p//PMyl9zMVNZj4uhFWNgJ+/uodjBBZZvba+WqI+e/wAxAlYM+QoBNgCJ9ppgAQRi9C0
9oXmdSevDr/qex8j4R1yURA+M0CaMR/gWJGZNhI2g6utsOIST4MM3Ie13vckXQnZIsh4GjPK+K/V
X03V2bc4vVZDnhcGMoUvl7H4XvD3fs6RkoS2wK6mbea+xutDiitCHxwWjHIwNG2N7yojImZbzg1N
ZtYQilJEOMa5lgAqzfPNKhG6xLkIT5lI3K0/wt8WT7xY7IuacLvXMbCLDOHzyE+GQmgv5Jn0qWc8
BNXNF8gPKF5K/KnphrjlNeODSQtXiGE+8Rq6bK/F1Tx/k6vljjhRPvMlyIAPcy6VbSrAJPAjkL8Z
PlkJeZvvsLWbgSxUuXayf+xSDHs6glOh9AZxfkhBnQ6BYCQruE22TCVJQWOlXbHgjyO+kFoi7lyy
IZFS5ZFJjdvwzXbnUixRvtJzjSRXV7MP/5oAuf+fRW56yz4ZECTT9hwd6Owqtku/k1mmXSgsR9+D
3ldpGUAGAnR2gPNd5n3FjuuUH6VQW9c8wT8DJCRFQbgl3lczWVxSyxC0rv6iDBAaqa1uC/J1+aSA
6EvXP3XgT1D49F+tfVSC69QO75Dkn5qERq7efzvqZ/WvRvFHjbRZfFCearjDHslQSklfxmgz5/gm
nJ34cc6BkoPIoeYhGsW48YkDNRLzvsjl4SmOw8kj6WRqsWRmOQcYqg13AR1/AFSsmWrAd+dmAV3w
gVRme+TgEkT83Vv56nPCaz1AvRL6jX900FrMlAwsK342DOyQN0r6s1Eq8iHsG1rG4fdkkQvvPEeH
wpmSfpyUHi85fmKb6ioVo5hblJyg30eQIBol4bzzHDlJ/jcF0s2PO9LbDirMjF/x6XH3En7XnL6q
U2V1CHO0wMBhtJUHHtZgAclxlACBEm4fAKsGG/tvEzfwL3EfZAqg8faCAsEiThmh7XAhOt2l4Af8
TgAD3Nkw4BOgjNa/8o061Rs0pMVzE4+f8YhL+MeHWWmjH+FgNvAh9hlW9hw3eoEQctyqaGgSU0Gf
gPUXhYMfFxmKtMbBw3qL2pQxTojaLonls976KooLpyOKN9j74lbmMaGKiTG3Q5a6c8Cidybp2qPM
89U2YMTNLpPNbTGPztJ8bUZ9IVfEGddh3dMJPeNjiGQrwb3Se4sklV80Ci/8PcKW5hvAWEgSYfC6
MagkZW18xP0Z0Wqc4Rh3UVUKncrdbNsZbLg4BIQ1g/5P+p4pDsQAudmctwRa6ZQjpLTkoweaEPMD
yfIbzHTqHCEapo8hc/zBEcMaBX6mW7RZJK0CGHyOhHEPRaDxHv3nJUH1syxFive6mJjXVzP+6noG
koWwadtHtrR5jpArUoz0qbH0ZwpIuhZsds/GHqUx1rUOj/EzDjGEkdNB68satn3Ey8nQ6lKCgAYw
qcPkcEu1TkVSkRWdwMFImJIF9bSxNvv3o9eSyNlqp4HRMi3rJ80CqCREMy8zNQtITlJqrXIAo0cb
f+2sv72/4zx1tpcQAGr49ejjNmBRor/ftIYPLk1Hu5+Gyx2mp7z65bxuV07ByyogjnmAZrmGZn+p
WMuDsybg3T81oNovTYPQ/1xLzf2XPKWBFMq8CczeKY801P4tuK5G8v9GEKrF9pUbDKapWp49aGtY
qzvTyPIh8iN6VoE0zRx/p4esGe1mjBr6DsRysWe5EawswqbEGMQzp3v+iSOdZuQRb0w6zVpEq14U
VHSTtdSbWfds3rxEfty/M6d7tv2yKixZ/jkMIfI4ZrV9l40faLW8ICZ1Fz8qPjZMst8nEzZYiXvV
9wRUdNZOdg5DQFc5UoEVNVJh7rkeiBgcxkzlPS+xYNe1GhsFLCADz18R7cY0RoP2qXf4eWveqwnw
aAn6z9a6Ce07mOmf/4vKhKehymCQoAOGnm9/36ZDscv5CR9KsMoKm9JuN07jpJjOr02xEU3BauQk
wKC+gta3erhE5RJEIh8TzIAr8wgE8qs7np8kVq9NYlcK5GiMBdsjVV9tv7wT5d7lE2uEzWZUw8l9
trEoAjtzlRTYX181um8/U8VNpLE+d8joIet4bGBdDj55dILUIreTz69OzH1YzTr+zVEOgr9oYcFp
33/H4J3fdaMCjvYNeE0NUspz4Wguz+sPp4nL4A/4YVMPPuiHSzAm1eunG44GemTzk2LOSNduGt5w
UnFcQ03xLwhd+rKn6R1l/IYDvPHvR+jfKCjkeIS3tFJY/q9Dw1rXRrSGx4f8SGWGlYLAxOwdKrf+
Fc2PO3xaSyailXLvh9rVBCMVODntuHUSE7vWidTreanfdSTN/G9Nal/zOXtLxvN1o3mP6EkgdS3b
7Qk+mzclvPTc4Qd3bBUQ52RTxozRgWkCM1hxV6I1IL+cHNfS1n+46BRo+No4G55kM0R2dmrk8/jK
VZMGtY9UjNa/X56LoKG8KqNJ9+EfLApcVsu5ic40dxS+SOVC8wDaGfU0/7clT+pRjtIHVg035B8F
N7d0M0LfghsX1ACWxfrfCw/0vGrF5v5uuxvYRtMl6/3fHhY50do44xT+2uaBqMQLKfrIV1kvZ2xg
ay5cyxaLHNGhzYECi933+SeIGJveFQgusMqJvyGGeWYOmAyMzrld/LbpRMg/1g+hVz54FaqgMnKd
q3+Gw4w3whJatbq+zsRMgAr59x1MekjTNQfyBzp0B7meSaoduBMgpJvoeN2zj4MKY0ig+Frwo4jh
5GaXfjBkxJr/WOqGDE9ai8nhIuFRTwDI0XlJnlwNTEM2M7Kjqqw6LHFRoFYM08askBM3ITPQfekE
/JbRxccq7NN/jVbiwr5zUOFJzdt3woFbvjgBzoxSVCyKonMc/KIKStbY0474y9e3AfuRepQapwGJ
yIizWk0TBJcnLwFWmcThBGptj/XSEqK793MgCyYMd0VlQ9tRLYID3qd+IjNs8KVqB/fyeBD0SeX3
8OAcegDHpFWz7H2K3wr5/VTCj93psmiHaiF8+/uWVW1CpIwgc1WEFEypNCUgM3SW5Tx+AR+HcmBM
Gx+Z4av5J3tQTivJE/UTXiuX7exaM6RXgfofx5F3FAYDwwJtKNs7xwMHMu9o5nbeYdlhgITzH1ZB
UoBOcz9hg3HiYCbpCeSh+PJrPYmWPZfVXlwN4h7bJjmYypfN//qXiQEgFnPm39E7agDynQyePP7G
5egPFQBfGRuuauLY8WCdqBUxNISBnYDhdgdgB6Rt7hAUfp5zAmulr9JkFR7wzU/Z6e5kMGVD0Q+C
lz84DycGYB73UL1o+vKokqj2C2SzWQwBBOK/jbczprtIeJZkDPrX2JYsXRH4aidJgM+88zC9gMIp
Hx6SfLPsqtU1JZvDvvDrq9ZpzMiwWX2D5Bxjc9c50PBFeFOO7PukK/R7iAisEhjEKJiT0RixUDqA
dnF+WapnSOcY7dsqeWLZD6VNFCYcmudkqjvah/DV4xkZ30YWU4WUyTSoNL+iV5Bsx+Lg4jzXhCmN
R2yRcpjQ4UB6ldCsHCZTXyQx27Of2QgUNabe0qqpUGCC6tkfYpM7504S0z/lpkClBBO0QzgEFN4y
Emyq+0whk2+GbcfCXJHTP2dTOqwxSQLwfwCy5ccHkjd55t/WC75fb3ZyyxJPlAv0GSjppzamUgX3
AQlc5cSGnRlSoSW5197KeOVKAL0OL+9zjk2IbZuSFxyIZ6teFNiL9dnh8qzbTkgCGmj5a1nN5d/m
GS9AYvakgeB6OJXWLBIXtoaJwlL/HU06dETIQ2K+t0qt2lz5Vd7gYyrIIseWfO8ICoUpF1JlgWS8
a13EiZTZ36tstOu915bRM8Pey9UwkQcMj+qHTNvwGmbzxtqnBATr34SmVoYaFBW9Q9ttA6nA+Tla
oy6AsnvXUa1G7AXIvtGo3YA4NbldIzzSik4zovd8IeaErUhQfPOt3L1sM23OgaACPDpifcKLesYp
ZJRLEWQfkefbpQnK5mBgd0IA9f0I5uMt0viNWActsYEMRw5lr146AjDlXI+WvxsW6YSQONwfFKi/
8+GvIcfCXUexWfj+RGIcK43SiCUkNOw7ksMMt2aSzUv3fd1FyuXg2bPIuEwI66ZSnTyS0feACDLg
tT/6WBMUURN0b/BZyka6FQFzyT+Mb6yo3oYG++hmZXFNNBEMeIIsn6qnUd2scJe8v+kVvduKe1Td
GVbAM70W/C3TrdmZ0Pygq/cL5SNILBxKEmoxevSnAjt7OG9CMZ6bHmie1gmCG2s1fXewojQx8trJ
lFMQrBaxjFFam/L1UdTSoRbN/EPL6oJq693Z9efHL/ryjz+CVOGtYwQZz+xxndkRxPj8uTliLSeD
aUgitsxU88XA2zq5oVBtRaABmkE9TKtgHgpz/Ej1req3vgNXs1OoTMwFIppcP9KtkeuTFSSzz15c
rfIJLlCNp75IkurJvW6HouLHxAYGYA9ADSANC5TMB7L2t59eulBgIcKZmvFuFpqxSbvTUhoa4dpY
I+r4aFmzkhWPLxNPRwa9j2qgznGVehsEy/vdn+RpOishcxTWGAcKD4ppcFJeuHaX9KjmxqxhXhbV
vM7sOf1H1x3WCtUWp5DOfH3BBUQI9hqBbn6koBiQxRtT+ZLYC2pUlL6veGYIbKPHfmpXMCQRnV5t
oeSDmzD5JC/3nst0qJOjpta2XLVYBVMQ/nB7AKxKhiSj9xSwyWZC23sGKHWPTnRsnbTCTJCin7Ii
v6e4/aoNRXUp/3Mlo1o+khZHKp1Ejy9uvL5BU+VZOV64w6JshNGzvKugO7M7LDhIsyhNdxP5iPsv
VsLYtWyit5gtDCFYm8B32bNGkyX5iir4nlaw1IdUINhNQmo6DC/2kvph1C+8H5ihuVBThsW2+Z4H
4p1ctmyjBOdcbBmBLZEau2OCxz86eKsEvN0PKgr/cMs170aHv7FGmRt0DAqhqzXztAjd4CJmne5x
l7alAVJlYI1ZZSIHso8Ev75pbPmmq9uV79YemvcDgOpc/JkDtHHJGPto4D90vpyAz87JBDtDdO0X
aF/UVwWMcezRYcXXLffWIZtCECc7Zb1KzXwXkqZ32s3RN66Su0UFB3v64ybD3CirAmcQtLk47o7u
8F3DbsNvJv3Ah39Yc1ssuyiMqMk4QMw6p96KOdg4WUcqnrULaUe60kyjG3Jt4sFeHG0xI5dF1Y73
1Tbxx65+fI+Wkqx5aG5dhaFuhWeuduW+zpPkY07mAEFoWqnTLhEERce48zpRuhyVAH9NAsfhGfAM
Ioqj81h2/to1t/oGfXM5YQJQgUNGl1UE9cO5J77TmDeaSkwHEEu8TysWnSiO2irV6U4wBPS640n8
mfo1ZhrfQcMOnjg7P/QTN/JyzPwyH46kNrL+/Ej7OEGVMkEnuw52AKXdBOREYxBrDHhBFb5VKZ3B
tl92fw+IoBkNbR6vPjT7b8T5QhkugBMSbyCJPbhALJDLRuK/tI1/B6eJtEwf7FyLzN/+2ycZPMTJ
tz2us8PCPKu8IDzhBY2nzztHCgmpCwWtM6RQa6jUCtsW3jcchIHpHboHRVUQPbJOanmBsTxlQLRc
pSSuC2GGazaRTl3qCtKLpOmO+pVDb1ZkR/wEUnvlrZU2AS68NCc+6k/I53o8UbgZR1qbYnAnpksD
2YzVUzZihSzRjGMAz1eryHXmnAK3lTiCY0ysfGezCNRmXQ0xOqd/RsFhNBNhZ1QVunmN1kVWxcdZ
QflJbEDTAqaOGTtz+BHR0fMHqNtvQurlkv9+JA52WZ6XDzhrYsr12QV4RbQ6Rc5DioU8xdopTV1b
DAe/zuVbgPQpD2KImGt7qjlFlaxD439/kFyIJoDx7GFYXUgJ7Xo2dYqnKZMrOAEscLTEA4QldQwQ
aGN/CRYW9Kp/KksiJ578RJSa2XGfQVSd+c6+guSx5vgiG6clzfuj46EayyioxSsN0N6uYMXB3iJs
ujd5LHPk+jSAeOPxEM49/1ZLQr7s4451NQXqUC6YXBCzexRVrFtUaKf9xlYc2NkVecXxxhYsNhCe
hxLUApnUihbyzKlDSJ/IHmAvdWNfUCVhRNGFdgrHndDGFX4oIS4uITMqCKwMv+3CJv9JjuO805mE
gS+Ylx1KGNErKYz8aadgsvlx98WgQEXSpnQwLhls9lYdmAeIFADd8PrrJzUw6t6SkC9wu7pDE8L3
hTLGztf+BkmBHiun/0i+LUQsuvoRLYUIckf9VmHPg4ZsEOmk8/zGfo3rpiBBTNfWyjJ+EZ6PBttG
Rkx8P7Av1YfOpk8bw774AuewkolPbSZD/Xwm+BJx3NAB4s7nUcIYeRSeU2+OsIoHlSx/4EONxEbw
ccPt/wLKiTNg4a5pw0U4EtEX8GcXjbPCsa7+Y0ZZ26xVIdkITq3BUorh9DL1OgLiBsixf+/fI0Xf
RB7wPZAxSPwxTlw/lq9MZnTSFdFJHGpsuj0xZn82Xsivjnmg8+zZO71kaTpWtdOlXHbwquIzo97S
A+PHe2ofMoL77Dk3CU9z5qrTaXZ0I5SGcoxSWUVyD+OefdKg6SM17juDjiVRouVrNAFqCF7cYthJ
FK0Ob6qWI3dXXQ/SzcDvW8d2On/wobRr51OciYzWPZ3Hvga3PnO12y8a/9fs45bYf1E8EvbVxgAd
/mMkQYhheaB4QwXjifmUFULLmC44wCcU2MelAvAu11452biIK/bJYuj1C5ErXm34gHjXvCqEEinE
TaD8FPhAYByfM4lQX7EmYwFT6zSQaiOeN6LWq/NWkqsGyNH6RNZ6NgLZ0/CidZkE0JFp4Yg0G1EG
wJMz7u82Oaf6nL3A7IJbi9FYLWV7FFzewDUhzakSNsNIrHgQZg8M2M2ZBFoMYcKnvRI7zZxSqUsB
FpeeNFHmEj0BOFfvyRbpLKqiSKQl68SlZOYIpqh2r5eg9cpmmnNzINhgQk/quk3A7l2Cbl2v0WQ6
/TJ/u+q/8vgStdeyGbihCJksYsn5cgzpsyIgJLTKDD/kwE+78Wuj3hup47Z9aB66m98EgoPPkKss
trRAQzwnZyjnkpRhMw/e9fL3gqQHwWweB3xG4T5BLHLaDx8LrCNc37ZZ1KsVvhlfSWG3rcB7kF8E
YoTUM2HVkIR5v4ZWtWz6iJzqqiFjDc82kV7qECLX+wVpse2FVoR95LLUGhXPtzG2R1wFIg89LgHl
xFkKHJTP0bTBP9Qa7dh4VUB1k9tBV3EJYqqYqDTY/AcM5/fD5zeeh6bvxtpKyzQ1imbHKKkFE9Gk
WnOgpD6apV+By0zeeYErIeyNudyIDas71edDNaA8kC+1UQFtKmPYCukQx6olp+o3CnRC715C1qAp
DuT984FyrVbX7GZQ+6QQb/3j5YCaCutnf2j+tEjyc3iKZMKpbp7LvXN0Lj58yOxxfJY7yfz1WvEP
5TMUhiMf5j5Rhn5lMtX5tNHzk6yvdskDvbxzGCXA9Ac3Xime1oecQiBTQ7DtDG/twMRcxSnFZ6IM
p6ApRJr8hThBtl2QK4iSPcDtp3KCWBU4o3PsmfJGRpE47SyxlZS4Qm1ZUV5CpKwXjrvvwV92zlLf
4HiXE/Pr1XzToAHFp1zKPKMzQPbA7fQqp6E74WJ2h5+I6/2yS/BDYMoriQBSBLSTNZUmcaFyyfr7
dwyV5nR6BYWAectSESzdOI5qBDitTdavs1+SkI5oBtIhUeDH8Ag+1x7NP/TQEEzneyPPhEaSZOvg
ILChYXYr36qlKTwUtUUgxJwH33vBl8SoUm+kG6lXSdQ3i8j+7Hechp8YsCpBjExOMUodOSmFbF9v
q0c9ILebI8Z2eBmrftru+95PdM3kwKtfIFB+oOapm8eF22qEotQwpgEs74ChgWCTHwQewK5CEy4d
wK/8b+Mba3ixqBhdPEi+EgdZ4yE07JaxMjNh7dOgIJXxBB4GDoDhNUWm5fWJrtTnm8T1LpVgUF7V
wDrGDDpKHegdoVQNGooJF/Q/UkM7/CY+EUAQAQfTAtcNb8dFc1v4aISXr91GajIs780AofGl1Pqi
3WTNk2JDXWkXhyZruX+IgmqMSyHB/HE4q+TahrJ1fufZV76G6cvEyMdDBWPaRRuozYX7korYVdXX
mC+XHvjN3wckmFh1Vwya9zMV+qlK6I36xQccIufWn9YpQm9nDLQoc5ruEMo/859KYyQShAhmis+X
RmsIkHbMo0XrVMe8l+sAFtOBCz5etSnZAbQzaM310lxdrDzSaTrU4IHWM3LwD0WOISnM1h0/mqp/
iAuwxPAdkS/fJdOuTC4/icW24rCpN4yuaXnL67+AGabXpp+GJv7weHmOoJcn/aBqAsxDvjkYn9rP
8FxOECvihmUxlpUUdzt+Q0tr9msvfY0Nw9G0j4H2b1D+4YfXQQqfMxevncgT1IstqujXWYbsiq6n
fiYqN5JsSmMwPRB59IVKkAbTGkfz/ZzfIIPhMdBv7VlqSLK62bFKT/PXeLIOtZSplBW9OUJJJD8S
+FDYRYN4w5h44rSAQ5hOTF2pyc7Oo4qcol6Z9OBn+7NyIzx9o7DEQqyUuVVZObfVUyFXeO0nSGUX
Q+ngdxkIa5+fhYz/Bb0uqb5hDtjSZGRJzkW0X2NRG5mdBa4Dx55YitfVDpXoeeAjMBqaOie6yCeL
ZVEEdcdaxWfDdcxRKLf0GIOgLO1JhiooQs38NjCnEELjs3JvmKJ6126mfT2I0n7hFVMMtB6tF9Wv
JZtmqk2nifLBZZV/VRoNBsZRD1J8PxLFEQx8rCj8NdQRKwQVoKfNtSIyiNhlAT2jW6O9zVAjcXbD
dC/vypW0Yc309RzxjTV6yRGAgtdt5Rvhxvc17k6tuFXY1LGf24NUA7tJRmstzVkZPMmd9A8lQ7zl
vYnGIFmwmYDKIGZ+oeDQWOJkccH0xdjje09wGJHNFttl09+dAcQd5EOOG3g6+iAfhOuR32TLvkZm
VNoOGBQVTRBXoT0Dc1jGGIZAOx0JwWfbiCOW8mEGcnc0DRig1pCq7dD3AXbw7Kgcq5Yto1vtEYBC
SOMvrkNedJTB1eyftq4lkEIp7kiwKeJFDicTNcAG0E3DyDPNv3M6XGZidwiWGVbARmV3OBGGDnxS
nPdwzyOJoiIfNPKPObuJL0/tlhHM4fK9T7fmzoqJ/4bzaCw7H4NDOGV1/bZMqXGTZMlqC5OXe0Vl
k63DzzIqp/Rp3PWZUFh5nhulgU3DFUxBA4mYqDxnd2K+y0QKv6cUGCQvQAUKewAZnEptoSZXWc3a
m2Z+t0Nx8HMjIlsTDpQwVhfydd7vX4/U0EDly0ZsQZVzf2Y8ObIbYfdDabyynce5mAXVauZAun64
AnQFcRLmTtaUlmrD5A8BnyUgqGx3xiLu+Pv2iRfN9jcH9AcBEfJKkoVpnMakiCr2tJgE8cSnZ6Ge
pZPNHNsscaCaatyXwg0hkCXpVFmyfXo3cz9+++KkgdTZyeoXEWeK1GiNF+wGAaLAXlPV3GQHd77H
+eRfXtKE3wvalcZW1G0OHE9rYhUMbEJvnM3FcfLJl4wxFSSm6t2pbRlXRCxll4+GpBajzeVcWwFA
/Sw9xtoCjrh70M6mjfHdNXlVpk++vvAygobP7n2/3JR+atfBFyNv4p6cq1TGi6NVtshI2sJKrhHV
4VXS9+mRuBsGhmtX755JZ6J7mD2/9m6bDElFmDhkdXK3/FE/AN6huObsoy8SRlgq2QLKiIC9Z7EY
KOJvCcb2jbCW8bw6SZh5LqLF5u7kd68g6mFgMdsy3fiY4DlgVD/SW9onyHjX6TwSPhGW47mnVkZO
OJupwM1yF8FYpcqj8+kiQJTRl0bao0yHnh/ppD95ex2xVH6cL5wU2mv71QQ8m3tp6GowVopNsLqS
QwaI/uicdwjwiqQ7oCvPsrw5+VFO0fbzWKyrkUuHPLMzeJROU8eRtmXnILMTnPGqmWoeIOmP4Zpr
SfkP5IPlRj/J2C8dYoteZhDYwk3Yiaet8M9iNUcSh43eNDt3sEa4o42bi85tIjJm40a8QQQDUv6s
YFxgtIVbTQXkb0lXUWKAU8t/tK0KVIu/hW5m9CiRaauLSj5sGcTqZwKJ/hqG1XtV3RFb8GfPqHW3
ZM9Lbiu8eQ2HTxVyUC+Q+4e+E/6VeoViCjSvjEGqxToHFKfC/euk2CP/4AvXr4hPMvqEGZusBDI+
lmt0Gj9hTJ3efY3USPOBoD35ZC2R9nlobrfqa/lLs90EAIZ9o+r2Jg2g78sOBtkvmpF8kSf++nFW
/EvsKPTfpT4nNed8LZ2sYNSJd5QMRTHyqd2BF0ESsL8RcOBM9H1XTbDP+ttFGV7vS28AOflRHQ9l
/KUdiZagrGVYX6a326lFuKk9uubXCVJGi4/y7X6xki9dqriARG1g/P8Way4wwyHVqLfSSFupcqkL
eiUHyC4V4cxI1eFKDza3f53IKW+mJB3QkXMHQX8q2VsYzGsQedjcvuDhUG0hEv1kUxhJezOwgHWJ
I1boMC1843I8HvhN5e6WXlJZiU9EFyEBljGav1AK4OQgctz27rGLNI+EzTwpzUKyi0iLuya3kIe5
FYa4J7Z7blpSiDnIo5F1gBT//E3dIsRcjpsVjnfOzdL4f/Vx357aTT8Qv8dfEaRL/he8CLF9w4rU
KuVNnh6hFDfdlZ1yHyW9n2qxmWMKiMR4F55helrjklkAdHqjrjXdI9KUrKuAq9J+0NSzxC9aNqJv
4orncF9tA5DDOtbVcMeefkTvfWuBwA92ld80H7PAqsFeR4WbD0PVLRNV46j0T/dihm3EDayZo8qG
OvXCpzEZ6T7vpTzzMULaOUACwTZylCeZR0+/e3fE687s6rzSK93/ZsHnn90lh3LUtFXAIcV11K6r
JGubI85qk6zgww5tOSmLDkJokklS+Et0T0cDrCcMnkPAVwcgu6llYNY4dmOkmQ3q30i4t+idzF3r
OA5urWUTzhiV9whXaIVmNouVPoCdeKPS2FVQbVNr3M4zG/zf7ok/+rnx3J5bd9r8rXKkh3jz82PL
zFAP2WVMKGBIn0ZctynjutcUGygdJYMcsZYhB30VDQy1ZSFCLLGRWdfJjfmim3jsZsoemt4FCfvv
7bZDbcBIm6NiA8Djl3m5P2rnL5Te9LK4p7x71HAHV/6J0j/Td1CnQrVD9g4aw76BqSiBcxebOR47
0nRLkmFT+j1+PfAk6QLFM/krM802ZMZWu9hfpAm2+QFwsD7WGmqkbrP+XWSFpLuNSXFkh+RZ6Els
cmseaimZwOUbcuCRfdTCMMOmfMBa1BPJxAj78fpFFIx7Cnrcs1PtKgwzTMHcYn8zqSONjuyDoA2w
ix84VNNYOnIovgr16Ww19pRXnWP0zcfE3Bxp22Zf4WodUZ7ZxuqSB9BdjpUus627GVhXu3t/sC6O
sHuT8Nh71nYPbEeCTmvJ1fX8fI0+oyXpAsqGlycv0hcF/0cNoO9S/tAmyiP5FrOeFEeYQF7CqQhj
vhvd0RLQxFHhDI6mWgrcdOTGdpSodxVF+Wa0CPnV/VZ2+87thkS5epAky3vAXl7PMYFc8hJiWj5u
unglIHXo3PrbIKmClhOD/ryvjgR8Dh5Hok13gf8rn9sFK2O9AWPpAYo5nBjeQldh7agt6nBgJ+PR
/8c516h0rN0tf1ErT/38f0/+pmBtLN8Xc6Q2iVXWtIp6hOf9TF73Ky8ExUVrFp7yNBUBnrxx3Ak3
LFArnIrv3W2NySYnP1ADdfAi+Gym4OXeocf7I9SaUE2t9Mo47xc1L7b6MbJVadDVfo3Xy+cgzEp+
9gZ1ZWF6zef3BDqGSc+Mb5+RfCPsCDt68Ljj7YG05b2ACaJOy0KEiZAYDLJzv24O8BZO8h/oSDxA
quVbglpobdI/tgnd6MB1IqRrSISUvayG0Ls8zdEN1JmvfvOY022AeHbAnJpTaEgZSEMYAh9Afsn6
TWMjmghEbNEa9YNokBbm7JcNLoNllfR46uWONYSZxBz5GMyv3y4T+O8f7r5bQy1uekab9WPJ7yXl
e/qZGlUQmj35yar3KaLHigM3xOsEmtGnu+bvGktTbZoFp/fdxotCMI8HrRkjJNTBu/Ac+gBNMaHN
BK6L0jzV07lULdAWW+21pQEvMDCcTB52StRAAlqEVxAu+K/XD6KqPRfGgHwORuC4FLDXrFPGElbq
BelBji/M9vT4rx3d+Qwng4u1DmMcRwAl0KSI+cPSB4U8VUil41NyFCCNo/NK+yfSkZ5U+Uav46Bh
OjkqdSU2Wzrc6htW2+skog8dJz8cwvLuIV2BThfqMO8KTIuBGthieDziTesius3VL1jd3Jq3/MA6
J2Csim+HGeSaFi/inpQgEUprNEVt6uweOxZaFRhIY8C6+RvXF+qFVRllER/59nlHrhT6MCUciFk5
je+WLVT5qsjmSmL58p0x8xKCBtdtZw75ukPcTjTgFqftq6rkEv5anBsedkFsUTz9llbUu5reZv7T
5VXqY+PF7/TngFK5BtenH47M4d1EsmcmimVkTS+O1eaIhp5gYgdBsapv2+HPrC6iZYRc4mtfpMW4
Boh2n698c9N6ZjtEs5qvMwtiTfmM0K7jgmicTE2RtKVE2SB2298DkgkkUY2enA+dET2200kULK7N
Ht1K5u++g7MJ8QmKmBOjc16Q/ShJfyeaWEGolv/dHJFgXHYWWMHcc0jk59fAWipiURZWqb16ndUN
z73mnkHTiuQzNELLkrZ6ieYcSDC2QMq4zAopssrnZQGLu+ufxPy8cTuNf9mqw8m/dh09NOuP13yD
uA4E4obEt1uXOssYWuhsJ8NILkSDntWbuZG3zP0ig9CjNk1x6YUzBqeJuRfFNrhfxe8YOtF0u9lO
DzJ4nd7UuKtHsC+v3mHavtu53DOTWkVUoStN+xPLypU3F33VhxVnF+GNyExEajKvFoC73KMTG4Ku
F3fKJX3CPgeA8N8ZhinTkRZnNKoo75xppzWgdGE7rArR8c8EMnQJZBuVMUZPpEGbYdqwfCPnoQ5k
a2nxGfsGOh6nu/rGSyIrfeWjLPOXjgnvHl4GJwrGws2Aod46H0C6pY4mZFyPD+nOFKsAm/0AFc0f
gBx+ueijTW6KmRSSNtS5DOgJ3rDWa8GDfXrk7Hzs63DjtgrIQeY26yGxoDyfE+wTnQYhX17Kifbh
n8UbBQbBpWQVO1iz/EjypPzhZlLGltsqtOVCMBQKakDwf6MCWLQaH43RxDuiYrxJeSicojhwHpPN
/Fy+il5vasWCro4x38euEwc4Wl5QD6RFQDJ/5cT0CNAccd/icz+FdfCvX0JfhmHugBVl4Zoiv1ZT
M3oiXF1GIHPF9RByrGoig1clD5swKG+OS4vy9N8LbxETGSGt5OsP5gfD92STq4LrH8RcK547RBa2
P5m3DqkvtNYt8I0uUYCXIHTRtTcD6uh3v3Rk6gF2WcOJecr9gb7w+G2SB+9n4/tzhwAmzar3uFz6
UO69iQZYe9kDxT57MKz8Mvl5i2Qq2D4a7qH3g4DKJ5hO7zBSRFjCggEkwqD+tm8TaIvai7Y43IE7
+uiFIOloOegBuUtUMPXrI4nsWXhPIRyG1WEVACqlLoCKG84de9pvI3koPbbJQOlBVm7TrhyP1j23
H8h9HCZr+WDMuzjW6BfoXTAtP9lbY13i0Sm1Oj1pketv34U9Z9ttxhGyj9XY/CNEZ1pOUOGB1YW3
NWddtMcP0u5shvwj98EKQGakFp983Fa6ta+xUniL1WP4ish8E+5pmncuZtbvzOzkIW1FFfjgXF9x
bYNHTM2A9dst2VIbgiASCI0eKmSbOc6gWdLwZdiaCm8ERzmNb0CR/aygp25GH/ytU9bGHUcDO1tP
bYUm/bFwxm2ZMGT7/j2P3ny5xRyQaaNoO7XksgT8lF00DJAkNw9ltKrsYCr5tunKorMP/PiC2MiL
+VpBDQfgI/XZ5gnbtz8C0vhdT+m2uTTsWCn1cZWK9SUga/ipiZ0vTHCCuGlbLoF7TVbK9WrfFLW9
L+vsifTQiR5zhYGC9UFXnM+TKxlVTJLsWOaOzUEpWn5TZWTQuQZSz86SU+Tx5aind9nMADFvyIQN
x3vHMoDHrHfcrn0rEvEprybB79dOiBYAAj9q1NMi8ynNiM0X67L+Xi35BuWRyJfPyopF2d+fgn+r
avpzYuxlKiTinK4Y8EBQkRXH7kwK8JQX4WTsU6L4Q4bxBzPoWBNe+J3+VSPKgB+h2lUq5TkDGwam
Cou/8O6PqYxGEQEp/Pe1gA6RrZF1lj2XkJLc1wbife3DvWFQbmDAZSi00Xj6U7ZxAPiZtdi+wCah
XgBhp/3B/RocbFCKVPzaPfCzlbdWS0ihxvCJzfhRQa4qBxdOeRBfdyxWhkNdFjYoZZFC6piI7Nta
op2aw9LDj1aOSiPFblDKG4iT/oRi5y7iQ6xNVfY33+oKoJd3LG28S214JUoDy3OL8e94KE59Vq5E
pa3jVs0RRYwZ0Uv9XV51AweSA/6Oq3msdfrVdM0p7LcEtpbm3HVIi2FMFuembP3jDBAv5X/x27vp
1e1hkkNta3UkEK6TIbiySIz3NO9CV52wdPvxd36vdR6DftUxQyoWuH7I42LNvO35XtDPVjopouxQ
FbxbX2J2g0/D8DvjlxXtZhbQot8srxJTr6W9coTM7WHGQ7VM4l6vMNTPSrRkNi+zVEKCni2GND4d
bcS62SdnafzLKwyDd1lCgS8d6prRjiOGY2PPbsQNVDbFhgUswPvFwfCpLG8rAXAGNVRtKQ89I4HI
AfMv/HEOP0bq+6m7/+5i5LGrgUcpa52XJwcs0mOMlsrfMqxvf+mQZQuY572QgUcufizomXt7y//K
WfvLePEFE5RZ4p9vkbexYdhyRZDePlzOVn8CVz9848V9wdkTOxyb64+7jWF+ddJ0mXqeef/KP3pm
bXJ6Je7WjUTJjcLlc93n4kQEEwrg12kNm24cM7q3IdFgorR+uyZn7+tVZve4JDd0fNTb9SylFkuA
qWh7v220F6xWBXD2WGhfxoiqflbFF1VO+8cYONuaVqoW9X2esjYMY4bivcRqImg+BcRoRhoNqOTD
+yARr2EuR1lY323L8GebfoIkdOOWni1wYfpoGRmHXr6MD+HgDsOoY2hqrgNy5vOyPEy8coEGDDvX
o8AetVD9HwXJnB2mbfLhQ3E8ltE7cFNpAeP1+nJm0+EWf2/he2kT5IaIcP0OfmboKmAPv9vhQ9mb
7gwDrVWGsaCCEoPsfUDm6bL9LyQlkAUpG44rh0vXX28fazDzk2p1RY1a/qkUToNO/V2JODVn/tiS
7S93lsM7t6q5l/TDe/0ut3gIf/YcS5n6yvZJjwmCPf4uzHtHKLXQ1EEU/+tXAI5bFbH1LhQ5hwFD
RwOMSP3+nkIIxWaPEHCJxlhZaANlJh6nMCvkGwWuXGzvm0xO5STbjlGEPqywxdmleg4kmdGUJvVs
f+ZXwrIqdU2iAtCVavPwpJC5anXrpl5QLXCRe62P6zbi/OG5QXEFfzCYAdw91bud4LdAoLiqD+pH
43bM8Ll4omb3Qnr/4fyLNFe0NXW3Ju2IwqXjEC9UTkpd9ob+MEtOejSnUc37qay/7OMi6+KWPLaI
Cg1LZRorpYofSa/d+dE+3fxEBRiFSiSEClty2+xv3m4iqODmHDa8UZ5UuGIfJzCHfCUZtWfZdz9I
sQ25Oxy2qNbbwL0dsYVaFypx9wQdrnUiKo85axv7Wx9Jh7wgQLdTLxCg5DWLfMVYsZGdaSKF9F+e
GXNUFMAkS8jFrc2HrFJC0MEJVKoG3hZ5qF0RhL9qQ/Md7acrF0/as3QGr6xm/jOPWJlfX0jDDChd
u1gnNzSYckiC2GKrTl0ERFtmOKgWGnpccZ6TPuFemMYOMpQES3UCzpwB30UESKjIDIQAfFVNgOe8
v6DLrcpJMSgE+0Xt196srUZyYlj2kHDz9ub1Z7g5hbQ9A8XDEsU/6uCpqllaPbR6QBdQimjG+/XW
9mJ68owgCOpCVC3BP/qt90VgyEEYv3v8jzj7hDXG1Q6sOMYvPedQqXV49sJ+/EqeATt7jrCcopD6
PqwVu2CsEn5vaS/i+qM/0WEQFeQY/os4TC7rmVIHBIQc2/3U73Zz9W6UJpKHEfhnbAexL5XNa04L
rxYSPJtu2egsYmoYVpesHOKfALreVltu0MnSb5e96datQesxUULvN2d8/ca7OhiZb99Q3l4jG5y4
CPpluoIuS/8j+2BEuVDyl8u4EhUj2o3ZBFfIxMIhqetsIyBi3EE/nxGVQYgr4pVahZAdrMWnWEfH
pfhcFZHvjZDGMNdTfT/hf8Kihq53jxFL7oraSDukg/sJET4j/eTM5BH2vL7tx3ZB2uSFj7rPDifA
oT+H4HKWcvs6JxIkRhhhSX8s8Hw5FuOd0upa5QVv8d/2rPm7ZBkp86GmcAAfDz296VjEAYgSyTVt
LEqzwhXU75K1gPTd+OfFDmmumSZPsE5eUVw7jeV9p9qK44A7y4NJgu4He6+D4JNrqnUdaOPnQ4jl
DlrpIubE/l4ht/VqLScuOL3kxLvTirywukz8Uk+66dr65ykKbMiaHr7Ckun/h6dH7tmJHsZ01Nfk
FVjpAsc6UFdyVxx4QmAYDu7tMMV6uo5CDeV6J7bEyJpUk+yFT6W1eKBD1JtEQj5BYu0MpYTem4DV
dFoHQMvdyOzoycmVUMZKCrDpjO4o54sJ69hkN7FJ+dEeS45fR93GOHb6vRwJ6UMtq/DQSGxvbFrj
SpnBExtXUVgvDu1DroyciJKmJpnRyzL56jaJq9sntMvvmxEY7xMzv6TDIAnT++bd2uXo+NaK7mty
vadRVT35YhyAYtf7GvK7dmSaVXPrRk2yZswk6oslkyntw+u6Ez+knk2d9i+2uHWeqoha5KqCUY1v
oXJEulsoGC/MuDDhbSzX318BZBwzLK7mABjHJDZ0BwWXL6LvvVO8On5LsaRyNKjvVGypEOi9iIAW
1BT3Kw+R6kUQgWViWrrd1XBqtmQUWWsvV7aAc7VIuMQ0nDONIyPbPykZ5l7R7JMHocE0CjzvHhUm
HjSeBShBocMY6T23wi3rFvcmsNOUUrIL+VyKIWQkek58OSM2R+5GVpzyyvAM6hmbICR3D64cjdfl
UnBUGC5evUDu7ZAIsYDKyF0mXYdW3LNxn0U3I2sU37UVtJZv0wjV3x1vst3BxswyqllCWQ8aWYQ6
n7ulacVp6RhJnVv1R07+emhUPIrBdZVxCHdaP+fglHc0K6hwDSgn1HdyWBVTPHERC6jbD20IB2qJ
iHCx8RSFv1gwgtqzaITvC7M5kSJAAcDtJWK2ixN9QF8YQ1XHNASSgnAr0+nWc8hgfdb3RYaeT4jf
kcKG7NmvFDBigkhMj5bjBcbvpen8EcVlf/SjR9cQ6PV9XUvU/ZQQFWpfOj9Y04+zRXtVEvkTQEjH
9jYZ65gWYbX0o3Yl68JE7l19sccHvuYaKDagvZAfNmbo1km8aVVm1Co5bdwNKjs3vq6Mb1B6tH7g
PywkDVyutOgqtlLDWjtyzMzKswl183qhdRtO3ny4pQac3c23oa2EiCVobsz6K5hJht1/wwdFC+57
dWd5wcWq1Ap9oqPggfUJY9jCFa0GvCcXBUa6yJGTUdCCZSO39jKNh5/xxrYGex7UFDQxW6kFvWl2
PNk3ViNDubkok/e1PeiGV3KaFe0z4Rh7vwd7CNFo21hkWYxg1sVenamJ5eyh8bYoin5DrJBG+gEt
hjPBAkGg4eT8ua8MjyM4vaVZ2smOTLiU4avGM0Jqug4GVbIeOrBuEbzNv9MEWoNl+dzIrQHajBke
kihVbimvNtcep41hNryeyar2Sx1hjZgjHu40P/q/HRe05g3L5uI77cVuZKs=
`pragma protect end_protected
